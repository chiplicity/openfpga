magic
tech sky130A
magscale 1 2
timestamp 1606227342
<< locali >>
rect 10057 19159 10091 19261
rect 13311 18785 13461 18819
rect 6101 18071 6135 18309
rect 15669 18275 15703 18377
rect 9873 18071 9907 18173
rect 4077 17119 4111 17221
rect 10057 17051 10091 17221
rect 10977 17187 11011 17289
rect 19809 17187 19843 17289
rect 7757 16575 7791 16745
rect 17877 15895 17911 16133
rect 3801 15351 3835 15589
rect 18705 15419 18739 15589
rect 9689 15011 9723 15113
rect 13277 14807 13311 15113
rect 17049 15011 17083 15113
rect 10517 14399 10551 14569
rect 15301 13243 15335 13345
rect 9045 12699 9079 12801
rect 15025 11611 15059 11781
rect 16037 11543 16071 11713
rect 14657 11135 14691 11305
rect 13921 10591 13955 10761
rect 14013 10591 14047 10693
rect 11621 9027 11655 9129
rect 17785 8891 17819 9129
rect 14231 7497 14323 7531
rect 6653 7191 6687 7497
rect 13277 7259 13311 7497
rect 13737 7259 13771 7429
rect 14289 7327 14323 7497
rect 14197 7191 14231 7293
rect 8861 6103 8895 6273
rect 12265 5015 12299 5253
rect 19257 5015 19291 5321
rect 10609 4471 10643 4573
rect 13093 4471 13127 4641
rect 3801 3383 3835 3553
rect 8217 3383 8251 3621
rect 17693 3519 17727 3621
rect 7849 2295 7883 2397
rect 10793 2363 10827 2601
<< viali >>
rect 1961 20009 1995 20043
rect 3065 20009 3099 20043
rect 3617 20009 3651 20043
rect 7941 20009 7975 20043
rect 8493 20009 8527 20043
rect 9781 20009 9815 20043
rect 13093 20009 13127 20043
rect 18981 20009 19015 20043
rect 19533 20009 19567 20043
rect 4712 19941 4746 19975
rect 11989 19941 12023 19975
rect 16313 19941 16347 19975
rect 1777 19873 1811 19907
rect 2329 19873 2363 19907
rect 2881 19873 2915 19907
rect 3433 19873 3467 19907
rect 6101 19873 6135 19907
rect 6929 19873 6963 19907
rect 7849 19873 7883 19907
rect 8861 19873 8895 19907
rect 10149 19873 10183 19907
rect 10793 19873 10827 19907
rect 11897 19873 11931 19907
rect 13461 19873 13495 19907
rect 14473 19873 14507 19907
rect 15485 19873 15519 19907
rect 16037 19873 16071 19907
rect 16773 19873 16807 19907
rect 17693 19873 17727 19907
rect 18797 19873 18831 19907
rect 19349 19873 19383 19907
rect 20269 19873 20303 19907
rect 4445 19805 4479 19839
rect 6377 19805 6411 19839
rect 8125 19805 8159 19839
rect 8953 19805 8987 19839
rect 9137 19805 9171 19839
rect 10241 19805 10275 19839
rect 10425 19805 10459 19839
rect 10977 19805 11011 19839
rect 12173 19805 12207 19839
rect 12633 19805 12667 19839
rect 13553 19805 13587 19839
rect 13737 19805 13771 19839
rect 14565 19805 14599 19839
rect 14657 19805 14691 19839
rect 17049 19805 17083 19839
rect 20361 19805 20395 19839
rect 20453 19805 20487 19839
rect 2513 19737 2547 19771
rect 7481 19737 7515 19771
rect 15669 19737 15703 19771
rect 5825 19669 5859 19703
rect 7113 19669 7147 19703
rect 11529 19669 11563 19703
rect 14105 19669 14139 19703
rect 17877 19669 17911 19703
rect 19901 19669 19935 19703
rect 3065 19465 3099 19499
rect 8217 19465 8251 19499
rect 13829 19465 13863 19499
rect 19349 19465 19383 19499
rect 10333 19397 10367 19431
rect 4353 19329 4387 19363
rect 14657 19329 14691 19363
rect 15761 19329 15795 19363
rect 17233 19329 17267 19363
rect 20361 19329 20395 19363
rect 1777 19261 1811 19295
rect 2329 19261 2363 19295
rect 2881 19261 2915 19295
rect 4721 19261 4755 19295
rect 4988 19261 5022 19295
rect 6837 19261 6871 19295
rect 7104 19261 7138 19295
rect 8493 19261 8527 19295
rect 10057 19261 10091 19295
rect 10149 19261 10183 19295
rect 10701 19261 10735 19295
rect 12449 19261 12483 19295
rect 14473 19261 14507 19295
rect 14565 19261 14599 19295
rect 15485 19261 15519 19295
rect 16129 19261 16163 19295
rect 17049 19261 17083 19295
rect 18061 19261 18095 19295
rect 18429 19261 18463 19295
rect 19165 19261 19199 19295
rect 20729 19261 20763 19295
rect 8760 19193 8794 19227
rect 10968 19193 11002 19227
rect 12694 19193 12728 19227
rect 16405 19193 16439 19227
rect 18981 19193 19015 19227
rect 1961 19125 1995 19159
rect 2513 19125 2547 19159
rect 3709 19125 3743 19159
rect 4077 19125 4111 19159
rect 4169 19125 4203 19159
rect 6101 19125 6135 19159
rect 9873 19125 9907 19159
rect 10057 19125 10091 19159
rect 12081 19125 12115 19159
rect 14105 19125 14139 19159
rect 15117 19125 15151 19159
rect 15577 19125 15611 19159
rect 18245 19125 18279 19159
rect 18613 19125 18647 19159
rect 19717 19125 19751 19159
rect 20085 19125 20119 19159
rect 20177 19125 20211 19159
rect 20913 19125 20947 19159
rect 1777 18921 1811 18955
rect 3433 18921 3467 18955
rect 4721 18921 4755 18955
rect 6101 18921 6135 18955
rect 8125 18921 8159 18955
rect 8585 18921 8619 18955
rect 11437 18921 11471 18955
rect 16681 18921 16715 18955
rect 18613 18921 18647 18955
rect 19441 18921 19475 18955
rect 2421 18853 2455 18887
rect 5089 18853 5123 18887
rect 10324 18853 10358 18887
rect 12173 18853 12207 18887
rect 13093 18853 13127 18887
rect 13809 18853 13843 18887
rect 17785 18853 17819 18887
rect 1593 18785 1627 18819
rect 2145 18785 2179 18819
rect 3341 18785 3375 18819
rect 4077 18785 4111 18819
rect 5181 18785 5215 18819
rect 6745 18785 6779 18819
rect 7012 18785 7046 18819
rect 8953 18785 8987 18819
rect 12081 18785 12115 18819
rect 12817 18785 12851 18819
rect 13277 18785 13311 18819
rect 13461 18785 13495 18819
rect 15669 18785 15703 18819
rect 17877 18785 17911 18819
rect 18429 18785 18463 18819
rect 19257 18785 19291 18819
rect 20177 18785 20211 18819
rect 3525 18717 3559 18751
rect 5365 18717 5399 18751
rect 6193 18717 6227 18751
rect 6377 18717 6411 18751
rect 9045 18717 9079 18751
rect 9137 18717 9171 18751
rect 10057 18717 10091 18751
rect 12265 18717 12299 18751
rect 13553 18717 13587 18751
rect 15761 18717 15795 18751
rect 15945 18717 15979 18751
rect 16773 18717 16807 18751
rect 16865 18717 16899 18751
rect 17969 18717 18003 18751
rect 20269 18717 20303 18751
rect 20361 18717 20395 18751
rect 4261 18649 4295 18683
rect 11713 18649 11747 18683
rect 2973 18581 3007 18615
rect 4537 18581 4571 18615
rect 5733 18581 5767 18615
rect 14933 18581 14967 18615
rect 15301 18581 15335 18615
rect 16313 18581 16347 18615
rect 17417 18581 17451 18615
rect 19809 18581 19843 18615
rect 2513 18377 2547 18411
rect 5181 18377 5215 18411
rect 7665 18377 7699 18411
rect 8953 18377 8987 18411
rect 9965 18377 9999 18411
rect 12449 18377 12483 18411
rect 15669 18377 15703 18411
rect 3157 18309 3191 18343
rect 6101 18309 6135 18343
rect 11345 18309 11379 18343
rect 14841 18309 14875 18343
rect 3709 18241 3743 18275
rect 4629 18241 4663 18275
rect 4721 18241 4755 18275
rect 5733 18241 5767 18275
rect 1777 18173 1811 18207
rect 2329 18173 2363 18207
rect 3525 18173 3559 18207
rect 3617 18105 3651 18139
rect 4537 18105 4571 18139
rect 5641 18105 5675 18139
rect 16865 18309 16899 18343
rect 6469 18241 6503 18275
rect 8217 18241 8251 18275
rect 9505 18241 9539 18275
rect 10425 18241 10459 18275
rect 10609 18241 10643 18275
rect 11989 18241 12023 18275
rect 13001 18241 13035 18275
rect 14381 18241 14415 18275
rect 15485 18241 15519 18275
rect 15669 18241 15703 18275
rect 16313 18241 16347 18275
rect 16497 18241 16531 18275
rect 17325 18241 17359 18275
rect 17417 18241 17451 18275
rect 18705 18241 18739 18275
rect 19993 18241 20027 18275
rect 6193 18173 6227 18207
rect 6837 18173 6871 18207
rect 9413 18173 9447 18207
rect 9873 18173 9907 18207
rect 11713 18173 11747 18207
rect 12817 18173 12851 18207
rect 16221 18173 16255 18207
rect 20453 18173 20487 18207
rect 15301 18105 15335 18139
rect 18429 18105 18463 18139
rect 19901 18105 19935 18139
rect 20729 18105 20763 18139
rect 1961 18037 1995 18071
rect 4169 18037 4203 18071
rect 5549 18037 5583 18071
rect 6101 18037 6135 18071
rect 7021 18037 7055 18071
rect 7481 18037 7515 18071
rect 8033 18037 8067 18071
rect 8125 18037 8159 18071
rect 9321 18037 9355 18071
rect 9873 18037 9907 18071
rect 10333 18037 10367 18071
rect 11805 18037 11839 18071
rect 12909 18037 12943 18071
rect 13829 18037 13863 18071
rect 14197 18037 14231 18071
rect 14289 18037 14323 18071
rect 15209 18037 15243 18071
rect 15853 18037 15887 18071
rect 17233 18037 17267 18071
rect 18061 18037 18095 18071
rect 18521 18037 18555 18071
rect 19441 18037 19475 18071
rect 19809 18037 19843 18071
rect 1685 17833 1719 17867
rect 3341 17833 3375 17867
rect 4077 17833 4111 17867
rect 4537 17833 4571 17867
rect 7297 17833 7331 17867
rect 7665 17833 7699 17867
rect 8493 17833 8527 17867
rect 8861 17833 8895 17867
rect 9689 17833 9723 17867
rect 12817 17833 12851 17867
rect 13185 17833 13219 17867
rect 14013 17833 14047 17867
rect 15301 17833 15335 17867
rect 16313 17833 16347 17867
rect 16773 17833 16807 17867
rect 17325 17833 17359 17867
rect 18705 17833 18739 17867
rect 19533 17833 19567 17867
rect 2329 17765 2363 17799
rect 3433 17765 3467 17799
rect 10701 17765 10735 17799
rect 13277 17765 13311 17799
rect 14473 17765 14507 17799
rect 17693 17765 17727 17799
rect 1501 17697 1535 17731
rect 2053 17697 2087 17731
rect 4445 17697 4479 17731
rect 5713 17697 5747 17731
rect 10057 17697 10091 17731
rect 11161 17697 11195 17731
rect 11428 17697 11462 17731
rect 14381 17697 14415 17731
rect 15669 17697 15703 17731
rect 15761 17697 15795 17731
rect 16681 17697 16715 17731
rect 19901 17697 19935 17731
rect 3617 17629 3651 17663
rect 4629 17629 4663 17663
rect 5089 17629 5123 17663
rect 5457 17629 5491 17663
rect 7757 17629 7791 17663
rect 7941 17629 7975 17663
rect 8953 17629 8987 17663
rect 9045 17629 9079 17663
rect 10149 17629 10183 17663
rect 10241 17629 10275 17663
rect 13369 17629 13403 17663
rect 14565 17629 14599 17663
rect 15853 17629 15887 17663
rect 16865 17629 16899 17663
rect 17785 17629 17819 17663
rect 17877 17629 17911 17663
rect 18797 17629 18831 17663
rect 18981 17629 19015 17663
rect 19993 17629 20027 17663
rect 20085 17629 20119 17663
rect 2973 17561 3007 17595
rect 6837 17561 6871 17595
rect 18337 17561 18371 17595
rect 7113 17493 7147 17527
rect 12541 17493 12575 17527
rect 1501 17289 1535 17323
rect 3893 17289 3927 17323
rect 5549 17289 5583 17323
rect 6377 17289 6411 17323
rect 7941 17289 7975 17323
rect 9137 17289 9171 17323
rect 10977 17289 11011 17323
rect 11161 17289 11195 17323
rect 13093 17289 13127 17323
rect 17601 17289 17635 17323
rect 19809 17289 19843 17323
rect 19901 17289 19935 17323
rect 4077 17221 4111 17255
rect 1961 17153 1995 17187
rect 2145 17153 2179 17187
rect 10057 17221 10091 17255
rect 10149 17221 10183 17255
rect 7757 17153 7791 17187
rect 8585 17153 8619 17187
rect 9689 17153 9723 17187
rect 2513 17085 2547 17119
rect 2780 17085 2814 17119
rect 4077 17085 4111 17119
rect 4169 17085 4203 17119
rect 4425 17085 4459 17119
rect 6193 17085 6227 17119
rect 18889 17221 18923 17255
rect 10701 17153 10735 17187
rect 10977 17153 11011 17187
rect 11805 17153 11839 17187
rect 13553 17153 13587 17187
rect 13737 17153 13771 17187
rect 18613 17153 18647 17187
rect 19441 17153 19475 17187
rect 19809 17153 19843 17187
rect 20361 17153 20395 17187
rect 20545 17153 20579 17187
rect 20913 17153 20947 17187
rect 11621 17085 11655 17119
rect 12541 17085 12575 17119
rect 14289 17085 14323 17119
rect 14545 17085 14579 17119
rect 16221 17085 16255 17119
rect 16488 17085 16522 17119
rect 20729 17085 20763 17119
rect 1869 17017 1903 17051
rect 7573 17017 7607 17051
rect 8309 17017 8343 17051
rect 9045 17017 9079 17051
rect 9597 17017 9631 17051
rect 10057 17017 10091 17051
rect 10609 17017 10643 17051
rect 11529 17017 11563 17051
rect 13461 17017 13495 17051
rect 18429 17017 18463 17051
rect 20269 17017 20303 17051
rect 7113 16949 7147 16983
rect 7481 16949 7515 16983
rect 8401 16949 8435 16983
rect 9505 16949 9539 16983
rect 10517 16949 10551 16983
rect 12725 16949 12759 16983
rect 15669 16949 15703 16983
rect 18061 16949 18095 16983
rect 18521 16949 18555 16983
rect 19257 16949 19291 16983
rect 19349 16949 19383 16983
rect 1593 16745 1627 16779
rect 1961 16745 1995 16779
rect 2329 16745 2363 16779
rect 3341 16745 3375 16779
rect 4077 16745 4111 16779
rect 4537 16745 4571 16779
rect 5457 16745 5491 16779
rect 5917 16745 5951 16779
rect 7481 16745 7515 16779
rect 7757 16745 7791 16779
rect 9321 16745 9355 16779
rect 9965 16745 9999 16779
rect 11713 16745 11747 16779
rect 12081 16745 12115 16779
rect 16681 16745 16715 16779
rect 18153 16745 18187 16779
rect 18613 16745 18647 16779
rect 19165 16745 19199 16779
rect 19993 16745 20027 16779
rect 21097 16745 21131 16779
rect 3433 16677 3467 16711
rect 5825 16677 5859 16711
rect 1409 16609 1443 16643
rect 4445 16609 4479 16643
rect 6837 16609 6871 16643
rect 17049 16677 17083 16711
rect 19533 16677 19567 16711
rect 20453 16677 20487 16711
rect 8197 16609 8231 16643
rect 9781 16609 9815 16643
rect 10333 16609 10367 16643
rect 10600 16609 10634 16643
rect 12449 16609 12483 16643
rect 13461 16609 13495 16643
rect 13728 16609 13762 16643
rect 15568 16609 15602 16643
rect 17509 16609 17543 16643
rect 17601 16609 17635 16643
rect 18521 16609 18555 16643
rect 20361 16609 20395 16643
rect 20913 16609 20947 16643
rect 2421 16541 2455 16575
rect 2605 16541 2639 16575
rect 3617 16541 3651 16575
rect 4629 16541 4663 16575
rect 6101 16541 6135 16575
rect 6929 16541 6963 16575
rect 7113 16541 7147 16575
rect 7757 16541 7791 16575
rect 7941 16541 7975 16575
rect 12541 16541 12575 16575
rect 12633 16541 12667 16575
rect 15301 16541 15335 16575
rect 17693 16541 17727 16575
rect 18797 16541 18831 16575
rect 19625 16541 19659 16575
rect 19809 16541 19843 16575
rect 20545 16541 20579 16575
rect 2973 16473 3007 16507
rect 14841 16473 14875 16507
rect 17141 16473 17175 16507
rect 6469 16405 6503 16439
rect 1685 16201 1719 16235
rect 4721 16201 4755 16235
rect 5733 16201 5767 16235
rect 8861 16201 8895 16235
rect 11345 16201 11379 16235
rect 15669 16201 15703 16235
rect 19073 16201 19107 16235
rect 2053 16133 2087 16167
rect 4445 16133 4479 16167
rect 11989 16133 12023 16167
rect 17877 16133 17911 16167
rect 2697 16065 2731 16099
rect 5273 16065 5307 16099
rect 6377 16065 6411 16099
rect 7481 16065 7515 16099
rect 13001 16065 13035 16099
rect 14013 16065 14047 16099
rect 15301 16065 15335 16099
rect 16221 16065 16255 16099
rect 17233 16065 17267 16099
rect 1501 15997 1535 16031
rect 3065 15997 3099 16031
rect 5089 15997 5123 16031
rect 6101 15997 6135 16031
rect 6929 15997 6963 16031
rect 7748 15997 7782 16031
rect 9413 15997 9447 16031
rect 9965 15997 9999 16031
rect 11805 15997 11839 16031
rect 13921 15997 13955 16031
rect 15117 15997 15151 16031
rect 2513 15929 2547 15963
rect 3332 15929 3366 15963
rect 5181 15929 5215 15963
rect 6193 15929 6227 15963
rect 10232 15929 10266 15963
rect 13829 15929 13863 15963
rect 16129 15929 16163 15963
rect 17049 15929 17083 15963
rect 19717 16065 19751 16099
rect 20453 16065 20487 16099
rect 18889 15997 18923 16031
rect 19533 15997 19567 16031
rect 20913 15929 20947 15963
rect 2421 15861 2455 15895
rect 7113 15861 7147 15895
rect 9597 15861 9631 15895
rect 12449 15861 12483 15895
rect 12817 15861 12851 15895
rect 12909 15861 12943 15895
rect 13461 15861 13495 15895
rect 14657 15861 14691 15895
rect 15025 15861 15059 15895
rect 16037 15861 16071 15895
rect 16681 15861 16715 15895
rect 17141 15861 17175 15895
rect 17877 15861 17911 15895
rect 19441 15861 19475 15895
rect 19901 15861 19935 15895
rect 20269 15861 20303 15895
rect 20361 15861 20395 15895
rect 1593 15657 1627 15691
rect 1961 15657 1995 15691
rect 3341 15657 3375 15691
rect 4077 15657 4111 15691
rect 4445 15657 4479 15691
rect 7021 15657 7055 15691
rect 8677 15657 8711 15691
rect 11805 15657 11839 15691
rect 13277 15657 13311 15691
rect 15945 15657 15979 15691
rect 3801 15589 3835 15623
rect 12265 15589 12299 15623
rect 14197 15589 14231 15623
rect 14289 15589 14323 15623
rect 16037 15589 16071 15623
rect 18705 15589 18739 15623
rect 19257 15589 19291 15623
rect 1409 15521 1443 15555
rect 2329 15521 2363 15555
rect 3433 15521 3467 15555
rect 2421 15453 2455 15487
rect 2605 15453 2639 15487
rect 3525 15453 3559 15487
rect 4537 15521 4571 15555
rect 5089 15521 5123 15555
rect 5641 15521 5675 15555
rect 5908 15521 5942 15555
rect 7553 15521 7587 15555
rect 9045 15521 9079 15555
rect 9689 15521 9723 15555
rect 9956 15521 9990 15555
rect 12173 15521 12207 15555
rect 13185 15521 13219 15555
rect 15025 15521 15059 15555
rect 17132 15521 17166 15555
rect 4629 15453 4663 15487
rect 7297 15453 7331 15487
rect 11345 15453 11379 15487
rect 12357 15453 12391 15487
rect 13369 15453 13403 15487
rect 14473 15453 14507 15487
rect 16129 15453 16163 15487
rect 16865 15453 16899 15487
rect 19165 15521 19199 15555
rect 19993 15521 20027 15555
rect 19349 15453 19383 15487
rect 20085 15453 20119 15487
rect 20177 15453 20211 15487
rect 5273 15385 5307 15419
rect 11069 15385 11103 15419
rect 18705 15385 18739 15419
rect 2973 15317 3007 15351
rect 3801 15317 3835 15351
rect 9229 15317 9263 15351
rect 12817 15317 12851 15351
rect 13829 15317 13863 15351
rect 14841 15317 14875 15351
rect 15577 15317 15611 15351
rect 18245 15317 18279 15351
rect 18797 15317 18831 15351
rect 19625 15317 19659 15351
rect 3433 15113 3467 15147
rect 6377 15113 6411 15147
rect 7665 15113 7699 15147
rect 9689 15113 9723 15147
rect 13001 15113 13035 15147
rect 13277 15113 13311 15147
rect 5181 15045 5215 15079
rect 1685 14977 1719 15011
rect 2789 14977 2823 15011
rect 4629 14977 4663 15011
rect 5825 14977 5859 15011
rect 7481 14977 7515 15011
rect 8217 14977 8251 15011
rect 8769 14977 8803 15011
rect 9505 14977 9539 15011
rect 9689 14977 9723 15011
rect 10425 14977 10459 15011
rect 11437 14977 11471 15011
rect 1501 14909 1535 14943
rect 3249 14909 3283 14943
rect 6193 14909 6227 14943
rect 7297 14909 7331 14943
rect 8033 14909 8067 14943
rect 11253 14909 11287 14943
rect 12817 14909 12851 14943
rect 4353 14841 4387 14875
rect 5549 14841 5583 14875
rect 7205 14841 7239 14875
rect 10333 14841 10367 14875
rect 11897 14841 11931 14875
rect 17049 15113 17083 15147
rect 19073 15113 19107 15147
rect 20085 15113 20119 15147
rect 14749 15045 14783 15079
rect 13369 14977 13403 15011
rect 17049 14977 17083 15011
rect 18521 14977 18555 15011
rect 18613 14977 18647 15011
rect 19625 14977 19659 15011
rect 20637 14977 20671 15011
rect 15025 14909 15059 14943
rect 15577 14909 15611 14943
rect 15844 14909 15878 14943
rect 17233 14909 17267 14943
rect 20545 14909 20579 14943
rect 13636 14841 13670 14875
rect 17509 14841 17543 14875
rect 18429 14841 18463 14875
rect 2237 14773 2271 14807
rect 2605 14773 2639 14807
rect 2697 14773 2731 14807
rect 3985 14773 4019 14807
rect 4445 14773 4479 14807
rect 4997 14773 5031 14807
rect 5641 14773 5675 14807
rect 6837 14773 6871 14807
rect 8125 14773 8159 14807
rect 8861 14773 8895 14807
rect 9229 14773 9263 14807
rect 9321 14773 9355 14807
rect 9873 14773 9907 14807
rect 10241 14773 10275 14807
rect 10885 14773 10919 14807
rect 11345 14773 11379 14807
rect 13277 14773 13311 14807
rect 15209 14773 15243 14807
rect 16957 14773 16991 14807
rect 18061 14773 18095 14807
rect 19441 14773 19475 14807
rect 19533 14773 19567 14807
rect 20453 14773 20487 14807
rect 6101 14569 6135 14603
rect 7389 14569 7423 14603
rect 8309 14569 8343 14603
rect 9689 14569 9723 14603
rect 10517 14569 10551 14603
rect 10701 14569 10735 14603
rect 11161 14569 11195 14603
rect 12173 14569 12207 14603
rect 14565 14569 14599 14603
rect 18613 14569 18647 14603
rect 2605 14501 2639 14535
rect 3525 14501 3559 14535
rect 4322 14501 4356 14535
rect 1501 14433 1535 14467
rect 3249 14433 3283 14467
rect 6837 14433 6871 14467
rect 7297 14433 7331 14467
rect 7849 14433 7883 14467
rect 9045 14433 9079 14467
rect 10057 14433 10091 14467
rect 11069 14501 11103 14535
rect 18981 14501 19015 14535
rect 20913 14501 20947 14535
rect 11989 14433 12023 14467
rect 12541 14433 12575 14467
rect 12808 14433 12842 14467
rect 15568 14433 15602 14467
rect 17408 14433 17442 14467
rect 20177 14433 20211 14467
rect 1777 14365 1811 14399
rect 2697 14365 2731 14399
rect 2881 14365 2915 14399
rect 4077 14365 4111 14399
rect 6193 14365 6227 14399
rect 6285 14365 6319 14399
rect 7481 14365 7515 14399
rect 8401 14365 8435 14399
rect 8493 14365 8527 14399
rect 10149 14365 10183 14399
rect 10333 14365 10367 14399
rect 10517 14365 10551 14399
rect 11253 14365 11287 14399
rect 14657 14365 14691 14399
rect 14749 14365 14783 14399
rect 15301 14365 15335 14399
rect 17141 14365 17175 14399
rect 19073 14365 19107 14399
rect 19165 14365 19199 14399
rect 20269 14365 20303 14399
rect 20361 14365 20395 14399
rect 7941 14297 7975 14331
rect 9229 14297 9263 14331
rect 18521 14297 18555 14331
rect 19625 14297 19659 14331
rect 2237 14229 2271 14263
rect 5457 14229 5491 14263
rect 5733 14229 5767 14263
rect 6929 14229 6963 14263
rect 13921 14229 13955 14263
rect 14197 14229 14231 14263
rect 16681 14229 16715 14263
rect 19809 14229 19843 14263
rect 6377 14025 6411 14059
rect 10057 14025 10091 14059
rect 12449 14025 12483 14059
rect 14933 14025 14967 14059
rect 19441 14025 19475 14059
rect 19717 14025 19751 14059
rect 9505 13957 9539 13991
rect 16957 13957 16991 13991
rect 2513 13889 2547 13923
rect 9045 13889 9079 13923
rect 13001 13889 13035 13923
rect 14013 13889 14047 13923
rect 17509 13889 17543 13923
rect 20269 13889 20303 13923
rect 2329 13821 2363 13855
rect 2881 13821 2915 13855
rect 4537 13821 4571 13855
rect 4804 13821 4838 13855
rect 6193 13821 6227 13855
rect 6837 13821 6871 13855
rect 7093 13821 7127 13855
rect 9689 13821 9723 13855
rect 9873 13821 9907 13855
rect 10425 13821 10459 13855
rect 10692 13821 10726 13855
rect 12817 13821 12851 13855
rect 12909 13821 12943 13855
rect 13921 13821 13955 13855
rect 14749 13821 14783 13855
rect 15301 13821 15335 13855
rect 17325 13821 17359 13855
rect 18061 13821 18095 13855
rect 20177 13821 20211 13855
rect 20729 13821 20763 13855
rect 3148 13753 3182 13787
rect 8861 13753 8895 13787
rect 15568 13753 15602 13787
rect 17417 13753 17451 13787
rect 18328 13753 18362 13787
rect 20085 13753 20119 13787
rect 1869 13685 1903 13719
rect 2237 13685 2271 13719
rect 4261 13685 4295 13719
rect 5917 13685 5951 13719
rect 8217 13685 8251 13719
rect 8493 13685 8527 13719
rect 8953 13685 8987 13719
rect 11805 13685 11839 13719
rect 13461 13685 13495 13719
rect 13829 13685 13863 13719
rect 16681 13685 16715 13719
rect 20913 13685 20947 13719
rect 4077 13481 4111 13515
rect 4537 13481 4571 13515
rect 5089 13481 5123 13515
rect 5549 13481 5583 13515
rect 6101 13481 6135 13515
rect 6561 13481 6595 13515
rect 8309 13481 8343 13515
rect 9229 13481 9263 13515
rect 16957 13481 16991 13515
rect 17325 13481 17359 13515
rect 18153 13481 18187 13515
rect 1777 13413 1811 13447
rect 5457 13413 5491 13447
rect 6469 13413 6503 13447
rect 17693 13413 17727 13447
rect 18613 13413 18647 13447
rect 1501 13345 1535 13379
rect 2237 13345 2271 13379
rect 2504 13345 2538 13379
rect 4445 13345 4479 13379
rect 7297 13345 7331 13379
rect 8217 13345 8251 13379
rect 9045 13345 9079 13379
rect 9781 13345 9815 13379
rect 10048 13345 10082 13379
rect 11621 13345 11655 13379
rect 11888 13345 11922 13379
rect 13185 13345 13219 13379
rect 13829 13345 13863 13379
rect 14289 13345 14323 13379
rect 15301 13345 15335 13379
rect 15853 13345 15887 13379
rect 15945 13345 15979 13379
rect 16681 13345 16715 13379
rect 16773 13345 16807 13379
rect 18521 13345 18555 13379
rect 19717 13345 19751 13379
rect 4721 13277 4755 13311
rect 5641 13277 5675 13311
rect 6653 13277 6687 13311
rect 8493 13277 8527 13311
rect 14381 13277 14415 13311
rect 14565 13277 14599 13311
rect 16037 13277 16071 13311
rect 17785 13277 17819 13311
rect 17969 13277 18003 13311
rect 18797 13277 18831 13311
rect 19809 13277 19843 13311
rect 19901 13277 19935 13311
rect 3617 13209 3651 13243
rect 15301 13209 15335 13243
rect 7113 13141 7147 13175
rect 7849 13141 7883 13175
rect 11161 13141 11195 13175
rect 13001 13141 13035 13175
rect 13369 13141 13403 13175
rect 13921 13141 13955 13175
rect 15485 13141 15519 13175
rect 16497 13141 16531 13175
rect 19257 13141 19291 13175
rect 19349 13141 19383 13175
rect 1869 12937 1903 12971
rect 4077 12937 4111 12971
rect 6285 12937 6319 12971
rect 7205 12937 7239 12971
rect 8953 12937 8987 12971
rect 9229 12937 9263 12971
rect 10517 12937 10551 12971
rect 14197 12937 14231 12971
rect 16221 12937 16255 12971
rect 19441 12937 19475 12971
rect 20913 12937 20947 12971
rect 2513 12801 2547 12835
rect 3709 12801 3743 12835
rect 4721 12801 4755 12835
rect 5641 12801 5675 12835
rect 9045 12801 9079 12835
rect 9781 12801 9815 12835
rect 11069 12801 11103 12835
rect 12541 12801 12575 12835
rect 14565 12801 14599 12835
rect 16773 12801 16807 12835
rect 18068 12801 18102 12835
rect 3433 12733 3467 12767
rect 5457 12733 5491 12767
rect 6101 12733 6135 12767
rect 7389 12733 7423 12767
rect 7573 12733 7607 12767
rect 11805 12733 11839 12767
rect 14381 12733 14415 12767
rect 17233 12733 17267 12767
rect 19533 12733 19567 12767
rect 19789 12733 19823 12767
rect 4445 12665 4479 12699
rect 7840 12665 7874 12699
rect 9045 12665 9079 12699
rect 9689 12665 9723 12699
rect 12808 12665 12842 12699
rect 14832 12665 14866 12699
rect 16681 12665 16715 12699
rect 17509 12665 17543 12699
rect 18328 12665 18362 12699
rect 2237 12597 2271 12631
rect 2329 12597 2363 12631
rect 3065 12597 3099 12631
rect 3525 12597 3559 12631
rect 4537 12597 4571 12631
rect 5089 12597 5123 12631
rect 5549 12597 5583 12631
rect 9597 12597 9631 12631
rect 10885 12597 10919 12631
rect 10977 12597 11011 12631
rect 11989 12597 12023 12631
rect 13921 12597 13955 12631
rect 15945 12597 15979 12631
rect 16589 12597 16623 12631
rect 2881 12393 2915 12427
rect 3341 12393 3375 12427
rect 4445 12393 4479 12427
rect 4537 12393 4571 12427
rect 10149 12393 10183 12427
rect 11805 12393 11839 12427
rect 12173 12393 12207 12427
rect 13001 12393 13035 12427
rect 17049 12393 17083 12427
rect 19441 12393 19475 12427
rect 11161 12325 11195 12359
rect 14565 12325 14599 12359
rect 19533 12325 19567 12359
rect 1501 12257 1535 12291
rect 1768 12257 1802 12291
rect 3157 12257 3191 12291
rect 5816 12257 5850 12291
rect 7205 12257 7239 12291
rect 7472 12257 7506 12291
rect 10057 12257 10091 12291
rect 11069 12257 11103 12291
rect 12265 12257 12299 12291
rect 13369 12257 13403 12291
rect 15301 12257 15335 12291
rect 15557 12257 15591 12291
rect 16865 12257 16899 12291
rect 17601 12257 17635 12291
rect 18061 12257 18095 12291
rect 18328 12257 18362 12291
rect 4629 12189 4663 12223
rect 5549 12189 5583 12223
rect 10241 12189 10275 12223
rect 11253 12189 11287 12223
rect 11529 12189 11563 12223
rect 12449 12189 12483 12223
rect 13461 12189 13495 12223
rect 13645 12189 13679 12223
rect 14657 12189 14691 12223
rect 14841 12189 14875 12223
rect 17693 12189 17727 12223
rect 17877 12189 17911 12223
rect 8585 12121 8619 12155
rect 10701 12121 10735 12155
rect 4077 12053 4111 12087
rect 6929 12053 6963 12087
rect 9689 12053 9723 12087
rect 12909 12053 12943 12087
rect 14197 12053 14231 12087
rect 16681 12053 16715 12087
rect 17233 12053 17267 12087
rect 3249 11849 3283 11883
rect 5733 11849 5767 11883
rect 7849 11849 7883 11883
rect 8033 11849 8067 11883
rect 11437 11849 11471 11883
rect 15209 11849 15243 11883
rect 16221 11849 16255 11883
rect 17601 11849 17635 11883
rect 20913 11849 20947 11883
rect 11345 11781 11379 11815
rect 14197 11781 14231 11815
rect 15025 11781 15059 11815
rect 19533 11781 19567 11815
rect 3801 11713 3835 11747
rect 4261 11713 4295 11747
rect 5365 11713 5399 11747
rect 6377 11713 6411 11747
rect 7481 11713 7515 11747
rect 7665 11713 7699 11747
rect 8585 11713 8619 11747
rect 9597 11713 9631 11747
rect 9781 11713 9815 11747
rect 9965 11713 9999 11747
rect 11989 11713 12023 11747
rect 14749 11713 14783 11747
rect 1593 11645 1627 11679
rect 1860 11645 1894 11679
rect 3617 11645 3651 11679
rect 6193 11645 6227 11679
rect 11805 11645 11839 11679
rect 12449 11645 12483 11679
rect 15669 11713 15703 11747
rect 15853 11713 15887 11747
rect 16037 11713 16071 11747
rect 16773 11713 16807 11747
rect 20269 11713 20303 11747
rect 15577 11645 15611 11679
rect 6101 11577 6135 11611
rect 10232 11577 10266 11611
rect 12716 11577 12750 11611
rect 14657 11577 14691 11611
rect 15025 11577 15059 11611
rect 17417 11645 17451 11679
rect 20729 11645 20763 11679
rect 20085 11577 20119 11611
rect 2973 11509 3007 11543
rect 3709 11509 3743 11543
rect 4721 11509 4755 11543
rect 5089 11509 5123 11543
rect 5181 11509 5215 11543
rect 7021 11509 7055 11543
rect 7389 11509 7423 11543
rect 8401 11509 8435 11543
rect 8493 11509 8527 11543
rect 9137 11509 9171 11543
rect 9505 11509 9539 11543
rect 11897 11509 11931 11543
rect 13829 11509 13863 11543
rect 14565 11509 14599 11543
rect 16037 11509 16071 11543
rect 16589 11509 16623 11543
rect 16681 11509 16715 11543
rect 19717 11509 19751 11543
rect 20177 11509 20211 11543
rect 1961 11305 1995 11339
rect 3709 11305 3743 11339
rect 4445 11305 4479 11339
rect 6469 11305 6503 11339
rect 8125 11305 8159 11339
rect 8401 11305 8435 11339
rect 13737 11305 13771 11339
rect 14105 11305 14139 11339
rect 14197 11305 14231 11339
rect 14657 11305 14691 11339
rect 15301 11305 15335 11339
rect 15669 11305 15703 11339
rect 16313 11305 16347 11339
rect 16681 11305 16715 11339
rect 17785 11305 17819 11339
rect 18797 11305 18831 11339
rect 20545 11305 20579 11339
rect 20913 11305 20947 11339
rect 4905 11237 4939 11271
rect 6990 11237 7024 11271
rect 8769 11237 8803 11271
rect 12265 11237 12299 11271
rect 1777 11169 1811 11203
rect 2329 11169 2363 11203
rect 2596 11169 2630 11203
rect 4813 11169 4847 11203
rect 5825 11169 5859 11203
rect 6653 11169 6687 11203
rect 8861 11169 8895 11203
rect 10517 11169 10551 11203
rect 13093 11169 13127 11203
rect 14749 11237 14783 11271
rect 19432 11237 19466 11271
rect 15761 11169 15795 11203
rect 17693 11169 17727 11203
rect 18613 11169 18647 11203
rect 4997 11101 5031 11135
rect 5917 11101 5951 11135
rect 6009 11101 6043 11135
rect 6745 11101 6779 11135
rect 8953 11101 8987 11135
rect 13185 11101 13219 11135
rect 13369 11101 13403 11135
rect 14289 11101 14323 11135
rect 14657 11101 14691 11135
rect 15853 11101 15887 11135
rect 16773 11101 16807 11135
rect 16957 11101 16991 11135
rect 17877 11101 17911 11135
rect 19165 11101 19199 11135
rect 5457 11033 5491 11067
rect 12725 11033 12759 11067
rect 17325 10965 17359 10999
rect 1685 10761 1719 10795
rect 4813 10761 4847 10795
rect 11529 10761 11563 10795
rect 13921 10761 13955 10795
rect 16865 10761 16899 10795
rect 20913 10761 20947 10795
rect 11253 10693 11287 10727
rect 2329 10625 2363 10659
rect 4077 10625 4111 10659
rect 4261 10625 4295 10659
rect 5457 10625 5491 10659
rect 5917 10625 5951 10659
rect 7481 10625 7515 10659
rect 8401 10625 8435 10659
rect 9413 10625 9447 10659
rect 12081 10625 12115 10659
rect 7205 10557 7239 10591
rect 8309 10557 8343 10591
rect 9229 10557 9263 10591
rect 9873 10557 9907 10591
rect 12449 10557 12483 10591
rect 12716 10557 12750 10591
rect 13921 10557 13955 10591
rect 14013 10693 14047 10727
rect 14105 10693 14139 10727
rect 14657 10625 14691 10659
rect 17417 10625 17451 10659
rect 18613 10625 18647 10659
rect 14013 10557 14047 10591
rect 14473 10557 14507 10591
rect 15209 10557 15243 10591
rect 15476 10557 15510 10591
rect 17325 10557 17359 10591
rect 18429 10557 18463 10591
rect 19533 10557 19567 10591
rect 3525 10489 3559 10523
rect 5273 10489 5307 10523
rect 7297 10489 7331 10523
rect 10140 10489 10174 10523
rect 19800 10489 19834 10523
rect 2053 10421 2087 10455
rect 2145 10421 2179 10455
rect 3617 10421 3651 10455
rect 3985 10421 4019 10455
rect 5181 10421 5215 10455
rect 6837 10421 6871 10455
rect 7849 10421 7883 10455
rect 8217 10421 8251 10455
rect 8861 10421 8895 10455
rect 9321 10421 9355 10455
rect 11897 10421 11931 10455
rect 11989 10421 12023 10455
rect 13829 10421 13863 10455
rect 14565 10421 14599 10455
rect 16589 10421 16623 10455
rect 17233 10421 17267 10455
rect 18061 10421 18095 10455
rect 18521 10421 18555 10455
rect 1777 10217 1811 10251
rect 2237 10217 2271 10251
rect 2973 10217 3007 10251
rect 3341 10217 3375 10251
rect 5733 10217 5767 10251
rect 6193 10217 6227 10251
rect 8769 10217 8803 10251
rect 11069 10217 11103 10251
rect 12357 10217 12391 10251
rect 16681 10217 16715 10251
rect 17693 10217 17727 10251
rect 18613 10217 18647 10251
rect 20361 10217 20395 10251
rect 3433 10149 3467 10183
rect 6101 10149 6135 10183
rect 7656 10149 7690 10183
rect 12725 10149 12759 10183
rect 13829 10149 13863 10183
rect 2145 10081 2179 10115
rect 4344 10081 4378 10115
rect 7297 10081 7331 10115
rect 7389 10081 7423 10115
rect 9689 10081 9723 10115
rect 9956 10081 9990 10115
rect 11713 10081 11747 10115
rect 13737 10081 13771 10115
rect 14565 10081 14599 10115
rect 15025 10081 15059 10115
rect 15669 10081 15703 10115
rect 17785 10081 17819 10115
rect 18429 10081 18463 10115
rect 18981 10081 19015 10115
rect 19248 10081 19282 10115
rect 2421 10013 2455 10047
rect 3617 10013 3651 10047
rect 4077 10013 4111 10047
rect 6285 10013 6319 10047
rect 11805 10013 11839 10047
rect 11989 10013 12023 10047
rect 12817 10013 12851 10047
rect 13001 10013 13035 10047
rect 13921 10013 13955 10047
rect 15761 10013 15795 10047
rect 15945 10013 15979 10047
rect 16773 10013 16807 10047
rect 16865 10013 16899 10047
rect 17877 10013 17911 10047
rect 5457 9945 5491 9979
rect 14381 9945 14415 9979
rect 15301 9945 15335 9979
rect 7113 9877 7147 9911
rect 11345 9877 11379 9911
rect 13369 9877 13403 9911
rect 14841 9877 14875 9911
rect 16313 9877 16347 9911
rect 17325 9877 17359 9911
rect 1869 9673 1903 9707
rect 2881 9673 2915 9707
rect 16313 9673 16347 9707
rect 10517 9605 10551 9639
rect 20913 9605 20947 9639
rect 2329 9537 2363 9571
rect 2513 9537 2547 9571
rect 3525 9537 3559 9571
rect 5917 9537 5951 9571
rect 11253 9537 11287 9571
rect 11345 9537 11379 9571
rect 14657 9537 14691 9571
rect 16773 9537 16807 9571
rect 16865 9537 16899 9571
rect 20361 9537 20395 9571
rect 2237 9469 2271 9503
rect 4261 9469 4295 9503
rect 4528 9469 4562 9503
rect 6837 9469 6871 9503
rect 7104 9469 7138 9503
rect 9137 9469 9171 9503
rect 12449 9469 12483 9503
rect 12716 9469 12750 9503
rect 17417 9469 17451 9503
rect 18061 9469 18095 9503
rect 20729 9469 20763 9503
rect 1409 9401 1443 9435
rect 3249 9401 3283 9435
rect 9404 9401 9438 9435
rect 11805 9401 11839 9435
rect 14924 9401 14958 9435
rect 18328 9401 18362 9435
rect 3341 9333 3375 9367
rect 5641 9333 5675 9367
rect 8217 9333 8251 9367
rect 10793 9333 10827 9367
rect 11161 9333 11195 9367
rect 13829 9333 13863 9367
rect 14197 9333 14231 9367
rect 16037 9333 16071 9367
rect 16681 9333 16715 9367
rect 17601 9333 17635 9367
rect 19441 9333 19475 9367
rect 19717 9333 19751 9367
rect 20085 9333 20119 9367
rect 20177 9333 20211 9367
rect 3709 9129 3743 9163
rect 5365 9129 5399 9163
rect 5917 9129 5951 9163
rect 6377 9129 6411 9163
rect 6929 9129 6963 9163
rect 7297 9129 7331 9163
rect 8309 9129 8343 9163
rect 10149 9129 10183 9163
rect 10793 9129 10827 9163
rect 11621 9129 11655 9163
rect 12173 9129 12207 9163
rect 16957 9129 16991 9163
rect 17325 9129 17359 9163
rect 17785 9129 17819 9163
rect 17969 9129 18003 9163
rect 18337 9129 18371 9163
rect 13636 9061 13670 9095
rect 2596 8993 2630 9027
rect 5273 8993 5307 9027
rect 6285 8993 6319 9027
rect 7389 8993 7423 9027
rect 8401 8993 8435 9027
rect 11161 8993 11195 9027
rect 11621 8993 11655 9027
rect 12265 8993 12299 9027
rect 15568 8993 15602 9027
rect 17417 8993 17451 9027
rect 2329 8925 2363 8959
rect 5549 8925 5583 8959
rect 6561 8925 6595 8959
rect 7481 8925 7515 8959
rect 8585 8925 8619 8959
rect 10241 8925 10275 8959
rect 10425 8925 10459 8959
rect 11253 8925 11287 8959
rect 11437 8925 11471 8959
rect 12357 8925 12391 8959
rect 13369 8925 13403 8959
rect 15301 8925 15335 8959
rect 17509 8925 17543 8959
rect 18429 9061 18463 9095
rect 19349 9061 19383 9095
rect 20269 9061 20303 9095
rect 19993 8993 20027 9027
rect 18613 8925 18647 8959
rect 19441 8925 19475 8959
rect 19625 8925 19659 8959
rect 4905 8857 4939 8891
rect 17785 8857 17819 8891
rect 18981 8857 19015 8891
rect 7941 8789 7975 8823
rect 9781 8789 9815 8823
rect 11805 8789 11839 8823
rect 14749 8789 14783 8823
rect 16681 8789 16715 8823
rect 6377 8585 6411 8619
rect 9689 8585 9723 8619
rect 11161 8585 11195 8619
rect 15117 8585 15151 8619
rect 18061 8585 18095 8619
rect 19073 8585 19107 8619
rect 2789 8517 2823 8551
rect 5089 8517 5123 8551
rect 10057 8517 10091 8551
rect 10149 8517 10183 8551
rect 14105 8517 14139 8551
rect 17325 8517 17359 8551
rect 17693 8517 17727 8551
rect 20085 8517 20119 8551
rect 5917 8449 5951 8483
rect 7297 8449 7331 8483
rect 7481 8449 7515 8483
rect 10701 8449 10735 8483
rect 11713 8449 11747 8483
rect 14565 8449 14599 8483
rect 14749 8449 14783 8483
rect 15669 8449 15703 8483
rect 16589 8449 16623 8483
rect 16773 8449 16807 8483
rect 18705 8449 18739 8483
rect 19533 8449 19567 8483
rect 19625 8449 19659 8483
rect 20637 8449 20671 8483
rect 1409 8381 1443 8415
rect 3709 8381 3743 8415
rect 6561 8381 6595 8415
rect 7205 8381 7239 8415
rect 8309 8381 8343 8415
rect 11529 8381 11563 8415
rect 12449 8381 12483 8415
rect 16497 8381 16531 8415
rect 17141 8381 17175 8415
rect 17877 8381 17911 8415
rect 19441 8381 19475 8415
rect 1676 8313 1710 8347
rect 3976 8313 4010 8347
rect 5825 8313 5859 8347
rect 8576 8313 8610 8347
rect 10517 8313 10551 8347
rect 10609 8313 10643 8347
rect 12716 8313 12750 8347
rect 15485 8313 15519 8347
rect 18521 8313 18555 8347
rect 20453 8313 20487 8347
rect 5365 8245 5399 8279
rect 5733 8245 5767 8279
rect 6837 8245 6871 8279
rect 11621 8245 11655 8279
rect 13829 8245 13863 8279
rect 14473 8245 14507 8279
rect 15577 8245 15611 8279
rect 16129 8245 16163 8279
rect 18429 8245 18463 8279
rect 20545 8245 20579 8279
rect 2973 8041 3007 8075
rect 6009 8041 6043 8075
rect 6377 8041 6411 8075
rect 7021 8041 7055 8075
rect 7389 8041 7423 8075
rect 8585 8041 8619 8075
rect 9045 8041 9079 8075
rect 9689 8041 9723 8075
rect 10057 8041 10091 8075
rect 10701 8041 10735 8075
rect 11161 8041 11195 8075
rect 11713 8041 11747 8075
rect 12173 8041 12207 8075
rect 12725 8041 12759 8075
rect 15301 8041 15335 8075
rect 18705 8041 18739 8075
rect 19165 8041 19199 8075
rect 19717 8041 19751 8075
rect 20913 8041 20947 8075
rect 6469 7973 6503 8007
rect 7481 7973 7515 8007
rect 12081 7973 12115 8007
rect 14197 7973 14231 8007
rect 15761 7973 15795 8007
rect 17294 7973 17328 8007
rect 1869 7905 1903 7939
rect 2881 7905 2915 7939
rect 3525 7905 3559 7939
rect 4353 7905 4387 7939
rect 4620 7905 4654 7939
rect 8401 7905 8435 7939
rect 8953 7905 8987 7939
rect 10149 7905 10183 7939
rect 11069 7905 11103 7939
rect 13093 7905 13127 7939
rect 14105 7905 14139 7939
rect 15669 7905 15703 7939
rect 16497 7905 16531 7939
rect 17049 7905 17083 7939
rect 19073 7905 19107 7939
rect 20085 7905 20119 7939
rect 1961 7837 1995 7871
rect 2145 7837 2179 7871
rect 3157 7837 3191 7871
rect 6653 7837 6687 7871
rect 7573 7837 7607 7871
rect 9229 7837 9263 7871
rect 10333 7837 10367 7871
rect 11345 7837 11379 7871
rect 12265 7837 12299 7871
rect 13185 7837 13219 7871
rect 13369 7837 13403 7871
rect 14289 7837 14323 7871
rect 14749 7837 14783 7871
rect 15945 7837 15979 7871
rect 19257 7837 19291 7871
rect 20177 7837 20211 7871
rect 20269 7837 20303 7871
rect 5733 7769 5767 7803
rect 18429 7769 18463 7803
rect 1501 7701 1535 7735
rect 2513 7701 2547 7735
rect 8217 7701 8251 7735
rect 13737 7701 13771 7735
rect 16681 7701 16715 7735
rect 4169 7497 4203 7531
rect 6653 7497 6687 7531
rect 12449 7497 12483 7531
rect 13277 7497 13311 7531
rect 13461 7497 13495 7531
rect 14197 7497 14231 7531
rect 14381 7497 14415 7531
rect 20729 7497 20763 7531
rect 3893 7429 3927 7463
rect 1961 7361 1995 7395
rect 2145 7361 2179 7395
rect 4813 7361 4847 7395
rect 6285 7361 6319 7395
rect 1869 7293 1903 7327
rect 2513 7293 2547 7327
rect 2780 7225 2814 7259
rect 4537 7225 4571 7259
rect 6101 7225 6135 7259
rect 8769 7429 8803 7463
rect 9505 7429 9539 7463
rect 9413 7361 9447 7395
rect 9965 7361 9999 7395
rect 10149 7361 10183 7395
rect 11161 7361 11195 7395
rect 13001 7361 13035 7395
rect 7389 7293 7423 7327
rect 9873 7293 9907 7327
rect 10977 7293 11011 7327
rect 11805 7293 11839 7327
rect 12817 7293 12851 7327
rect 13737 7429 13771 7463
rect 14013 7429 14047 7463
rect 13645 7293 13679 7327
rect 7634 7225 7668 7259
rect 8861 7225 8895 7259
rect 10885 7225 10919 7259
rect 12909 7225 12943 7259
rect 13277 7225 13311 7259
rect 15025 7361 15059 7395
rect 16037 7361 16071 7395
rect 17601 7361 17635 7395
rect 18613 7361 18647 7395
rect 13829 7293 13863 7327
rect 14197 7293 14231 7327
rect 14289 7293 14323 7327
rect 14841 7293 14875 7327
rect 16221 7293 16255 7327
rect 17325 7293 17359 7327
rect 19349 7293 19383 7327
rect 19605 7293 19639 7327
rect 13737 7225 13771 7259
rect 15853 7225 15887 7259
rect 17417 7225 17451 7259
rect 18429 7225 18463 7259
rect 1501 7157 1535 7191
rect 4629 7157 4663 7191
rect 5733 7157 5767 7191
rect 6193 7157 6227 7191
rect 6653 7157 6687 7191
rect 10517 7157 10551 7191
rect 11989 7157 12023 7191
rect 14197 7157 14231 7191
rect 14749 7157 14783 7191
rect 15393 7157 15427 7191
rect 15761 7157 15795 7191
rect 16405 7157 16439 7191
rect 16773 7157 16807 7191
rect 16957 7157 16991 7191
rect 18061 7157 18095 7191
rect 18521 7157 18555 7191
rect 4905 6953 4939 6987
rect 5917 6953 5951 6987
rect 14657 6953 14691 6987
rect 17969 6953 18003 6987
rect 20545 6953 20579 6987
rect 2421 6885 2455 6919
rect 13369 6885 13403 6919
rect 13461 6885 13495 6919
rect 14565 6885 14599 6919
rect 3065 6817 3099 6851
rect 7297 6817 7331 6851
rect 8309 6817 8343 6851
rect 8401 6817 8435 6851
rect 10057 6817 10091 6851
rect 10149 6817 10183 6851
rect 11345 6817 11379 6851
rect 11612 6817 11646 6851
rect 15761 6817 15795 6851
rect 16845 6817 16879 6851
rect 18521 6817 18555 6851
rect 19432 6817 19466 6851
rect 2513 6749 2547 6783
rect 2697 6749 2731 6783
rect 3249 6749 3283 6783
rect 4445 6749 4479 6783
rect 4997 6749 5031 6783
rect 5089 6749 5123 6783
rect 6009 6749 6043 6783
rect 6193 6749 6227 6783
rect 7389 6749 7423 6783
rect 7573 6749 7607 6783
rect 8493 6749 8527 6783
rect 10241 6749 10275 6783
rect 10885 6749 10919 6783
rect 13599 6749 13633 6783
rect 14841 6749 14875 6783
rect 15853 6749 15887 6783
rect 16037 6749 16071 6783
rect 16589 6749 16623 6783
rect 19165 6749 19199 6783
rect 2053 6681 2087 6715
rect 9689 6681 9723 6715
rect 12725 6681 12759 6715
rect 4537 6613 4571 6647
rect 5549 6613 5583 6647
rect 6929 6613 6963 6647
rect 7941 6613 7975 6647
rect 13001 6613 13035 6647
rect 14197 6613 14231 6647
rect 15393 6613 15427 6647
rect 18705 6613 18739 6647
rect 2881 6409 2915 6443
rect 3525 6409 3559 6443
rect 10701 6409 10735 6443
rect 14197 6409 14231 6443
rect 16589 6409 16623 6443
rect 16865 6409 16899 6443
rect 20361 6409 20395 6443
rect 4077 6273 4111 6307
rect 5089 6273 5123 6307
rect 5181 6273 5215 6307
rect 6101 6273 6135 6307
rect 6193 6273 6227 6307
rect 7389 6273 7423 6307
rect 7573 6273 7607 6307
rect 8585 6273 8619 6307
rect 8861 6273 8895 6307
rect 11161 6273 11195 6307
rect 11345 6273 11379 6307
rect 14841 6273 14875 6307
rect 15209 6273 15243 6307
rect 17417 6273 17451 6307
rect 20913 6273 20947 6307
rect 1501 6205 1535 6239
rect 4997 6205 5031 6239
rect 8493 6205 8527 6239
rect 1768 6137 1802 6171
rect 3893 6137 3927 6171
rect 6009 6137 6043 6171
rect 8401 6137 8435 6171
rect 9045 6205 9079 6239
rect 11805 6205 11839 6239
rect 12449 6205 12483 6239
rect 12716 6205 12750 6239
rect 17325 6205 17359 6239
rect 18429 6205 18463 6239
rect 18981 6205 19015 6239
rect 20637 6205 20671 6239
rect 9312 6137 9346 6171
rect 14657 6137 14691 6171
rect 15476 6137 15510 6171
rect 19248 6137 19282 6171
rect 3985 6069 4019 6103
rect 4629 6069 4663 6103
rect 5641 6069 5675 6103
rect 6929 6069 6963 6103
rect 7297 6069 7331 6103
rect 8033 6069 8067 6103
rect 8861 6069 8895 6103
rect 10425 6069 10459 6103
rect 11069 6069 11103 6103
rect 11989 6069 12023 6103
rect 13829 6069 13863 6103
rect 14565 6069 14599 6103
rect 17233 6069 17267 6103
rect 18613 6069 18647 6103
rect 3157 5865 3191 5899
rect 5457 5865 5491 5899
rect 6653 5865 6687 5899
rect 6745 5865 6779 5899
rect 8953 5865 8987 5899
rect 11805 5865 11839 5899
rect 16681 5865 16715 5899
rect 16957 5865 16991 5899
rect 18429 5865 18463 5899
rect 19165 5865 19199 5899
rect 2044 5797 2078 5831
rect 11713 5797 11747 5831
rect 12624 5797 12658 5831
rect 14105 5797 14139 5831
rect 15546 5797 15580 5831
rect 17325 5797 17359 5831
rect 1777 5729 1811 5763
rect 4344 5729 4378 5763
rect 7297 5729 7331 5763
rect 7564 5729 7598 5763
rect 9956 5729 9990 5763
rect 12357 5729 12391 5763
rect 14565 5729 14599 5763
rect 14657 5729 14691 5763
rect 15301 5729 15335 5763
rect 17417 5729 17451 5763
rect 18337 5729 18371 5763
rect 18981 5729 19015 5763
rect 19901 5729 19935 5763
rect 3433 5661 3467 5695
rect 4077 5661 4111 5695
rect 6837 5661 6871 5695
rect 9689 5661 9723 5695
rect 11897 5661 11931 5695
rect 14749 5661 14783 5695
rect 17509 5661 17543 5695
rect 18613 5661 18647 5695
rect 19993 5661 20027 5695
rect 20177 5661 20211 5695
rect 8677 5593 8711 5627
rect 11345 5593 11379 5627
rect 14197 5593 14231 5627
rect 17969 5593 18003 5627
rect 6285 5525 6319 5559
rect 11069 5525 11103 5559
rect 13737 5525 13771 5559
rect 19533 5525 19567 5559
rect 2053 5321 2087 5355
rect 12449 5321 12483 5355
rect 14289 5321 14323 5355
rect 15301 5321 15335 5355
rect 16957 5321 16991 5355
rect 18061 5321 18095 5355
rect 19257 5321 19291 5355
rect 20729 5321 20763 5355
rect 6837 5253 6871 5287
rect 9597 5253 9631 5287
rect 12265 5253 12299 5287
rect 2605 5185 2639 5219
rect 3709 5185 3743 5219
rect 7481 5185 7515 5219
rect 8769 5185 8803 5219
rect 10149 5185 10183 5219
rect 11161 5185 11195 5219
rect 11897 5185 11931 5219
rect 4353 5117 4387 5151
rect 4620 5117 4654 5151
rect 8493 5117 8527 5151
rect 10977 5117 11011 5151
rect 11621 5117 11655 5151
rect 8585 5049 8619 5083
rect 11069 5049 11103 5083
rect 13001 5185 13035 5219
rect 13645 5185 13679 5219
rect 14933 5185 14967 5219
rect 15853 5185 15887 5219
rect 17509 5185 17543 5219
rect 18613 5185 18647 5219
rect 13461 5117 13495 5151
rect 15669 5117 15703 5151
rect 16405 5117 16439 5151
rect 14749 5049 14783 5083
rect 15761 5049 15795 5083
rect 17325 5049 17359 5083
rect 19349 5117 19383 5151
rect 19605 5117 19639 5151
rect 2421 4981 2455 5015
rect 2513 4981 2547 5015
rect 3065 4981 3099 5015
rect 3433 4981 3467 5015
rect 3525 4981 3559 5015
rect 5733 4981 5767 5015
rect 7205 4981 7239 5015
rect 7297 4981 7331 5015
rect 8125 4981 8159 5015
rect 9965 4981 9999 5015
rect 10057 4981 10091 5015
rect 10609 4981 10643 5015
rect 12265 4981 12299 5015
rect 12817 4981 12851 5015
rect 12909 4981 12943 5015
rect 14657 4981 14691 5015
rect 16589 4981 16623 5015
rect 17417 4981 17451 5015
rect 18429 4981 18463 5015
rect 18521 4981 18555 5015
rect 19257 4981 19291 5015
rect 2053 4777 2087 4811
rect 4997 4777 5031 4811
rect 5549 4777 5583 4811
rect 7665 4777 7699 4811
rect 8401 4777 8435 4811
rect 9229 4777 9263 4811
rect 9689 4777 9723 4811
rect 10057 4777 10091 4811
rect 11529 4777 11563 4811
rect 14197 4777 14231 4811
rect 16681 4777 16715 4811
rect 18797 4777 18831 4811
rect 19625 4777 19659 4811
rect 8309 4709 8343 4743
rect 12633 4709 12667 4743
rect 14657 4709 14691 4743
rect 15568 4709 15602 4743
rect 17684 4709 17718 4743
rect 2421 4641 2455 4675
rect 3525 4641 3559 4675
rect 5457 4641 5491 4675
rect 6285 4641 6319 4675
rect 6552 4641 6586 4675
rect 9045 4641 9079 4675
rect 10701 4641 10735 4675
rect 11437 4641 11471 4675
rect 13093 4641 13127 4675
rect 13277 4641 13311 4675
rect 14565 4641 14599 4675
rect 15301 4641 15335 4675
rect 17417 4641 17451 4675
rect 19073 4641 19107 4675
rect 19993 4641 20027 4675
rect 2513 4573 2547 4607
rect 2697 4573 2731 4607
rect 2881 4573 2915 4607
rect 3617 4573 3651 4607
rect 3801 4573 3835 4607
rect 5733 4573 5767 4607
rect 8493 4573 8527 4607
rect 10149 4573 10183 4607
rect 10333 4573 10367 4607
rect 10609 4573 10643 4607
rect 11713 4573 11747 4607
rect 12173 4573 12207 4607
rect 12725 4573 12759 4607
rect 12817 4573 12851 4607
rect 3157 4505 3191 4539
rect 11069 4505 11103 4539
rect 13553 4573 13587 4607
rect 14841 4573 14875 4607
rect 20085 4573 20119 4607
rect 20177 4573 20211 4607
rect 20913 4573 20947 4607
rect 5089 4437 5123 4471
rect 7941 4437 7975 4471
rect 10609 4437 10643 4471
rect 10885 4437 10919 4471
rect 12265 4437 12299 4471
rect 13093 4437 13127 4471
rect 19257 4437 19291 4471
rect 4077 4233 4111 4267
rect 4905 4233 4939 4267
rect 7021 4233 7055 4267
rect 10149 4233 10183 4267
rect 18061 4233 18095 4267
rect 19717 4233 19751 4267
rect 19901 4233 19935 4267
rect 11161 4165 11195 4199
rect 13829 4165 13863 4199
rect 15301 4165 15335 4199
rect 4629 4097 4663 4131
rect 5549 4097 5583 4131
rect 6377 4097 6411 4131
rect 7573 4097 7607 4131
rect 10609 4097 10643 4131
rect 10701 4097 10735 4131
rect 11713 4097 11747 4131
rect 14565 4097 14599 4131
rect 14657 4097 14691 4131
rect 15853 4097 15887 4131
rect 16865 4097 16899 4131
rect 18613 4097 18647 4131
rect 19165 4097 19199 4131
rect 20453 4097 20487 4131
rect 2053 4029 2087 4063
rect 5365 4029 5399 4063
rect 6101 4029 6135 4063
rect 7481 4029 7515 4063
rect 8493 4029 8527 4063
rect 8760 4029 8794 4063
rect 12449 4029 12483 4063
rect 16773 4029 16807 4063
rect 17417 4029 17451 4063
rect 18981 4029 19015 4063
rect 20269 4029 20303 4063
rect 2320 3961 2354 3995
rect 4445 3961 4479 3995
rect 5273 3961 5307 3995
rect 12716 3961 12750 3995
rect 20361 3961 20395 3995
rect 3433 3893 3467 3927
rect 4537 3893 4571 3927
rect 5733 3893 5767 3927
rect 6193 3893 6227 3927
rect 7389 3893 7423 3927
rect 9873 3893 9907 3927
rect 10517 3893 10551 3927
rect 11529 3893 11563 3927
rect 11621 3893 11655 3927
rect 14105 3893 14139 3927
rect 14473 3893 14507 3927
rect 15669 3893 15703 3927
rect 15761 3893 15795 3927
rect 16313 3893 16347 3927
rect 16681 3893 16715 3927
rect 17601 3893 17635 3927
rect 18429 3893 18463 3927
rect 18521 3893 18555 3927
rect 1961 3689 1995 3723
rect 2329 3689 2363 3723
rect 2973 3689 3007 3723
rect 3433 3689 3467 3723
rect 4077 3689 4111 3723
rect 4445 3689 4479 3723
rect 7113 3689 7147 3723
rect 7389 3689 7423 3723
rect 7757 3689 7791 3723
rect 8585 3689 8619 3723
rect 11529 3689 11563 3723
rect 11897 3689 11931 3723
rect 11989 3689 12023 3723
rect 14013 3689 14047 3723
rect 15393 3689 15427 3723
rect 17325 3689 17359 3723
rect 17877 3689 17911 3723
rect 18245 3689 18279 3723
rect 19625 3689 19659 3723
rect 3341 3621 3375 3655
rect 8217 3621 8251 3655
rect 11069 3621 11103 3655
rect 12909 3621 12943 3655
rect 16405 3621 16439 3655
rect 17233 3621 17267 3655
rect 17693 3621 17727 3655
rect 19165 3621 19199 3655
rect 2421 3553 2455 3587
rect 3801 3553 3835 3587
rect 4537 3553 4571 3587
rect 5733 3553 5767 3587
rect 6000 3553 6034 3587
rect 2605 3485 2639 3519
rect 3525 3485 3559 3519
rect 4629 3485 4663 3519
rect 7849 3485 7883 3519
rect 7941 3485 7975 3519
rect 3801 3349 3835 3383
rect 8953 3553 8987 3587
rect 9045 3553 9079 3587
rect 10057 3553 10091 3587
rect 10793 3553 10827 3587
rect 13001 3553 13035 3587
rect 13921 3553 13955 3587
rect 14565 3553 14599 3587
rect 15761 3553 15795 3587
rect 15853 3553 15887 3587
rect 18889 3553 18923 3587
rect 19993 3553 20027 3587
rect 8493 3485 8527 3519
rect 9229 3485 9263 3519
rect 10149 3485 10183 3519
rect 10333 3485 10367 3519
rect 10517 3485 10551 3519
rect 12173 3485 12207 3519
rect 13093 3485 13127 3519
rect 14105 3485 14139 3519
rect 16037 3485 16071 3519
rect 17509 3485 17543 3519
rect 17693 3485 17727 3519
rect 18337 3485 18371 3519
rect 18521 3485 18555 3519
rect 20085 3485 20119 3519
rect 20269 3485 20303 3519
rect 9689 3417 9723 3451
rect 12541 3417 12575 3451
rect 13553 3417 13587 3451
rect 8217 3349 8251 3383
rect 14749 3349 14783 3383
rect 16865 3349 16899 3383
rect 2145 3145 2179 3179
rect 4537 3145 4571 3179
rect 6193 3145 6227 3179
rect 8217 3145 8251 3179
rect 10149 3145 10183 3179
rect 11805 3145 11839 3179
rect 12449 3145 12483 3179
rect 14473 3145 14507 3179
rect 15485 3145 15519 3179
rect 18429 3145 18463 3179
rect 16957 3077 16991 3111
rect 2697 3009 2731 3043
rect 6837 3009 6871 3043
rect 13001 3009 13035 3043
rect 14013 3009 14047 3043
rect 15117 3009 15151 3043
rect 16129 3009 16163 3043
rect 17509 3009 17543 3043
rect 18889 3009 18923 3043
rect 19073 3009 19107 3043
rect 19901 3009 19935 3043
rect 19993 3009 20027 3043
rect 2513 2941 2547 2975
rect 3157 2941 3191 2975
rect 4813 2941 4847 2975
rect 8769 2941 8803 2975
rect 10425 2941 10459 2975
rect 10692 2941 10726 2975
rect 12909 2941 12943 2975
rect 14841 2941 14875 2975
rect 15853 2941 15887 2975
rect 17417 2941 17451 2975
rect 19809 2941 19843 2975
rect 20545 2941 20579 2975
rect 3424 2873 3458 2907
rect 5058 2873 5092 2907
rect 7104 2873 7138 2907
rect 9036 2873 9070 2907
rect 12817 2873 12851 2907
rect 14933 2873 14967 2907
rect 15945 2873 15979 2907
rect 17325 2873 17359 2907
rect 18797 2873 18831 2907
rect 2605 2805 2639 2839
rect 13461 2805 13495 2839
rect 13829 2805 13863 2839
rect 13921 2805 13955 2839
rect 19441 2805 19475 2839
rect 20729 2805 20763 2839
rect 2237 2601 2271 2635
rect 2789 2601 2823 2635
rect 3341 2601 3375 2635
rect 4629 2601 4663 2635
rect 5089 2601 5123 2635
rect 5825 2601 5859 2635
rect 6193 2601 6227 2635
rect 6929 2601 6963 2635
rect 7389 2601 7423 2635
rect 7941 2601 7975 2635
rect 9321 2601 9355 2635
rect 10241 2601 10275 2635
rect 10333 2601 10367 2635
rect 10793 2601 10827 2635
rect 12265 2601 12299 2635
rect 12725 2601 12759 2635
rect 13185 2601 13219 2635
rect 13737 2601 13771 2635
rect 14105 2601 14139 2635
rect 14197 2601 14231 2635
rect 15485 2601 15519 2635
rect 15945 2601 15979 2635
rect 16497 2601 16531 2635
rect 16957 2601 16991 2635
rect 19073 2601 19107 2635
rect 19533 2601 19567 2635
rect 20085 2601 20119 2635
rect 20453 2601 20487 2635
rect 2145 2533 2179 2567
rect 3433 2533 3467 2567
rect 4537 2533 4571 2567
rect 7297 2533 7331 2567
rect 8309 2533 8343 2567
rect 4997 2465 5031 2499
rect 9137 2465 9171 2499
rect 2421 2397 2455 2431
rect 3525 2397 3559 2431
rect 5273 2397 5307 2431
rect 6285 2397 6319 2431
rect 6469 2397 6503 2431
rect 7573 2397 7607 2431
rect 7849 2397 7883 2431
rect 8401 2397 8435 2431
rect 8493 2397 8527 2431
rect 10517 2397 10551 2431
rect 11152 2533 11186 2567
rect 19441 2533 19475 2567
rect 13093 2465 13127 2499
rect 14841 2465 14875 2499
rect 15853 2465 15887 2499
rect 16865 2465 16899 2499
rect 17509 2465 17543 2499
rect 18521 2465 18555 2499
rect 10885 2397 10919 2431
rect 13369 2397 13403 2431
rect 14289 2397 14323 2431
rect 16037 2397 16071 2431
rect 17049 2397 17083 2431
rect 17693 2397 17727 2431
rect 19625 2397 19659 2431
rect 20545 2397 20579 2431
rect 20637 2397 20671 2431
rect 9873 2329 9907 2363
rect 10793 2329 10827 2363
rect 1777 2261 1811 2295
rect 2973 2261 3007 2295
rect 7849 2261 7883 2295
rect 15025 2261 15059 2295
rect 18705 2261 18739 2295
<< metal1 >>
rect 3050 22176 3056 22228
rect 3108 22216 3114 22228
rect 3694 22216 3700 22228
rect 3108 22188 3700 22216
rect 3108 22176 3114 22188
rect 3694 22176 3700 22188
rect 3752 22176 3758 22228
rect 9674 20408 9680 20460
rect 9732 20448 9738 20460
rect 10870 20448 10876 20460
rect 9732 20420 10876 20448
rect 9732 20408 9738 20420
rect 10870 20408 10876 20420
rect 10928 20448 10934 20460
rect 16666 20448 16672 20460
rect 10928 20420 16672 20448
rect 10928 20408 10934 20420
rect 16666 20408 16672 20420
rect 16724 20408 16730 20460
rect 7374 20340 7380 20392
rect 7432 20380 7438 20392
rect 8202 20380 8208 20392
rect 7432 20352 8208 20380
rect 7432 20340 7438 20352
rect 8202 20340 8208 20352
rect 8260 20340 8266 20392
rect 10226 20340 10232 20392
rect 10284 20380 10290 20392
rect 17770 20380 17776 20392
rect 10284 20352 17776 20380
rect 10284 20340 10290 20352
rect 17770 20340 17776 20352
rect 17828 20340 17834 20392
rect 3602 20272 3608 20324
rect 3660 20312 3666 20324
rect 16298 20312 16304 20324
rect 3660 20284 16304 20312
rect 3660 20272 3666 20284
rect 16298 20272 16304 20284
rect 16356 20272 16362 20324
rect 3326 20204 3332 20256
rect 3384 20244 3390 20256
rect 15378 20244 15384 20256
rect 3384 20216 15384 20244
rect 3384 20204 3390 20216
rect 15378 20204 15384 20216
rect 15436 20204 15442 20256
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 1949 20043 2007 20049
rect 1949 20009 1961 20043
rect 1995 20040 2007 20043
rect 2866 20040 2872 20052
rect 1995 20012 2872 20040
rect 1995 20009 2007 20012
rect 1949 20003 2007 20009
rect 2866 20000 2872 20012
rect 2924 20000 2930 20052
rect 3053 20043 3111 20049
rect 3053 20009 3065 20043
rect 3099 20040 3111 20043
rect 3326 20040 3332 20052
rect 3099 20012 3332 20040
rect 3099 20009 3111 20012
rect 3053 20003 3111 20009
rect 3326 20000 3332 20012
rect 3384 20000 3390 20052
rect 3602 20040 3608 20052
rect 3563 20012 3608 20040
rect 3602 20000 3608 20012
rect 3660 20000 3666 20052
rect 5718 20040 5724 20052
rect 3988 20012 5724 20040
rect 1765 19907 1823 19913
rect 1765 19873 1777 19907
rect 1811 19904 1823 19907
rect 1854 19904 1860 19916
rect 1811 19876 1860 19904
rect 1811 19873 1823 19876
rect 1765 19867 1823 19873
rect 1854 19864 1860 19876
rect 1912 19864 1918 19916
rect 2130 19864 2136 19916
rect 2188 19904 2194 19916
rect 2317 19907 2375 19913
rect 2317 19904 2329 19907
rect 2188 19876 2329 19904
rect 2188 19864 2194 19876
rect 2317 19873 2329 19876
rect 2363 19873 2375 19907
rect 2317 19867 2375 19873
rect 2869 19907 2927 19913
rect 2869 19873 2881 19907
rect 2915 19904 2927 19907
rect 3326 19904 3332 19916
rect 2915 19876 3332 19904
rect 2915 19873 2927 19876
rect 2869 19867 2927 19873
rect 3326 19864 3332 19876
rect 3384 19864 3390 19916
rect 3421 19907 3479 19913
rect 3421 19873 3433 19907
rect 3467 19904 3479 19907
rect 3988 19904 4016 20012
rect 5718 20000 5724 20012
rect 5776 20000 5782 20052
rect 7929 20043 7987 20049
rect 7929 20009 7941 20043
rect 7975 20040 7987 20043
rect 8481 20043 8539 20049
rect 8481 20040 8493 20043
rect 7975 20012 8493 20040
rect 7975 20009 7987 20012
rect 7929 20003 7987 20009
rect 8481 20009 8493 20012
rect 8527 20009 8539 20043
rect 9766 20040 9772 20052
rect 9727 20012 9772 20040
rect 8481 20003 8539 20009
rect 9766 20000 9772 20012
rect 9824 20000 9830 20052
rect 13081 20043 13139 20049
rect 13081 20009 13093 20043
rect 13127 20009 13139 20043
rect 13081 20003 13139 20009
rect 4700 19975 4758 19981
rect 4700 19941 4712 19975
rect 4746 19972 4758 19975
rect 8018 19972 8024 19984
rect 4746 19944 8024 19972
rect 4746 19941 4758 19944
rect 4700 19935 4758 19941
rect 8018 19932 8024 19944
rect 8076 19932 8082 19984
rect 9858 19972 9864 19984
rect 8680 19944 9864 19972
rect 3467 19876 4016 19904
rect 3467 19873 3479 19876
rect 3421 19867 3479 19873
rect 5166 19864 5172 19916
rect 5224 19904 5230 19916
rect 6089 19907 6147 19913
rect 6089 19904 6101 19907
rect 5224 19876 6101 19904
rect 5224 19864 5230 19876
rect 6089 19873 6101 19876
rect 6135 19873 6147 19907
rect 6914 19904 6920 19916
rect 6875 19876 6920 19904
rect 6089 19867 6147 19873
rect 6914 19864 6920 19876
rect 6972 19864 6978 19916
rect 7742 19864 7748 19916
rect 7800 19904 7806 19916
rect 7837 19907 7895 19913
rect 7837 19904 7849 19907
rect 7800 19876 7849 19904
rect 7800 19864 7806 19876
rect 7837 19873 7849 19876
rect 7883 19873 7895 19907
rect 8680 19904 8708 19944
rect 9858 19932 9864 19944
rect 9916 19932 9922 19984
rect 9950 19932 9956 19984
rect 10008 19972 10014 19984
rect 11977 19975 12035 19981
rect 11977 19972 11989 19975
rect 10008 19944 11989 19972
rect 10008 19932 10014 19944
rect 11977 19941 11989 19944
rect 12023 19941 12035 19975
rect 13096 19972 13124 20003
rect 13262 20000 13268 20052
rect 13320 20040 13326 20052
rect 14458 20040 14464 20052
rect 13320 20012 14464 20040
rect 13320 20000 13326 20012
rect 14458 20000 14464 20012
rect 14516 20000 14522 20052
rect 18966 20040 18972 20052
rect 18927 20012 18972 20040
rect 18966 20000 18972 20012
rect 19024 20000 19030 20052
rect 19242 20000 19248 20052
rect 19300 20040 19306 20052
rect 19521 20043 19579 20049
rect 19521 20040 19533 20043
rect 19300 20012 19533 20040
rect 19300 20000 19306 20012
rect 19521 20009 19533 20012
rect 19567 20009 19579 20043
rect 19521 20003 19579 20009
rect 16301 19975 16359 19981
rect 13096 19944 16160 19972
rect 11977 19935 12035 19941
rect 8846 19904 8852 19916
rect 7837 19867 7895 19873
rect 8036 19876 8708 19904
rect 8807 19876 8852 19904
rect 4433 19839 4491 19845
rect 4433 19805 4445 19839
rect 4479 19805 4491 19839
rect 4433 19799 4491 19805
rect 6365 19839 6423 19845
rect 6365 19805 6377 19839
rect 6411 19836 6423 19839
rect 8036 19836 8064 19876
rect 8846 19864 8852 19876
rect 8904 19864 8910 19916
rect 9674 19864 9680 19916
rect 9732 19904 9738 19916
rect 10137 19907 10195 19913
rect 10137 19904 10149 19907
rect 9732 19876 10149 19904
rect 9732 19864 9738 19876
rect 10137 19873 10149 19876
rect 10183 19873 10195 19907
rect 10137 19867 10195 19873
rect 10502 19864 10508 19916
rect 10560 19904 10566 19916
rect 10781 19907 10839 19913
rect 10781 19904 10793 19907
rect 10560 19876 10793 19904
rect 10560 19864 10566 19876
rect 10781 19873 10793 19876
rect 10827 19873 10839 19907
rect 11882 19904 11888 19916
rect 11843 19876 11888 19904
rect 10781 19867 10839 19873
rect 11882 19864 11888 19876
rect 11940 19864 11946 19916
rect 13446 19904 13452 19916
rect 13407 19876 13452 19904
rect 13446 19864 13452 19876
rect 13504 19864 13510 19916
rect 14274 19864 14280 19916
rect 14332 19904 14338 19916
rect 14461 19907 14519 19913
rect 14461 19904 14473 19907
rect 14332 19876 14473 19904
rect 14332 19864 14338 19876
rect 14461 19873 14473 19876
rect 14507 19873 14519 19907
rect 14461 19867 14519 19873
rect 15194 19864 15200 19916
rect 15252 19904 15258 19916
rect 15473 19907 15531 19913
rect 15473 19904 15485 19907
rect 15252 19876 15485 19904
rect 15252 19864 15258 19876
rect 15473 19873 15485 19876
rect 15519 19873 15531 19907
rect 15473 19867 15531 19873
rect 16025 19907 16083 19913
rect 16025 19873 16037 19907
rect 16071 19873 16083 19907
rect 16132 19904 16160 19944
rect 16301 19941 16313 19975
rect 16347 19972 16359 19975
rect 17954 19972 17960 19984
rect 16347 19944 17960 19972
rect 16347 19941 16359 19944
rect 16301 19935 16359 19941
rect 17954 19932 17960 19944
rect 18012 19932 18018 19984
rect 16761 19907 16819 19913
rect 16761 19904 16773 19907
rect 16132 19876 16773 19904
rect 16025 19867 16083 19873
rect 16761 19873 16773 19876
rect 16807 19873 16819 19907
rect 16761 19867 16819 19873
rect 6411 19808 8064 19836
rect 8113 19839 8171 19845
rect 6411 19805 6423 19808
rect 6365 19799 6423 19805
rect 8113 19805 8125 19839
rect 8159 19836 8171 19839
rect 8202 19836 8208 19848
rect 8159 19808 8208 19836
rect 8159 19805 8171 19808
rect 8113 19799 8171 19805
rect 2501 19771 2559 19777
rect 2501 19737 2513 19771
rect 2547 19768 2559 19771
rect 2774 19768 2780 19780
rect 2547 19740 2780 19768
rect 2547 19737 2559 19740
rect 2501 19731 2559 19737
rect 2774 19728 2780 19740
rect 2832 19728 2838 19780
rect 4448 19700 4476 19799
rect 8202 19796 8208 19808
rect 8260 19796 8266 19848
rect 8938 19836 8944 19848
rect 8899 19808 8944 19836
rect 8938 19796 8944 19808
rect 8996 19796 9002 19848
rect 9125 19839 9183 19845
rect 9125 19805 9137 19839
rect 9171 19836 9183 19839
rect 9214 19836 9220 19848
rect 9171 19808 9220 19836
rect 9171 19805 9183 19808
rect 9125 19799 9183 19805
rect 9214 19796 9220 19808
rect 9272 19796 9278 19848
rect 10229 19839 10287 19845
rect 10229 19805 10241 19839
rect 10275 19836 10287 19839
rect 10275 19808 10364 19836
rect 10275 19805 10287 19808
rect 10229 19799 10287 19805
rect 7469 19771 7527 19777
rect 7469 19737 7481 19771
rect 7515 19768 7527 19771
rect 10336 19768 10364 19808
rect 10410 19796 10416 19848
rect 10468 19836 10474 19848
rect 10468 19808 10513 19836
rect 10468 19796 10474 19808
rect 10686 19796 10692 19848
rect 10744 19836 10750 19848
rect 10965 19839 11023 19845
rect 10965 19836 10977 19839
rect 10744 19808 10977 19836
rect 10744 19796 10750 19808
rect 10965 19805 10977 19808
rect 11011 19805 11023 19839
rect 10965 19799 11023 19805
rect 11698 19796 11704 19848
rect 11756 19836 11762 19848
rect 12161 19839 12219 19845
rect 12161 19836 12173 19839
rect 11756 19808 12173 19836
rect 11756 19796 11762 19808
rect 12161 19805 12173 19808
rect 12207 19836 12219 19839
rect 12434 19836 12440 19848
rect 12207 19808 12440 19836
rect 12207 19805 12219 19808
rect 12161 19799 12219 19805
rect 12434 19796 12440 19808
rect 12492 19796 12498 19848
rect 12621 19839 12679 19845
rect 12621 19805 12633 19839
rect 12667 19805 12679 19839
rect 13538 19836 13544 19848
rect 13499 19808 13544 19836
rect 12621 19799 12679 19805
rect 7515 19740 10364 19768
rect 12636 19768 12664 19799
rect 13538 19796 13544 19808
rect 13596 19796 13602 19848
rect 13722 19836 13728 19848
rect 13683 19808 13728 19836
rect 13722 19796 13728 19808
rect 13780 19796 13786 19848
rect 14366 19796 14372 19848
rect 14424 19836 14430 19848
rect 14553 19839 14611 19845
rect 14553 19836 14565 19839
rect 14424 19808 14565 19836
rect 14424 19796 14430 19808
rect 14553 19805 14565 19808
rect 14599 19805 14611 19839
rect 14553 19799 14611 19805
rect 14642 19796 14648 19848
rect 14700 19836 14706 19848
rect 14700 19808 14745 19836
rect 14700 19796 14706 19808
rect 15378 19796 15384 19848
rect 15436 19836 15442 19848
rect 16040 19836 16068 19867
rect 17402 19864 17408 19916
rect 17460 19904 17466 19916
rect 17681 19907 17739 19913
rect 17681 19904 17693 19907
rect 17460 19876 17693 19904
rect 17460 19864 17466 19876
rect 17681 19873 17693 19876
rect 17727 19873 17739 19907
rect 17681 19867 17739 19873
rect 18785 19907 18843 19913
rect 18785 19873 18797 19907
rect 18831 19904 18843 19907
rect 18874 19904 18880 19916
rect 18831 19876 18880 19904
rect 18831 19873 18843 19876
rect 18785 19867 18843 19873
rect 18874 19864 18880 19876
rect 18932 19864 18938 19916
rect 19337 19907 19395 19913
rect 19337 19873 19349 19907
rect 19383 19904 19395 19907
rect 20070 19904 20076 19916
rect 19383 19876 20076 19904
rect 19383 19873 19395 19876
rect 19337 19867 19395 19873
rect 20070 19864 20076 19876
rect 20128 19864 20134 19916
rect 20257 19907 20315 19913
rect 20257 19873 20269 19907
rect 20303 19904 20315 19907
rect 20990 19904 20996 19916
rect 20303 19876 20996 19904
rect 20303 19873 20315 19876
rect 20257 19867 20315 19873
rect 20990 19864 20996 19876
rect 21048 19864 21054 19916
rect 17034 19836 17040 19848
rect 15436 19808 16068 19836
rect 16995 19808 17040 19836
rect 15436 19796 15442 19808
rect 17034 19796 17040 19808
rect 17092 19796 17098 19848
rect 20088 19836 20116 19864
rect 20349 19839 20407 19845
rect 20349 19836 20361 19839
rect 20088 19808 20361 19836
rect 20349 19805 20361 19808
rect 20395 19805 20407 19839
rect 20349 19799 20407 19805
rect 20438 19796 20444 19848
rect 20496 19836 20502 19848
rect 20496 19808 20541 19836
rect 20496 19796 20502 19808
rect 14458 19768 14464 19780
rect 12636 19740 14464 19768
rect 7515 19737 7527 19740
rect 7469 19731 7527 19737
rect 14458 19728 14464 19740
rect 14516 19728 14522 19780
rect 15657 19771 15715 19777
rect 15657 19737 15669 19771
rect 15703 19768 15715 19771
rect 18966 19768 18972 19780
rect 15703 19740 18972 19768
rect 15703 19737 15715 19740
rect 15657 19731 15715 19737
rect 18966 19728 18972 19740
rect 19024 19728 19030 19780
rect 4706 19700 4712 19712
rect 4448 19672 4712 19700
rect 4706 19660 4712 19672
rect 4764 19660 4770 19712
rect 5350 19660 5356 19712
rect 5408 19700 5414 19712
rect 5813 19703 5871 19709
rect 5813 19700 5825 19703
rect 5408 19672 5825 19700
rect 5408 19660 5414 19672
rect 5813 19669 5825 19672
rect 5859 19669 5871 19703
rect 5813 19663 5871 19669
rect 7101 19703 7159 19709
rect 7101 19669 7113 19703
rect 7147 19700 7159 19703
rect 8110 19700 8116 19712
rect 7147 19672 8116 19700
rect 7147 19669 7159 19672
rect 7101 19663 7159 19669
rect 8110 19660 8116 19672
rect 8168 19660 8174 19712
rect 8294 19660 8300 19712
rect 8352 19700 8358 19712
rect 10410 19700 10416 19712
rect 8352 19672 10416 19700
rect 8352 19660 8358 19672
rect 10410 19660 10416 19672
rect 10468 19660 10474 19712
rect 11517 19703 11575 19709
rect 11517 19669 11529 19703
rect 11563 19700 11575 19703
rect 12894 19700 12900 19712
rect 11563 19672 12900 19700
rect 11563 19669 11575 19672
rect 11517 19663 11575 19669
rect 12894 19660 12900 19672
rect 12952 19660 12958 19712
rect 14093 19703 14151 19709
rect 14093 19669 14105 19703
rect 14139 19700 14151 19703
rect 14182 19700 14188 19712
rect 14139 19672 14188 19700
rect 14139 19669 14151 19672
rect 14093 19663 14151 19669
rect 14182 19660 14188 19672
rect 14240 19660 14246 19712
rect 17865 19703 17923 19709
rect 17865 19669 17877 19703
rect 17911 19700 17923 19703
rect 18782 19700 18788 19712
rect 17911 19672 18788 19700
rect 17911 19669 17923 19672
rect 17865 19663 17923 19669
rect 18782 19660 18788 19672
rect 18840 19660 18846 19712
rect 19886 19700 19892 19712
rect 19847 19672 19892 19700
rect 19886 19660 19892 19672
rect 19944 19660 19950 19712
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 3053 19499 3111 19505
rect 3053 19465 3065 19499
rect 3099 19496 3111 19499
rect 3142 19496 3148 19508
rect 3099 19468 3148 19496
rect 3099 19465 3111 19468
rect 3053 19459 3111 19465
rect 3142 19456 3148 19468
rect 3200 19456 3206 19508
rect 3326 19456 3332 19508
rect 3384 19496 3390 19508
rect 3384 19468 7972 19496
rect 3384 19456 3390 19468
rect 7944 19428 7972 19468
rect 8018 19456 8024 19508
rect 8076 19496 8082 19508
rect 8205 19499 8263 19505
rect 8205 19496 8217 19499
rect 8076 19468 8217 19496
rect 8076 19456 8082 19468
rect 8205 19465 8217 19468
rect 8251 19496 8263 19499
rect 8294 19496 8300 19508
rect 8251 19468 8300 19496
rect 8251 19465 8263 19468
rect 8205 19459 8263 19465
rect 8294 19456 8300 19468
rect 8352 19456 8358 19508
rect 12342 19496 12348 19508
rect 8496 19468 12348 19496
rect 8496 19428 8524 19468
rect 12342 19456 12348 19468
rect 12400 19456 12406 19508
rect 12434 19456 12440 19508
rect 12492 19496 12498 19508
rect 12492 19468 13400 19496
rect 12492 19456 12498 19468
rect 2240 19400 3188 19428
rect 7944 19400 8524 19428
rect 1670 19252 1676 19304
rect 1728 19292 1734 19304
rect 1765 19295 1823 19301
rect 1765 19292 1777 19295
rect 1728 19264 1777 19292
rect 1728 19252 1734 19264
rect 1765 19261 1777 19264
rect 1811 19261 1823 19295
rect 2240 19292 2268 19400
rect 1765 19255 1823 19261
rect 1863 19264 2268 19292
rect 2317 19295 2375 19301
rect 1118 19184 1124 19236
rect 1176 19224 1182 19236
rect 1863 19224 1891 19264
rect 2317 19261 2329 19295
rect 2363 19292 2375 19295
rect 2682 19292 2688 19304
rect 2363 19264 2688 19292
rect 2363 19261 2375 19264
rect 2317 19255 2375 19261
rect 2682 19252 2688 19264
rect 2740 19252 2746 19304
rect 2866 19292 2872 19304
rect 2827 19264 2872 19292
rect 2866 19252 2872 19264
rect 2924 19252 2930 19304
rect 3050 19252 3056 19304
rect 3108 19252 3114 19304
rect 3068 19224 3096 19252
rect 1176 19196 1891 19224
rect 1964 19196 3096 19224
rect 3160 19224 3188 19400
rect 10226 19388 10232 19440
rect 10284 19428 10290 19440
rect 10321 19431 10379 19437
rect 10321 19428 10333 19431
rect 10284 19400 10333 19428
rect 10284 19388 10290 19400
rect 10321 19397 10333 19400
rect 10367 19397 10379 19431
rect 13372 19428 13400 19468
rect 13722 19456 13728 19508
rect 13780 19496 13786 19508
rect 13817 19499 13875 19505
rect 13817 19496 13829 19499
rect 13780 19468 13829 19496
rect 13780 19456 13786 19468
rect 13817 19465 13829 19468
rect 13863 19465 13875 19499
rect 19334 19496 19340 19508
rect 19295 19468 19340 19496
rect 13817 19459 13875 19465
rect 19334 19456 19340 19468
rect 19392 19456 19398 19508
rect 18874 19428 18880 19440
rect 13372 19400 14688 19428
rect 10321 19391 10379 19397
rect 14660 19369 14688 19400
rect 15304 19400 18880 19428
rect 4341 19363 4399 19369
rect 4341 19360 4353 19363
rect 4251 19332 4353 19360
rect 4341 19329 4353 19332
rect 4387 19360 4399 19363
rect 14645 19363 14703 19369
rect 4387 19332 4844 19360
rect 4387 19329 4399 19332
rect 4341 19323 4399 19329
rect 3510 19252 3516 19304
rect 3568 19292 3574 19304
rect 4356 19292 4384 19323
rect 4706 19292 4712 19304
rect 3568 19264 4384 19292
rect 4667 19264 4712 19292
rect 3568 19252 3574 19264
rect 4706 19252 4712 19264
rect 4764 19252 4770 19304
rect 3160 19196 4016 19224
rect 1176 19184 1182 19196
rect 1964 19165 1992 19196
rect 3988 19168 4016 19196
rect 1949 19159 2007 19165
rect 1949 19125 1961 19159
rect 1995 19125 2007 19159
rect 1949 19119 2007 19125
rect 2501 19159 2559 19165
rect 2501 19125 2513 19159
rect 2547 19156 2559 19159
rect 2958 19156 2964 19168
rect 2547 19128 2964 19156
rect 2547 19125 2559 19128
rect 2501 19119 2559 19125
rect 2958 19116 2964 19128
rect 3016 19116 3022 19168
rect 3697 19159 3755 19165
rect 3697 19125 3709 19159
rect 3743 19156 3755 19159
rect 3878 19156 3884 19168
rect 3743 19128 3884 19156
rect 3743 19125 3755 19128
rect 3697 19119 3755 19125
rect 3878 19116 3884 19128
rect 3936 19116 3942 19168
rect 3970 19116 3976 19168
rect 4028 19156 4034 19168
rect 4065 19159 4123 19165
rect 4065 19156 4077 19159
rect 4028 19128 4077 19156
rect 4028 19116 4034 19128
rect 4065 19125 4077 19128
rect 4111 19125 4123 19159
rect 4065 19119 4123 19125
rect 4157 19159 4215 19165
rect 4157 19125 4169 19159
rect 4203 19156 4215 19159
rect 4706 19156 4712 19168
rect 4203 19128 4712 19156
rect 4203 19125 4215 19128
rect 4157 19119 4215 19125
rect 4706 19116 4712 19128
rect 4764 19116 4770 19168
rect 4816 19156 4844 19332
rect 6748 19332 6960 19360
rect 4976 19295 5034 19301
rect 4976 19261 4988 19295
rect 5022 19292 5034 19295
rect 5350 19292 5356 19304
rect 5022 19264 5356 19292
rect 5022 19261 5034 19264
rect 4976 19255 5034 19261
rect 5350 19252 5356 19264
rect 5408 19252 5414 19304
rect 6454 19252 6460 19304
rect 6512 19292 6518 19304
rect 6748 19292 6776 19332
rect 6512 19264 6776 19292
rect 6825 19295 6883 19301
rect 6512 19252 6518 19264
rect 6825 19261 6837 19295
rect 6871 19261 6883 19295
rect 6932 19292 6960 19332
rect 12268 19332 12572 19360
rect 7092 19295 7150 19301
rect 7092 19292 7104 19295
rect 6932 19264 7104 19292
rect 6825 19255 6883 19261
rect 7092 19261 7104 19264
rect 7138 19292 7150 19295
rect 7650 19292 7656 19304
rect 7138 19264 7656 19292
rect 7138 19261 7150 19264
rect 7092 19255 7150 19261
rect 6730 19184 6736 19236
rect 6788 19224 6794 19236
rect 6840 19224 6868 19255
rect 7650 19252 7656 19264
rect 7708 19252 7714 19304
rect 8481 19295 8539 19301
rect 8481 19292 8493 19295
rect 7760 19264 8493 19292
rect 7558 19224 7564 19236
rect 6788 19196 7564 19224
rect 6788 19184 6794 19196
rect 7558 19184 7564 19196
rect 7616 19224 7622 19236
rect 7760 19224 7788 19264
rect 8481 19261 8493 19264
rect 8527 19261 8539 19295
rect 10045 19295 10103 19301
rect 10045 19292 10057 19295
rect 8481 19255 8539 19261
rect 8680 19264 10057 19292
rect 7616 19196 7788 19224
rect 7616 19184 7622 19196
rect 8110 19184 8116 19236
rect 8168 19224 8174 19236
rect 8680 19224 8708 19264
rect 10045 19261 10057 19264
rect 10091 19261 10103 19295
rect 10045 19255 10103 19261
rect 10137 19295 10195 19301
rect 10137 19261 10149 19295
rect 10183 19292 10195 19295
rect 10410 19292 10416 19304
rect 10183 19264 10416 19292
rect 10183 19261 10195 19264
rect 10137 19255 10195 19261
rect 10410 19252 10416 19264
rect 10468 19252 10474 19304
rect 10689 19295 10747 19301
rect 10689 19261 10701 19295
rect 10735 19292 10747 19295
rect 10778 19292 10784 19304
rect 10735 19264 10784 19292
rect 10735 19261 10747 19264
rect 10689 19255 10747 19261
rect 10778 19252 10784 19264
rect 10836 19252 10842 19304
rect 11238 19252 11244 19304
rect 11296 19292 11302 19304
rect 12268 19292 12296 19332
rect 11296 19264 12296 19292
rect 11296 19252 11302 19264
rect 12342 19252 12348 19304
rect 12400 19292 12406 19304
rect 12437 19295 12495 19301
rect 12437 19292 12449 19295
rect 12400 19264 12449 19292
rect 12400 19252 12406 19264
rect 12437 19261 12449 19264
rect 12483 19261 12495 19295
rect 12544 19292 12572 19332
rect 14645 19329 14657 19363
rect 14691 19329 14703 19363
rect 14645 19323 14703 19329
rect 12544 19264 12839 19292
rect 12437 19255 12495 19261
rect 8168 19196 8708 19224
rect 8748 19227 8806 19233
rect 8168 19184 8174 19196
rect 8748 19193 8760 19227
rect 8794 19224 8806 19227
rect 9122 19224 9128 19236
rect 8794 19196 9128 19224
rect 8794 19193 8806 19196
rect 8748 19187 8806 19193
rect 9122 19184 9128 19196
rect 9180 19184 9186 19236
rect 10956 19227 11014 19233
rect 10956 19193 10968 19227
rect 11002 19224 11014 19227
rect 11422 19224 11428 19236
rect 11002 19196 11428 19224
rect 11002 19193 11014 19196
rect 10956 19187 11014 19193
rect 11422 19184 11428 19196
rect 11480 19224 11486 19236
rect 11698 19224 11704 19236
rect 11480 19196 11704 19224
rect 11480 19184 11486 19196
rect 11698 19184 11704 19196
rect 11756 19184 11762 19236
rect 12682 19227 12740 19233
rect 12682 19224 12694 19227
rect 12084 19196 12694 19224
rect 6089 19159 6147 19165
rect 6089 19156 6101 19159
rect 4816 19128 6101 19156
rect 6089 19125 6101 19128
rect 6135 19125 6147 19159
rect 6089 19119 6147 19125
rect 7282 19116 7288 19168
rect 7340 19156 7346 19168
rect 8662 19156 8668 19168
rect 7340 19128 8668 19156
rect 7340 19116 7346 19128
rect 8662 19116 8668 19128
rect 8720 19116 8726 19168
rect 9214 19116 9220 19168
rect 9272 19156 9278 19168
rect 9861 19159 9919 19165
rect 9861 19156 9873 19159
rect 9272 19128 9873 19156
rect 9272 19116 9278 19128
rect 9861 19125 9873 19128
rect 9907 19125 9919 19159
rect 9861 19119 9919 19125
rect 10045 19159 10103 19165
rect 10045 19125 10057 19159
rect 10091 19156 10103 19159
rect 10226 19156 10232 19168
rect 10091 19128 10232 19156
rect 10091 19125 10103 19128
rect 10045 19119 10103 19125
rect 10226 19116 10232 19128
rect 10284 19116 10290 19168
rect 12084 19165 12112 19196
rect 12682 19193 12694 19196
rect 12728 19193 12740 19227
rect 12811 19224 12839 19264
rect 13078 19252 13084 19304
rect 13136 19292 13142 19304
rect 14458 19292 14464 19304
rect 13136 19264 14320 19292
rect 14419 19264 14464 19292
rect 13136 19252 13142 19264
rect 13170 19224 13176 19236
rect 12811 19196 13176 19224
rect 12682 19187 12740 19193
rect 13170 19184 13176 19196
rect 13228 19184 13234 19236
rect 14292 19224 14320 19264
rect 14458 19252 14464 19264
rect 14516 19252 14522 19304
rect 14553 19295 14611 19301
rect 14553 19261 14565 19295
rect 14599 19292 14611 19295
rect 15010 19292 15016 19304
rect 14599 19264 15016 19292
rect 14599 19261 14611 19264
rect 14553 19255 14611 19261
rect 15010 19252 15016 19264
rect 15068 19292 15074 19304
rect 15304 19292 15332 19400
rect 18874 19388 18880 19400
rect 18932 19388 18938 19440
rect 15749 19363 15807 19369
rect 15749 19329 15761 19363
rect 15795 19360 15807 19363
rect 16206 19360 16212 19372
rect 15795 19332 16212 19360
rect 15795 19329 15807 19332
rect 15749 19323 15807 19329
rect 16206 19320 16212 19332
rect 16264 19320 16270 19372
rect 17126 19320 17132 19372
rect 17184 19360 17190 19372
rect 17221 19363 17279 19369
rect 17221 19360 17233 19363
rect 17184 19332 17233 19360
rect 17184 19320 17190 19332
rect 17221 19329 17233 19332
rect 17267 19329 17279 19363
rect 20346 19360 20352 19372
rect 20307 19332 20352 19360
rect 17221 19323 17279 19329
rect 20346 19320 20352 19332
rect 20404 19320 20410 19372
rect 15068 19264 15332 19292
rect 15473 19295 15531 19301
rect 15068 19252 15074 19264
rect 15473 19261 15485 19295
rect 15519 19292 15531 19295
rect 15930 19292 15936 19304
rect 15519 19264 15936 19292
rect 15519 19261 15531 19264
rect 15473 19255 15531 19261
rect 15930 19252 15936 19264
rect 15988 19252 15994 19304
rect 16114 19292 16120 19304
rect 16075 19264 16120 19292
rect 16114 19252 16120 19264
rect 16172 19252 16178 19304
rect 16574 19252 16580 19304
rect 16632 19292 16638 19304
rect 17037 19295 17095 19301
rect 17037 19292 17049 19295
rect 16632 19264 17049 19292
rect 16632 19252 16638 19264
rect 17037 19261 17049 19264
rect 17083 19261 17095 19295
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 17037 19255 17095 19261
rect 17144 19264 18061 19292
rect 16393 19227 16451 19233
rect 14292 19196 16344 19224
rect 12069 19159 12127 19165
rect 12069 19125 12081 19159
rect 12115 19156 12127 19159
rect 12250 19156 12256 19168
rect 12115 19128 12256 19156
rect 12115 19125 12127 19128
rect 12069 19119 12127 19125
rect 12250 19116 12256 19128
rect 12308 19116 12314 19168
rect 12986 19116 12992 19168
rect 13044 19156 13050 19168
rect 14093 19159 14151 19165
rect 14093 19156 14105 19159
rect 13044 19128 14105 19156
rect 13044 19116 13050 19128
rect 14093 19125 14105 19128
rect 14139 19125 14151 19159
rect 15102 19156 15108 19168
rect 15063 19128 15108 19156
rect 14093 19119 14151 19125
rect 15102 19116 15108 19128
rect 15160 19116 15166 19168
rect 15470 19116 15476 19168
rect 15528 19156 15534 19168
rect 15565 19159 15623 19165
rect 15565 19156 15577 19159
rect 15528 19128 15577 19156
rect 15528 19116 15534 19128
rect 15565 19125 15577 19128
rect 15611 19125 15623 19159
rect 16316 19156 16344 19196
rect 16393 19193 16405 19227
rect 16439 19224 16451 19227
rect 17144 19224 17172 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18414 19292 18420 19304
rect 18375 19264 18420 19292
rect 18049 19255 18107 19261
rect 18414 19252 18420 19264
rect 18472 19252 18478 19304
rect 19153 19295 19211 19301
rect 19153 19261 19165 19295
rect 19199 19261 19211 19295
rect 20162 19292 20168 19304
rect 19153 19255 19211 19261
rect 19260 19264 20168 19292
rect 18969 19227 19027 19233
rect 18969 19224 18981 19227
rect 16439 19196 17172 19224
rect 17420 19196 18981 19224
rect 16439 19193 16451 19196
rect 16393 19187 16451 19193
rect 17420 19156 17448 19196
rect 18969 19193 18981 19196
rect 19015 19224 19027 19227
rect 19168 19224 19196 19255
rect 19015 19196 19196 19224
rect 19015 19193 19027 19196
rect 18969 19187 19027 19193
rect 16316 19128 17448 19156
rect 18233 19159 18291 19165
rect 15565 19119 15623 19125
rect 18233 19125 18245 19159
rect 18279 19156 18291 19159
rect 18506 19156 18512 19168
rect 18279 19128 18512 19156
rect 18279 19125 18291 19128
rect 18233 19119 18291 19125
rect 18506 19116 18512 19128
rect 18564 19116 18570 19168
rect 18601 19159 18659 19165
rect 18601 19125 18613 19159
rect 18647 19156 18659 19159
rect 18690 19156 18696 19168
rect 18647 19128 18696 19156
rect 18647 19125 18659 19128
rect 18601 19119 18659 19125
rect 18690 19116 18696 19128
rect 18748 19116 18754 19168
rect 18874 19116 18880 19168
rect 18932 19156 18938 19168
rect 19260 19156 19288 19264
rect 20162 19252 20168 19264
rect 20220 19252 20226 19304
rect 20717 19295 20775 19301
rect 20717 19261 20729 19295
rect 20763 19292 20775 19295
rect 21266 19292 21272 19304
rect 20763 19264 21272 19292
rect 20763 19261 20775 19264
rect 20717 19255 20775 19261
rect 21266 19252 21272 19264
rect 21324 19252 21330 19304
rect 19334 19184 19340 19236
rect 19392 19224 19398 19236
rect 20622 19224 20628 19236
rect 19392 19196 20628 19224
rect 19392 19184 19398 19196
rect 20622 19184 20628 19196
rect 20680 19184 20686 19236
rect 19702 19156 19708 19168
rect 18932 19128 19288 19156
rect 19663 19128 19708 19156
rect 18932 19116 18938 19128
rect 19702 19116 19708 19128
rect 19760 19116 19766 19168
rect 19886 19116 19892 19168
rect 19944 19156 19950 19168
rect 20073 19159 20131 19165
rect 20073 19156 20085 19159
rect 19944 19128 20085 19156
rect 19944 19116 19950 19128
rect 20073 19125 20085 19128
rect 20119 19125 20131 19159
rect 20073 19119 20131 19125
rect 20162 19116 20168 19168
rect 20220 19156 20226 19168
rect 20898 19156 20904 19168
rect 20220 19128 20265 19156
rect 20859 19128 20904 19156
rect 20220 19116 20226 19128
rect 20898 19116 20904 19128
rect 20956 19116 20962 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 1762 18952 1768 18964
rect 1723 18924 1768 18952
rect 1762 18912 1768 18924
rect 1820 18912 1826 18964
rect 2498 18912 2504 18964
rect 2556 18952 2562 18964
rect 3421 18955 3479 18961
rect 3421 18952 3433 18955
rect 2556 18924 3433 18952
rect 2556 18912 2562 18924
rect 3421 18921 3433 18924
rect 3467 18952 3479 18955
rect 4062 18952 4068 18964
rect 3467 18924 4068 18952
rect 3467 18921 3479 18924
rect 3421 18915 3479 18921
rect 4062 18912 4068 18924
rect 4120 18912 4126 18964
rect 4706 18952 4712 18964
rect 4667 18924 4712 18952
rect 4706 18912 4712 18924
rect 4764 18912 4770 18964
rect 6089 18955 6147 18961
rect 6089 18921 6101 18955
rect 6135 18952 6147 18955
rect 7282 18952 7288 18964
rect 6135 18924 7288 18952
rect 6135 18921 6147 18924
rect 6089 18915 6147 18921
rect 7282 18912 7288 18924
rect 7340 18912 7346 18964
rect 7650 18912 7656 18964
rect 7708 18952 7714 18964
rect 8113 18955 8171 18961
rect 8113 18952 8125 18955
rect 7708 18924 8125 18952
rect 7708 18912 7714 18924
rect 8113 18921 8125 18924
rect 8159 18952 8171 18955
rect 8202 18952 8208 18964
rect 8159 18924 8208 18952
rect 8159 18921 8171 18924
rect 8113 18915 8171 18921
rect 8202 18912 8208 18924
rect 8260 18912 8266 18964
rect 8573 18955 8631 18961
rect 8573 18921 8585 18955
rect 8619 18952 8631 18955
rect 8938 18952 8944 18964
rect 8619 18924 8944 18952
rect 8619 18921 8631 18924
rect 8573 18915 8631 18921
rect 8938 18912 8944 18924
rect 8996 18912 9002 18964
rect 10962 18952 10968 18964
rect 10336 18924 10968 18952
rect 1854 18844 1860 18896
rect 1912 18884 1918 18896
rect 10336 18893 10364 18924
rect 10962 18912 10968 18924
rect 11020 18912 11026 18964
rect 11422 18952 11428 18964
rect 11383 18924 11428 18952
rect 11422 18912 11428 18924
rect 11480 18952 11486 18964
rect 12066 18952 12072 18964
rect 11480 18924 12072 18952
rect 11480 18912 11486 18924
rect 12066 18912 12072 18924
rect 12124 18912 12130 18964
rect 12434 18912 12440 18964
rect 12492 18952 12498 18964
rect 16666 18952 16672 18964
rect 12492 18924 12572 18952
rect 16627 18924 16672 18952
rect 12492 18912 12498 18924
rect 2409 18887 2467 18893
rect 2409 18884 2421 18887
rect 1912 18856 2421 18884
rect 1912 18844 1918 18856
rect 2409 18853 2421 18856
rect 2455 18853 2467 18887
rect 5077 18887 5135 18893
rect 5077 18884 5089 18887
rect 2409 18847 2467 18853
rect 3252 18856 5089 18884
rect 1578 18816 1584 18828
rect 1539 18788 1584 18816
rect 1578 18776 1584 18788
rect 1636 18776 1642 18828
rect 2133 18819 2191 18825
rect 2133 18785 2145 18819
rect 2179 18816 2191 18819
rect 2222 18816 2228 18828
rect 2179 18788 2228 18816
rect 2179 18785 2191 18788
rect 2133 18779 2191 18785
rect 2222 18776 2228 18788
rect 2280 18776 2286 18828
rect 3252 18816 3280 18856
rect 5077 18853 5089 18856
rect 5123 18884 5135 18887
rect 10312 18887 10370 18893
rect 5123 18856 8616 18884
rect 5123 18853 5135 18856
rect 5077 18847 5135 18853
rect 2700 18788 3280 18816
rect 3329 18819 3387 18825
rect 658 18708 664 18760
rect 716 18748 722 18760
rect 2700 18748 2728 18788
rect 3329 18785 3341 18819
rect 3375 18785 3387 18819
rect 3329 18779 3387 18785
rect 716 18720 2728 18748
rect 716 18708 722 18720
rect 2038 18640 2044 18692
rect 2096 18680 2102 18692
rect 3050 18680 3056 18692
rect 2096 18652 3056 18680
rect 2096 18640 2102 18652
rect 3050 18640 3056 18652
rect 3108 18640 3114 18692
rect 3344 18680 3372 18779
rect 3418 18776 3424 18828
rect 3476 18816 3482 18828
rect 4065 18819 4123 18825
rect 3476 18788 4016 18816
rect 3476 18776 3482 18788
rect 3510 18748 3516 18760
rect 3471 18720 3516 18748
rect 3510 18708 3516 18720
rect 3568 18708 3574 18760
rect 3988 18748 4016 18788
rect 4065 18785 4077 18819
rect 4111 18816 4123 18819
rect 4338 18816 4344 18828
rect 4111 18788 4344 18816
rect 4111 18785 4123 18788
rect 4065 18779 4123 18785
rect 4338 18776 4344 18788
rect 4396 18776 4402 18828
rect 5169 18819 5227 18825
rect 5169 18785 5181 18819
rect 5215 18816 5227 18819
rect 5258 18816 5264 18828
rect 5215 18788 5264 18816
rect 5215 18785 5227 18788
rect 5169 18779 5227 18785
rect 5258 18776 5264 18788
rect 5316 18776 5322 18828
rect 6730 18816 6736 18828
rect 6691 18788 6736 18816
rect 6730 18776 6736 18788
rect 6788 18776 6794 18828
rect 7000 18819 7058 18825
rect 7000 18785 7012 18819
rect 7046 18816 7058 18819
rect 8294 18816 8300 18828
rect 7046 18788 8300 18816
rect 7046 18785 7058 18788
rect 7000 18779 7058 18785
rect 8294 18776 8300 18788
rect 8352 18776 8358 18828
rect 5350 18748 5356 18760
rect 3988 18720 5212 18748
rect 5311 18720 5356 18748
rect 3418 18680 3424 18692
rect 3344 18652 3424 18680
rect 3418 18640 3424 18652
rect 3476 18640 3482 18692
rect 3602 18640 3608 18692
rect 3660 18680 3666 18692
rect 4249 18683 4307 18689
rect 4249 18680 4261 18683
rect 3660 18652 4261 18680
rect 3660 18640 3666 18652
rect 4249 18649 4261 18652
rect 4295 18649 4307 18683
rect 4249 18643 4307 18649
rect 4338 18640 4344 18692
rect 4396 18680 4402 18692
rect 5184 18680 5212 18720
rect 5350 18708 5356 18720
rect 5408 18708 5414 18760
rect 6178 18748 6184 18760
rect 6139 18720 6184 18748
rect 6178 18708 6184 18720
rect 6236 18708 6242 18760
rect 6365 18751 6423 18757
rect 6365 18717 6377 18751
rect 6411 18748 6423 18751
rect 6454 18748 6460 18760
rect 6411 18720 6460 18748
rect 6411 18717 6423 18720
rect 6365 18711 6423 18717
rect 6454 18708 6460 18720
rect 6512 18708 6518 18760
rect 8588 18748 8616 18856
rect 10312 18853 10324 18887
rect 10358 18853 10370 18887
rect 10312 18847 10370 18853
rect 11146 18844 11152 18896
rect 11204 18884 11210 18896
rect 12161 18887 12219 18893
rect 12161 18884 12173 18887
rect 11204 18856 12173 18884
rect 11204 18844 11210 18856
rect 12161 18853 12173 18856
rect 12207 18853 12219 18887
rect 12544 18884 12572 18924
rect 16666 18912 16672 18924
rect 16724 18912 16730 18964
rect 18598 18952 18604 18964
rect 16776 18924 18092 18952
rect 18559 18924 18604 18952
rect 13814 18893 13820 18896
rect 13081 18887 13139 18893
rect 13081 18884 13093 18887
rect 12161 18847 12219 18853
rect 12268 18856 12480 18884
rect 12544 18856 13093 18884
rect 8662 18776 8668 18828
rect 8720 18816 8726 18828
rect 8941 18819 8999 18825
rect 8941 18816 8953 18819
rect 8720 18788 8953 18816
rect 8720 18776 8726 18788
rect 8941 18785 8953 18788
rect 8987 18816 8999 18819
rect 11698 18816 11704 18828
rect 8987 18788 11704 18816
rect 8987 18785 8999 18788
rect 8941 18779 8999 18785
rect 11698 18776 11704 18788
rect 11756 18776 11762 18828
rect 12069 18819 12127 18825
rect 12069 18785 12081 18819
rect 12115 18816 12127 18819
rect 12268 18816 12296 18856
rect 12115 18788 12296 18816
rect 12452 18816 12480 18856
rect 13081 18853 13093 18856
rect 13127 18853 13139 18887
rect 13081 18847 13139 18853
rect 13797 18887 13820 18893
rect 13797 18853 13809 18887
rect 13797 18847 13820 18853
rect 13814 18844 13820 18847
rect 13872 18844 13878 18896
rect 14090 18844 14096 18896
rect 14148 18884 14154 18896
rect 16776 18884 16804 18924
rect 17770 18884 17776 18896
rect 14148 18856 16804 18884
rect 17731 18856 17776 18884
rect 14148 18844 14154 18856
rect 17770 18844 17776 18856
rect 17828 18844 17834 18896
rect 17954 18844 17960 18896
rect 18012 18844 18018 18896
rect 18064 18884 18092 18924
rect 18598 18912 18604 18924
rect 18656 18912 18662 18964
rect 19426 18952 19432 18964
rect 19387 18924 19432 18952
rect 19426 18912 19432 18924
rect 19484 18912 19490 18964
rect 19610 18884 19616 18896
rect 18064 18856 19616 18884
rect 19610 18844 19616 18856
rect 19668 18844 19674 18896
rect 12805 18819 12863 18825
rect 12452 18788 12756 18816
rect 12115 18785 12127 18788
rect 12069 18779 12127 18785
rect 9033 18751 9091 18757
rect 9033 18748 9045 18751
rect 8588 18720 9045 18748
rect 9033 18717 9045 18720
rect 9079 18717 9091 18751
rect 9033 18711 9091 18717
rect 6730 18680 6736 18692
rect 4396 18652 4568 18680
rect 5184 18652 6736 18680
rect 4396 18640 4402 18652
rect 2961 18615 3019 18621
rect 2961 18581 2973 18615
rect 3007 18612 3019 18615
rect 4154 18612 4160 18624
rect 3007 18584 4160 18612
rect 3007 18581 3019 18584
rect 2961 18575 3019 18581
rect 4154 18572 4160 18584
rect 4212 18572 4218 18624
rect 4540 18621 4568 18652
rect 6730 18640 6736 18652
rect 6788 18640 6794 18692
rect 9048 18680 9076 18711
rect 9122 18708 9128 18760
rect 9180 18748 9186 18760
rect 10045 18751 10103 18757
rect 9180 18720 9225 18748
rect 9180 18708 9186 18720
rect 10045 18717 10057 18751
rect 10091 18717 10103 18751
rect 12250 18748 12256 18760
rect 12211 18720 12256 18748
rect 10045 18711 10103 18717
rect 9490 18680 9496 18692
rect 9048 18652 9496 18680
rect 9490 18640 9496 18652
rect 9548 18640 9554 18692
rect 9582 18640 9588 18692
rect 9640 18680 9646 18692
rect 10060 18680 10088 18711
rect 12250 18708 12256 18720
rect 12308 18708 12314 18760
rect 12728 18748 12756 18788
rect 12805 18785 12817 18819
rect 12851 18816 12863 18819
rect 13265 18819 13323 18825
rect 13265 18816 13277 18819
rect 12851 18788 13277 18816
rect 12851 18785 12863 18788
rect 12805 18779 12863 18785
rect 13265 18785 13277 18788
rect 13311 18785 13323 18819
rect 13265 18779 13323 18785
rect 13449 18819 13507 18825
rect 13449 18785 13461 18819
rect 13495 18816 13507 18819
rect 15286 18816 15292 18828
rect 13495 18788 15292 18816
rect 13495 18785 13507 18788
rect 13449 18779 13507 18785
rect 15286 18776 15292 18788
rect 15344 18776 15350 18828
rect 15654 18816 15660 18828
rect 15615 18788 15660 18816
rect 15654 18776 15660 18788
rect 15712 18776 15718 18828
rect 17862 18816 17868 18828
rect 16224 18788 16896 18816
rect 17823 18788 17868 18816
rect 16224 18760 16252 18788
rect 12986 18748 12992 18760
rect 12728 18720 12992 18748
rect 12986 18708 12992 18720
rect 13044 18708 13050 18760
rect 13354 18708 13360 18760
rect 13412 18748 13418 18760
rect 13541 18751 13599 18757
rect 13541 18748 13553 18751
rect 13412 18720 13553 18748
rect 13412 18708 13418 18720
rect 13541 18717 13553 18720
rect 13587 18717 13599 18751
rect 15746 18748 15752 18760
rect 15707 18720 15752 18748
rect 13541 18711 13599 18717
rect 15746 18708 15752 18720
rect 15804 18708 15810 18760
rect 15933 18751 15991 18757
rect 15933 18717 15945 18751
rect 15979 18748 15991 18751
rect 16206 18748 16212 18760
rect 15979 18720 16212 18748
rect 15979 18717 15991 18720
rect 15933 18711 15991 18717
rect 16206 18708 16212 18720
rect 16264 18708 16270 18760
rect 16666 18708 16672 18760
rect 16724 18748 16730 18760
rect 16868 18757 16896 18788
rect 17862 18776 17868 18788
rect 17920 18776 17926 18828
rect 17972 18816 18000 18844
rect 18417 18819 18475 18825
rect 18417 18816 18429 18819
rect 17972 18788 18429 18816
rect 18417 18785 18429 18788
rect 18463 18785 18475 18819
rect 18417 18779 18475 18785
rect 18598 18776 18604 18828
rect 18656 18816 18662 18828
rect 19245 18819 19303 18825
rect 19245 18816 19257 18819
rect 18656 18788 19257 18816
rect 18656 18776 18662 18788
rect 19245 18785 19257 18788
rect 19291 18785 19303 18819
rect 19245 18779 19303 18785
rect 19978 18776 19984 18828
rect 20036 18816 20042 18828
rect 20165 18819 20223 18825
rect 20165 18816 20177 18819
rect 20036 18788 20177 18816
rect 20036 18776 20042 18788
rect 20165 18785 20177 18788
rect 20211 18785 20223 18819
rect 20165 18779 20223 18785
rect 16761 18751 16819 18757
rect 16761 18748 16773 18751
rect 16724 18720 16773 18748
rect 16724 18708 16730 18720
rect 16761 18717 16773 18720
rect 16807 18717 16819 18751
rect 16761 18711 16819 18717
rect 16853 18751 16911 18757
rect 16853 18717 16865 18751
rect 16899 18717 16911 18751
rect 16853 18711 16911 18717
rect 17586 18708 17592 18760
rect 17644 18748 17650 18760
rect 17957 18751 18015 18757
rect 17957 18748 17969 18751
rect 17644 18720 17969 18748
rect 17644 18708 17650 18720
rect 17957 18717 17969 18720
rect 18003 18717 18015 18751
rect 17957 18711 18015 18717
rect 18506 18708 18512 18760
rect 18564 18748 18570 18760
rect 20257 18751 20315 18757
rect 20257 18748 20269 18751
rect 18564 18720 20269 18748
rect 18564 18708 18570 18720
rect 20257 18717 20269 18720
rect 20303 18717 20315 18751
rect 20257 18711 20315 18717
rect 20346 18708 20352 18760
rect 20404 18748 20410 18760
rect 20404 18720 20449 18748
rect 20404 18708 20410 18720
rect 9640 18652 10088 18680
rect 11701 18683 11759 18689
rect 9640 18640 9646 18652
rect 11701 18649 11713 18683
rect 11747 18680 11759 18683
rect 13446 18680 13452 18692
rect 11747 18652 13452 18680
rect 11747 18649 11759 18652
rect 11701 18643 11759 18649
rect 13446 18640 13452 18652
rect 13504 18640 13510 18692
rect 21542 18680 21548 18692
rect 14476 18652 21548 18680
rect 4525 18615 4583 18621
rect 4525 18581 4537 18615
rect 4571 18612 4583 18615
rect 5350 18612 5356 18624
rect 4571 18584 5356 18612
rect 4571 18581 4583 18584
rect 4525 18575 4583 18581
rect 5350 18572 5356 18584
rect 5408 18572 5414 18624
rect 5721 18615 5779 18621
rect 5721 18581 5733 18615
rect 5767 18612 5779 18615
rect 9674 18612 9680 18624
rect 5767 18584 9680 18612
rect 5767 18581 5779 18584
rect 5721 18575 5779 18581
rect 9674 18572 9680 18584
rect 9732 18572 9738 18624
rect 13170 18572 13176 18624
rect 13228 18612 13234 18624
rect 14476 18612 14504 18652
rect 21542 18640 21548 18652
rect 21600 18640 21606 18692
rect 13228 18584 14504 18612
rect 14921 18615 14979 18621
rect 13228 18572 13234 18584
rect 14921 18581 14933 18615
rect 14967 18612 14979 18615
rect 15010 18612 15016 18624
rect 14967 18584 15016 18612
rect 14967 18581 14979 18584
rect 14921 18575 14979 18581
rect 15010 18572 15016 18584
rect 15068 18572 15074 18624
rect 15289 18615 15347 18621
rect 15289 18581 15301 18615
rect 15335 18612 15347 18615
rect 16022 18612 16028 18624
rect 15335 18584 16028 18612
rect 15335 18581 15347 18584
rect 15289 18575 15347 18581
rect 16022 18572 16028 18584
rect 16080 18572 16086 18624
rect 16298 18612 16304 18624
rect 16259 18584 16304 18612
rect 16298 18572 16304 18584
rect 16356 18572 16362 18624
rect 17405 18615 17463 18621
rect 17405 18581 17417 18615
rect 17451 18612 17463 18615
rect 17678 18612 17684 18624
rect 17451 18584 17684 18612
rect 17451 18581 17463 18584
rect 17405 18575 17463 18581
rect 17678 18572 17684 18584
rect 17736 18572 17742 18624
rect 19794 18612 19800 18624
rect 19755 18584 19800 18612
rect 19794 18572 19800 18584
rect 19852 18572 19858 18624
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 2501 18411 2559 18417
rect 2501 18377 2513 18411
rect 2547 18408 2559 18411
rect 2774 18408 2780 18420
rect 2547 18380 2780 18408
rect 2547 18377 2559 18380
rect 2501 18371 2559 18377
rect 2774 18368 2780 18380
rect 2832 18368 2838 18420
rect 3050 18368 3056 18420
rect 3108 18408 3114 18420
rect 3108 18380 3372 18408
rect 3108 18368 3114 18380
rect 3145 18343 3203 18349
rect 3145 18309 3157 18343
rect 3191 18309 3203 18343
rect 3344 18340 3372 18380
rect 3418 18368 3424 18420
rect 3476 18408 3482 18420
rect 3694 18408 3700 18420
rect 3476 18380 3700 18408
rect 3476 18368 3482 18380
rect 3694 18368 3700 18380
rect 3752 18408 3758 18420
rect 4982 18408 4988 18420
rect 3752 18380 4988 18408
rect 3752 18368 3758 18380
rect 4982 18368 4988 18380
rect 5040 18368 5046 18420
rect 5166 18408 5172 18420
rect 5127 18380 5172 18408
rect 5166 18368 5172 18380
rect 5224 18368 5230 18420
rect 6178 18368 6184 18420
rect 6236 18408 6242 18420
rect 7653 18411 7711 18417
rect 7653 18408 7665 18411
rect 6236 18380 7665 18408
rect 6236 18368 6242 18380
rect 7653 18377 7665 18380
rect 7699 18377 7711 18411
rect 7653 18371 7711 18377
rect 8110 18368 8116 18420
rect 8168 18408 8174 18420
rect 8662 18408 8668 18420
rect 8168 18380 8668 18408
rect 8168 18368 8174 18380
rect 8662 18368 8668 18380
rect 8720 18368 8726 18420
rect 8846 18368 8852 18420
rect 8904 18408 8910 18420
rect 8941 18411 8999 18417
rect 8941 18408 8953 18411
rect 8904 18380 8953 18408
rect 8904 18368 8910 18380
rect 8941 18377 8953 18380
rect 8987 18377 8999 18411
rect 8941 18371 8999 18377
rect 9030 18368 9036 18420
rect 9088 18408 9094 18420
rect 9398 18408 9404 18420
rect 9088 18380 9404 18408
rect 9088 18368 9094 18380
rect 9398 18368 9404 18380
rect 9456 18368 9462 18420
rect 9490 18368 9496 18420
rect 9548 18408 9554 18420
rect 9674 18408 9680 18420
rect 9548 18380 9680 18408
rect 9548 18368 9554 18380
rect 9674 18368 9680 18380
rect 9732 18368 9738 18420
rect 9950 18408 9956 18420
rect 9911 18380 9956 18408
rect 9950 18368 9956 18380
rect 10008 18368 10014 18420
rect 10410 18368 10416 18420
rect 10468 18408 10474 18420
rect 12437 18411 12495 18417
rect 10468 18380 10548 18408
rect 10468 18368 10474 18380
rect 6089 18343 6147 18349
rect 6089 18340 6101 18343
rect 3344 18312 6101 18340
rect 3145 18303 3203 18309
rect 1762 18204 1768 18216
rect 1723 18176 1768 18204
rect 1762 18164 1768 18176
rect 1820 18164 1826 18216
rect 2314 18204 2320 18216
rect 2275 18176 2320 18204
rect 2314 18164 2320 18176
rect 2372 18164 2378 18216
rect 3050 18164 3056 18216
rect 3108 18204 3114 18216
rect 3160 18204 3188 18303
rect 3528 18213 3556 18312
rect 6089 18309 6101 18312
rect 6135 18309 6147 18343
rect 9766 18340 9772 18352
rect 6089 18303 6147 18309
rect 6196 18312 9772 18340
rect 3602 18232 3608 18284
rect 3660 18272 3666 18284
rect 3697 18275 3755 18281
rect 3697 18272 3709 18275
rect 3660 18244 3709 18272
rect 3660 18232 3666 18244
rect 3697 18241 3709 18244
rect 3743 18241 3755 18275
rect 3697 18235 3755 18241
rect 3878 18232 3884 18284
rect 3936 18272 3942 18284
rect 4617 18275 4675 18281
rect 4617 18272 4629 18275
rect 3936 18244 4629 18272
rect 3936 18232 3942 18244
rect 4617 18241 4629 18244
rect 4663 18241 4675 18275
rect 4617 18235 4675 18241
rect 4706 18232 4712 18284
rect 4764 18272 4770 18284
rect 4764 18244 4809 18272
rect 4764 18232 4770 18244
rect 5534 18232 5540 18284
rect 5592 18272 5598 18284
rect 5721 18275 5779 18281
rect 5721 18272 5733 18275
rect 5592 18244 5733 18272
rect 5592 18232 5598 18244
rect 5721 18241 5733 18244
rect 5767 18241 5779 18275
rect 5721 18235 5779 18241
rect 3108 18176 3188 18204
rect 3513 18207 3571 18213
rect 3108 18164 3114 18176
rect 3513 18173 3525 18207
rect 3559 18173 3571 18207
rect 3513 18167 3571 18173
rect 4062 18164 4068 18216
rect 4120 18204 4126 18216
rect 6196 18213 6224 18312
rect 9766 18300 9772 18312
rect 9824 18300 9830 18352
rect 6457 18275 6515 18281
rect 6457 18241 6469 18275
rect 6503 18272 6515 18275
rect 8110 18272 8116 18284
rect 6503 18244 8116 18272
rect 6503 18241 6515 18244
rect 6457 18235 6515 18241
rect 8110 18232 8116 18244
rect 8168 18232 8174 18284
rect 8205 18275 8263 18281
rect 8205 18241 8217 18275
rect 8251 18272 8263 18275
rect 8294 18272 8300 18284
rect 8251 18244 8300 18272
rect 8251 18241 8263 18244
rect 8205 18235 8263 18241
rect 8294 18232 8300 18244
rect 8352 18272 8358 18284
rect 9030 18272 9036 18284
rect 8352 18244 9036 18272
rect 8352 18232 8358 18244
rect 9030 18232 9036 18244
rect 9088 18232 9094 18284
rect 9122 18232 9128 18284
rect 9180 18272 9186 18284
rect 9493 18275 9551 18281
rect 9493 18272 9505 18275
rect 9180 18244 9505 18272
rect 9180 18232 9186 18244
rect 9493 18241 9505 18244
rect 9539 18241 9551 18275
rect 9493 18235 9551 18241
rect 9674 18232 9680 18284
rect 9732 18272 9738 18284
rect 10413 18275 10471 18281
rect 10413 18272 10425 18275
rect 9732 18244 10425 18272
rect 9732 18232 9738 18244
rect 10413 18241 10425 18244
rect 10459 18241 10471 18275
rect 10413 18235 10471 18241
rect 6181 18207 6239 18213
rect 4120 18176 6132 18204
rect 4120 18164 4126 18176
rect 1486 18096 1492 18148
rect 1544 18136 1550 18148
rect 3605 18139 3663 18145
rect 3605 18136 3617 18139
rect 1544 18108 3617 18136
rect 1544 18096 1550 18108
rect 3605 18105 3617 18108
rect 3651 18136 3663 18139
rect 3786 18136 3792 18148
rect 3651 18108 3792 18136
rect 3651 18105 3663 18108
rect 3605 18099 3663 18105
rect 3786 18096 3792 18108
rect 3844 18096 3850 18148
rect 4522 18136 4528 18148
rect 4483 18108 4528 18136
rect 4522 18096 4528 18108
rect 4580 18096 4586 18148
rect 4706 18096 4712 18148
rect 4764 18136 4770 18148
rect 5629 18139 5687 18145
rect 5629 18136 5641 18139
rect 4764 18108 5641 18136
rect 4764 18096 4770 18108
rect 5629 18105 5641 18108
rect 5675 18105 5687 18139
rect 6104 18136 6132 18176
rect 6181 18173 6193 18207
rect 6227 18173 6239 18207
rect 6181 18167 6239 18173
rect 6270 18164 6276 18216
rect 6328 18204 6334 18216
rect 6825 18207 6883 18213
rect 6825 18204 6837 18207
rect 6328 18176 6837 18204
rect 6328 18164 6334 18176
rect 6825 18173 6837 18176
rect 6871 18173 6883 18207
rect 9401 18207 9459 18213
rect 9401 18204 9413 18207
rect 6825 18167 6883 18173
rect 6932 18176 9413 18204
rect 6932 18136 6960 18176
rect 9401 18173 9413 18176
rect 9447 18204 9459 18207
rect 9861 18207 9919 18213
rect 9861 18204 9873 18207
rect 9447 18176 9873 18204
rect 9447 18173 9459 18176
rect 9401 18167 9459 18173
rect 9861 18173 9873 18176
rect 9907 18173 9919 18207
rect 10520 18204 10548 18380
rect 12437 18377 12449 18411
rect 12483 18408 12495 18411
rect 13538 18408 13544 18420
rect 12483 18380 13544 18408
rect 12483 18377 12495 18380
rect 12437 18371 12495 18377
rect 13538 18368 13544 18380
rect 13596 18368 13602 18420
rect 13722 18368 13728 18420
rect 13780 18408 13786 18420
rect 15657 18411 15715 18417
rect 15657 18408 15669 18411
rect 13780 18380 15669 18408
rect 13780 18368 13786 18380
rect 15657 18377 15669 18380
rect 15703 18377 15715 18411
rect 15657 18371 15715 18377
rect 15746 18368 15752 18420
rect 15804 18408 15810 18420
rect 16942 18408 16948 18420
rect 15804 18380 16948 18408
rect 15804 18368 15810 18380
rect 16942 18368 16948 18380
rect 17000 18368 17006 18420
rect 18690 18408 18696 18420
rect 18248 18380 18696 18408
rect 18248 18352 18276 18380
rect 18690 18368 18696 18380
rect 18748 18368 18754 18420
rect 19242 18368 19248 18420
rect 19300 18408 19306 18420
rect 19334 18408 19340 18420
rect 19300 18380 19340 18408
rect 19300 18368 19306 18380
rect 19334 18368 19340 18380
rect 19392 18368 19398 18420
rect 19610 18368 19616 18420
rect 19668 18408 19674 18420
rect 22002 18408 22008 18420
rect 19668 18380 22008 18408
rect 19668 18368 19674 18380
rect 22002 18368 22008 18380
rect 22060 18368 22066 18420
rect 11333 18343 11391 18349
rect 11333 18309 11345 18343
rect 11379 18340 11391 18343
rect 13262 18340 13268 18352
rect 11379 18312 13268 18340
rect 11379 18309 11391 18312
rect 11333 18303 11391 18309
rect 13262 18300 13268 18312
rect 13320 18300 13326 18352
rect 13446 18300 13452 18352
rect 13504 18340 13510 18352
rect 14829 18343 14887 18349
rect 13504 18312 14228 18340
rect 13504 18300 13510 18312
rect 10597 18275 10655 18281
rect 10597 18241 10609 18275
rect 10643 18272 10655 18275
rect 10962 18272 10968 18284
rect 10643 18244 10968 18272
rect 10643 18241 10655 18244
rect 10597 18235 10655 18241
rect 10962 18232 10968 18244
rect 11020 18272 11026 18284
rect 11977 18275 12035 18281
rect 11977 18272 11989 18275
rect 11020 18244 11989 18272
rect 11020 18232 11026 18244
rect 11977 18241 11989 18244
rect 12023 18241 12035 18275
rect 11977 18235 12035 18241
rect 11701 18207 11759 18213
rect 11701 18204 11713 18207
rect 10520 18176 11713 18204
rect 9861 18167 9919 18173
rect 11701 18173 11713 18176
rect 11747 18204 11759 18207
rect 11790 18204 11796 18216
rect 11747 18176 11796 18204
rect 11747 18173 11759 18176
rect 11701 18167 11759 18173
rect 11790 18164 11796 18176
rect 11848 18164 11854 18216
rect 11992 18204 12020 18235
rect 12250 18232 12256 18284
rect 12308 18272 12314 18284
rect 12989 18275 13047 18281
rect 12989 18272 13001 18275
rect 12308 18244 13001 18272
rect 12308 18232 12314 18244
rect 12989 18241 13001 18244
rect 13035 18241 13047 18275
rect 12989 18235 13047 18241
rect 13906 18232 13912 18284
rect 13964 18272 13970 18284
rect 14090 18272 14096 18284
rect 13964 18244 14096 18272
rect 13964 18232 13970 18244
rect 14090 18232 14096 18244
rect 14148 18232 14154 18284
rect 12618 18204 12624 18216
rect 11992 18176 12624 18204
rect 12618 18164 12624 18176
rect 12676 18164 12682 18216
rect 12805 18207 12863 18213
rect 12805 18173 12817 18207
rect 12851 18173 12863 18207
rect 14200 18204 14228 18312
rect 14829 18309 14841 18343
rect 14875 18340 14887 18343
rect 16758 18340 16764 18352
rect 14875 18312 16764 18340
rect 14875 18309 14887 18312
rect 14829 18303 14887 18309
rect 16758 18300 16764 18312
rect 16816 18300 16822 18352
rect 16853 18343 16911 18349
rect 16853 18309 16865 18343
rect 16899 18340 16911 18343
rect 17494 18340 17500 18352
rect 16899 18312 17500 18340
rect 16899 18309 16911 18312
rect 16853 18303 16911 18309
rect 17494 18300 17500 18312
rect 17552 18300 17558 18352
rect 18230 18300 18236 18352
rect 18288 18300 18294 18352
rect 20346 18340 20352 18352
rect 18708 18312 20352 18340
rect 14366 18272 14372 18284
rect 14327 18244 14372 18272
rect 14366 18232 14372 18244
rect 14424 18232 14430 18284
rect 15473 18275 15531 18281
rect 15473 18241 15485 18275
rect 15519 18272 15531 18275
rect 15562 18272 15568 18284
rect 15519 18244 15568 18272
rect 15519 18241 15531 18244
rect 15473 18235 15531 18241
rect 15562 18232 15568 18244
rect 15620 18232 15626 18284
rect 15657 18275 15715 18281
rect 15657 18241 15669 18275
rect 15703 18272 15715 18275
rect 16301 18275 16359 18281
rect 16301 18272 16313 18275
rect 15703 18244 16313 18272
rect 15703 18241 15715 18244
rect 15657 18235 15715 18241
rect 16301 18241 16313 18244
rect 16347 18241 16359 18275
rect 16301 18235 16359 18241
rect 16485 18275 16543 18281
rect 16485 18241 16497 18275
rect 16531 18272 16543 18275
rect 16942 18272 16948 18284
rect 16531 18244 16948 18272
rect 16531 18241 16543 18244
rect 16485 18235 16543 18241
rect 16942 18232 16948 18244
rect 17000 18232 17006 18284
rect 17310 18272 17316 18284
rect 17271 18244 17316 18272
rect 17310 18232 17316 18244
rect 17368 18232 17374 18284
rect 18708 18281 18736 18312
rect 20346 18300 20352 18312
rect 20404 18300 20410 18352
rect 17405 18275 17463 18281
rect 17405 18241 17417 18275
rect 17451 18272 17463 18275
rect 18693 18275 18751 18281
rect 18693 18272 18705 18275
rect 17451 18244 18705 18272
rect 17451 18241 17463 18244
rect 17405 18235 17463 18241
rect 18693 18241 18705 18244
rect 18739 18241 18751 18275
rect 18693 18235 18751 18241
rect 19518 18232 19524 18284
rect 19576 18272 19582 18284
rect 19981 18275 20039 18281
rect 19981 18272 19993 18275
rect 19576 18244 19993 18272
rect 19576 18232 19582 18244
rect 19981 18241 19993 18244
rect 20027 18241 20039 18275
rect 19981 18235 20039 18241
rect 16209 18207 16267 18213
rect 16209 18204 16221 18207
rect 14200 18176 16221 18204
rect 12805 18167 12863 18173
rect 16209 18173 16221 18176
rect 16255 18173 16267 18207
rect 18598 18204 18604 18216
rect 16209 18167 16267 18173
rect 16500 18176 18604 18204
rect 12526 18136 12532 18148
rect 6104 18108 6960 18136
rect 7024 18108 12532 18136
rect 5629 18099 5687 18105
rect 1949 18071 2007 18077
rect 1949 18037 1961 18071
rect 1995 18068 2007 18071
rect 3234 18068 3240 18080
rect 1995 18040 3240 18068
rect 1995 18037 2007 18040
rect 1949 18031 2007 18037
rect 3234 18028 3240 18040
rect 3292 18028 3298 18080
rect 4154 18068 4160 18080
rect 4115 18040 4160 18068
rect 4154 18028 4160 18040
rect 4212 18028 4218 18080
rect 4890 18028 4896 18080
rect 4948 18068 4954 18080
rect 5537 18071 5595 18077
rect 5537 18068 5549 18071
rect 4948 18040 5549 18068
rect 4948 18028 4954 18040
rect 5537 18037 5549 18040
rect 5583 18037 5595 18071
rect 5537 18031 5595 18037
rect 6089 18071 6147 18077
rect 6089 18037 6101 18071
rect 6135 18068 6147 18071
rect 6454 18068 6460 18080
rect 6135 18040 6460 18068
rect 6135 18037 6147 18040
rect 6089 18031 6147 18037
rect 6454 18028 6460 18040
rect 6512 18028 6518 18080
rect 7024 18077 7052 18108
rect 12526 18096 12532 18108
rect 12584 18096 12590 18148
rect 12820 18080 12848 18167
rect 16500 18148 16528 18176
rect 18598 18164 18604 18176
rect 18656 18164 18662 18216
rect 19150 18164 19156 18216
rect 19208 18204 19214 18216
rect 20441 18207 20499 18213
rect 20441 18204 20453 18207
rect 19208 18176 20453 18204
rect 19208 18164 19214 18176
rect 20441 18173 20453 18176
rect 20487 18173 20499 18207
rect 20441 18167 20499 18173
rect 15289 18139 15347 18145
rect 15289 18136 15301 18139
rect 13832 18108 15301 18136
rect 7009 18071 7067 18077
rect 7009 18037 7021 18071
rect 7055 18037 7067 18071
rect 7466 18068 7472 18080
rect 7427 18040 7472 18068
rect 7009 18031 7067 18037
rect 7466 18028 7472 18040
rect 7524 18068 7530 18080
rect 7650 18068 7656 18080
rect 7524 18040 7656 18068
rect 7524 18028 7530 18040
rect 7650 18028 7656 18040
rect 7708 18068 7714 18080
rect 8021 18071 8079 18077
rect 8021 18068 8033 18071
rect 7708 18040 8033 18068
rect 7708 18028 7714 18040
rect 8021 18037 8033 18040
rect 8067 18037 8079 18071
rect 8021 18031 8079 18037
rect 8113 18071 8171 18077
rect 8113 18037 8125 18071
rect 8159 18068 8171 18071
rect 8202 18068 8208 18080
rect 8159 18040 8208 18068
rect 8159 18037 8171 18040
rect 8113 18031 8171 18037
rect 8202 18028 8208 18040
rect 8260 18028 8266 18080
rect 9309 18071 9367 18077
rect 9309 18037 9321 18071
rect 9355 18068 9367 18071
rect 9490 18068 9496 18080
rect 9355 18040 9496 18068
rect 9355 18037 9367 18040
rect 9309 18031 9367 18037
rect 9490 18028 9496 18040
rect 9548 18028 9554 18080
rect 9861 18071 9919 18077
rect 9861 18037 9873 18071
rect 9907 18068 9919 18071
rect 10321 18071 10379 18077
rect 10321 18068 10333 18071
rect 9907 18040 10333 18068
rect 9907 18037 9919 18040
rect 9861 18031 9919 18037
rect 10321 18037 10333 18040
rect 10367 18037 10379 18071
rect 10321 18031 10379 18037
rect 10410 18028 10416 18080
rect 10468 18068 10474 18080
rect 11793 18071 11851 18077
rect 11793 18068 11805 18071
rect 10468 18040 11805 18068
rect 10468 18028 10474 18040
rect 11793 18037 11805 18040
rect 11839 18037 11851 18071
rect 11793 18031 11851 18037
rect 12793 18028 12799 18080
rect 12851 18028 12857 18080
rect 12897 18071 12955 18077
rect 12897 18037 12909 18071
rect 12943 18068 12955 18071
rect 13078 18068 13084 18080
rect 12943 18040 13084 18068
rect 12943 18037 12955 18040
rect 12897 18031 12955 18037
rect 13078 18028 13084 18040
rect 13136 18028 13142 18080
rect 13832 18077 13860 18108
rect 15289 18105 15301 18108
rect 15335 18105 15347 18139
rect 15289 18099 15347 18105
rect 16482 18096 16488 18148
rect 16540 18096 16546 18148
rect 18417 18139 18475 18145
rect 18417 18105 18429 18139
rect 18463 18136 18475 18139
rect 18690 18136 18696 18148
rect 18463 18108 18696 18136
rect 18463 18105 18475 18108
rect 18417 18099 18475 18105
rect 18690 18096 18696 18108
rect 18748 18096 18754 18148
rect 19334 18096 19340 18148
rect 19392 18136 19398 18148
rect 19889 18139 19947 18145
rect 19889 18136 19901 18139
rect 19392 18108 19901 18136
rect 19392 18096 19398 18108
rect 19889 18105 19901 18108
rect 19935 18105 19947 18139
rect 20714 18136 20720 18148
rect 20675 18108 20720 18136
rect 19889 18099 19947 18105
rect 20714 18096 20720 18108
rect 20772 18096 20778 18148
rect 13817 18071 13875 18077
rect 13817 18037 13829 18071
rect 13863 18037 13875 18071
rect 14182 18068 14188 18080
rect 14143 18040 14188 18068
rect 13817 18031 13875 18037
rect 14182 18028 14188 18040
rect 14240 18028 14246 18080
rect 14274 18028 14280 18080
rect 14332 18068 14338 18080
rect 15194 18068 15200 18080
rect 14332 18040 14377 18068
rect 15155 18040 15200 18068
rect 14332 18028 14338 18040
rect 15194 18028 15200 18040
rect 15252 18028 15258 18080
rect 15470 18028 15476 18080
rect 15528 18068 15534 18080
rect 15841 18071 15899 18077
rect 15841 18068 15853 18071
rect 15528 18040 15853 18068
rect 15528 18028 15534 18040
rect 15841 18037 15853 18040
rect 15887 18037 15899 18071
rect 17218 18068 17224 18080
rect 17179 18040 17224 18068
rect 15841 18031 15899 18037
rect 17218 18028 17224 18040
rect 17276 18028 17282 18080
rect 18046 18068 18052 18080
rect 18007 18040 18052 18068
rect 18046 18028 18052 18040
rect 18104 18028 18110 18080
rect 18509 18071 18567 18077
rect 18509 18037 18521 18071
rect 18555 18068 18567 18071
rect 18598 18068 18604 18080
rect 18555 18040 18604 18068
rect 18555 18037 18567 18040
rect 18509 18031 18567 18037
rect 18598 18028 18604 18040
rect 18656 18028 18662 18080
rect 19426 18068 19432 18080
rect 19387 18040 19432 18068
rect 19426 18028 19432 18040
rect 19484 18028 19490 18080
rect 19794 18068 19800 18080
rect 19755 18040 19800 18068
rect 19794 18028 19800 18040
rect 19852 18028 19858 18080
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 1670 17864 1676 17876
rect 1631 17836 1676 17864
rect 1670 17824 1676 17836
rect 1728 17824 1734 17876
rect 1946 17824 1952 17876
rect 2004 17864 2010 17876
rect 3234 17864 3240 17876
rect 2004 17836 3240 17864
rect 2004 17824 2010 17836
rect 3234 17824 3240 17836
rect 3292 17824 3298 17876
rect 3329 17867 3387 17873
rect 3329 17833 3341 17867
rect 3375 17864 3387 17867
rect 4065 17867 4123 17873
rect 4065 17864 4077 17867
rect 3375 17836 4077 17864
rect 3375 17833 3387 17836
rect 3329 17827 3387 17833
rect 4065 17833 4077 17836
rect 4111 17833 4123 17867
rect 4065 17827 4123 17833
rect 4246 17824 4252 17876
rect 4304 17864 4310 17876
rect 4525 17867 4583 17873
rect 4525 17864 4537 17867
rect 4304 17836 4537 17864
rect 4304 17824 4310 17836
rect 4525 17833 4537 17836
rect 4571 17833 4583 17867
rect 4525 17827 4583 17833
rect 4982 17824 4988 17876
rect 5040 17864 5046 17876
rect 6822 17864 6828 17876
rect 5040 17836 6828 17864
rect 5040 17824 5046 17836
rect 6822 17824 6828 17836
rect 6880 17824 6886 17876
rect 7282 17864 7288 17876
rect 7243 17836 7288 17864
rect 7282 17824 7288 17836
rect 7340 17824 7346 17876
rect 7653 17867 7711 17873
rect 7653 17864 7665 17867
rect 7576 17836 7665 17864
rect 2314 17796 2320 17808
rect 2275 17768 2320 17796
rect 2314 17756 2320 17768
rect 2372 17756 2378 17808
rect 3421 17799 3479 17805
rect 3421 17765 3433 17799
rect 3467 17796 3479 17799
rect 4154 17796 4160 17808
rect 3467 17768 4160 17796
rect 3467 17765 3479 17768
rect 3421 17759 3479 17765
rect 4154 17756 4160 17768
rect 4212 17756 4218 17808
rect 1489 17731 1547 17737
rect 1489 17697 1501 17731
rect 1535 17697 1547 17731
rect 1489 17691 1547 17697
rect 2041 17731 2099 17737
rect 2041 17697 2053 17731
rect 2087 17728 2099 17731
rect 3050 17728 3056 17740
rect 2087 17700 3056 17728
rect 2087 17697 2099 17700
rect 2041 17691 2099 17697
rect 1504 17660 1532 17691
rect 3050 17688 3056 17700
rect 3108 17688 3114 17740
rect 3510 17688 3516 17740
rect 3568 17728 3574 17740
rect 4433 17731 4491 17737
rect 4433 17728 4445 17731
rect 3568 17700 4445 17728
rect 3568 17688 3574 17700
rect 4433 17697 4445 17700
rect 4479 17697 4491 17731
rect 4433 17691 4491 17697
rect 4798 17688 4804 17740
rect 4856 17728 4862 17740
rect 4856 17700 5212 17728
rect 4856 17688 4862 17700
rect 5184 17672 5212 17700
rect 5534 17688 5540 17740
rect 5592 17728 5598 17740
rect 5701 17731 5759 17737
rect 5701 17728 5713 17731
rect 5592 17700 5713 17728
rect 5592 17688 5598 17700
rect 5701 17697 5713 17700
rect 5747 17697 5759 17731
rect 5701 17691 5759 17697
rect 7466 17688 7472 17740
rect 7524 17728 7530 17740
rect 7576 17728 7604 17836
rect 7653 17833 7665 17836
rect 7699 17833 7711 17867
rect 7653 17827 7711 17833
rect 7742 17824 7748 17876
rect 7800 17864 7806 17876
rect 8481 17867 8539 17873
rect 8481 17864 8493 17867
rect 7800 17836 8493 17864
rect 7800 17824 7806 17836
rect 8481 17833 8493 17836
rect 8527 17833 8539 17867
rect 8481 17827 8539 17833
rect 8849 17867 8907 17873
rect 8849 17833 8861 17867
rect 8895 17864 8907 17867
rect 9677 17867 9735 17873
rect 9677 17864 9689 17867
rect 8895 17836 9689 17864
rect 8895 17833 8907 17836
rect 8849 17827 8907 17833
rect 9677 17833 9689 17836
rect 9723 17833 9735 17867
rect 12158 17864 12164 17876
rect 9677 17827 9735 17833
rect 9784 17836 12164 17864
rect 7834 17756 7840 17808
rect 7892 17796 7898 17808
rect 9784 17796 9812 17836
rect 12158 17824 12164 17836
rect 12216 17824 12222 17876
rect 12802 17864 12808 17876
rect 12763 17836 12808 17864
rect 12802 17824 12808 17836
rect 12860 17824 12866 17876
rect 13173 17867 13231 17873
rect 13173 17833 13185 17867
rect 13219 17864 13231 17867
rect 13446 17864 13452 17876
rect 13219 17836 13452 17864
rect 13219 17833 13231 17836
rect 13173 17827 13231 17833
rect 13446 17824 13452 17836
rect 13504 17824 13510 17876
rect 14001 17867 14059 17873
rect 14001 17833 14013 17867
rect 14047 17864 14059 17867
rect 14182 17864 14188 17876
rect 14047 17836 14188 17864
rect 14047 17833 14059 17836
rect 14001 17827 14059 17833
rect 14182 17824 14188 17836
rect 14240 17824 14246 17876
rect 15286 17864 15292 17876
rect 15247 17836 15292 17864
rect 15286 17824 15292 17836
rect 15344 17824 15350 17876
rect 16301 17867 16359 17873
rect 16301 17833 16313 17867
rect 16347 17864 16359 17867
rect 16574 17864 16580 17876
rect 16347 17836 16580 17864
rect 16347 17833 16359 17836
rect 16301 17827 16359 17833
rect 16574 17824 16580 17836
rect 16632 17824 16638 17876
rect 16758 17864 16764 17876
rect 16719 17836 16764 17864
rect 16758 17824 16764 17836
rect 16816 17824 16822 17876
rect 17313 17867 17371 17873
rect 17313 17833 17325 17867
rect 17359 17864 17371 17867
rect 18693 17867 18751 17873
rect 18693 17864 18705 17867
rect 17359 17836 18705 17864
rect 17359 17833 17371 17836
rect 17313 17827 17371 17833
rect 18693 17833 18705 17836
rect 18739 17833 18751 17867
rect 18693 17827 18751 17833
rect 19521 17867 19579 17873
rect 19521 17833 19533 17867
rect 19567 17864 19579 17867
rect 19794 17864 19800 17876
rect 19567 17836 19800 17864
rect 19567 17833 19579 17836
rect 19521 17827 19579 17833
rect 19794 17824 19800 17836
rect 19852 17824 19858 17876
rect 10502 17796 10508 17808
rect 7892 17768 9812 17796
rect 9876 17768 10508 17796
rect 7892 17756 7898 17768
rect 9876 17728 9904 17768
rect 10502 17756 10508 17768
rect 10560 17756 10566 17808
rect 10689 17799 10747 17805
rect 10689 17765 10701 17799
rect 10735 17796 10747 17799
rect 13078 17796 13084 17808
rect 10735 17768 13084 17796
rect 10735 17765 10747 17768
rect 10689 17759 10747 17765
rect 13078 17756 13084 17768
rect 13136 17756 13142 17808
rect 13262 17756 13268 17808
rect 13320 17796 13326 17808
rect 13320 17768 13365 17796
rect 13320 17756 13326 17768
rect 13538 17756 13544 17808
rect 13596 17796 13602 17808
rect 14461 17799 14519 17805
rect 14461 17796 14473 17799
rect 13596 17768 14473 17796
rect 13596 17756 13602 17768
rect 14461 17765 14473 17768
rect 14507 17765 14519 17799
rect 14461 17759 14519 17765
rect 15102 17756 15108 17808
rect 15160 17796 15166 17808
rect 17681 17799 17739 17805
rect 17681 17796 17693 17799
rect 15160 17768 16528 17796
rect 15160 17756 15166 17768
rect 10042 17728 10048 17740
rect 7524 17700 7604 17728
rect 7668 17700 9904 17728
rect 10003 17700 10048 17728
rect 7524 17688 7530 17700
rect 2774 17660 2780 17672
rect 1504 17632 2780 17660
rect 2774 17620 2780 17632
rect 2832 17620 2838 17672
rect 3602 17660 3608 17672
rect 3563 17632 3608 17660
rect 3602 17620 3608 17632
rect 3660 17620 3666 17672
rect 4154 17620 4160 17672
rect 4212 17660 4218 17672
rect 4614 17660 4620 17672
rect 4212 17632 4620 17660
rect 4212 17620 4218 17632
rect 4614 17620 4620 17632
rect 4672 17620 4678 17672
rect 5074 17660 5080 17672
rect 5035 17632 5080 17660
rect 5074 17620 5080 17632
rect 5132 17620 5138 17672
rect 5166 17620 5172 17672
rect 5224 17660 5230 17672
rect 5445 17663 5503 17669
rect 5445 17660 5457 17663
rect 5224 17632 5457 17660
rect 5224 17620 5230 17632
rect 5445 17629 5457 17632
rect 5491 17629 5503 17663
rect 7668 17660 7696 17700
rect 10042 17688 10048 17700
rect 10100 17688 10106 17740
rect 10778 17688 10784 17740
rect 10836 17728 10842 17740
rect 11149 17731 11207 17737
rect 11149 17728 11161 17731
rect 10836 17700 11161 17728
rect 10836 17688 10842 17700
rect 11149 17697 11161 17700
rect 11195 17697 11207 17731
rect 11149 17691 11207 17697
rect 11416 17731 11474 17737
rect 11416 17697 11428 17731
rect 11462 17728 11474 17731
rect 11698 17728 11704 17740
rect 11462 17700 11704 17728
rect 11462 17697 11474 17700
rect 11416 17691 11474 17697
rect 11698 17688 11704 17700
rect 11756 17728 11762 17740
rect 11756 17700 13492 17728
rect 11756 17688 11762 17700
rect 5445 17623 5503 17629
rect 6472 17632 7696 17660
rect 2961 17595 3019 17601
rect 2961 17561 2973 17595
rect 3007 17592 3019 17595
rect 4706 17592 4712 17604
rect 3007 17564 4712 17592
rect 3007 17561 3019 17564
rect 2961 17555 3019 17561
rect 4706 17552 4712 17564
rect 4764 17552 4770 17604
rect 2866 17484 2872 17536
rect 2924 17524 2930 17536
rect 5258 17524 5264 17536
rect 2924 17496 5264 17524
rect 2924 17484 2930 17496
rect 5258 17484 5264 17496
rect 5316 17484 5322 17536
rect 5442 17484 5448 17536
rect 5500 17524 5506 17536
rect 6472 17524 6500 17632
rect 7742 17620 7748 17672
rect 7800 17660 7806 17672
rect 7929 17663 7987 17669
rect 7800 17632 7845 17660
rect 7800 17620 7806 17632
rect 7929 17629 7941 17663
rect 7975 17629 7987 17663
rect 8938 17660 8944 17672
rect 8899 17632 8944 17660
rect 7929 17623 7987 17629
rect 6825 17595 6883 17601
rect 6825 17561 6837 17595
rect 6871 17592 6883 17595
rect 7944 17592 7972 17623
rect 8938 17620 8944 17632
rect 8996 17620 9002 17672
rect 9030 17620 9036 17672
rect 9088 17660 9094 17672
rect 9214 17660 9220 17672
rect 9088 17632 9220 17660
rect 9088 17620 9094 17632
rect 9214 17620 9220 17632
rect 9272 17620 9278 17672
rect 9398 17620 9404 17672
rect 9456 17660 9462 17672
rect 10137 17663 10195 17669
rect 10137 17660 10149 17663
rect 9456 17632 10149 17660
rect 9456 17620 9462 17632
rect 10137 17629 10149 17632
rect 10183 17629 10195 17663
rect 10137 17623 10195 17629
rect 10229 17663 10287 17669
rect 10229 17629 10241 17663
rect 10275 17629 10287 17663
rect 10229 17623 10287 17629
rect 9048 17592 9076 17620
rect 6871 17564 7880 17592
rect 7944 17564 9076 17592
rect 6871 17561 6883 17564
rect 6825 17555 6883 17561
rect 5500 17496 6500 17524
rect 5500 17484 5506 17496
rect 6638 17484 6644 17536
rect 6696 17524 6702 17536
rect 7101 17527 7159 17533
rect 7101 17524 7113 17527
rect 6696 17496 7113 17524
rect 6696 17484 6702 17496
rect 7101 17493 7113 17496
rect 7147 17524 7159 17527
rect 7742 17524 7748 17536
rect 7147 17496 7748 17524
rect 7147 17493 7159 17496
rect 7101 17487 7159 17493
rect 7742 17484 7748 17496
rect 7800 17484 7806 17536
rect 7852 17524 7880 17564
rect 9122 17552 9128 17604
rect 9180 17592 9186 17604
rect 10244 17592 10272 17623
rect 12250 17620 12256 17672
rect 12308 17660 12314 17672
rect 13357 17663 13415 17669
rect 13357 17660 13369 17663
rect 12308 17632 13369 17660
rect 12308 17620 12314 17632
rect 13357 17629 13369 17632
rect 13403 17629 13415 17663
rect 13357 17623 13415 17629
rect 9180 17564 10272 17592
rect 13464 17592 13492 17700
rect 13906 17688 13912 17740
rect 13964 17728 13970 17740
rect 14369 17731 14427 17737
rect 14369 17728 14381 17731
rect 13964 17700 14381 17728
rect 13964 17688 13970 17700
rect 14369 17697 14381 17700
rect 14415 17697 14427 17731
rect 15654 17728 15660 17740
rect 15615 17700 15660 17728
rect 14369 17691 14427 17697
rect 15654 17688 15660 17700
rect 15712 17688 15718 17740
rect 15749 17731 15807 17737
rect 15749 17697 15761 17731
rect 15795 17728 15807 17731
rect 15930 17728 15936 17740
rect 15795 17700 15936 17728
rect 15795 17697 15807 17700
rect 15749 17691 15807 17697
rect 15930 17688 15936 17700
rect 15988 17688 15994 17740
rect 13814 17620 13820 17672
rect 13872 17660 13878 17672
rect 14553 17663 14611 17669
rect 14553 17660 14565 17663
rect 13872 17632 14565 17660
rect 13872 17620 13878 17632
rect 14553 17629 14565 17632
rect 14599 17660 14611 17663
rect 15010 17660 15016 17672
rect 14599 17632 15016 17660
rect 14599 17629 14611 17632
rect 14553 17623 14611 17629
rect 15010 17620 15016 17632
rect 15068 17620 15074 17672
rect 15841 17663 15899 17669
rect 15841 17629 15853 17663
rect 15887 17629 15899 17663
rect 15841 17623 15899 17629
rect 15856 17592 15884 17623
rect 13464 17564 15884 17592
rect 16500 17592 16528 17768
rect 16592 17768 17693 17796
rect 16592 17740 16620 17768
rect 17681 17765 17693 17768
rect 17727 17765 17739 17799
rect 19610 17796 19616 17808
rect 17681 17759 17739 17765
rect 17788 17768 19616 17796
rect 16574 17688 16580 17740
rect 16632 17688 16638 17740
rect 16669 17731 16727 17737
rect 16669 17697 16681 17731
rect 16715 17728 16727 17731
rect 16758 17728 16764 17740
rect 16715 17700 16764 17728
rect 16715 17697 16727 17700
rect 16669 17691 16727 17697
rect 16758 17688 16764 17700
rect 16816 17688 16822 17740
rect 17126 17688 17132 17740
rect 17184 17728 17190 17740
rect 17788 17728 17816 17768
rect 19610 17756 19616 17768
rect 19668 17756 19674 17808
rect 19978 17796 19984 17808
rect 19812 17768 19984 17796
rect 19812 17740 19840 17768
rect 19978 17756 19984 17768
rect 20036 17756 20042 17808
rect 19702 17728 19708 17740
rect 17184 17700 17816 17728
rect 17880 17700 19708 17728
rect 17184 17688 17190 17700
rect 16850 17620 16856 17672
rect 16908 17660 16914 17672
rect 17770 17660 17776 17672
rect 16908 17632 16953 17660
rect 17731 17632 17776 17660
rect 16908 17620 16914 17632
rect 17770 17620 17776 17632
rect 17828 17620 17834 17672
rect 17880 17669 17908 17700
rect 19702 17688 19708 17700
rect 19760 17688 19766 17740
rect 19794 17688 19800 17740
rect 19852 17688 19858 17740
rect 19889 17731 19947 17737
rect 19889 17697 19901 17731
rect 19935 17728 19947 17731
rect 20162 17728 20168 17740
rect 19935 17700 20168 17728
rect 19935 17697 19947 17700
rect 19889 17691 19947 17697
rect 20162 17688 20168 17700
rect 20220 17688 20226 17740
rect 17865 17663 17923 17669
rect 17865 17629 17877 17663
rect 17911 17629 17923 17663
rect 18782 17660 18788 17672
rect 18743 17632 18788 17660
rect 17865 17623 17923 17629
rect 18782 17620 18788 17632
rect 18840 17620 18846 17672
rect 18966 17660 18972 17672
rect 18927 17632 18972 17660
rect 18966 17620 18972 17632
rect 19024 17660 19030 17672
rect 19978 17660 19984 17672
rect 19024 17632 19840 17660
rect 19939 17632 19984 17660
rect 19024 17620 19030 17632
rect 18325 17595 18383 17601
rect 16500 17564 16804 17592
rect 9180 17552 9186 17564
rect 10502 17524 10508 17536
rect 7852 17496 10508 17524
rect 10502 17484 10508 17496
rect 10560 17484 10566 17536
rect 12529 17527 12587 17533
rect 12529 17493 12541 17527
rect 12575 17524 12587 17527
rect 12618 17524 12624 17536
rect 12575 17496 12624 17524
rect 12575 17493 12587 17496
rect 12529 17487 12587 17493
rect 12618 17484 12624 17496
rect 12676 17484 12682 17536
rect 16776 17524 16804 17564
rect 18325 17561 18337 17595
rect 18371 17592 18383 17595
rect 19334 17592 19340 17604
rect 18371 17564 19340 17592
rect 18371 17561 18383 17564
rect 18325 17555 18383 17561
rect 19334 17552 19340 17564
rect 19392 17552 19398 17604
rect 19812 17592 19840 17632
rect 19978 17620 19984 17632
rect 20036 17620 20042 17672
rect 20073 17663 20131 17669
rect 20073 17629 20085 17663
rect 20119 17629 20131 17663
rect 20073 17623 20131 17629
rect 20088 17592 20116 17623
rect 19812 17564 20116 17592
rect 20898 17524 20904 17536
rect 16776 17496 20904 17524
rect 20898 17484 20904 17496
rect 20956 17484 20962 17536
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 1489 17323 1547 17329
rect 1489 17289 1501 17323
rect 1535 17320 1547 17323
rect 3510 17320 3516 17332
rect 1535 17292 3516 17320
rect 1535 17289 1547 17292
rect 1489 17283 1547 17289
rect 3510 17280 3516 17292
rect 3568 17280 3574 17332
rect 3602 17280 3608 17332
rect 3660 17320 3666 17332
rect 3881 17323 3939 17329
rect 3881 17320 3893 17323
rect 3660 17292 3893 17320
rect 3660 17280 3666 17292
rect 3881 17289 3893 17292
rect 3927 17289 3939 17323
rect 5534 17320 5540 17332
rect 5495 17292 5540 17320
rect 3881 17283 3939 17289
rect 1946 17184 1952 17196
rect 1907 17156 1952 17184
rect 1946 17144 1952 17156
rect 2004 17144 2010 17196
rect 2130 17184 2136 17196
rect 2091 17156 2136 17184
rect 2130 17144 2136 17156
rect 2188 17144 2194 17196
rect 3896 17184 3924 17283
rect 5534 17280 5540 17292
rect 5592 17280 5598 17332
rect 6365 17323 6423 17329
rect 6365 17289 6377 17323
rect 6411 17320 6423 17323
rect 7834 17320 7840 17332
rect 6411 17292 7840 17320
rect 6411 17289 6423 17292
rect 6365 17283 6423 17289
rect 7834 17280 7840 17292
rect 7892 17280 7898 17332
rect 7929 17323 7987 17329
rect 7929 17289 7941 17323
rect 7975 17320 7987 17323
rect 8202 17320 8208 17332
rect 7975 17292 8208 17320
rect 7975 17289 7987 17292
rect 7929 17283 7987 17289
rect 8202 17280 8208 17292
rect 8260 17280 8266 17332
rect 8938 17280 8944 17332
rect 8996 17320 9002 17332
rect 9125 17323 9183 17329
rect 9125 17320 9137 17323
rect 8996 17292 9137 17320
rect 8996 17280 9002 17292
rect 9125 17289 9137 17292
rect 9171 17289 9183 17323
rect 9125 17283 9183 17289
rect 9214 17280 9220 17332
rect 9272 17320 9278 17332
rect 10965 17323 11023 17329
rect 10965 17320 10977 17323
rect 9272 17292 10977 17320
rect 9272 17280 9278 17292
rect 10965 17289 10977 17292
rect 11011 17289 11023 17323
rect 11146 17320 11152 17332
rect 11107 17292 11152 17320
rect 10965 17283 11023 17289
rect 11146 17280 11152 17292
rect 11204 17280 11210 17332
rect 13081 17323 13139 17329
rect 13081 17289 13093 17323
rect 13127 17320 13139 17323
rect 14182 17320 14188 17332
rect 13127 17292 14188 17320
rect 13127 17289 13139 17292
rect 13081 17283 13139 17289
rect 14182 17280 14188 17292
rect 14240 17280 14246 17332
rect 17310 17320 17316 17332
rect 14292 17292 17316 17320
rect 4065 17255 4123 17261
rect 4065 17221 4077 17255
rect 4111 17252 4123 17255
rect 4154 17252 4160 17264
rect 4111 17224 4160 17252
rect 4111 17221 4123 17224
rect 4065 17215 4123 17221
rect 4154 17212 4160 17224
rect 4212 17212 4218 17264
rect 5258 17212 5264 17264
rect 5316 17252 5322 17264
rect 10045 17255 10103 17261
rect 10045 17252 10057 17255
rect 5316 17224 10057 17252
rect 5316 17212 5322 17224
rect 10045 17221 10057 17224
rect 10091 17221 10103 17255
rect 10045 17215 10103 17221
rect 10137 17255 10195 17261
rect 10137 17221 10149 17255
rect 10183 17252 10195 17255
rect 11422 17252 11428 17264
rect 10183 17224 11428 17252
rect 10183 17221 10195 17224
rect 10137 17215 10195 17221
rect 11422 17212 11428 17224
rect 11480 17212 11486 17264
rect 11606 17212 11612 17264
rect 11664 17252 11670 17264
rect 14292 17252 14320 17292
rect 17310 17280 17316 17292
rect 17368 17280 17374 17332
rect 17589 17323 17647 17329
rect 17589 17289 17601 17323
rect 17635 17320 17647 17323
rect 17862 17320 17868 17332
rect 17635 17292 17868 17320
rect 17635 17289 17647 17292
rect 17589 17283 17647 17289
rect 17862 17280 17868 17292
rect 17920 17280 17926 17332
rect 17954 17280 17960 17332
rect 18012 17320 18018 17332
rect 19797 17323 19855 17329
rect 19797 17320 19809 17323
rect 18012 17292 19809 17320
rect 18012 17280 18018 17292
rect 19797 17289 19809 17292
rect 19843 17289 19855 17323
rect 19797 17283 19855 17289
rect 19889 17323 19947 17329
rect 19889 17289 19901 17323
rect 19935 17320 19947 17323
rect 20162 17320 20168 17332
rect 19935 17292 20168 17320
rect 19935 17289 19947 17292
rect 19889 17283 19947 17289
rect 20162 17280 20168 17292
rect 20220 17280 20226 17332
rect 11664 17224 14320 17252
rect 11664 17212 11670 17224
rect 18414 17212 18420 17264
rect 18472 17252 18478 17264
rect 18877 17255 18935 17261
rect 18472 17224 18644 17252
rect 18472 17212 18478 17224
rect 3896 17156 4292 17184
rect 1394 17076 1400 17128
rect 1452 17116 1458 17128
rect 1452 17088 2452 17116
rect 1452 17076 1458 17088
rect 1857 17051 1915 17057
rect 1857 17017 1869 17051
rect 1903 17048 1915 17051
rect 2424 17048 2452 17088
rect 2498 17076 2504 17128
rect 2556 17116 2562 17128
rect 2768 17119 2826 17125
rect 2556 17088 2601 17116
rect 2556 17076 2562 17088
rect 2768 17085 2780 17119
rect 2814 17116 2826 17119
rect 4065 17119 4123 17125
rect 4065 17116 4077 17119
rect 2814 17088 4077 17116
rect 2814 17085 2826 17088
rect 2768 17079 2826 17085
rect 4065 17085 4077 17088
rect 4111 17085 4123 17119
rect 4065 17079 4123 17085
rect 4157 17119 4215 17125
rect 4157 17085 4169 17119
rect 4203 17085 4215 17119
rect 4264 17116 4292 17156
rect 6546 17144 6552 17196
rect 6604 17184 6610 17196
rect 6914 17184 6920 17196
rect 6604 17156 6920 17184
rect 6604 17144 6610 17156
rect 6914 17144 6920 17156
rect 6972 17144 6978 17196
rect 7745 17187 7803 17193
rect 7745 17153 7757 17187
rect 7791 17153 7803 17187
rect 7745 17147 7803 17153
rect 8573 17187 8631 17193
rect 8573 17153 8585 17187
rect 8619 17184 8631 17187
rect 9122 17184 9128 17196
rect 8619 17156 9128 17184
rect 8619 17153 8631 17156
rect 8573 17147 8631 17153
rect 4413 17119 4471 17125
rect 4413 17116 4425 17119
rect 4264 17088 4425 17116
rect 4157 17079 4215 17085
rect 4413 17085 4425 17088
rect 4459 17085 4471 17119
rect 4413 17079 4471 17085
rect 6181 17119 6239 17125
rect 6181 17085 6193 17119
rect 6227 17116 6239 17119
rect 7006 17116 7012 17128
rect 6227 17088 7012 17116
rect 6227 17085 6239 17088
rect 6181 17079 6239 17085
rect 2958 17048 2964 17060
rect 1903 17020 2360 17048
rect 2424 17020 2964 17048
rect 1903 17017 1915 17020
rect 1857 17011 1915 17017
rect 2332 16980 2360 17020
rect 2958 17008 2964 17020
rect 3016 17008 3022 17060
rect 3142 17008 3148 17060
rect 3200 17048 3206 17060
rect 4172 17048 4200 17079
rect 7006 17076 7012 17088
rect 7064 17076 7070 17128
rect 7760 17060 7788 17147
rect 9122 17144 9128 17156
rect 9180 17184 9186 17196
rect 9677 17187 9735 17193
rect 9677 17184 9689 17187
rect 9180 17156 9689 17184
rect 9180 17144 9186 17156
rect 9677 17153 9689 17156
rect 9723 17153 9735 17187
rect 9677 17147 9735 17153
rect 10502 17144 10508 17196
rect 10560 17184 10566 17196
rect 10689 17187 10747 17193
rect 10689 17184 10701 17187
rect 10560 17156 10701 17184
rect 10560 17144 10566 17156
rect 10689 17153 10701 17156
rect 10735 17153 10747 17187
rect 10689 17147 10747 17153
rect 10965 17187 11023 17193
rect 10965 17153 10977 17187
rect 11011 17184 11023 17187
rect 11793 17187 11851 17193
rect 11011 17156 11744 17184
rect 11011 17153 11023 17156
rect 10965 17147 11023 17153
rect 9858 17116 9864 17128
rect 8220 17088 9864 17116
rect 5166 17048 5172 17060
rect 3200 17020 5172 17048
rect 3200 17008 3206 17020
rect 5166 17008 5172 17020
rect 5224 17008 5230 17060
rect 6914 17008 6920 17060
rect 6972 17048 6978 17060
rect 7561 17051 7619 17057
rect 7561 17048 7573 17051
rect 6972 17020 7573 17048
rect 6972 17008 6978 17020
rect 7561 17017 7573 17020
rect 7607 17017 7619 17051
rect 7561 17011 7619 17017
rect 7742 17008 7748 17060
rect 7800 17008 7806 17060
rect 2866 16980 2872 16992
rect 2332 16952 2872 16980
rect 2866 16940 2872 16952
rect 2924 16940 2930 16992
rect 3326 16940 3332 16992
rect 3384 16980 3390 16992
rect 4890 16980 4896 16992
rect 3384 16952 4896 16980
rect 3384 16940 3390 16952
rect 4890 16940 4896 16952
rect 4948 16940 4954 16992
rect 7098 16980 7104 16992
rect 7059 16952 7104 16980
rect 7098 16940 7104 16952
rect 7156 16940 7162 16992
rect 7469 16983 7527 16989
rect 7469 16949 7481 16983
rect 7515 16980 7527 16983
rect 8220 16980 8248 17088
rect 9858 17076 9864 17088
rect 9916 17076 9922 17128
rect 9950 17076 9956 17128
rect 10008 17116 10014 17128
rect 11609 17119 11667 17125
rect 11609 17116 11621 17119
rect 10008 17088 11621 17116
rect 10008 17076 10014 17088
rect 11609 17085 11621 17088
rect 11655 17085 11667 17119
rect 11716 17116 11744 17156
rect 11793 17153 11805 17187
rect 11839 17184 11851 17187
rect 12250 17184 12256 17196
rect 11839 17156 12256 17184
rect 11839 17153 11851 17156
rect 11793 17147 11851 17153
rect 12250 17144 12256 17156
rect 12308 17144 12314 17196
rect 13541 17187 13599 17193
rect 13541 17184 13553 17187
rect 12360 17156 13553 17184
rect 12360 17116 12388 17156
rect 13541 17153 13553 17156
rect 13587 17153 13599 17187
rect 13541 17147 13599 17153
rect 13725 17187 13783 17193
rect 13725 17153 13737 17187
rect 13771 17184 13783 17187
rect 13814 17184 13820 17196
rect 13771 17156 13820 17184
rect 13771 17153 13783 17156
rect 13725 17147 13783 17153
rect 13814 17144 13820 17156
rect 13872 17184 13878 17196
rect 14182 17184 14188 17196
rect 13872 17156 14188 17184
rect 13872 17144 13878 17156
rect 14182 17144 14188 17156
rect 14240 17144 14246 17196
rect 18616 17193 18644 17224
rect 18877 17221 18889 17255
rect 18923 17252 18935 17255
rect 18923 17224 20760 17252
rect 18923 17221 18935 17224
rect 18877 17215 18935 17221
rect 18601 17187 18659 17193
rect 18601 17153 18613 17187
rect 18647 17153 18659 17187
rect 18601 17147 18659 17153
rect 19334 17144 19340 17196
rect 19392 17184 19398 17196
rect 19429 17187 19487 17193
rect 19429 17184 19441 17187
rect 19392 17156 19441 17184
rect 19392 17144 19398 17156
rect 19429 17153 19441 17156
rect 19475 17153 19487 17187
rect 19429 17147 19487 17153
rect 19797 17187 19855 17193
rect 19797 17153 19809 17187
rect 19843 17184 19855 17187
rect 20349 17187 20407 17193
rect 20349 17184 20361 17187
rect 19843 17156 20361 17184
rect 19843 17153 19855 17156
rect 19797 17147 19855 17153
rect 20349 17153 20361 17156
rect 20395 17153 20407 17187
rect 20530 17184 20536 17196
rect 20491 17156 20536 17184
rect 20349 17147 20407 17153
rect 20530 17144 20536 17156
rect 20588 17144 20594 17196
rect 12526 17116 12532 17128
rect 11716 17088 12388 17116
rect 12487 17088 12532 17116
rect 11609 17079 11667 17085
rect 12526 17076 12532 17088
rect 12584 17076 12590 17128
rect 13354 17076 13360 17128
rect 13412 17116 13418 17128
rect 14274 17116 14280 17128
rect 13412 17088 14280 17116
rect 13412 17076 13418 17088
rect 14274 17076 14280 17088
rect 14332 17076 14338 17128
rect 14366 17076 14372 17128
rect 14424 17116 14430 17128
rect 14533 17119 14591 17125
rect 14533 17116 14545 17119
rect 14424 17088 14545 17116
rect 14424 17076 14430 17088
rect 14533 17085 14545 17088
rect 14579 17085 14591 17119
rect 14533 17079 14591 17085
rect 15010 17076 15016 17128
rect 15068 17116 15074 17128
rect 16206 17116 16212 17128
rect 15068 17088 15875 17116
rect 16167 17088 16212 17116
rect 15068 17076 15074 17088
rect 8297 17051 8355 17057
rect 8297 17017 8309 17051
rect 8343 17048 8355 17051
rect 8846 17048 8852 17060
rect 8343 17020 8852 17048
rect 8343 17017 8355 17020
rect 8297 17011 8355 17017
rect 8846 17008 8852 17020
rect 8904 17008 8910 17060
rect 9033 17051 9091 17057
rect 9033 17017 9045 17051
rect 9079 17048 9091 17051
rect 9398 17048 9404 17060
rect 9079 17020 9404 17048
rect 9079 17017 9091 17020
rect 9033 17011 9091 17017
rect 9398 17008 9404 17020
rect 9456 17048 9462 17060
rect 9585 17051 9643 17057
rect 9585 17048 9597 17051
rect 9456 17020 9597 17048
rect 9456 17008 9462 17020
rect 9585 17017 9597 17020
rect 9631 17017 9643 17051
rect 9585 17011 9643 17017
rect 10045 17051 10103 17057
rect 10045 17017 10057 17051
rect 10091 17048 10103 17051
rect 10597 17051 10655 17057
rect 10597 17048 10609 17051
rect 10091 17020 10609 17048
rect 10091 17017 10103 17020
rect 10045 17011 10103 17017
rect 10597 17017 10609 17020
rect 10643 17017 10655 17051
rect 10597 17011 10655 17017
rect 11517 17051 11575 17057
rect 11517 17017 11529 17051
rect 11563 17048 11575 17051
rect 13446 17048 13452 17060
rect 11563 17020 12020 17048
rect 13407 17020 13452 17048
rect 11563 17017 11575 17020
rect 11517 17011 11575 17017
rect 7515 16952 8248 16980
rect 8389 16983 8447 16989
rect 7515 16949 7527 16952
rect 7469 16943 7527 16949
rect 8389 16949 8401 16983
rect 8435 16980 8447 16983
rect 8478 16980 8484 16992
rect 8435 16952 8484 16980
rect 8435 16949 8447 16952
rect 8389 16943 8447 16949
rect 8478 16940 8484 16952
rect 8536 16940 8542 16992
rect 9490 16980 9496 16992
rect 9451 16952 9496 16980
rect 9490 16940 9496 16952
rect 9548 16940 9554 16992
rect 9674 16940 9680 16992
rect 9732 16980 9738 16992
rect 10505 16983 10563 16989
rect 10505 16980 10517 16983
rect 9732 16952 10517 16980
rect 9732 16940 9738 16952
rect 10505 16949 10517 16952
rect 10551 16949 10563 16983
rect 11992 16980 12020 17020
rect 13446 17008 13452 17020
rect 13504 17008 13510 17060
rect 15847 17048 15875 17088
rect 16206 17076 16212 17088
rect 16264 17076 16270 17128
rect 16476 17119 16534 17125
rect 16476 17085 16488 17119
rect 16522 17116 16534 17119
rect 16850 17116 16856 17128
rect 16522 17088 16856 17116
rect 16522 17085 16534 17088
rect 16476 17079 16534 17085
rect 16850 17076 16856 17088
rect 16908 17076 16914 17128
rect 16942 17076 16948 17128
rect 17000 17116 17006 17128
rect 19242 17116 19248 17128
rect 17000 17088 19248 17116
rect 17000 17076 17006 17088
rect 19242 17076 19248 17088
rect 19300 17076 19306 17128
rect 20732 17125 20760 17224
rect 20898 17184 20904 17196
rect 20859 17156 20904 17184
rect 20898 17144 20904 17156
rect 20956 17144 20962 17196
rect 20717 17119 20775 17125
rect 20717 17085 20729 17119
rect 20763 17085 20775 17119
rect 20717 17079 20775 17085
rect 18322 17048 18328 17060
rect 15488 17020 15792 17048
rect 15847 17020 18328 17048
rect 12434 16980 12440 16992
rect 11992 16952 12440 16980
rect 10505 16943 10563 16949
rect 12434 16940 12440 16952
rect 12492 16940 12498 16992
rect 12713 16983 12771 16989
rect 12713 16949 12725 16983
rect 12759 16980 12771 16983
rect 15488 16980 15516 17020
rect 12759 16952 15516 16980
rect 12759 16949 12771 16952
rect 12713 16943 12771 16949
rect 15562 16940 15568 16992
rect 15620 16980 15626 16992
rect 15657 16983 15715 16989
rect 15657 16980 15669 16983
rect 15620 16952 15669 16980
rect 15620 16940 15626 16952
rect 15657 16949 15669 16952
rect 15703 16949 15715 16983
rect 15764 16980 15792 17020
rect 18322 17008 18328 17020
rect 18380 17008 18386 17060
rect 18417 17051 18475 17057
rect 18417 17017 18429 17051
rect 18463 17048 18475 17051
rect 20257 17051 20315 17057
rect 18463 17020 18644 17048
rect 18463 17017 18475 17020
rect 18417 17011 18475 17017
rect 17126 16980 17132 16992
rect 15764 16952 17132 16980
rect 15657 16943 15715 16949
rect 17126 16940 17132 16952
rect 17184 16940 17190 16992
rect 18046 16980 18052 16992
rect 18007 16952 18052 16980
rect 18046 16940 18052 16952
rect 18104 16940 18110 16992
rect 18138 16940 18144 16992
rect 18196 16980 18202 16992
rect 18509 16983 18567 16989
rect 18509 16980 18521 16983
rect 18196 16952 18521 16980
rect 18196 16940 18202 16952
rect 18509 16949 18521 16952
rect 18555 16949 18567 16983
rect 18616 16980 18644 17020
rect 20257 17017 20269 17051
rect 20303 17048 20315 17051
rect 20806 17048 20812 17060
rect 20303 17020 20812 17048
rect 20303 17017 20315 17020
rect 20257 17011 20315 17017
rect 20806 17008 20812 17020
rect 20864 17008 20870 17060
rect 18874 16980 18880 16992
rect 18616 16952 18880 16980
rect 18509 16943 18567 16949
rect 18874 16940 18880 16952
rect 18932 16940 18938 16992
rect 19242 16980 19248 16992
rect 19203 16952 19248 16980
rect 19242 16940 19248 16952
rect 19300 16940 19306 16992
rect 19334 16940 19340 16992
rect 19392 16980 19398 16992
rect 19392 16952 19437 16980
rect 19392 16940 19398 16952
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 1578 16776 1584 16788
rect 1539 16748 1584 16776
rect 1578 16736 1584 16748
rect 1636 16736 1642 16788
rect 1949 16779 2007 16785
rect 1949 16745 1961 16779
rect 1995 16745 2007 16779
rect 2314 16776 2320 16788
rect 2275 16748 2320 16776
rect 1949 16739 2007 16745
rect 198 16668 204 16720
rect 256 16708 262 16720
rect 1964 16708 1992 16739
rect 2314 16736 2320 16748
rect 2372 16736 2378 16788
rect 2406 16736 2412 16788
rect 2464 16776 2470 16788
rect 2774 16776 2780 16788
rect 2464 16748 2780 16776
rect 2464 16736 2470 16748
rect 2774 16736 2780 16748
rect 2832 16736 2838 16788
rect 3329 16779 3387 16785
rect 3329 16745 3341 16779
rect 3375 16776 3387 16779
rect 4065 16779 4123 16785
rect 4065 16776 4077 16779
rect 3375 16748 4077 16776
rect 3375 16745 3387 16748
rect 3329 16739 3387 16745
rect 4065 16745 4077 16748
rect 4111 16745 4123 16779
rect 4065 16739 4123 16745
rect 4246 16736 4252 16788
rect 4304 16776 4310 16788
rect 4525 16779 4583 16785
rect 4525 16776 4537 16779
rect 4304 16748 4537 16776
rect 4304 16736 4310 16748
rect 4525 16745 4537 16748
rect 4571 16745 4583 16779
rect 5442 16776 5448 16788
rect 5403 16748 5448 16776
rect 4525 16739 4583 16745
rect 5442 16736 5448 16748
rect 5500 16736 5506 16788
rect 5905 16779 5963 16785
rect 5905 16745 5917 16779
rect 5951 16776 5963 16779
rect 7098 16776 7104 16788
rect 5951 16748 7104 16776
rect 5951 16745 5963 16748
rect 5905 16739 5963 16745
rect 7098 16736 7104 16748
rect 7156 16736 7162 16788
rect 7466 16776 7472 16788
rect 7427 16748 7472 16776
rect 7466 16736 7472 16748
rect 7524 16736 7530 16788
rect 7745 16779 7803 16785
rect 7745 16745 7757 16779
rect 7791 16776 7803 16779
rect 8570 16776 8576 16788
rect 7791 16748 8576 16776
rect 7791 16745 7803 16748
rect 7745 16739 7803 16745
rect 8570 16736 8576 16748
rect 8628 16736 8634 16788
rect 9122 16736 9128 16788
rect 9180 16776 9186 16788
rect 9309 16779 9367 16785
rect 9309 16776 9321 16779
rect 9180 16748 9321 16776
rect 9180 16736 9186 16748
rect 9309 16745 9321 16748
rect 9355 16745 9367 16779
rect 9309 16739 9367 16745
rect 9953 16779 10011 16785
rect 9953 16745 9965 16779
rect 9999 16745 10011 16779
rect 11698 16776 11704 16788
rect 11659 16748 11704 16776
rect 9953 16739 10011 16745
rect 3421 16711 3479 16717
rect 256 16680 1900 16708
rect 1964 16680 3372 16708
rect 256 16668 262 16680
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 1872 16640 1900 16680
rect 3344 16640 3372 16680
rect 3421 16677 3433 16711
rect 3467 16708 3479 16711
rect 4706 16708 4712 16720
rect 3467 16680 4712 16708
rect 3467 16677 3479 16680
rect 3421 16671 3479 16677
rect 4706 16668 4712 16680
rect 4764 16668 4770 16720
rect 5813 16711 5871 16717
rect 5813 16677 5825 16711
rect 5859 16708 5871 16711
rect 7650 16708 7656 16720
rect 5859 16680 7656 16708
rect 5859 16677 5871 16680
rect 5813 16671 5871 16677
rect 7650 16668 7656 16680
rect 7708 16668 7714 16720
rect 9674 16708 9680 16720
rect 7751 16680 9680 16708
rect 1872 16612 2268 16640
rect 3344 16612 4108 16640
rect 2240 16572 2268 16612
rect 2406 16572 2412 16584
rect 2240 16544 2412 16572
rect 2406 16532 2412 16544
rect 2464 16532 2470 16584
rect 2593 16575 2651 16581
rect 2593 16541 2605 16575
rect 2639 16572 2651 16575
rect 3602 16572 3608 16584
rect 2639 16544 3464 16572
rect 3563 16544 3608 16572
rect 2639 16541 2651 16544
rect 2593 16535 2651 16541
rect 2961 16507 3019 16513
rect 2961 16473 2973 16507
rect 3007 16504 3019 16507
rect 3326 16504 3332 16516
rect 3007 16476 3332 16504
rect 3007 16473 3019 16476
rect 2961 16467 3019 16473
rect 3326 16464 3332 16476
rect 3384 16464 3390 16516
rect 3436 16436 3464 16544
rect 3602 16532 3608 16544
rect 3660 16532 3666 16584
rect 4080 16504 4108 16612
rect 4154 16600 4160 16652
rect 4212 16640 4218 16652
rect 4433 16643 4491 16649
rect 4433 16640 4445 16643
rect 4212 16612 4445 16640
rect 4212 16600 4218 16612
rect 4433 16609 4445 16612
rect 4479 16609 4491 16643
rect 4433 16603 4491 16609
rect 6730 16600 6736 16652
rect 6788 16640 6794 16652
rect 6825 16643 6883 16649
rect 6825 16640 6837 16643
rect 6788 16612 6837 16640
rect 6788 16600 6794 16612
rect 6825 16609 6837 16612
rect 6871 16609 6883 16643
rect 7751 16640 7779 16680
rect 9674 16668 9680 16680
rect 9732 16668 9738 16720
rect 9968 16708 9996 16739
rect 11698 16736 11704 16748
rect 11756 16736 11762 16788
rect 11882 16736 11888 16788
rect 11940 16776 11946 16788
rect 12069 16779 12127 16785
rect 12069 16776 12081 16779
rect 11940 16748 12081 16776
rect 11940 16736 11946 16748
rect 12069 16745 12081 16748
rect 12115 16745 12127 16779
rect 15010 16776 15016 16788
rect 12069 16739 12127 16745
rect 12176 16748 15016 16776
rect 11514 16708 11520 16720
rect 9968 16680 11520 16708
rect 11514 16668 11520 16680
rect 11572 16668 11578 16720
rect 8202 16649 8208 16652
rect 8185 16643 8208 16649
rect 8185 16640 8197 16643
rect 6825 16603 6883 16609
rect 6932 16612 7779 16640
rect 7852 16612 8197 16640
rect 4338 16532 4344 16584
rect 4396 16572 4402 16584
rect 4617 16575 4675 16581
rect 4617 16572 4629 16575
rect 4396 16544 4629 16572
rect 4396 16532 4402 16544
rect 4617 16541 4629 16544
rect 4663 16572 4675 16575
rect 5258 16572 5264 16584
rect 4663 16544 5264 16572
rect 4663 16541 4675 16544
rect 4617 16535 4675 16541
rect 5258 16532 5264 16544
rect 5316 16532 5322 16584
rect 6089 16575 6147 16581
rect 6089 16541 6101 16575
rect 6135 16541 6147 16575
rect 6089 16535 6147 16541
rect 5534 16504 5540 16516
rect 4080 16476 5540 16504
rect 5534 16464 5540 16476
rect 5592 16464 5598 16516
rect 6104 16504 6132 16535
rect 6454 16532 6460 16584
rect 6512 16572 6518 16584
rect 6932 16581 6960 16612
rect 6917 16575 6975 16581
rect 6917 16572 6929 16575
rect 6512 16544 6929 16572
rect 6512 16532 6518 16544
rect 6917 16541 6929 16544
rect 6963 16541 6975 16575
rect 7098 16572 7104 16584
rect 7011 16544 7104 16572
rect 6917 16535 6975 16541
rect 7098 16532 7104 16544
rect 7156 16572 7162 16584
rect 7745 16575 7803 16581
rect 7745 16572 7757 16575
rect 7156 16544 7757 16572
rect 7156 16532 7162 16544
rect 7745 16541 7757 16544
rect 7791 16541 7803 16575
rect 7745 16535 7803 16541
rect 7852 16504 7880 16612
rect 8185 16609 8197 16612
rect 8260 16640 8266 16652
rect 8260 16612 8333 16640
rect 8185 16603 8208 16609
rect 8202 16600 8208 16603
rect 8260 16600 8266 16612
rect 8478 16600 8484 16652
rect 8536 16640 8542 16652
rect 9122 16640 9128 16652
rect 8536 16612 9128 16640
rect 8536 16600 8542 16612
rect 9122 16600 9128 16612
rect 9180 16640 9186 16652
rect 9769 16643 9827 16649
rect 9769 16640 9781 16643
rect 9180 16612 9781 16640
rect 9180 16600 9186 16612
rect 9769 16609 9781 16612
rect 9815 16609 9827 16643
rect 9769 16603 9827 16609
rect 10321 16643 10379 16649
rect 10321 16609 10333 16643
rect 10367 16640 10379 16643
rect 10410 16640 10416 16652
rect 10367 16612 10416 16640
rect 10367 16609 10379 16612
rect 10321 16603 10379 16609
rect 10410 16600 10416 16612
rect 10468 16600 10474 16652
rect 10588 16643 10646 16649
rect 10588 16609 10600 16643
rect 10634 16640 10646 16643
rect 11146 16640 11152 16652
rect 10634 16612 11152 16640
rect 10634 16609 10646 16612
rect 10588 16603 10646 16609
rect 11146 16600 11152 16612
rect 11204 16600 11210 16652
rect 12066 16600 12072 16652
rect 12124 16640 12130 16652
rect 12176 16640 12204 16748
rect 15010 16736 15016 16748
rect 15068 16736 15074 16788
rect 16669 16779 16727 16785
rect 16669 16745 16681 16779
rect 16715 16776 16727 16779
rect 16850 16776 16856 16788
rect 16715 16748 16856 16776
rect 16715 16745 16727 16748
rect 16669 16739 16727 16745
rect 16850 16736 16856 16748
rect 16908 16736 16914 16788
rect 17402 16736 17408 16788
rect 17460 16776 17466 16788
rect 17460 16748 17540 16776
rect 17460 16736 17466 16748
rect 14366 16668 14372 16720
rect 14424 16668 14430 16720
rect 15838 16708 15844 16720
rect 14844 16680 15844 16708
rect 12124 16612 12204 16640
rect 12437 16643 12495 16649
rect 12124 16600 12130 16612
rect 12437 16609 12449 16643
rect 12483 16640 12495 16643
rect 13262 16640 13268 16652
rect 12483 16612 13268 16640
rect 12483 16609 12495 16612
rect 12437 16603 12495 16609
rect 13262 16600 13268 16612
rect 13320 16600 13326 16652
rect 13354 16600 13360 16652
rect 13412 16640 13418 16652
rect 13449 16643 13507 16649
rect 13449 16640 13461 16643
rect 13412 16612 13461 16640
rect 13412 16600 13418 16612
rect 13449 16609 13461 16612
rect 13495 16609 13507 16643
rect 13449 16603 13507 16609
rect 13716 16643 13774 16649
rect 13716 16609 13728 16643
rect 13762 16640 13774 16643
rect 14182 16640 14188 16652
rect 13762 16612 14188 16640
rect 13762 16609 13774 16612
rect 13716 16603 13774 16609
rect 14182 16600 14188 16612
rect 14240 16600 14246 16652
rect 14384 16640 14412 16668
rect 14844 16640 14872 16680
rect 15838 16668 15844 16680
rect 15896 16668 15902 16720
rect 17037 16711 17095 16717
rect 17037 16677 17049 16711
rect 17083 16708 17095 16711
rect 17126 16708 17132 16720
rect 17083 16680 17132 16708
rect 17083 16677 17095 16680
rect 17037 16671 17095 16677
rect 17126 16668 17132 16680
rect 17184 16668 17190 16720
rect 15562 16649 15568 16652
rect 14384 16612 14872 16640
rect 7929 16575 7987 16581
rect 7929 16541 7941 16575
rect 7975 16541 7987 16575
rect 12526 16572 12532 16584
rect 12487 16544 12532 16572
rect 7929 16535 7987 16541
rect 6104 16476 7880 16504
rect 6178 16436 6184 16448
rect 3436 16408 6184 16436
rect 6178 16396 6184 16408
rect 6236 16396 6242 16448
rect 6454 16436 6460 16448
rect 6415 16408 6460 16436
rect 6454 16396 6460 16408
rect 6512 16396 6518 16448
rect 7558 16396 7564 16448
rect 7616 16436 7622 16448
rect 7944 16436 7972 16535
rect 12526 16532 12532 16544
rect 12584 16532 12590 16584
rect 12618 16532 12624 16584
rect 12676 16572 12682 16584
rect 12676 16544 12721 16572
rect 12676 16532 12682 16544
rect 11422 16464 11428 16516
rect 11480 16504 11486 16516
rect 12434 16504 12440 16516
rect 11480 16476 12440 16504
rect 11480 16464 11486 16476
rect 12434 16464 12440 16476
rect 12492 16464 12498 16516
rect 14844 16513 14872 16612
rect 15556 16603 15568 16649
rect 15620 16640 15626 16652
rect 17512 16649 17540 16748
rect 17770 16736 17776 16788
rect 17828 16776 17834 16788
rect 18141 16779 18199 16785
rect 18141 16776 18153 16779
rect 17828 16748 18153 16776
rect 17828 16736 17834 16748
rect 18141 16745 18153 16748
rect 18187 16745 18199 16779
rect 18141 16739 18199 16745
rect 18230 16736 18236 16788
rect 18288 16776 18294 16788
rect 18506 16776 18512 16788
rect 18288 16748 18512 16776
rect 18288 16736 18294 16748
rect 18506 16736 18512 16748
rect 18564 16776 18570 16788
rect 18601 16779 18659 16785
rect 18601 16776 18613 16779
rect 18564 16748 18613 16776
rect 18564 16736 18570 16748
rect 18601 16745 18613 16748
rect 18647 16745 18659 16779
rect 18601 16739 18659 16745
rect 18782 16736 18788 16788
rect 18840 16776 18846 16788
rect 19153 16779 19211 16785
rect 19153 16776 19165 16779
rect 18840 16748 19165 16776
rect 18840 16736 18846 16748
rect 19153 16745 19165 16748
rect 19199 16745 19211 16779
rect 19978 16776 19984 16788
rect 19939 16748 19984 16776
rect 19153 16739 19211 16745
rect 19978 16736 19984 16748
rect 20036 16736 20042 16788
rect 21085 16779 21143 16785
rect 21085 16776 21097 16779
rect 20272 16748 21097 16776
rect 18046 16668 18052 16720
rect 18104 16708 18110 16720
rect 19521 16711 19579 16717
rect 19521 16708 19533 16711
rect 18104 16680 19533 16708
rect 18104 16668 18110 16680
rect 19521 16677 19533 16680
rect 19567 16677 19579 16711
rect 19521 16671 19579 16677
rect 17497 16643 17555 16649
rect 15620 16612 15656 16640
rect 15562 16600 15568 16603
rect 15620 16600 15626 16612
rect 17497 16609 17509 16643
rect 17543 16609 17555 16643
rect 17497 16603 17555 16609
rect 17589 16643 17647 16649
rect 17589 16609 17601 16643
rect 17635 16640 17647 16643
rect 17770 16640 17776 16652
rect 17635 16612 17776 16640
rect 17635 16609 17647 16612
rect 17589 16603 17647 16609
rect 15289 16575 15347 16581
rect 15289 16541 15301 16575
rect 15335 16541 15347 16575
rect 15289 16535 15347 16541
rect 14829 16507 14887 16513
rect 14829 16473 14841 16507
rect 14875 16473 14887 16507
rect 14829 16467 14887 16473
rect 9674 16436 9680 16448
rect 7616 16408 9680 16436
rect 7616 16396 7622 16408
rect 9674 16396 9680 16408
rect 9732 16396 9738 16448
rect 11882 16396 11888 16448
rect 11940 16436 11946 16448
rect 14918 16436 14924 16448
rect 11940 16408 14924 16436
rect 11940 16396 11946 16408
rect 14918 16396 14924 16408
rect 14976 16396 14982 16448
rect 15304 16436 15332 16535
rect 17310 16532 17316 16584
rect 17368 16572 17374 16584
rect 17512 16572 17540 16603
rect 17770 16600 17776 16612
rect 17828 16600 17834 16652
rect 18506 16640 18512 16652
rect 18467 16612 18512 16640
rect 18506 16600 18512 16612
rect 18564 16600 18570 16652
rect 19058 16600 19064 16652
rect 19116 16640 19122 16652
rect 20272 16640 20300 16748
rect 21085 16745 21097 16748
rect 21131 16745 21143 16779
rect 21085 16739 21143 16745
rect 20441 16711 20499 16717
rect 20441 16677 20453 16711
rect 20487 16708 20499 16711
rect 21358 16708 21364 16720
rect 20487 16680 21364 16708
rect 20487 16677 20499 16680
rect 20441 16671 20499 16677
rect 21358 16668 21364 16680
rect 21416 16668 21422 16720
rect 19116 16612 20300 16640
rect 20349 16643 20407 16649
rect 19116 16600 19122 16612
rect 20349 16609 20361 16643
rect 20395 16640 20407 16643
rect 20898 16640 20904 16652
rect 20395 16612 20668 16640
rect 20859 16612 20904 16640
rect 20395 16609 20407 16612
rect 20349 16603 20407 16609
rect 17368 16544 17540 16572
rect 17681 16575 17739 16581
rect 17368 16532 17374 16544
rect 17681 16541 17693 16575
rect 17727 16572 17739 16575
rect 17727 16544 17816 16572
rect 17727 16541 17739 16544
rect 17681 16535 17739 16541
rect 17788 16516 17816 16544
rect 18414 16532 18420 16584
rect 18472 16572 18478 16584
rect 18782 16572 18788 16584
rect 18472 16544 18788 16572
rect 18472 16532 18478 16544
rect 18782 16532 18788 16544
rect 18840 16532 18846 16584
rect 19610 16572 19616 16584
rect 19571 16544 19616 16572
rect 19610 16532 19616 16544
rect 19668 16532 19674 16584
rect 19702 16532 19708 16584
rect 19760 16572 19766 16584
rect 19797 16575 19855 16581
rect 19797 16572 19809 16575
rect 19760 16544 19809 16572
rect 19760 16532 19766 16544
rect 19797 16541 19809 16544
rect 19843 16572 19855 16575
rect 20530 16572 20536 16584
rect 19843 16544 20536 16572
rect 19843 16541 19855 16544
rect 19797 16535 19855 16541
rect 20530 16532 20536 16544
rect 20588 16532 20594 16584
rect 16574 16464 16580 16516
rect 16632 16504 16638 16516
rect 17129 16507 17187 16513
rect 17129 16504 17141 16507
rect 16632 16476 17141 16504
rect 16632 16464 16638 16476
rect 17129 16473 17141 16476
rect 17175 16473 17187 16507
rect 17129 16467 17187 16473
rect 17770 16464 17776 16516
rect 17828 16464 17834 16516
rect 16206 16436 16212 16448
rect 15304 16408 16212 16436
rect 16206 16396 16212 16408
rect 16264 16396 16270 16448
rect 16850 16396 16856 16448
rect 16908 16436 16914 16448
rect 20640 16436 20668 16612
rect 20898 16600 20904 16612
rect 20956 16600 20962 16652
rect 16908 16408 20668 16436
rect 16908 16396 16914 16408
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 1670 16232 1676 16244
rect 1631 16204 1676 16232
rect 1670 16192 1676 16204
rect 1728 16192 1734 16244
rect 2498 16192 2504 16244
rect 2556 16232 2562 16244
rect 4706 16232 4712 16244
rect 2556 16204 3096 16232
rect 4667 16204 4712 16232
rect 2556 16192 2562 16204
rect 2041 16167 2099 16173
rect 2041 16133 2053 16167
rect 2087 16164 2099 16167
rect 2087 16136 2636 16164
rect 2087 16133 2099 16136
rect 2041 16127 2099 16133
rect 1489 16031 1547 16037
rect 1489 15997 1501 16031
rect 1535 16028 1547 16031
rect 1670 16028 1676 16040
rect 1535 16000 1676 16028
rect 1535 15997 1547 16000
rect 1489 15991 1547 15997
rect 1670 15988 1676 16000
rect 1728 15988 1734 16040
rect 2498 15960 2504 15972
rect 2459 15932 2504 15960
rect 2498 15920 2504 15932
rect 2556 15920 2562 15972
rect 2608 15960 2636 16136
rect 2685 16099 2743 16105
rect 2685 16065 2697 16099
rect 2731 16096 2743 16099
rect 2774 16096 2780 16108
rect 2731 16068 2780 16096
rect 2731 16065 2743 16068
rect 2685 16059 2743 16065
rect 2774 16056 2780 16068
rect 2832 16056 2838 16108
rect 3068 16037 3096 16204
rect 4706 16192 4712 16204
rect 4764 16192 4770 16244
rect 5721 16235 5779 16241
rect 5721 16201 5733 16235
rect 5767 16232 5779 16235
rect 6914 16232 6920 16244
rect 5767 16204 6920 16232
rect 5767 16201 5779 16204
rect 5721 16195 5779 16201
rect 6914 16192 6920 16204
rect 6972 16192 6978 16244
rect 7006 16192 7012 16244
rect 7064 16232 7070 16244
rect 7466 16232 7472 16244
rect 7064 16204 7472 16232
rect 7064 16192 7070 16204
rect 7466 16192 7472 16204
rect 7524 16232 7530 16244
rect 8110 16232 8116 16244
rect 7524 16204 8116 16232
rect 7524 16192 7530 16204
rect 8110 16192 8116 16204
rect 8168 16192 8174 16244
rect 8202 16192 8208 16244
rect 8260 16232 8266 16244
rect 8849 16235 8907 16241
rect 8849 16232 8861 16235
rect 8260 16204 8861 16232
rect 8260 16192 8266 16204
rect 8849 16201 8861 16204
rect 8895 16201 8907 16235
rect 8849 16195 8907 16201
rect 8938 16192 8944 16244
rect 8996 16232 9002 16244
rect 8996 16204 10916 16232
rect 8996 16192 9002 16204
rect 4433 16167 4491 16173
rect 4433 16133 4445 16167
rect 4479 16164 4491 16167
rect 4479 16136 5304 16164
rect 4479 16133 4491 16136
rect 4433 16127 4491 16133
rect 5276 16108 5304 16136
rect 6178 16124 6184 16176
rect 6236 16164 6242 16176
rect 7098 16164 7104 16176
rect 6236 16136 7104 16164
rect 6236 16124 6242 16136
rect 7098 16124 7104 16136
rect 7156 16124 7162 16176
rect 10888 16164 10916 16204
rect 11146 16192 11152 16244
rect 11204 16232 11210 16244
rect 11333 16235 11391 16241
rect 11333 16232 11345 16235
rect 11204 16204 11345 16232
rect 11204 16192 11210 16204
rect 11333 16201 11345 16204
rect 11379 16232 11391 16235
rect 12618 16232 12624 16244
rect 11379 16204 12624 16232
rect 11379 16201 11391 16204
rect 11333 16195 11391 16201
rect 12618 16192 12624 16204
rect 12676 16192 12682 16244
rect 12802 16192 12808 16244
rect 12860 16232 12866 16244
rect 14458 16232 14464 16244
rect 12860 16204 14464 16232
rect 12860 16192 12866 16204
rect 14458 16192 14464 16204
rect 14516 16192 14522 16244
rect 14642 16192 14648 16244
rect 14700 16232 14706 16244
rect 14700 16204 15148 16232
rect 14700 16192 14706 16204
rect 11977 16167 12035 16173
rect 10888 16136 11836 16164
rect 5258 16056 5264 16108
rect 5316 16096 5322 16108
rect 6365 16099 6423 16105
rect 5316 16068 5361 16096
rect 5316 16056 5322 16068
rect 6365 16065 6377 16099
rect 6411 16096 6423 16099
rect 6822 16096 6828 16108
rect 6411 16068 6828 16096
rect 6411 16065 6423 16068
rect 6365 16059 6423 16065
rect 6822 16056 6828 16068
rect 6880 16056 6886 16108
rect 7006 16056 7012 16108
rect 7064 16096 7070 16108
rect 7469 16099 7527 16105
rect 7469 16096 7481 16099
rect 7064 16068 7481 16096
rect 7064 16056 7070 16068
rect 7469 16065 7481 16068
rect 7515 16065 7527 16099
rect 7469 16059 7527 16065
rect 3053 16031 3111 16037
rect 3053 15997 3065 16031
rect 3099 16028 3111 16031
rect 3142 16028 3148 16040
rect 3099 16000 3148 16028
rect 3099 15997 3111 16000
rect 3053 15991 3111 15997
rect 3142 15988 3148 16000
rect 3200 15988 3206 16040
rect 5077 16031 5135 16037
rect 5077 16028 5089 16031
rect 3252 16000 5089 16028
rect 3252 15960 3280 16000
rect 5077 15997 5089 16000
rect 5123 15997 5135 16031
rect 5077 15991 5135 15997
rect 6089 16031 6147 16037
rect 6089 15997 6101 16031
rect 6135 16028 6147 16031
rect 6454 16028 6460 16040
rect 6135 16000 6460 16028
rect 6135 15997 6147 16000
rect 6089 15991 6147 15997
rect 6454 15988 6460 16000
rect 6512 15988 6518 16040
rect 6917 16031 6975 16037
rect 6917 15997 6929 16031
rect 6963 16028 6975 16031
rect 7282 16028 7288 16040
rect 6963 16000 7288 16028
rect 6963 15997 6975 16000
rect 6917 15991 6975 15997
rect 7282 15988 7288 16000
rect 7340 15988 7346 16040
rect 7484 16028 7512 16059
rect 7558 16028 7564 16040
rect 7484 16000 7564 16028
rect 7558 15988 7564 16000
rect 7616 15988 7622 16040
rect 7742 16037 7748 16040
rect 7736 16028 7748 16037
rect 7703 16000 7748 16028
rect 7736 15991 7748 16000
rect 7742 15988 7748 15991
rect 7800 15988 7806 16040
rect 9401 16031 9459 16037
rect 9401 15997 9413 16031
rect 9447 16028 9459 16031
rect 9582 16028 9588 16040
rect 9447 16000 9588 16028
rect 9447 15997 9459 16000
rect 9401 15991 9459 15997
rect 9582 15988 9588 16000
rect 9640 15988 9646 16040
rect 9674 15988 9680 16040
rect 9732 16028 9738 16040
rect 11808 16037 11836 16136
rect 11977 16133 11989 16167
rect 12023 16164 12035 16167
rect 15120 16164 15148 16204
rect 15194 16192 15200 16244
rect 15252 16232 15258 16244
rect 15657 16235 15715 16241
rect 15657 16232 15669 16235
rect 15252 16204 15669 16232
rect 15252 16192 15258 16204
rect 15657 16201 15669 16204
rect 15703 16201 15715 16235
rect 15657 16195 15715 16201
rect 17126 16192 17132 16244
rect 17184 16232 17190 16244
rect 18506 16232 18512 16244
rect 17184 16204 18512 16232
rect 17184 16192 17190 16204
rect 18506 16192 18512 16204
rect 18564 16192 18570 16244
rect 19061 16235 19119 16241
rect 19061 16201 19073 16235
rect 19107 16232 19119 16235
rect 19610 16232 19616 16244
rect 19107 16204 19616 16232
rect 19107 16201 19119 16204
rect 19061 16195 19119 16201
rect 19610 16192 19616 16204
rect 19668 16192 19674 16244
rect 17865 16167 17923 16173
rect 12023 16136 15056 16164
rect 15120 16136 15332 16164
rect 12023 16133 12035 16136
rect 11977 16127 12035 16133
rect 12250 16056 12256 16108
rect 12308 16096 12314 16108
rect 12989 16099 13047 16105
rect 12989 16096 13001 16099
rect 12308 16068 13001 16096
rect 12308 16056 12314 16068
rect 12989 16065 13001 16068
rect 13035 16065 13047 16099
rect 12989 16059 13047 16065
rect 13354 16056 13360 16108
rect 13412 16096 13418 16108
rect 13630 16096 13636 16108
rect 13412 16068 13636 16096
rect 13412 16056 13418 16068
rect 13630 16056 13636 16068
rect 13688 16056 13694 16108
rect 14001 16099 14059 16105
rect 14001 16065 14013 16099
rect 14047 16065 14059 16099
rect 15028 16096 15056 16136
rect 15304 16105 15332 16136
rect 17865 16133 17877 16167
rect 17911 16164 17923 16167
rect 20898 16164 20904 16176
rect 17911 16136 20904 16164
rect 17911 16133 17923 16136
rect 17865 16127 17923 16133
rect 20898 16124 20904 16136
rect 20956 16164 20962 16176
rect 21174 16164 21180 16176
rect 20956 16136 21180 16164
rect 20956 16124 20962 16136
rect 21174 16124 21180 16136
rect 21232 16124 21238 16176
rect 15289 16099 15347 16105
rect 15028 16068 15240 16096
rect 14001 16059 14059 16065
rect 9953 16031 10011 16037
rect 9953 16028 9965 16031
rect 9732 16000 9965 16028
rect 9732 15988 9738 16000
rect 9953 15997 9965 16000
rect 9999 15997 10011 16031
rect 9953 15991 10011 15997
rect 11793 16031 11851 16037
rect 11793 15997 11805 16031
rect 11839 15997 11851 16031
rect 11793 15991 11851 15997
rect 12434 15988 12440 16040
rect 12492 16028 12498 16040
rect 13909 16031 13967 16037
rect 13909 16028 13921 16031
rect 12492 16000 13921 16028
rect 12492 15988 12498 16000
rect 13909 15997 13921 16000
rect 13955 15997 13967 16031
rect 13909 15991 13967 15997
rect 2608 15932 3280 15960
rect 3320 15963 3378 15969
rect 3320 15929 3332 15963
rect 3366 15960 3378 15963
rect 3510 15960 3516 15972
rect 3366 15932 3516 15960
rect 3366 15929 3378 15932
rect 3320 15923 3378 15929
rect 3510 15920 3516 15932
rect 3568 15920 3574 15972
rect 5169 15963 5227 15969
rect 5169 15960 5181 15963
rect 3620 15932 5181 15960
rect 2406 15892 2412 15904
rect 2367 15864 2412 15892
rect 2406 15852 2412 15864
rect 2464 15852 2470 15904
rect 2590 15852 2596 15904
rect 2648 15892 2654 15904
rect 3620 15892 3648 15932
rect 5169 15929 5181 15932
rect 5215 15929 5227 15963
rect 5169 15923 5227 15929
rect 5534 15920 5540 15972
rect 5592 15960 5598 15972
rect 6181 15963 6239 15969
rect 6181 15960 6193 15963
rect 5592 15932 6193 15960
rect 5592 15920 5598 15932
rect 6181 15929 6193 15932
rect 6227 15929 6239 15963
rect 7300 15960 7328 15988
rect 14016 15972 14044 16059
rect 14458 15988 14464 16040
rect 14516 16028 14522 16040
rect 15105 16031 15163 16037
rect 15105 16028 15117 16031
rect 14516 16000 15117 16028
rect 14516 15988 14522 16000
rect 15105 15997 15117 16000
rect 15151 15997 15163 16031
rect 15212 16028 15240 16068
rect 15289 16065 15301 16099
rect 15335 16065 15347 16099
rect 15289 16059 15347 16065
rect 15838 16056 15844 16108
rect 15896 16096 15902 16108
rect 16209 16099 16267 16105
rect 16209 16096 16221 16099
rect 15896 16068 16221 16096
rect 15896 16056 15902 16068
rect 16209 16065 16221 16068
rect 16255 16096 16267 16099
rect 17221 16099 17279 16105
rect 17221 16096 17233 16099
rect 16255 16068 17233 16096
rect 16255 16065 16267 16068
rect 16209 16059 16267 16065
rect 17221 16065 17233 16068
rect 17267 16096 17279 16099
rect 17770 16096 17776 16108
rect 17267 16068 17776 16096
rect 17267 16065 17279 16068
rect 17221 16059 17279 16065
rect 17770 16056 17776 16068
rect 17828 16056 17834 16108
rect 18782 16056 18788 16108
rect 18840 16096 18846 16108
rect 19705 16099 19763 16105
rect 19705 16096 19717 16099
rect 18840 16068 19717 16096
rect 18840 16056 18846 16068
rect 19705 16065 19717 16068
rect 19751 16065 19763 16099
rect 20438 16096 20444 16108
rect 20399 16068 20444 16096
rect 19705 16059 19763 16065
rect 15378 16028 15384 16040
rect 15212 16000 15384 16028
rect 15105 15991 15163 15997
rect 15378 15988 15384 16000
rect 15436 15988 15442 16040
rect 16666 15988 16672 16040
rect 16724 16028 16730 16040
rect 18877 16031 18935 16037
rect 18877 16028 18889 16031
rect 16724 16000 18889 16028
rect 16724 15988 16730 16000
rect 18877 15997 18889 16000
rect 18923 16028 18935 16031
rect 19521 16031 19579 16037
rect 19521 16028 19533 16031
rect 18923 16000 19533 16028
rect 18923 15997 18935 16000
rect 18877 15991 18935 15997
rect 19521 15997 19533 16000
rect 19567 15997 19579 16031
rect 19720 16028 19748 16059
rect 20438 16056 20444 16068
rect 20496 16056 20502 16108
rect 20622 16028 20628 16040
rect 19720 16000 20628 16028
rect 19521 15991 19579 15997
rect 20622 15988 20628 16000
rect 20680 15988 20686 16040
rect 10042 15960 10048 15972
rect 7300 15932 10048 15960
rect 6181 15923 6239 15929
rect 10042 15920 10048 15932
rect 10100 15920 10106 15972
rect 10220 15963 10278 15969
rect 10220 15929 10232 15963
rect 10266 15960 10278 15963
rect 10870 15960 10876 15972
rect 10266 15932 10876 15960
rect 10266 15929 10278 15932
rect 10220 15923 10278 15929
rect 10870 15920 10876 15932
rect 10928 15920 10934 15972
rect 13814 15960 13820 15972
rect 13775 15932 13820 15960
rect 13814 15920 13820 15932
rect 13872 15920 13878 15972
rect 13998 15960 14004 15972
rect 13911 15932 14004 15960
rect 2648 15864 3648 15892
rect 2648 15852 2654 15864
rect 3694 15852 3700 15904
rect 3752 15892 3758 15904
rect 6914 15892 6920 15904
rect 3752 15864 6920 15892
rect 3752 15852 3758 15864
rect 6914 15852 6920 15864
rect 6972 15852 6978 15904
rect 7098 15892 7104 15904
rect 7059 15864 7104 15892
rect 7098 15852 7104 15864
rect 7156 15852 7162 15904
rect 9585 15895 9643 15901
rect 9585 15861 9597 15895
rect 9631 15892 9643 15895
rect 12342 15892 12348 15904
rect 9631 15864 12348 15892
rect 9631 15861 9643 15864
rect 9585 15855 9643 15861
rect 12342 15852 12348 15864
rect 12400 15852 12406 15904
rect 12437 15895 12495 15901
rect 12437 15861 12449 15895
rect 12483 15892 12495 15895
rect 12526 15892 12532 15904
rect 12483 15864 12532 15892
rect 12483 15861 12495 15864
rect 12437 15855 12495 15861
rect 12526 15852 12532 15864
rect 12584 15852 12590 15904
rect 12710 15852 12716 15904
rect 12768 15892 12774 15904
rect 12805 15895 12863 15901
rect 12805 15892 12817 15895
rect 12768 15864 12817 15892
rect 12768 15852 12774 15864
rect 12805 15861 12817 15864
rect 12851 15861 12863 15895
rect 12805 15855 12863 15861
rect 12897 15895 12955 15901
rect 12897 15861 12909 15895
rect 12943 15892 12955 15895
rect 13170 15892 13176 15904
rect 12943 15864 13176 15892
rect 12943 15861 12955 15864
rect 12897 15855 12955 15861
rect 13170 15852 13176 15864
rect 13228 15852 13234 15904
rect 13446 15892 13452 15904
rect 13407 15864 13452 15892
rect 13446 15852 13452 15864
rect 13504 15852 13510 15904
rect 13538 15852 13544 15904
rect 13596 15892 13602 15904
rect 13924 15892 13952 15932
rect 13998 15920 14004 15932
rect 14056 15920 14062 15972
rect 16117 15963 16175 15969
rect 16117 15960 16129 15963
rect 14660 15932 16129 15960
rect 14660 15901 14688 15932
rect 16117 15929 16129 15932
rect 16163 15929 16175 15963
rect 16117 15923 16175 15929
rect 17037 15963 17095 15969
rect 17037 15929 17049 15963
rect 17083 15960 17095 15963
rect 20901 15963 20959 15969
rect 20901 15960 20913 15963
rect 17083 15932 20913 15960
rect 17083 15929 17095 15932
rect 17037 15923 17095 15929
rect 20901 15929 20913 15932
rect 20947 15929 20959 15963
rect 20901 15923 20959 15929
rect 13596 15864 13952 15892
rect 14645 15895 14703 15901
rect 13596 15852 13602 15864
rect 14645 15861 14657 15895
rect 14691 15861 14703 15895
rect 14645 15855 14703 15861
rect 15013 15895 15071 15901
rect 15013 15861 15025 15895
rect 15059 15892 15071 15895
rect 15838 15892 15844 15904
rect 15059 15864 15844 15892
rect 15059 15861 15071 15864
rect 15013 15855 15071 15861
rect 15838 15852 15844 15864
rect 15896 15852 15902 15904
rect 16025 15895 16083 15901
rect 16025 15861 16037 15895
rect 16071 15892 16083 15895
rect 16482 15892 16488 15904
rect 16071 15864 16488 15892
rect 16071 15861 16083 15864
rect 16025 15855 16083 15861
rect 16482 15852 16488 15864
rect 16540 15852 16546 15904
rect 16666 15892 16672 15904
rect 16627 15864 16672 15892
rect 16666 15852 16672 15864
rect 16724 15852 16730 15904
rect 17129 15895 17187 15901
rect 17129 15861 17141 15895
rect 17175 15892 17187 15895
rect 17865 15895 17923 15901
rect 17865 15892 17877 15895
rect 17175 15864 17877 15892
rect 17175 15861 17187 15864
rect 17129 15855 17187 15861
rect 17865 15861 17877 15864
rect 17911 15861 17923 15895
rect 17865 15855 17923 15861
rect 19429 15895 19487 15901
rect 19429 15861 19441 15895
rect 19475 15892 19487 15895
rect 19610 15892 19616 15904
rect 19475 15864 19616 15892
rect 19475 15861 19487 15864
rect 19429 15855 19487 15861
rect 19610 15852 19616 15864
rect 19668 15852 19674 15904
rect 19889 15895 19947 15901
rect 19889 15861 19901 15895
rect 19935 15892 19947 15895
rect 19978 15892 19984 15904
rect 19935 15864 19984 15892
rect 19935 15861 19947 15864
rect 19889 15855 19947 15861
rect 19978 15852 19984 15864
rect 20036 15852 20042 15904
rect 20254 15892 20260 15904
rect 20215 15864 20260 15892
rect 20254 15852 20260 15864
rect 20312 15852 20318 15904
rect 20346 15852 20352 15904
rect 20404 15892 20410 15904
rect 20404 15864 20449 15892
rect 20404 15852 20410 15864
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 1486 15648 1492 15700
rect 1544 15688 1550 15700
rect 1581 15691 1639 15697
rect 1581 15688 1593 15691
rect 1544 15660 1593 15688
rect 1544 15648 1550 15660
rect 1581 15657 1593 15660
rect 1627 15657 1639 15691
rect 1581 15651 1639 15657
rect 1949 15691 2007 15697
rect 1949 15657 1961 15691
rect 1995 15688 2007 15691
rect 2590 15688 2596 15700
rect 1995 15660 2596 15688
rect 1995 15657 2007 15660
rect 1949 15651 2007 15657
rect 2590 15648 2596 15660
rect 2648 15648 2654 15700
rect 3326 15688 3332 15700
rect 3287 15660 3332 15688
rect 3326 15648 3332 15660
rect 3384 15648 3390 15700
rect 4065 15691 4123 15697
rect 4065 15657 4077 15691
rect 4111 15688 4123 15691
rect 4154 15688 4160 15700
rect 4111 15660 4160 15688
rect 4111 15657 4123 15660
rect 4065 15651 4123 15657
rect 4154 15648 4160 15660
rect 4212 15648 4218 15700
rect 4433 15691 4491 15697
rect 4433 15657 4445 15691
rect 4479 15688 4491 15691
rect 5074 15688 5080 15700
rect 4479 15660 5080 15688
rect 4479 15657 4491 15660
rect 4433 15651 4491 15657
rect 5074 15648 5080 15660
rect 5132 15648 5138 15700
rect 6822 15648 6828 15700
rect 6880 15688 6886 15700
rect 7009 15691 7067 15697
rect 7009 15688 7021 15691
rect 6880 15660 7021 15688
rect 6880 15648 6886 15660
rect 7009 15657 7021 15660
rect 7055 15657 7067 15691
rect 7009 15651 7067 15657
rect 3694 15620 3700 15632
rect 1504 15592 3700 15620
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15552 1455 15555
rect 1504 15552 1532 15592
rect 3694 15580 3700 15592
rect 3752 15580 3758 15632
rect 3789 15623 3847 15629
rect 3789 15589 3801 15623
rect 3835 15620 3847 15623
rect 4246 15620 4252 15632
rect 3835 15592 4252 15620
rect 3835 15589 3847 15592
rect 3789 15583 3847 15589
rect 4246 15580 4252 15592
rect 4304 15580 4310 15632
rect 4448 15592 5028 15620
rect 1443 15524 1532 15552
rect 1443 15521 1455 15524
rect 1397 15515 1455 15521
rect 1578 15512 1584 15564
rect 1636 15552 1642 15564
rect 2038 15552 2044 15564
rect 1636 15524 2044 15552
rect 1636 15512 1642 15524
rect 2038 15512 2044 15524
rect 2096 15552 2102 15564
rect 2317 15555 2375 15561
rect 2317 15552 2329 15555
rect 2096 15524 2329 15552
rect 2096 15512 2102 15524
rect 2317 15521 2329 15524
rect 2363 15521 2375 15555
rect 2317 15515 2375 15521
rect 3421 15555 3479 15561
rect 3421 15521 3433 15555
rect 3467 15552 3479 15555
rect 4448 15552 4476 15592
rect 3467 15524 4476 15552
rect 4525 15555 4583 15561
rect 3467 15521 3479 15524
rect 3421 15515 3479 15521
rect 4525 15521 4537 15555
rect 4571 15552 4583 15555
rect 4890 15552 4896 15564
rect 4571 15524 4896 15552
rect 4571 15521 4583 15524
rect 4525 15515 4583 15521
rect 4890 15512 4896 15524
rect 4948 15512 4954 15564
rect 2409 15487 2467 15493
rect 2409 15453 2421 15487
rect 2455 15484 2467 15487
rect 2498 15484 2504 15496
rect 2455 15456 2504 15484
rect 2455 15453 2467 15456
rect 2409 15447 2467 15453
rect 2498 15444 2504 15456
rect 2556 15444 2562 15496
rect 2593 15487 2651 15493
rect 2593 15453 2605 15487
rect 2639 15484 2651 15487
rect 2774 15484 2780 15496
rect 2639 15456 2780 15484
rect 2639 15453 2651 15456
rect 2593 15447 2651 15453
rect 2774 15444 2780 15456
rect 2832 15484 2838 15496
rect 3510 15484 3516 15496
rect 2832 15456 3516 15484
rect 2832 15444 2838 15456
rect 3510 15444 3516 15456
rect 3568 15484 3574 15496
rect 4617 15487 4675 15493
rect 4617 15484 4629 15487
rect 3568 15456 4629 15484
rect 3568 15444 3574 15456
rect 4617 15453 4629 15456
rect 4663 15453 4675 15487
rect 5000 15484 5028 15592
rect 5092 15592 6960 15620
rect 5092 15561 5120 15592
rect 5077 15555 5135 15561
rect 5077 15521 5089 15555
rect 5123 15521 5135 15555
rect 5077 15515 5135 15521
rect 5442 15512 5448 15564
rect 5500 15552 5506 15564
rect 5629 15555 5687 15561
rect 5629 15552 5641 15555
rect 5500 15524 5641 15552
rect 5500 15512 5506 15524
rect 5629 15521 5641 15524
rect 5675 15521 5687 15555
rect 5629 15515 5687 15521
rect 5896 15555 5954 15561
rect 5896 15521 5908 15555
rect 5942 15552 5954 15555
rect 6178 15552 6184 15564
rect 5942 15524 6184 15552
rect 5942 15521 5954 15524
rect 5896 15515 5954 15521
rect 6178 15512 6184 15524
rect 6236 15512 6242 15564
rect 5534 15484 5540 15496
rect 5000 15456 5540 15484
rect 4617 15447 4675 15453
rect 5534 15444 5540 15456
rect 5592 15444 5598 15496
rect 3970 15376 3976 15428
rect 4028 15416 4034 15428
rect 5261 15419 5319 15425
rect 5261 15416 5273 15419
rect 4028 15388 5273 15416
rect 4028 15376 4034 15388
rect 5261 15385 5273 15388
rect 5307 15385 5319 15419
rect 5261 15379 5319 15385
rect 2961 15351 3019 15357
rect 2961 15317 2973 15351
rect 3007 15348 3019 15351
rect 3789 15351 3847 15357
rect 3789 15348 3801 15351
rect 3007 15320 3801 15348
rect 3007 15317 3019 15320
rect 2961 15311 3019 15317
rect 3789 15317 3801 15320
rect 3835 15317 3847 15351
rect 3789 15311 3847 15317
rect 4062 15308 4068 15360
rect 4120 15348 4126 15360
rect 6362 15348 6368 15360
rect 4120 15320 6368 15348
rect 4120 15308 4126 15320
rect 6362 15308 6368 15320
rect 6420 15308 6426 15360
rect 6932 15348 6960 15592
rect 7024 15552 7052 15651
rect 7742 15648 7748 15700
rect 7800 15688 7806 15700
rect 8202 15688 8208 15700
rect 7800 15660 8208 15688
rect 7800 15648 7806 15660
rect 8202 15648 8208 15660
rect 8260 15688 8266 15700
rect 8665 15691 8723 15697
rect 8665 15688 8677 15691
rect 8260 15660 8677 15688
rect 8260 15648 8266 15660
rect 8665 15657 8677 15660
rect 8711 15657 8723 15691
rect 8665 15651 8723 15657
rect 9674 15648 9680 15700
rect 9732 15688 9738 15700
rect 10410 15688 10416 15700
rect 9732 15660 10416 15688
rect 9732 15648 9738 15660
rect 10410 15648 10416 15660
rect 10468 15648 10474 15700
rect 11793 15691 11851 15697
rect 11793 15657 11805 15691
rect 11839 15688 11851 15691
rect 11882 15688 11888 15700
rect 11839 15660 11888 15688
rect 11839 15657 11851 15660
rect 11793 15651 11851 15657
rect 11882 15648 11888 15660
rect 11940 15648 11946 15700
rect 11992 15660 12388 15688
rect 7098 15580 7104 15632
rect 7156 15620 7162 15632
rect 11992 15620 12020 15660
rect 12253 15623 12311 15629
rect 12253 15620 12265 15623
rect 7156 15592 12020 15620
rect 12084 15592 12265 15620
rect 7156 15580 7162 15592
rect 7541 15555 7599 15561
rect 7541 15552 7553 15555
rect 7024 15524 7553 15552
rect 7541 15521 7553 15524
rect 7587 15552 7599 15555
rect 9030 15552 9036 15564
rect 7587 15524 8892 15552
rect 8991 15524 9036 15552
rect 7587 15521 7599 15524
rect 7541 15515 7599 15521
rect 7006 15444 7012 15496
rect 7064 15484 7070 15496
rect 7285 15487 7343 15493
rect 7285 15484 7297 15487
rect 7064 15456 7297 15484
rect 7064 15444 7070 15456
rect 7285 15453 7297 15456
rect 7331 15453 7343 15487
rect 8864 15484 8892 15524
rect 9030 15512 9036 15524
rect 9088 15512 9094 15564
rect 9674 15552 9680 15564
rect 9635 15524 9680 15552
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 9944 15555 10002 15561
rect 9944 15521 9956 15555
rect 9990 15552 10002 15555
rect 10502 15552 10508 15564
rect 9990 15524 10508 15552
rect 9990 15521 10002 15524
rect 9944 15515 10002 15521
rect 10502 15512 10508 15524
rect 10560 15512 10566 15564
rect 10962 15512 10968 15564
rect 11020 15552 11026 15564
rect 12084 15552 12112 15592
rect 12253 15589 12265 15592
rect 12299 15589 12311 15623
rect 12360 15620 12388 15660
rect 12526 15648 12532 15700
rect 12584 15688 12590 15700
rect 13265 15691 13323 15697
rect 13265 15688 13277 15691
rect 12584 15660 13277 15688
rect 12584 15648 12590 15660
rect 13265 15657 13277 15660
rect 13311 15657 13323 15691
rect 13265 15651 13323 15657
rect 13630 15648 13636 15700
rect 13688 15688 13694 15700
rect 15838 15688 15844 15700
rect 13688 15660 15844 15688
rect 13688 15648 13694 15660
rect 15838 15648 15844 15660
rect 15896 15648 15902 15700
rect 15933 15691 15991 15697
rect 15933 15657 15945 15691
rect 15979 15688 15991 15691
rect 16666 15688 16672 15700
rect 15979 15660 16672 15688
rect 15979 15657 15991 15660
rect 15933 15651 15991 15657
rect 16666 15648 16672 15660
rect 16724 15648 16730 15700
rect 21358 15688 21364 15700
rect 16776 15660 21364 15688
rect 12802 15620 12808 15632
rect 12360 15592 12808 15620
rect 12253 15583 12311 15589
rect 12802 15580 12808 15592
rect 12860 15580 12866 15632
rect 13078 15580 13084 15632
rect 13136 15620 13142 15632
rect 14185 15623 14243 15629
rect 14185 15620 14197 15623
rect 13136 15592 14197 15620
rect 13136 15580 13142 15592
rect 14185 15589 14197 15592
rect 14231 15589 14243 15623
rect 14185 15583 14243 15589
rect 14277 15623 14335 15629
rect 14277 15589 14289 15623
rect 14323 15620 14335 15623
rect 14366 15620 14372 15632
rect 14323 15592 14372 15620
rect 14323 15589 14335 15592
rect 14277 15583 14335 15589
rect 14366 15580 14372 15592
rect 14424 15580 14430 15632
rect 16025 15623 16083 15629
rect 14476 15592 15148 15620
rect 11020 15524 12112 15552
rect 12161 15555 12219 15561
rect 11020 15512 11026 15524
rect 12161 15521 12173 15555
rect 12207 15521 12219 15555
rect 12161 15515 12219 15521
rect 9214 15484 9220 15496
rect 8864 15456 9220 15484
rect 7285 15447 7343 15453
rect 9214 15444 9220 15456
rect 9272 15444 9278 15496
rect 11146 15444 11152 15496
rect 11204 15484 11210 15496
rect 11333 15487 11391 15493
rect 11333 15484 11345 15487
rect 11204 15456 11345 15484
rect 11204 15444 11210 15456
rect 11333 15453 11345 15456
rect 11379 15453 11391 15487
rect 11333 15447 11391 15453
rect 11882 15444 11888 15496
rect 11940 15484 11946 15496
rect 12176 15484 12204 15515
rect 12434 15512 12440 15564
rect 12492 15552 12498 15564
rect 13173 15555 13231 15561
rect 13173 15552 13185 15555
rect 12492 15524 13185 15552
rect 12492 15512 12498 15524
rect 13173 15521 13185 15524
rect 13219 15552 13231 15555
rect 14476 15552 14504 15592
rect 15010 15552 15016 15564
rect 13219 15524 14504 15552
rect 14971 15524 15016 15552
rect 13219 15521 13231 15524
rect 13173 15515 13231 15521
rect 15010 15512 15016 15524
rect 15068 15512 15074 15564
rect 15120 15552 15148 15592
rect 16025 15589 16037 15623
rect 16071 15620 16083 15623
rect 16574 15620 16580 15632
rect 16071 15592 16580 15620
rect 16071 15589 16083 15592
rect 16025 15583 16083 15589
rect 16574 15580 16580 15592
rect 16632 15580 16638 15632
rect 16776 15552 16804 15660
rect 21358 15648 21364 15660
rect 21416 15648 21422 15700
rect 17402 15580 17408 15632
rect 17460 15620 17466 15632
rect 18693 15623 18751 15629
rect 18693 15620 18705 15623
rect 17460 15592 18705 15620
rect 17460 15580 17466 15592
rect 18693 15589 18705 15592
rect 18739 15589 18751 15623
rect 18693 15583 18751 15589
rect 19245 15623 19303 15629
rect 19245 15589 19257 15623
rect 19291 15620 19303 15623
rect 19702 15620 19708 15632
rect 19291 15592 19708 15620
rect 19291 15589 19303 15592
rect 19245 15583 19303 15589
rect 19702 15580 19708 15592
rect 19760 15580 19766 15632
rect 15120 15524 16804 15552
rect 17120 15555 17178 15561
rect 17120 15521 17132 15555
rect 17166 15552 17178 15555
rect 19150 15552 19156 15564
rect 17166 15524 18828 15552
rect 19111 15524 19156 15552
rect 17166 15521 17178 15524
rect 17120 15515 17178 15521
rect 18800 15496 18828 15524
rect 19150 15512 19156 15524
rect 19208 15512 19214 15564
rect 19426 15512 19432 15564
rect 19484 15552 19490 15564
rect 19981 15555 20039 15561
rect 19981 15552 19993 15555
rect 19484 15524 19993 15552
rect 19484 15512 19490 15524
rect 19981 15521 19993 15524
rect 20027 15521 20039 15555
rect 19981 15515 20039 15521
rect 11940 15456 12204 15484
rect 11940 15444 11946 15456
rect 12250 15444 12256 15496
rect 12308 15484 12314 15496
rect 12345 15487 12403 15493
rect 12345 15484 12357 15487
rect 12308 15456 12357 15484
rect 12308 15444 12314 15456
rect 12345 15453 12357 15456
rect 12391 15453 12403 15487
rect 12345 15447 12403 15453
rect 13357 15487 13415 15493
rect 13357 15453 13369 15487
rect 13403 15484 13415 15487
rect 13538 15484 13544 15496
rect 13403 15456 13544 15484
rect 13403 15453 13415 15456
rect 13357 15447 13415 15453
rect 9490 15416 9496 15428
rect 8220 15388 9496 15416
rect 8220 15348 8248 15388
rect 9490 15376 9496 15388
rect 9548 15376 9554 15428
rect 10870 15376 10876 15428
rect 10928 15416 10934 15428
rect 11057 15419 11115 15425
rect 11057 15416 11069 15419
rect 10928 15388 11069 15416
rect 10928 15376 10934 15388
rect 11057 15385 11069 15388
rect 11103 15416 11115 15419
rect 13372 15416 13400 15447
rect 13538 15444 13544 15456
rect 13596 15444 13602 15496
rect 14461 15487 14519 15493
rect 14461 15453 14473 15487
rect 14507 15453 14519 15487
rect 14461 15447 14519 15453
rect 11103 15388 13400 15416
rect 11103 15385 11115 15388
rect 11057 15379 11115 15385
rect 13998 15376 14004 15428
rect 14056 15416 14062 15428
rect 14476 15416 14504 15447
rect 15562 15444 15568 15496
rect 15620 15484 15626 15496
rect 16117 15487 16175 15493
rect 16117 15484 16129 15487
rect 15620 15456 16129 15484
rect 15620 15444 15626 15456
rect 16117 15453 16129 15456
rect 16163 15453 16175 15487
rect 16117 15447 16175 15453
rect 16853 15487 16911 15493
rect 16853 15453 16865 15487
rect 16899 15453 16911 15487
rect 18782 15484 18788 15496
rect 18695 15456 18788 15484
rect 16853 15447 16911 15453
rect 14056 15388 14504 15416
rect 14056 15376 14062 15388
rect 16206 15376 16212 15428
rect 16264 15416 16270 15428
rect 16868 15416 16896 15447
rect 18782 15444 18788 15456
rect 18840 15484 18846 15496
rect 19337 15487 19395 15493
rect 19337 15484 19349 15487
rect 18840 15456 19349 15484
rect 18840 15444 18846 15456
rect 19337 15453 19349 15456
rect 19383 15453 19395 15487
rect 20070 15484 20076 15496
rect 20031 15456 20076 15484
rect 19337 15447 19395 15453
rect 16264 15388 16896 15416
rect 16264 15376 16270 15388
rect 6932 15320 8248 15348
rect 9217 15351 9275 15357
rect 9217 15317 9229 15351
rect 9263 15348 9275 15351
rect 12434 15348 12440 15360
rect 9263 15320 12440 15348
rect 9263 15317 9275 15320
rect 9217 15311 9275 15317
rect 12434 15308 12440 15320
rect 12492 15308 12498 15360
rect 12802 15348 12808 15360
rect 12763 15320 12808 15348
rect 12802 15308 12808 15320
rect 12860 15308 12866 15360
rect 13814 15348 13820 15360
rect 13775 15320 13820 15348
rect 13814 15308 13820 15320
rect 13872 15308 13878 15360
rect 14274 15308 14280 15360
rect 14332 15348 14338 15360
rect 14829 15351 14887 15357
rect 14829 15348 14841 15351
rect 14332 15320 14841 15348
rect 14332 15308 14338 15320
rect 14829 15317 14841 15320
rect 14875 15317 14887 15351
rect 14829 15311 14887 15317
rect 15565 15351 15623 15357
rect 15565 15317 15577 15351
rect 15611 15348 15623 15351
rect 16758 15348 16764 15360
rect 15611 15320 16764 15348
rect 15611 15317 15623 15320
rect 15565 15311 15623 15317
rect 16758 15308 16764 15320
rect 16816 15308 16822 15360
rect 16868 15348 16896 15388
rect 18693 15419 18751 15425
rect 18693 15385 18705 15419
rect 18739 15416 18751 15419
rect 19352 15416 19380 15447
rect 20070 15444 20076 15456
rect 20128 15444 20134 15496
rect 20165 15487 20223 15493
rect 20165 15453 20177 15487
rect 20211 15453 20223 15487
rect 20165 15447 20223 15453
rect 20180 15416 20208 15447
rect 18739 15388 18920 15416
rect 19352 15388 20208 15416
rect 18739 15385 18751 15388
rect 18693 15379 18751 15385
rect 17034 15348 17040 15360
rect 16868 15320 17040 15348
rect 17034 15308 17040 15320
rect 17092 15308 17098 15360
rect 17954 15308 17960 15360
rect 18012 15348 18018 15360
rect 18233 15351 18291 15357
rect 18233 15348 18245 15351
rect 18012 15320 18245 15348
rect 18012 15308 18018 15320
rect 18233 15317 18245 15320
rect 18279 15317 18291 15351
rect 18233 15311 18291 15317
rect 18506 15308 18512 15360
rect 18564 15348 18570 15360
rect 18785 15351 18843 15357
rect 18785 15348 18797 15351
rect 18564 15320 18797 15348
rect 18564 15308 18570 15320
rect 18785 15317 18797 15320
rect 18831 15317 18843 15351
rect 18892 15348 18920 15388
rect 19334 15348 19340 15360
rect 18892 15320 19340 15348
rect 18785 15311 18843 15317
rect 19334 15308 19340 15320
rect 19392 15308 19398 15360
rect 19610 15348 19616 15360
rect 19571 15320 19616 15348
rect 19610 15308 19616 15320
rect 19668 15308 19674 15360
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 3418 15144 3424 15156
rect 3379 15116 3424 15144
rect 3418 15104 3424 15116
rect 3476 15104 3482 15156
rect 3970 15104 3976 15156
rect 4028 15144 4034 15156
rect 5442 15144 5448 15156
rect 4028 15116 5448 15144
rect 4028 15104 4034 15116
rect 5442 15104 5448 15116
rect 5500 15104 5506 15156
rect 6362 15144 6368 15156
rect 6323 15116 6368 15144
rect 6362 15104 6368 15116
rect 6420 15104 6426 15156
rect 7190 15104 7196 15156
rect 7248 15144 7254 15156
rect 7466 15144 7472 15156
rect 7248 15116 7472 15144
rect 7248 15104 7254 15116
rect 7466 15104 7472 15116
rect 7524 15104 7530 15156
rect 7650 15144 7656 15156
rect 7611 15116 7656 15144
rect 7650 15104 7656 15116
rect 7708 15104 7714 15156
rect 8570 15104 8576 15156
rect 8628 15144 8634 15156
rect 8938 15144 8944 15156
rect 8628 15116 8944 15144
rect 8628 15104 8634 15116
rect 8938 15104 8944 15116
rect 8996 15144 9002 15156
rect 9677 15147 9735 15153
rect 9677 15144 9689 15147
rect 8996 15116 9689 15144
rect 8996 15104 9002 15116
rect 9677 15113 9689 15116
rect 9723 15144 9735 15147
rect 10318 15144 10324 15156
rect 9723 15116 10324 15144
rect 9723 15113 9735 15116
rect 9677 15107 9735 15113
rect 10318 15104 10324 15116
rect 10376 15104 10382 15156
rect 12710 15104 12716 15156
rect 12768 15144 12774 15156
rect 12989 15147 13047 15153
rect 12989 15144 13001 15147
rect 12768 15116 13001 15144
rect 12768 15104 12774 15116
rect 12989 15113 13001 15116
rect 13035 15113 13047 15147
rect 12989 15107 13047 15113
rect 13265 15147 13323 15153
rect 13265 15113 13277 15147
rect 13311 15144 13323 15147
rect 14274 15144 14280 15156
rect 13311 15116 14280 15144
rect 13311 15113 13323 15116
rect 13265 15107 13323 15113
rect 3142 15036 3148 15088
rect 3200 15076 3206 15088
rect 3988 15076 4016 15104
rect 5166 15076 5172 15088
rect 3200 15048 4016 15076
rect 5127 15048 5172 15076
rect 3200 15036 3206 15048
rect 5166 15036 5172 15048
rect 5224 15036 5230 15088
rect 6178 15036 6184 15088
rect 6236 15076 6242 15088
rect 6546 15076 6552 15088
rect 6236 15048 6552 15076
rect 6236 15036 6242 15048
rect 6546 15036 6552 15048
rect 6604 15036 6610 15088
rect 7558 15036 7564 15088
rect 7616 15076 7622 15088
rect 13170 15076 13176 15088
rect 7616 15048 13176 15076
rect 7616 15036 7622 15048
rect 13170 15036 13176 15048
rect 13228 15036 13234 15088
rect 1670 15008 1676 15020
rect 1631 14980 1676 15008
rect 1670 14968 1676 14980
rect 1728 14968 1734 15020
rect 2777 15011 2835 15017
rect 2777 14977 2789 15011
rect 2823 15008 2835 15011
rect 2958 15008 2964 15020
rect 2823 14980 2964 15008
rect 2823 14977 2835 14980
rect 2777 14971 2835 14977
rect 2958 14968 2964 14980
rect 3016 15008 3022 15020
rect 4617 15011 4675 15017
rect 4617 15008 4629 15011
rect 3016 14980 4629 15008
rect 3016 14968 3022 14980
rect 4617 14977 4629 14980
rect 4663 15008 4675 15011
rect 5813 15011 5871 15017
rect 5813 15008 5825 15011
rect 4663 14980 5825 15008
rect 4663 14977 4675 14980
rect 4617 14971 4675 14977
rect 5813 14977 5825 14980
rect 5859 14977 5871 15011
rect 7466 15008 7472 15020
rect 7427 14980 7472 15008
rect 5813 14971 5871 14977
rect 7466 14968 7472 14980
rect 7524 14968 7530 15020
rect 8202 15008 8208 15020
rect 8163 14980 8208 15008
rect 8202 14968 8208 14980
rect 8260 14968 8266 15020
rect 8757 15011 8815 15017
rect 8757 14977 8769 15011
rect 8803 15008 8815 15011
rect 9306 15008 9312 15020
rect 8803 14980 9312 15008
rect 8803 14977 8815 14980
rect 8757 14971 8815 14977
rect 9306 14968 9312 14980
rect 9364 14968 9370 15020
rect 9493 15011 9551 15017
rect 9493 14977 9505 15011
rect 9539 15008 9551 15011
rect 9677 15011 9735 15017
rect 9677 15008 9689 15011
rect 9539 14980 9689 15008
rect 9539 14977 9551 14980
rect 9493 14971 9551 14977
rect 9677 14977 9689 14980
rect 9723 14977 9735 15011
rect 9677 14971 9735 14977
rect 9766 14968 9772 15020
rect 9824 15008 9830 15020
rect 10413 15011 10471 15017
rect 10413 15008 10425 15011
rect 9824 14980 10425 15008
rect 9824 14968 9830 14980
rect 10413 14977 10425 14980
rect 10459 15008 10471 15011
rect 10962 15008 10968 15020
rect 10459 14980 10968 15008
rect 10459 14977 10471 14980
rect 10413 14971 10471 14977
rect 10962 14968 10968 14980
rect 11020 15008 11026 15020
rect 11425 15011 11483 15017
rect 11425 15008 11437 15011
rect 11020 14980 11437 15008
rect 11020 14968 11026 14980
rect 11425 14977 11437 14980
rect 11471 14977 11483 15011
rect 11425 14971 11483 14977
rect 12434 14968 12440 15020
rect 12492 15008 12498 15020
rect 13262 15008 13268 15020
rect 12492 14980 13268 15008
rect 12492 14968 12498 14980
rect 13262 14968 13268 14980
rect 13320 14968 13326 15020
rect 13372 15017 13400 15116
rect 14274 15104 14280 15116
rect 14332 15104 14338 15156
rect 16850 15144 16856 15156
rect 15479 15116 16856 15144
rect 14737 15079 14795 15085
rect 14737 15045 14749 15079
rect 14783 15076 14795 15079
rect 15378 15076 15384 15088
rect 14783 15048 15384 15076
rect 14783 15045 14795 15048
rect 14737 15039 14795 15045
rect 15378 15036 15384 15048
rect 15436 15036 15442 15088
rect 13357 15011 13415 15017
rect 13357 14977 13369 15011
rect 13403 14977 13415 15011
rect 13357 14971 13415 14977
rect 1486 14940 1492 14952
rect 1447 14912 1492 14940
rect 1486 14900 1492 14912
rect 1544 14900 1550 14952
rect 2866 14900 2872 14952
rect 2924 14940 2930 14952
rect 3237 14943 3295 14949
rect 3237 14940 3249 14943
rect 2924 14912 3249 14940
rect 2924 14900 2930 14912
rect 3237 14909 3249 14912
rect 3283 14940 3295 14943
rect 3418 14940 3424 14952
rect 3283 14912 3424 14940
rect 3283 14909 3295 14912
rect 3237 14903 3295 14909
rect 3418 14900 3424 14912
rect 3476 14900 3482 14952
rect 3510 14900 3516 14952
rect 3568 14940 3574 14952
rect 6181 14943 6239 14949
rect 6181 14940 6193 14943
rect 3568 14912 6193 14940
rect 3568 14900 3574 14912
rect 6181 14909 6193 14912
rect 6227 14909 6239 14943
rect 6181 14903 6239 14909
rect 7285 14943 7343 14949
rect 7285 14909 7297 14943
rect 7331 14940 7343 14943
rect 7650 14940 7656 14952
rect 7331 14912 7656 14940
rect 7331 14909 7343 14912
rect 7285 14903 7343 14909
rect 7650 14900 7656 14912
rect 7708 14900 7714 14952
rect 8021 14943 8079 14949
rect 8021 14909 8033 14943
rect 8067 14940 8079 14943
rect 8067 14912 10916 14940
rect 8067 14909 8079 14912
rect 8021 14903 8079 14909
rect 4341 14875 4399 14881
rect 4341 14841 4353 14875
rect 4387 14872 4399 14875
rect 5442 14872 5448 14884
rect 4387 14844 5448 14872
rect 4387 14841 4399 14844
rect 4341 14835 4399 14841
rect 5442 14832 5448 14844
rect 5500 14832 5506 14884
rect 5537 14875 5595 14881
rect 5537 14841 5549 14875
rect 5583 14872 5595 14875
rect 6086 14872 6092 14884
rect 5583 14844 6092 14872
rect 5583 14841 5595 14844
rect 5537 14835 5595 14841
rect 6086 14832 6092 14844
rect 6144 14832 6150 14884
rect 6914 14832 6920 14884
rect 6972 14872 6978 14884
rect 7193 14875 7251 14881
rect 7193 14872 7205 14875
rect 6972 14844 7205 14872
rect 6972 14832 6978 14844
rect 7193 14841 7205 14844
rect 7239 14872 7251 14875
rect 7926 14872 7932 14884
rect 7239 14844 7932 14872
rect 7239 14841 7251 14844
rect 7193 14835 7251 14841
rect 7926 14832 7932 14844
rect 7984 14832 7990 14884
rect 10321 14875 10379 14881
rect 10321 14872 10333 14875
rect 8864 14844 10333 14872
rect 2038 14764 2044 14816
rect 2096 14804 2102 14816
rect 2225 14807 2283 14813
rect 2225 14804 2237 14807
rect 2096 14776 2237 14804
rect 2096 14764 2102 14776
rect 2225 14773 2237 14776
rect 2271 14773 2283 14807
rect 2590 14804 2596 14816
rect 2551 14776 2596 14804
rect 2225 14767 2283 14773
rect 2590 14764 2596 14776
rect 2648 14764 2654 14816
rect 2685 14807 2743 14813
rect 2685 14773 2697 14807
rect 2731 14804 2743 14807
rect 3878 14804 3884 14816
rect 2731 14776 3884 14804
rect 2731 14773 2743 14776
rect 2685 14767 2743 14773
rect 3878 14764 3884 14776
rect 3936 14764 3942 14816
rect 3973 14807 4031 14813
rect 3973 14773 3985 14807
rect 4019 14804 4031 14807
rect 4154 14804 4160 14816
rect 4019 14776 4160 14804
rect 4019 14773 4031 14776
rect 3973 14767 4031 14773
rect 4154 14764 4160 14776
rect 4212 14764 4218 14816
rect 4433 14807 4491 14813
rect 4433 14773 4445 14807
rect 4479 14804 4491 14807
rect 4614 14804 4620 14816
rect 4479 14776 4620 14804
rect 4479 14773 4491 14776
rect 4433 14767 4491 14773
rect 4614 14764 4620 14776
rect 4672 14764 4678 14816
rect 4985 14807 5043 14813
rect 4985 14773 4997 14807
rect 5031 14804 5043 14807
rect 5629 14807 5687 14813
rect 5629 14804 5641 14807
rect 5031 14776 5641 14804
rect 5031 14773 5043 14776
rect 4985 14767 5043 14773
rect 5629 14773 5641 14776
rect 5675 14804 5687 14807
rect 6546 14804 6552 14816
rect 5675 14776 6552 14804
rect 5675 14773 5687 14776
rect 5629 14767 5687 14773
rect 6546 14764 6552 14776
rect 6604 14764 6610 14816
rect 6822 14804 6828 14816
rect 6783 14776 6828 14804
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 8113 14807 8171 14813
rect 8113 14773 8125 14807
rect 8159 14804 8171 14807
rect 8570 14804 8576 14816
rect 8159 14776 8576 14804
rect 8159 14773 8171 14776
rect 8113 14767 8171 14773
rect 8570 14764 8576 14776
rect 8628 14764 8634 14816
rect 8864 14813 8892 14844
rect 10321 14841 10333 14844
rect 10367 14841 10379 14875
rect 10321 14835 10379 14841
rect 8849 14807 8907 14813
rect 8849 14773 8861 14807
rect 8895 14773 8907 14807
rect 9214 14804 9220 14816
rect 9175 14776 9220 14804
rect 8849 14767 8907 14773
rect 9214 14764 9220 14776
rect 9272 14764 9278 14816
rect 9306 14764 9312 14816
rect 9364 14804 9370 14816
rect 9364 14776 9409 14804
rect 9364 14764 9370 14776
rect 9766 14764 9772 14816
rect 9824 14804 9830 14816
rect 9861 14807 9919 14813
rect 9861 14804 9873 14807
rect 9824 14776 9873 14804
rect 9824 14764 9830 14776
rect 9861 14773 9873 14776
rect 9907 14773 9919 14807
rect 10226 14804 10232 14816
rect 10187 14776 10232 14804
rect 9861 14767 9919 14773
rect 10226 14764 10232 14776
rect 10284 14764 10290 14816
rect 10888 14813 10916 14912
rect 11146 14900 11152 14952
rect 11204 14940 11210 14952
rect 11241 14943 11299 14949
rect 11241 14940 11253 14943
rect 11204 14912 11253 14940
rect 11204 14900 11210 14912
rect 11241 14909 11253 14912
rect 11287 14909 11299 14943
rect 12526 14940 12532 14952
rect 11241 14903 11299 14909
rect 11348 14912 12532 14940
rect 10873 14807 10931 14813
rect 10873 14773 10885 14807
rect 10919 14773 10931 14807
rect 10873 14767 10931 14773
rect 11146 14764 11152 14816
rect 11204 14804 11210 14816
rect 11348 14813 11376 14912
rect 12526 14900 12532 14912
rect 12584 14900 12590 14952
rect 12805 14943 12863 14949
rect 12805 14909 12817 14943
rect 12851 14940 12863 14943
rect 12851 14912 13860 14940
rect 12851 14909 12863 14912
rect 12805 14903 12863 14909
rect 11885 14875 11943 14881
rect 11885 14841 11897 14875
rect 11931 14872 11943 14875
rect 13624 14875 13682 14881
rect 11931 14844 13584 14872
rect 11931 14841 11943 14844
rect 11885 14835 11943 14841
rect 11333 14807 11391 14813
rect 11333 14804 11345 14807
rect 11204 14776 11345 14804
rect 11204 14764 11210 14776
rect 11333 14773 11345 14776
rect 11379 14773 11391 14807
rect 11333 14767 11391 14773
rect 11974 14764 11980 14816
rect 12032 14804 12038 14816
rect 12250 14804 12256 14816
rect 12032 14776 12256 14804
rect 12032 14764 12038 14776
rect 12250 14764 12256 14776
rect 12308 14764 12314 14816
rect 12526 14764 12532 14816
rect 12584 14804 12590 14816
rect 13265 14807 13323 14813
rect 13265 14804 13277 14807
rect 12584 14776 13277 14804
rect 12584 14764 12590 14776
rect 13265 14773 13277 14776
rect 13311 14773 13323 14807
rect 13556 14804 13584 14844
rect 13624 14841 13636 14875
rect 13670 14872 13682 14875
rect 13722 14872 13728 14884
rect 13670 14844 13728 14872
rect 13670 14841 13682 14844
rect 13624 14835 13682 14841
rect 13722 14832 13728 14844
rect 13780 14832 13786 14884
rect 13832 14872 13860 14912
rect 13906 14900 13912 14952
rect 13964 14940 13970 14952
rect 15013 14943 15071 14949
rect 15013 14940 15025 14943
rect 13964 14912 15025 14940
rect 13964 14900 13970 14912
rect 15013 14909 15025 14912
rect 15059 14940 15071 14943
rect 15479 14940 15507 15116
rect 16850 15104 16856 15116
rect 16908 15104 16914 15156
rect 17037 15147 17095 15153
rect 17037 15113 17049 15147
rect 17083 15144 17095 15147
rect 19061 15147 19119 15153
rect 17083 15116 18828 15144
rect 17083 15113 17095 15116
rect 17037 15107 17095 15113
rect 16666 15036 16672 15088
rect 16724 15076 16730 15088
rect 17218 15076 17224 15088
rect 16724 15048 17224 15076
rect 16724 15036 16730 15048
rect 17218 15036 17224 15048
rect 17276 15036 17282 15088
rect 18046 15036 18052 15088
rect 18104 15076 18110 15088
rect 18800 15076 18828 15116
rect 19061 15113 19073 15147
rect 19107 15144 19119 15147
rect 19426 15144 19432 15156
rect 19107 15116 19432 15144
rect 19107 15113 19119 15116
rect 19061 15107 19119 15113
rect 19426 15104 19432 15116
rect 19484 15104 19490 15156
rect 20070 15144 20076 15156
rect 20031 15116 20076 15144
rect 20070 15104 20076 15116
rect 20128 15104 20134 15156
rect 19242 15076 19248 15088
rect 18104 15048 18736 15076
rect 18800 15048 19248 15076
rect 18104 15036 18110 15048
rect 16758 14968 16764 15020
rect 16816 15008 16822 15020
rect 17037 15011 17095 15017
rect 17037 15008 17049 15011
rect 16816 14980 17049 15008
rect 16816 14968 16822 14980
rect 17037 14977 17049 14980
rect 17083 14977 17095 15011
rect 17954 15008 17960 15020
rect 17037 14971 17095 14977
rect 17144 14980 17960 15008
rect 15059 14912 15507 14940
rect 15565 14943 15623 14949
rect 15059 14909 15071 14912
rect 15013 14903 15071 14909
rect 15565 14909 15577 14943
rect 15611 14909 15623 14943
rect 15565 14903 15623 14909
rect 15832 14943 15890 14949
rect 15832 14909 15844 14943
rect 15878 14940 15890 14943
rect 17144 14940 17172 14980
rect 17954 14968 17960 14980
rect 18012 14968 18018 15020
rect 18506 15008 18512 15020
rect 18467 14980 18512 15008
rect 18506 14968 18512 14980
rect 18564 14968 18570 15020
rect 18601 15011 18659 15017
rect 18601 14977 18613 15011
rect 18647 14977 18659 15011
rect 18601 14971 18659 14977
rect 15878 14912 17172 14940
rect 17221 14943 17279 14949
rect 15878 14909 15890 14912
rect 15832 14903 15890 14909
rect 17221 14909 17233 14943
rect 17267 14940 17279 14943
rect 17402 14940 17408 14952
rect 17267 14912 17408 14940
rect 17267 14909 17279 14912
rect 17221 14903 17279 14909
rect 15102 14872 15108 14884
rect 13832 14844 15108 14872
rect 15102 14832 15108 14844
rect 15160 14832 15166 14884
rect 15580 14872 15608 14903
rect 17402 14900 17408 14912
rect 17460 14900 17466 14952
rect 17972 14940 18000 14968
rect 18616 14940 18644 14971
rect 17972 14912 18644 14940
rect 18708 14940 18736 15048
rect 19242 15036 19248 15048
rect 19300 15036 19306 15088
rect 19334 14968 19340 15020
rect 19392 15008 19398 15020
rect 19613 15011 19671 15017
rect 19613 15008 19625 15011
rect 19392 14980 19625 15008
rect 19392 14968 19398 14980
rect 19613 14977 19625 14980
rect 19659 15008 19671 15011
rect 20625 15011 20683 15017
rect 20625 15008 20637 15011
rect 19659 14980 20637 15008
rect 19659 14977 19671 14980
rect 19613 14971 19671 14977
rect 20625 14977 20637 14980
rect 20671 14977 20683 15011
rect 20625 14971 20683 14977
rect 20533 14943 20591 14949
rect 20533 14940 20545 14943
rect 18708 14912 20545 14940
rect 20533 14909 20545 14912
rect 20579 14909 20591 14943
rect 20533 14903 20591 14909
rect 16206 14872 16212 14884
rect 15580 14844 16212 14872
rect 16206 14832 16212 14844
rect 16264 14832 16270 14884
rect 16850 14832 16856 14884
rect 16908 14872 16914 14884
rect 17497 14875 17555 14881
rect 17497 14872 17509 14875
rect 16908 14844 17509 14872
rect 16908 14832 16914 14844
rect 17497 14841 17509 14844
rect 17543 14841 17555 14875
rect 17497 14835 17555 14841
rect 18417 14875 18475 14881
rect 18417 14841 18429 14875
rect 18463 14872 18475 14875
rect 19610 14872 19616 14884
rect 18463 14844 19616 14872
rect 18463 14841 18475 14844
rect 18417 14835 18475 14841
rect 19610 14832 19616 14844
rect 19668 14832 19674 14884
rect 14274 14804 14280 14816
rect 13556 14776 14280 14804
rect 13265 14767 13323 14773
rect 14274 14764 14280 14776
rect 14332 14764 14338 14816
rect 15197 14807 15255 14813
rect 15197 14773 15209 14807
rect 15243 14804 15255 14807
rect 15286 14804 15292 14816
rect 15243 14776 15292 14804
rect 15243 14773 15255 14776
rect 15197 14767 15255 14773
rect 15286 14764 15292 14776
rect 15344 14764 15350 14816
rect 15746 14764 15752 14816
rect 15804 14804 15810 14816
rect 16945 14807 17003 14813
rect 16945 14804 16957 14807
rect 15804 14776 16957 14804
rect 15804 14764 15810 14776
rect 16945 14773 16957 14776
rect 16991 14804 17003 14807
rect 17402 14804 17408 14816
rect 16991 14776 17408 14804
rect 16991 14773 17003 14776
rect 16945 14767 17003 14773
rect 17402 14764 17408 14776
rect 17460 14764 17466 14816
rect 18049 14807 18107 14813
rect 18049 14773 18061 14807
rect 18095 14804 18107 14807
rect 19058 14804 19064 14816
rect 18095 14776 19064 14804
rect 18095 14773 18107 14776
rect 18049 14767 18107 14773
rect 19058 14764 19064 14776
rect 19116 14764 19122 14816
rect 19426 14804 19432 14816
rect 19387 14776 19432 14804
rect 19426 14764 19432 14776
rect 19484 14764 19490 14816
rect 19521 14807 19579 14813
rect 19521 14773 19533 14807
rect 19567 14804 19579 14807
rect 19886 14804 19892 14816
rect 19567 14776 19892 14804
rect 19567 14773 19579 14776
rect 19521 14767 19579 14773
rect 19886 14764 19892 14776
rect 19944 14764 19950 14816
rect 20162 14764 20168 14816
rect 20220 14804 20226 14816
rect 20441 14807 20499 14813
rect 20441 14804 20453 14807
rect 20220 14776 20453 14804
rect 20220 14764 20226 14776
rect 20441 14773 20453 14776
rect 20487 14773 20499 14807
rect 20441 14767 20499 14773
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 1486 14560 1492 14612
rect 1544 14600 1550 14612
rect 5350 14600 5356 14612
rect 1544 14572 5356 14600
rect 1544 14560 1550 14572
rect 5350 14560 5356 14572
rect 5408 14560 5414 14612
rect 6089 14603 6147 14609
rect 6089 14569 6101 14603
rect 6135 14600 6147 14603
rect 6822 14600 6828 14612
rect 6135 14572 6828 14600
rect 6135 14569 6147 14572
rect 6089 14563 6147 14569
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 6914 14560 6920 14612
rect 6972 14600 6978 14612
rect 7377 14603 7435 14609
rect 7377 14600 7389 14603
rect 6972 14572 7389 14600
rect 6972 14560 6978 14572
rect 7377 14569 7389 14572
rect 7423 14600 7435 14603
rect 7558 14600 7564 14612
rect 7423 14572 7564 14600
rect 7423 14569 7435 14572
rect 7377 14563 7435 14569
rect 7558 14560 7564 14572
rect 7616 14560 7622 14612
rect 8297 14603 8355 14609
rect 8297 14569 8309 14603
rect 8343 14600 8355 14603
rect 9122 14600 9128 14612
rect 8343 14572 9128 14600
rect 8343 14569 8355 14572
rect 8297 14563 8355 14569
rect 9122 14560 9128 14572
rect 9180 14560 9186 14612
rect 9677 14603 9735 14609
rect 9677 14569 9689 14603
rect 9723 14600 9735 14603
rect 10226 14600 10232 14612
rect 9723 14572 10232 14600
rect 9723 14569 9735 14572
rect 9677 14563 9735 14569
rect 10226 14560 10232 14572
rect 10284 14560 10290 14612
rect 10318 14560 10324 14612
rect 10376 14600 10382 14612
rect 10505 14603 10563 14609
rect 10505 14600 10517 14603
rect 10376 14572 10517 14600
rect 10376 14560 10382 14572
rect 10505 14569 10517 14572
rect 10551 14569 10563 14603
rect 10505 14563 10563 14569
rect 10689 14603 10747 14609
rect 10689 14569 10701 14603
rect 10735 14569 10747 14603
rect 10689 14563 10747 14569
rect 11149 14603 11207 14609
rect 11149 14569 11161 14603
rect 11195 14600 11207 14603
rect 11974 14600 11980 14612
rect 11195 14572 11980 14600
rect 11195 14569 11207 14572
rect 11149 14563 11207 14569
rect 2593 14535 2651 14541
rect 2593 14501 2605 14535
rect 2639 14532 2651 14535
rect 3142 14532 3148 14544
rect 2639 14504 3148 14532
rect 2639 14501 2651 14504
rect 2593 14495 2651 14501
rect 3142 14492 3148 14504
rect 3200 14492 3206 14544
rect 3510 14532 3516 14544
rect 3471 14504 3516 14532
rect 3510 14492 3516 14504
rect 3568 14492 3574 14544
rect 4246 14492 4252 14544
rect 4304 14541 4310 14544
rect 4304 14535 4368 14541
rect 4304 14501 4322 14535
rect 4356 14501 4368 14535
rect 4304 14495 4368 14501
rect 5552 14504 7972 14532
rect 4304 14492 4310 14495
rect 5552 14476 5580 14504
rect 1486 14464 1492 14476
rect 1447 14436 1492 14464
rect 1486 14424 1492 14436
rect 1544 14424 1550 14476
rect 3234 14464 3240 14476
rect 3195 14436 3240 14464
rect 3234 14424 3240 14436
rect 3292 14424 3298 14476
rect 4890 14464 4896 14476
rect 3620 14436 4896 14464
rect 1762 14396 1768 14408
rect 1723 14368 1768 14396
rect 1762 14356 1768 14368
rect 1820 14356 1826 14408
rect 2685 14399 2743 14405
rect 2685 14365 2697 14399
rect 2731 14365 2743 14399
rect 2685 14359 2743 14365
rect 2869 14399 2927 14405
rect 2869 14365 2881 14399
rect 2915 14396 2927 14399
rect 2958 14396 2964 14408
rect 2915 14368 2964 14396
rect 2915 14365 2927 14368
rect 2869 14359 2927 14365
rect 2700 14328 2728 14359
rect 2958 14356 2964 14368
rect 3016 14356 3022 14408
rect 3510 14328 3516 14340
rect 2700 14300 3516 14328
rect 3510 14288 3516 14300
rect 3568 14288 3574 14340
rect 2222 14260 2228 14272
rect 2183 14232 2228 14260
rect 2222 14220 2228 14232
rect 2280 14220 2286 14272
rect 2590 14220 2596 14272
rect 2648 14260 2654 14272
rect 3620 14260 3648 14436
rect 4890 14424 4896 14436
rect 4948 14424 4954 14476
rect 5534 14424 5540 14476
rect 5592 14424 5598 14476
rect 5626 14424 5632 14476
rect 5684 14464 5690 14476
rect 5684 14436 6316 14464
rect 5684 14424 5690 14436
rect 3970 14356 3976 14408
rect 4028 14396 4034 14408
rect 6288 14405 6316 14436
rect 6454 14424 6460 14476
rect 6512 14464 6518 14476
rect 6825 14467 6883 14473
rect 6825 14464 6837 14467
rect 6512 14436 6837 14464
rect 6512 14424 6518 14436
rect 6825 14433 6837 14436
rect 6871 14464 6883 14467
rect 7285 14467 7343 14473
rect 7285 14464 7297 14467
rect 6871 14436 7297 14464
rect 6871 14433 6883 14436
rect 6825 14427 6883 14433
rect 7285 14433 7297 14436
rect 7331 14464 7343 14467
rect 7834 14464 7840 14476
rect 7331 14436 7840 14464
rect 7331 14433 7343 14436
rect 7285 14427 7343 14433
rect 7834 14424 7840 14436
rect 7892 14424 7898 14476
rect 7944 14464 7972 14504
rect 8570 14492 8576 14544
rect 8628 14532 8634 14544
rect 10704 14532 10732 14563
rect 11974 14560 11980 14572
rect 12032 14560 12038 14612
rect 12158 14600 12164 14612
rect 12119 14572 12164 14600
rect 12158 14560 12164 14572
rect 12216 14560 12222 14612
rect 12710 14560 12716 14612
rect 12768 14560 12774 14612
rect 13814 14560 13820 14612
rect 13872 14600 13878 14612
rect 14553 14603 14611 14609
rect 14553 14600 14565 14603
rect 13872 14572 14565 14600
rect 13872 14560 13878 14572
rect 14553 14569 14565 14572
rect 14599 14569 14611 14603
rect 14553 14563 14611 14569
rect 15286 14560 15292 14612
rect 15344 14600 15350 14612
rect 17862 14600 17868 14612
rect 15344 14572 17868 14600
rect 15344 14560 15350 14572
rect 17862 14560 17868 14572
rect 17920 14560 17926 14612
rect 18601 14603 18659 14609
rect 18601 14569 18613 14603
rect 18647 14600 18659 14603
rect 19150 14600 19156 14612
rect 18647 14572 19156 14600
rect 18647 14569 18659 14572
rect 18601 14563 18659 14569
rect 19150 14560 19156 14572
rect 19208 14560 19214 14612
rect 19426 14560 19432 14612
rect 19484 14560 19490 14612
rect 8628 14504 10732 14532
rect 11057 14535 11115 14541
rect 8628 14492 8634 14504
rect 11057 14501 11069 14535
rect 11103 14532 11115 14535
rect 11330 14532 11336 14544
rect 11103 14504 11336 14532
rect 11103 14501 11115 14504
rect 11057 14495 11115 14501
rect 11330 14492 11336 14504
rect 11388 14492 11394 14544
rect 12728 14532 12756 14560
rect 11992 14504 12756 14532
rect 7944 14436 8616 14464
rect 4065 14399 4123 14405
rect 4065 14396 4077 14399
rect 4028 14368 4077 14396
rect 4028 14356 4034 14368
rect 4065 14365 4077 14368
rect 4111 14365 4123 14399
rect 4065 14359 4123 14365
rect 6181 14399 6239 14405
rect 6181 14365 6193 14399
rect 6227 14365 6239 14399
rect 6181 14359 6239 14365
rect 6273 14399 6331 14405
rect 6273 14365 6285 14399
rect 6319 14365 6331 14399
rect 7466 14396 7472 14408
rect 7427 14368 7472 14396
rect 6273 14359 6331 14365
rect 6196 14328 6224 14359
rect 7466 14356 7472 14368
rect 7524 14396 7530 14408
rect 8386 14396 8392 14408
rect 7524 14368 8248 14396
rect 8347 14368 8392 14396
rect 7524 14356 7530 14368
rect 7929 14331 7987 14337
rect 7929 14328 7941 14331
rect 6196 14300 7941 14328
rect 7929 14297 7941 14300
rect 7975 14297 7987 14331
rect 8220 14328 8248 14368
rect 8386 14356 8392 14368
rect 8444 14356 8450 14408
rect 8481 14399 8539 14405
rect 8481 14365 8493 14399
rect 8527 14365 8539 14399
rect 8481 14359 8539 14365
rect 8496 14328 8524 14359
rect 8220 14300 8524 14328
rect 7929 14291 7987 14297
rect 2648 14232 3648 14260
rect 2648 14220 2654 14232
rect 4798 14220 4804 14272
rect 4856 14260 4862 14272
rect 5445 14263 5503 14269
rect 5445 14260 5457 14263
rect 4856 14232 5457 14260
rect 4856 14220 4862 14232
rect 5445 14229 5457 14232
rect 5491 14229 5503 14263
rect 5445 14223 5503 14229
rect 5534 14220 5540 14272
rect 5592 14260 5598 14272
rect 5721 14263 5779 14269
rect 5721 14260 5733 14263
rect 5592 14232 5733 14260
rect 5592 14220 5598 14232
rect 5721 14229 5733 14232
rect 5767 14229 5779 14263
rect 6914 14260 6920 14272
rect 6875 14232 6920 14260
rect 5721 14223 5779 14229
rect 6914 14220 6920 14232
rect 6972 14220 6978 14272
rect 8588 14260 8616 14436
rect 8662 14424 8668 14476
rect 8720 14464 8726 14476
rect 9033 14467 9091 14473
rect 9033 14464 9045 14467
rect 8720 14436 9045 14464
rect 8720 14424 8726 14436
rect 9033 14433 9045 14436
rect 9079 14433 9091 14467
rect 10042 14464 10048 14476
rect 10003 14436 10048 14464
rect 9033 14427 9091 14433
rect 10042 14424 10048 14436
rect 10100 14424 10106 14476
rect 11992 14473 12020 14504
rect 12986 14492 12992 14544
rect 13044 14532 13050 14544
rect 18969 14535 19027 14541
rect 18969 14532 18981 14535
rect 13044 14504 18981 14532
rect 13044 14492 13050 14504
rect 18969 14501 18981 14504
rect 19015 14501 19027 14535
rect 18969 14495 19027 14501
rect 11977 14467 12035 14473
rect 11977 14433 11989 14467
rect 12023 14433 12035 14467
rect 12526 14464 12532 14476
rect 12487 14436 12532 14464
rect 11977 14427 12035 14433
rect 12526 14424 12532 14436
rect 12584 14424 12590 14476
rect 12796 14467 12854 14473
rect 12796 14433 12808 14467
rect 12842 14464 12854 14467
rect 14918 14464 14924 14476
rect 12842 14436 14924 14464
rect 12842 14433 12854 14436
rect 12796 14427 12854 14433
rect 14918 14424 14924 14436
rect 14976 14424 14982 14476
rect 15378 14424 15384 14476
rect 15436 14464 15442 14476
rect 15556 14467 15614 14473
rect 15556 14464 15568 14467
rect 15436 14436 15568 14464
rect 15436 14424 15442 14436
rect 15556 14433 15568 14436
rect 15602 14464 15614 14467
rect 16942 14464 16948 14476
rect 15602 14436 16948 14464
rect 15602 14433 15614 14436
rect 15556 14427 15614 14433
rect 16942 14424 16948 14436
rect 17000 14424 17006 14476
rect 17396 14467 17454 14473
rect 17396 14433 17408 14467
rect 17442 14464 17454 14467
rect 19444 14464 19472 14560
rect 20901 14535 20959 14541
rect 20901 14532 20913 14535
rect 19996 14504 20913 14532
rect 19996 14464 20024 14504
rect 20901 14501 20913 14504
rect 20947 14501 20959 14535
rect 20901 14495 20959 14501
rect 20162 14464 20168 14476
rect 17442 14436 19196 14464
rect 19444 14436 20024 14464
rect 20123 14436 20168 14464
rect 17442 14433 17454 14436
rect 17396 14427 17454 14433
rect 10137 14399 10195 14405
rect 10137 14365 10149 14399
rect 10183 14396 10195 14399
rect 10226 14396 10232 14408
rect 10183 14368 10232 14396
rect 10183 14365 10195 14368
rect 10137 14359 10195 14365
rect 10226 14356 10232 14368
rect 10284 14356 10290 14408
rect 10321 14399 10379 14405
rect 10321 14365 10333 14399
rect 10367 14396 10379 14399
rect 10505 14399 10563 14405
rect 10505 14396 10517 14399
rect 10367 14368 10517 14396
rect 10367 14365 10379 14368
rect 10321 14359 10379 14365
rect 10505 14365 10517 14368
rect 10551 14365 10563 14399
rect 10505 14359 10563 14365
rect 10962 14356 10968 14408
rect 11020 14396 11026 14408
rect 11241 14399 11299 14405
rect 11241 14396 11253 14399
rect 11020 14368 11253 14396
rect 11020 14356 11026 14368
rect 11241 14365 11253 14368
rect 11287 14365 11299 14399
rect 11241 14359 11299 14365
rect 13998 14356 14004 14408
rect 14056 14396 14062 14408
rect 14645 14399 14703 14405
rect 14645 14396 14657 14399
rect 14056 14368 14657 14396
rect 14056 14356 14062 14368
rect 14645 14365 14657 14368
rect 14691 14365 14703 14399
rect 14645 14359 14703 14365
rect 14737 14399 14795 14405
rect 14737 14365 14749 14399
rect 14783 14365 14795 14399
rect 15286 14396 15292 14408
rect 15247 14368 15292 14396
rect 14737 14359 14795 14365
rect 9217 14331 9275 14337
rect 9217 14297 9229 14331
rect 9263 14328 9275 14331
rect 11698 14328 11704 14340
rect 9263 14300 11704 14328
rect 9263 14297 9275 14300
rect 9217 14291 9275 14297
rect 11698 14288 11704 14300
rect 11756 14288 11762 14340
rect 14752 14328 14780 14359
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 17034 14356 17040 14408
rect 17092 14396 17098 14408
rect 17129 14399 17187 14405
rect 17129 14396 17141 14399
rect 17092 14368 17141 14396
rect 17092 14356 17098 14368
rect 17129 14365 17141 14368
rect 17175 14365 17187 14399
rect 19058 14396 19064 14408
rect 19019 14368 19064 14396
rect 17129 14359 17187 14365
rect 13648 14300 14780 14328
rect 11606 14260 11612 14272
rect 8588 14232 11612 14260
rect 11606 14220 11612 14232
rect 11664 14220 11670 14272
rect 12710 14220 12716 14272
rect 12768 14260 12774 14272
rect 13648 14260 13676 14300
rect 12768 14232 13676 14260
rect 12768 14220 12774 14232
rect 13722 14220 13728 14272
rect 13780 14260 13786 14272
rect 13909 14263 13967 14269
rect 13909 14260 13921 14263
rect 13780 14232 13921 14260
rect 13780 14220 13786 14232
rect 13909 14229 13921 14232
rect 13955 14229 13967 14263
rect 13909 14223 13967 14229
rect 14185 14263 14243 14269
rect 14185 14229 14197 14263
rect 14231 14260 14243 14263
rect 15654 14260 15660 14272
rect 14231 14232 15660 14260
rect 14231 14229 14243 14232
rect 14185 14223 14243 14229
rect 15654 14220 15660 14232
rect 15712 14220 15718 14272
rect 16669 14263 16727 14269
rect 16669 14229 16681 14263
rect 16715 14260 16727 14263
rect 17034 14260 17040 14272
rect 16715 14232 17040 14260
rect 16715 14229 16727 14232
rect 16669 14223 16727 14229
rect 17034 14220 17040 14232
rect 17092 14220 17098 14272
rect 17144 14260 17172 14359
rect 19058 14356 19064 14368
rect 19116 14356 19122 14408
rect 19168 14405 19196 14436
rect 20162 14424 20168 14436
rect 20220 14424 20226 14476
rect 19153 14399 19211 14405
rect 19153 14365 19165 14399
rect 19199 14396 19211 14399
rect 19426 14396 19432 14408
rect 19199 14368 19432 14396
rect 19199 14365 19211 14368
rect 19153 14359 19211 14365
rect 19426 14356 19432 14368
rect 19484 14356 19490 14408
rect 20257 14399 20315 14405
rect 20257 14365 20269 14399
rect 20303 14365 20315 14399
rect 20257 14359 20315 14365
rect 18509 14331 18567 14337
rect 18509 14297 18521 14331
rect 18555 14328 18567 14331
rect 18782 14328 18788 14340
rect 18555 14300 18788 14328
rect 18555 14297 18567 14300
rect 18509 14291 18567 14297
rect 18782 14288 18788 14300
rect 18840 14288 18846 14340
rect 19610 14328 19616 14340
rect 19571 14300 19616 14328
rect 19610 14288 19616 14300
rect 19668 14328 19674 14340
rect 20272 14328 20300 14359
rect 20346 14356 20352 14408
rect 20404 14396 20410 14408
rect 20404 14368 20449 14396
rect 20404 14356 20410 14368
rect 19668 14300 20300 14328
rect 19668 14288 19674 14300
rect 17862 14260 17868 14272
rect 17144 14232 17868 14260
rect 17862 14220 17868 14232
rect 17920 14220 17926 14272
rect 19242 14220 19248 14272
rect 19300 14260 19306 14272
rect 19797 14263 19855 14269
rect 19797 14260 19809 14263
rect 19300 14232 19809 14260
rect 19300 14220 19306 14232
rect 19797 14229 19809 14232
rect 19843 14229 19855 14263
rect 19797 14223 19855 14229
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 2866 14056 2872 14068
rect 2608 14028 2872 14056
rect 2501 13923 2559 13929
rect 2501 13889 2513 13923
rect 2547 13920 2559 13923
rect 2608 13920 2636 14028
rect 2866 14016 2872 14028
rect 2924 14056 2930 14068
rect 3786 14056 3792 14068
rect 2924 14028 3792 14056
rect 2924 14016 2930 14028
rect 3786 14016 3792 14028
rect 3844 14016 3850 14068
rect 4062 14016 4068 14068
rect 4120 14056 4126 14068
rect 6365 14059 6423 14065
rect 6365 14056 6377 14059
rect 4120 14028 6377 14056
rect 4120 14016 4126 14028
rect 6365 14025 6377 14028
rect 6411 14025 6423 14059
rect 9214 14056 9220 14068
rect 6365 14019 6423 14025
rect 6472 14028 9220 14056
rect 2547 13892 2636 13920
rect 2547 13889 2559 13892
rect 2501 13883 2559 13889
rect 4062 13880 4068 13932
rect 4120 13920 4126 13932
rect 4120 13892 4660 13920
rect 4120 13880 4126 13892
rect 2317 13855 2375 13861
rect 2317 13821 2329 13855
rect 2363 13852 2375 13855
rect 2406 13852 2412 13864
rect 2363 13824 2412 13852
rect 2363 13821 2375 13824
rect 2317 13815 2375 13821
rect 2406 13812 2412 13824
rect 2464 13812 2470 13864
rect 2869 13855 2927 13861
rect 2869 13821 2881 13855
rect 2915 13852 2927 13855
rect 3970 13852 3976 13864
rect 2915 13824 3976 13852
rect 2915 13821 2927 13824
rect 2869 13815 2927 13821
rect 2130 13744 2136 13796
rect 2188 13784 2194 13796
rect 2884 13784 2912 13815
rect 3970 13812 3976 13824
rect 4028 13852 4034 13864
rect 4522 13852 4528 13864
rect 4028 13824 4528 13852
rect 4028 13812 4034 13824
rect 4522 13812 4528 13824
rect 4580 13812 4586 13864
rect 2188 13756 2912 13784
rect 3136 13787 3194 13793
rect 2188 13744 2194 13756
rect 3136 13753 3148 13787
rect 3182 13784 3194 13787
rect 3602 13784 3608 13796
rect 3182 13756 3608 13784
rect 3182 13753 3194 13756
rect 3136 13747 3194 13753
rect 3602 13744 3608 13756
rect 3660 13744 3666 13796
rect 4632 13784 4660 13892
rect 4798 13861 4804 13864
rect 4792 13852 4804 13861
rect 4759 13824 4804 13852
rect 4792 13815 4804 13824
rect 4798 13812 4804 13815
rect 4856 13812 4862 13864
rect 6086 13852 6092 13864
rect 4908 13824 6092 13852
rect 4908 13784 4936 13824
rect 6086 13812 6092 13824
rect 6144 13812 6150 13864
rect 6181 13855 6239 13861
rect 6181 13821 6193 13855
rect 6227 13852 6239 13855
rect 6270 13852 6276 13864
rect 6227 13824 6276 13852
rect 6227 13821 6239 13824
rect 6181 13815 6239 13821
rect 6270 13812 6276 13824
rect 6328 13852 6334 13864
rect 6472 13852 6500 14028
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 10045 14059 10103 14065
rect 10045 14025 10057 14059
rect 10091 14056 10103 14059
rect 12437 14059 12495 14065
rect 10091 14028 11376 14056
rect 10091 14025 10103 14028
rect 10045 14019 10103 14025
rect 9493 13991 9551 13997
rect 9493 13957 9505 13991
rect 9539 13988 9551 13991
rect 9858 13988 9864 14000
rect 9539 13960 9864 13988
rect 9539 13957 9551 13960
rect 9493 13951 9551 13957
rect 9858 13948 9864 13960
rect 9916 13948 9922 14000
rect 11348 13988 11376 14028
rect 12437 14025 12449 14059
rect 12483 14056 12495 14059
rect 14182 14056 14188 14068
rect 12483 14028 14188 14056
rect 12483 14025 12495 14028
rect 12437 14019 12495 14025
rect 14182 14016 14188 14028
rect 14240 14016 14246 14068
rect 14921 14059 14979 14065
rect 14921 14025 14933 14059
rect 14967 14056 14979 14059
rect 17954 14056 17960 14068
rect 14967 14028 17960 14056
rect 14967 14025 14979 14028
rect 14921 14019 14979 14025
rect 17954 14016 17960 14028
rect 18012 14016 18018 14068
rect 19426 14056 19432 14068
rect 19387 14028 19432 14056
rect 19426 14016 19432 14028
rect 19484 14016 19490 14068
rect 19702 14056 19708 14068
rect 19663 14028 19708 14056
rect 19702 14016 19708 14028
rect 19760 14016 19766 14068
rect 11348 13960 12480 13988
rect 8202 13880 8208 13932
rect 8260 13920 8266 13932
rect 9033 13923 9091 13929
rect 9033 13920 9045 13923
rect 8260 13892 9045 13920
rect 8260 13880 8266 13892
rect 9033 13889 9045 13892
rect 9079 13889 9091 13923
rect 9876 13920 9904 13948
rect 12452 13932 12480 13960
rect 13538 13948 13544 14000
rect 13596 13988 13602 14000
rect 13596 13960 14136 13988
rect 13596 13948 13602 13960
rect 9876 13892 10180 13920
rect 9033 13883 9091 13889
rect 6822 13852 6828 13864
rect 6328 13824 6500 13852
rect 6783 13824 6828 13852
rect 6328 13812 6334 13824
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 7081 13855 7139 13861
rect 7081 13852 7093 13855
rect 6932 13824 7093 13852
rect 6932 13784 6960 13824
rect 7081 13821 7093 13824
rect 7127 13821 7139 13855
rect 7081 13815 7139 13821
rect 8386 13812 8392 13864
rect 8444 13852 8450 13864
rect 9677 13855 9735 13861
rect 9677 13852 9689 13855
rect 8444 13824 9689 13852
rect 8444 13812 8450 13824
rect 9677 13821 9689 13824
rect 9723 13821 9735 13855
rect 9677 13815 9735 13821
rect 9766 13812 9772 13864
rect 9824 13852 9830 13864
rect 9861 13855 9919 13861
rect 9861 13852 9873 13855
rect 9824 13824 9873 13852
rect 9824 13812 9830 13824
rect 9861 13821 9873 13824
rect 9907 13821 9919 13855
rect 10152 13852 10180 13892
rect 12434 13880 12440 13932
rect 12492 13880 12498 13932
rect 12618 13880 12624 13932
rect 12676 13920 12682 13932
rect 12989 13923 13047 13929
rect 12989 13920 13001 13923
rect 12676 13892 13001 13920
rect 12676 13880 12682 13892
rect 12989 13889 13001 13892
rect 13035 13889 13047 13923
rect 12989 13883 13047 13889
rect 13262 13880 13268 13932
rect 13320 13920 13326 13932
rect 14001 13923 14059 13929
rect 14001 13920 14013 13923
rect 13320 13892 14013 13920
rect 13320 13880 13326 13892
rect 14001 13889 14013 13892
rect 14047 13889 14059 13923
rect 14001 13883 14059 13889
rect 10410 13852 10416 13864
rect 10152 13824 10416 13852
rect 9861 13815 9919 13821
rect 10410 13812 10416 13824
rect 10468 13812 10474 13864
rect 10680 13855 10738 13861
rect 10680 13821 10692 13855
rect 10726 13852 10738 13855
rect 11146 13852 11152 13864
rect 10726 13824 11152 13852
rect 10726 13821 10738 13824
rect 10680 13815 10738 13821
rect 11146 13812 11152 13824
rect 11204 13812 11210 13864
rect 12802 13852 12808 13864
rect 12763 13824 12808 13852
rect 12802 13812 12808 13824
rect 12860 13812 12866 13864
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13852 12955 13855
rect 13446 13852 13452 13864
rect 12943 13824 13452 13852
rect 12943 13821 12955 13824
rect 12897 13815 12955 13821
rect 13446 13812 13452 13824
rect 13504 13812 13510 13864
rect 13630 13812 13636 13864
rect 13688 13852 13694 13864
rect 13909 13855 13967 13861
rect 13909 13852 13921 13855
rect 13688 13824 13921 13852
rect 13688 13812 13694 13824
rect 13909 13821 13921 13824
rect 13955 13821 13967 13855
rect 14108 13852 14136 13960
rect 16574 13948 16580 14000
rect 16632 13988 16638 14000
rect 16945 13991 17003 13997
rect 16945 13988 16957 13991
rect 16632 13960 16957 13988
rect 16632 13948 16638 13960
rect 16945 13957 16957 13960
rect 16991 13957 17003 13991
rect 16945 13951 17003 13957
rect 14182 13880 14188 13932
rect 14240 13920 14246 13932
rect 14240 13892 15424 13920
rect 14240 13880 14246 13892
rect 14737 13855 14795 13861
rect 14737 13852 14749 13855
rect 14108 13824 14749 13852
rect 13909 13815 13967 13821
rect 14737 13821 14749 13824
rect 14783 13821 14795 13855
rect 15286 13852 15292 13864
rect 15247 13824 15292 13852
rect 14737 13815 14795 13821
rect 15286 13812 15292 13824
rect 15344 13812 15350 13864
rect 15396 13852 15424 13892
rect 17402 13880 17408 13932
rect 17460 13920 17466 13932
rect 17497 13923 17555 13929
rect 17497 13920 17509 13923
rect 17460 13892 17509 13920
rect 17460 13880 17466 13892
rect 17497 13889 17509 13892
rect 17543 13889 17555 13923
rect 19444 13920 19472 14016
rect 20257 13923 20315 13929
rect 20257 13920 20269 13923
rect 19444 13892 20269 13920
rect 17497 13883 17555 13889
rect 20257 13889 20269 13892
rect 20303 13889 20315 13923
rect 20257 13883 20315 13889
rect 17313 13855 17371 13861
rect 17313 13852 17325 13855
rect 15396 13824 17325 13852
rect 17313 13821 17325 13824
rect 17359 13821 17371 13855
rect 17313 13815 17371 13821
rect 17862 13812 17868 13864
rect 17920 13852 17926 13864
rect 18049 13855 18107 13861
rect 18049 13852 18061 13855
rect 17920 13824 18061 13852
rect 17920 13812 17926 13824
rect 18049 13821 18061 13824
rect 18095 13821 18107 13855
rect 20165 13855 20223 13861
rect 20165 13852 20177 13855
rect 18049 13815 18107 13821
rect 18156 13824 20177 13852
rect 4632 13756 4936 13784
rect 5920 13756 6960 13784
rect 1854 13716 1860 13728
rect 1815 13688 1860 13716
rect 1854 13676 1860 13688
rect 1912 13676 1918 13728
rect 2225 13719 2283 13725
rect 2225 13685 2237 13719
rect 2271 13716 2283 13719
rect 2498 13716 2504 13728
rect 2271 13688 2504 13716
rect 2271 13685 2283 13688
rect 2225 13679 2283 13685
rect 2498 13676 2504 13688
rect 2556 13676 2562 13728
rect 3694 13676 3700 13728
rect 3752 13716 3758 13728
rect 4246 13716 4252 13728
rect 3752 13688 4252 13716
rect 3752 13676 3758 13688
rect 4246 13676 4252 13688
rect 4304 13716 4310 13728
rect 5626 13716 5632 13728
rect 4304 13688 5632 13716
rect 4304 13676 4310 13688
rect 5626 13676 5632 13688
rect 5684 13676 5690 13728
rect 5810 13676 5816 13728
rect 5868 13716 5874 13728
rect 5920 13725 5948 13756
rect 7374 13744 7380 13796
rect 7432 13784 7438 13796
rect 8849 13787 8907 13793
rect 8849 13784 8861 13787
rect 7432 13756 8861 13784
rect 7432 13744 7438 13756
rect 8849 13753 8861 13756
rect 8895 13784 8907 13787
rect 13078 13784 13084 13796
rect 8895 13756 13084 13784
rect 8895 13753 8907 13756
rect 8849 13747 8907 13753
rect 13078 13744 13084 13756
rect 13136 13744 13142 13796
rect 15556 13787 15614 13793
rect 13464 13756 15516 13784
rect 5905 13719 5963 13725
rect 5905 13716 5917 13719
rect 5868 13688 5917 13716
rect 5868 13676 5874 13688
rect 5905 13685 5917 13688
rect 5951 13685 5963 13719
rect 8202 13716 8208 13728
rect 8163 13688 8208 13716
rect 5905 13679 5963 13685
rect 8202 13676 8208 13688
rect 8260 13676 8266 13728
rect 8294 13676 8300 13728
rect 8352 13716 8358 13728
rect 8481 13719 8539 13725
rect 8481 13716 8493 13719
rect 8352 13688 8493 13716
rect 8352 13676 8358 13688
rect 8481 13685 8493 13688
rect 8527 13685 8539 13719
rect 8481 13679 8539 13685
rect 8570 13676 8576 13728
rect 8628 13716 8634 13728
rect 8941 13719 8999 13725
rect 8941 13716 8953 13719
rect 8628 13688 8953 13716
rect 8628 13676 8634 13688
rect 8941 13685 8953 13688
rect 8987 13685 8999 13719
rect 8941 13679 8999 13685
rect 9122 13676 9128 13728
rect 9180 13716 9186 13728
rect 9490 13716 9496 13728
rect 9180 13688 9496 13716
rect 9180 13676 9186 13688
rect 9490 13676 9496 13688
rect 9548 13676 9554 13728
rect 11793 13719 11851 13725
rect 11793 13685 11805 13719
rect 11839 13716 11851 13719
rect 12342 13716 12348 13728
rect 11839 13688 12348 13716
rect 11839 13685 11851 13688
rect 11793 13679 11851 13685
rect 12342 13676 12348 13688
rect 12400 13676 12406 13728
rect 12434 13676 12440 13728
rect 12492 13716 12498 13728
rect 13354 13716 13360 13728
rect 12492 13688 13360 13716
rect 12492 13676 12498 13688
rect 13354 13676 13360 13688
rect 13412 13676 13418 13728
rect 13464 13725 13492 13756
rect 13449 13719 13507 13725
rect 13449 13685 13461 13719
rect 13495 13685 13507 13719
rect 13814 13716 13820 13728
rect 13775 13688 13820 13716
rect 13449 13679 13507 13685
rect 13814 13676 13820 13688
rect 13872 13676 13878 13728
rect 15488 13716 15516 13756
rect 15556 13753 15568 13787
rect 15602 13784 15614 13787
rect 15746 13784 15752 13796
rect 15602 13756 15752 13784
rect 15602 13753 15614 13756
rect 15556 13747 15614 13753
rect 15746 13744 15752 13756
rect 15804 13744 15810 13796
rect 16758 13784 16764 13796
rect 16316 13756 16764 13784
rect 16316 13716 16344 13756
rect 16758 13744 16764 13756
rect 16816 13744 16822 13796
rect 16942 13744 16948 13796
rect 17000 13784 17006 13796
rect 17405 13787 17463 13793
rect 17405 13784 17417 13787
rect 17000 13756 17417 13784
rect 17000 13744 17006 13756
rect 17405 13753 17417 13756
rect 17451 13753 17463 13787
rect 17405 13747 17463 13753
rect 17954 13744 17960 13796
rect 18012 13784 18018 13796
rect 18156 13784 18184 13824
rect 20165 13821 20177 13824
rect 20211 13821 20223 13855
rect 20165 13815 20223 13821
rect 20717 13855 20775 13861
rect 20717 13821 20729 13855
rect 20763 13852 20775 13855
rect 21082 13852 21088 13864
rect 20763 13824 21088 13852
rect 20763 13821 20775 13824
rect 20717 13815 20775 13821
rect 21082 13812 21088 13824
rect 21140 13812 21146 13864
rect 18322 13793 18328 13796
rect 18316 13784 18328 13793
rect 18012 13756 18184 13784
rect 18283 13756 18328 13784
rect 18012 13744 18018 13756
rect 18316 13747 18328 13756
rect 18322 13744 18328 13747
rect 18380 13744 18386 13796
rect 19426 13784 19432 13796
rect 18892 13756 19432 13784
rect 16666 13716 16672 13728
rect 15488 13688 16344 13716
rect 16627 13688 16672 13716
rect 16666 13676 16672 13688
rect 16724 13676 16730 13728
rect 17218 13676 17224 13728
rect 17276 13716 17282 13728
rect 18892 13716 18920 13756
rect 19426 13744 19432 13756
rect 19484 13744 19490 13796
rect 19610 13744 19616 13796
rect 19668 13784 19674 13796
rect 20073 13787 20131 13793
rect 20073 13784 20085 13787
rect 19668 13756 20085 13784
rect 19668 13744 19674 13756
rect 20073 13753 20085 13756
rect 20119 13753 20131 13787
rect 20073 13747 20131 13753
rect 17276 13688 18920 13716
rect 17276 13676 17282 13688
rect 18966 13676 18972 13728
rect 19024 13716 19030 13728
rect 19886 13716 19892 13728
rect 19024 13688 19892 13716
rect 19024 13676 19030 13688
rect 19886 13676 19892 13688
rect 19944 13676 19950 13728
rect 20898 13716 20904 13728
rect 20859 13688 20904 13716
rect 20898 13676 20904 13688
rect 20956 13676 20962 13728
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 3234 13472 3240 13524
rect 3292 13512 3298 13524
rect 4065 13515 4123 13521
rect 4065 13512 4077 13515
rect 3292 13484 4077 13512
rect 3292 13472 3298 13484
rect 4065 13481 4077 13484
rect 4111 13481 4123 13515
rect 4065 13475 4123 13481
rect 4525 13515 4583 13521
rect 4525 13481 4537 13515
rect 4571 13512 4583 13515
rect 5077 13515 5135 13521
rect 5077 13512 5089 13515
rect 4571 13484 5089 13512
rect 4571 13481 4583 13484
rect 4525 13475 4583 13481
rect 5077 13481 5089 13484
rect 5123 13481 5135 13515
rect 5534 13512 5540 13524
rect 5495 13484 5540 13512
rect 5077 13475 5135 13481
rect 5534 13472 5540 13484
rect 5592 13472 5598 13524
rect 6089 13515 6147 13521
rect 6089 13481 6101 13515
rect 6135 13481 6147 13515
rect 6089 13475 6147 13481
rect 6549 13515 6607 13521
rect 6549 13481 6561 13515
rect 6595 13512 6607 13515
rect 6914 13512 6920 13524
rect 6595 13484 6920 13512
rect 6595 13481 6607 13484
rect 6549 13475 6607 13481
rect 1765 13447 1823 13453
rect 1765 13413 1777 13447
rect 1811 13444 1823 13447
rect 5166 13444 5172 13456
rect 1811 13416 5172 13444
rect 1811 13413 1823 13416
rect 1765 13407 1823 13413
rect 5166 13404 5172 13416
rect 5224 13404 5230 13456
rect 5445 13447 5503 13453
rect 5445 13413 5457 13447
rect 5491 13444 5503 13447
rect 6104 13444 6132 13475
rect 6914 13472 6920 13484
rect 6972 13472 6978 13524
rect 7190 13472 7196 13524
rect 7248 13512 7254 13524
rect 7742 13512 7748 13524
rect 7248 13484 7748 13512
rect 7248 13472 7254 13484
rect 7742 13472 7748 13484
rect 7800 13472 7806 13524
rect 8294 13512 8300 13524
rect 8255 13484 8300 13512
rect 8294 13472 8300 13484
rect 8352 13472 8358 13524
rect 9217 13515 9275 13521
rect 9217 13481 9229 13515
rect 9263 13512 9275 13515
rect 12434 13512 12440 13524
rect 9263 13484 12440 13512
rect 9263 13481 9275 13484
rect 9217 13475 9275 13481
rect 12434 13472 12440 13484
rect 12492 13472 12498 13524
rect 13078 13472 13084 13524
rect 13136 13512 13142 13524
rect 16945 13515 17003 13521
rect 13136 13484 16804 13512
rect 13136 13472 13142 13484
rect 5491 13416 6132 13444
rect 6457 13447 6515 13453
rect 5491 13413 5503 13416
rect 5445 13407 5503 13413
rect 6457 13413 6469 13447
rect 6503 13444 6515 13447
rect 7208 13444 7236 13472
rect 8386 13444 8392 13456
rect 6503 13416 7236 13444
rect 7300 13416 8392 13444
rect 6503 13413 6515 13416
rect 6457 13407 6515 13413
rect 1489 13379 1547 13385
rect 1489 13345 1501 13379
rect 1535 13376 1547 13379
rect 1946 13376 1952 13388
rect 1535 13348 1952 13376
rect 1535 13345 1547 13348
rect 1489 13339 1547 13345
rect 1946 13336 1952 13348
rect 2004 13336 2010 13388
rect 2130 13336 2136 13388
rect 2188 13376 2194 13388
rect 2225 13379 2283 13385
rect 2225 13376 2237 13379
rect 2188 13348 2237 13376
rect 2188 13336 2194 13348
rect 2225 13345 2237 13348
rect 2271 13345 2283 13379
rect 2225 13339 2283 13345
rect 2492 13379 2550 13385
rect 2492 13345 2504 13379
rect 2538 13376 2550 13379
rect 2866 13376 2872 13388
rect 2538 13348 2872 13376
rect 2538 13345 2550 13348
rect 2492 13339 2550 13345
rect 2866 13336 2872 13348
rect 2924 13336 2930 13388
rect 4062 13336 4068 13388
rect 4120 13376 4126 13388
rect 4433 13379 4491 13385
rect 4433 13376 4445 13379
rect 4120 13348 4445 13376
rect 4120 13336 4126 13348
rect 4433 13345 4445 13348
rect 4479 13345 4491 13379
rect 5810 13376 5816 13388
rect 4433 13339 4491 13345
rect 4724 13348 5816 13376
rect 4724 13317 4752 13348
rect 5810 13336 5816 13348
rect 5868 13336 5874 13388
rect 7190 13336 7196 13388
rect 7248 13376 7254 13388
rect 7300 13385 7328 13416
rect 8386 13404 8392 13416
rect 8444 13404 8450 13456
rect 10686 13444 10692 13456
rect 9048 13416 10692 13444
rect 9048 13385 9076 13416
rect 10686 13404 10692 13416
rect 10744 13404 10750 13456
rect 12618 13444 12624 13456
rect 11624 13416 12624 13444
rect 7285 13379 7343 13385
rect 7285 13376 7297 13379
rect 7248 13348 7297 13376
rect 7248 13336 7254 13348
rect 7285 13345 7297 13348
rect 7331 13345 7343 13379
rect 7285 13339 7343 13345
rect 8205 13379 8263 13385
rect 8205 13345 8217 13379
rect 8251 13376 8263 13379
rect 9033 13379 9091 13385
rect 8251 13348 8984 13376
rect 8251 13345 8263 13348
rect 8205 13339 8263 13345
rect 4709 13311 4767 13317
rect 4709 13277 4721 13311
rect 4755 13277 4767 13311
rect 4709 13271 4767 13277
rect 4798 13268 4804 13320
rect 4856 13308 4862 13320
rect 5629 13311 5687 13317
rect 5629 13308 5641 13311
rect 4856 13280 5641 13308
rect 4856 13268 4862 13280
rect 5629 13277 5641 13280
rect 5675 13277 5687 13311
rect 5629 13271 5687 13277
rect 5718 13268 5724 13320
rect 5776 13308 5782 13320
rect 6641 13311 6699 13317
rect 6641 13308 6653 13311
rect 5776 13280 6653 13308
rect 5776 13268 5782 13280
rect 6641 13277 6653 13280
rect 6687 13277 6699 13311
rect 8478 13308 8484 13320
rect 8439 13280 8484 13308
rect 6641 13271 6699 13277
rect 8478 13268 8484 13280
rect 8536 13268 8542 13320
rect 8956 13308 8984 13348
rect 9033 13345 9045 13379
rect 9079 13345 9091 13379
rect 9033 13339 9091 13345
rect 9769 13379 9827 13385
rect 9769 13345 9781 13379
rect 9815 13376 9827 13379
rect 9858 13376 9864 13388
rect 9815 13348 9864 13376
rect 9815 13345 9827 13348
rect 9769 13339 9827 13345
rect 9858 13336 9864 13348
rect 9916 13336 9922 13388
rect 10036 13379 10094 13385
rect 10036 13345 10048 13379
rect 10082 13376 10094 13379
rect 10962 13376 10968 13388
rect 10082 13348 10968 13376
rect 10082 13345 10094 13348
rect 10036 13339 10094 13345
rect 10962 13336 10968 13348
rect 11020 13336 11026 13388
rect 11624 13385 11652 13416
rect 12618 13404 12624 13416
rect 12676 13404 12682 13456
rect 13722 13444 13728 13456
rect 12728 13416 13728 13444
rect 11609 13379 11667 13385
rect 11609 13345 11621 13379
rect 11655 13345 11667 13379
rect 11609 13339 11667 13345
rect 11876 13379 11934 13385
rect 11876 13345 11888 13379
rect 11922 13376 11934 13379
rect 12342 13376 12348 13388
rect 11922 13348 12348 13376
rect 11922 13345 11934 13348
rect 11876 13339 11934 13345
rect 12342 13336 12348 13348
rect 12400 13336 12406 13388
rect 12434 13336 12440 13388
rect 12492 13376 12498 13388
rect 12728 13376 12756 13416
rect 13722 13404 13728 13416
rect 13780 13404 13786 13456
rect 14182 13404 14188 13456
rect 14240 13444 14246 13456
rect 15010 13444 15016 13456
rect 14240 13416 15016 13444
rect 14240 13404 14246 13416
rect 15010 13404 15016 13416
rect 15068 13444 15074 13456
rect 16776 13444 16804 13484
rect 16945 13481 16957 13515
rect 16991 13512 17003 13515
rect 17126 13512 17132 13524
rect 16991 13484 17132 13512
rect 16991 13481 17003 13484
rect 16945 13475 17003 13481
rect 17126 13472 17132 13484
rect 17184 13472 17190 13524
rect 17313 13515 17371 13521
rect 17313 13481 17325 13515
rect 17359 13512 17371 13515
rect 17954 13512 17960 13524
rect 17359 13484 17960 13512
rect 17359 13481 17371 13484
rect 17313 13475 17371 13481
rect 17954 13472 17960 13484
rect 18012 13472 18018 13524
rect 18141 13515 18199 13521
rect 18141 13481 18153 13515
rect 18187 13512 18199 13515
rect 18782 13512 18788 13524
rect 18187 13484 18788 13512
rect 18187 13481 18199 13484
rect 18141 13475 18199 13481
rect 18782 13472 18788 13484
rect 18840 13472 18846 13524
rect 17681 13447 17739 13453
rect 17681 13444 17693 13447
rect 15068 13416 16712 13444
rect 16776 13416 17693 13444
rect 15068 13404 15074 13416
rect 12492 13348 12756 13376
rect 13173 13379 13231 13385
rect 12492 13336 12498 13348
rect 13173 13345 13185 13379
rect 13219 13376 13231 13379
rect 13446 13376 13452 13388
rect 13219 13348 13452 13376
rect 13219 13345 13231 13348
rect 13173 13339 13231 13345
rect 13446 13336 13452 13348
rect 13504 13336 13510 13388
rect 13817 13379 13875 13385
rect 13817 13345 13829 13379
rect 13863 13376 13875 13379
rect 13906 13376 13912 13388
rect 13863 13348 13912 13376
rect 13863 13345 13875 13348
rect 13817 13339 13875 13345
rect 13906 13336 13912 13348
rect 13964 13376 13970 13388
rect 14277 13379 14335 13385
rect 14277 13376 14289 13379
rect 13964 13348 14289 13376
rect 13964 13336 13970 13348
rect 14277 13345 14289 13348
rect 14323 13376 14335 13379
rect 15102 13376 15108 13388
rect 14323 13348 15108 13376
rect 14323 13345 14335 13348
rect 14277 13339 14335 13345
rect 15102 13336 15108 13348
rect 15160 13336 15166 13388
rect 15289 13379 15347 13385
rect 15289 13345 15301 13379
rect 15335 13376 15347 13379
rect 15378 13376 15384 13388
rect 15335 13348 15384 13376
rect 15335 13345 15347 13348
rect 15289 13339 15347 13345
rect 15378 13336 15384 13348
rect 15436 13336 15442 13388
rect 15562 13336 15568 13388
rect 15620 13376 15626 13388
rect 15841 13379 15899 13385
rect 15841 13376 15853 13379
rect 15620 13348 15853 13376
rect 15620 13336 15626 13348
rect 15841 13345 15853 13348
rect 15887 13345 15899 13379
rect 15841 13339 15899 13345
rect 15930 13336 15936 13388
rect 15988 13376 15994 13388
rect 16684 13385 16712 13416
rect 16960 13388 16988 13416
rect 17681 13413 17693 13416
rect 17727 13413 17739 13447
rect 17681 13407 17739 13413
rect 18414 13404 18420 13456
rect 18472 13444 18478 13456
rect 18601 13447 18659 13453
rect 18601 13444 18613 13447
rect 18472 13416 18613 13444
rect 18472 13404 18478 13416
rect 18601 13413 18613 13416
rect 18647 13413 18659 13447
rect 20898 13444 20904 13456
rect 18601 13407 18659 13413
rect 19076 13416 20904 13444
rect 16669 13379 16727 13385
rect 15988 13348 16033 13376
rect 15988 13336 15994 13348
rect 16669 13345 16681 13379
rect 16715 13345 16727 13379
rect 16669 13339 16727 13345
rect 16758 13336 16764 13388
rect 16816 13376 16822 13388
rect 16816 13348 16861 13376
rect 16816 13336 16822 13348
rect 16942 13336 16948 13388
rect 17000 13336 17006 13388
rect 18509 13379 18567 13385
rect 18509 13345 18521 13379
rect 18555 13376 18567 13379
rect 18966 13376 18972 13388
rect 18555 13348 18972 13376
rect 18555 13345 18567 13348
rect 18509 13339 18567 13345
rect 18966 13336 18972 13348
rect 19024 13336 19030 13388
rect 9214 13308 9220 13320
rect 8956 13280 9220 13308
rect 9214 13268 9220 13280
rect 9272 13268 9278 13320
rect 13354 13268 13360 13320
rect 13412 13308 13418 13320
rect 14369 13311 14427 13317
rect 14369 13308 14381 13311
rect 13412 13280 14381 13308
rect 13412 13268 13418 13280
rect 14369 13277 14381 13280
rect 14415 13277 14427 13311
rect 14369 13271 14427 13277
rect 14553 13311 14611 13317
rect 14553 13277 14565 13311
rect 14599 13308 14611 13311
rect 14642 13308 14648 13320
rect 14599 13280 14648 13308
rect 14599 13277 14611 13280
rect 14553 13271 14611 13277
rect 14642 13268 14648 13280
rect 14700 13308 14706 13320
rect 15470 13308 15476 13320
rect 14700 13280 15476 13308
rect 14700 13268 14706 13280
rect 15470 13268 15476 13280
rect 15528 13268 15534 13320
rect 16022 13308 16028 13320
rect 15983 13280 16028 13308
rect 16022 13268 16028 13280
rect 16080 13268 16086 13320
rect 17773 13311 17831 13317
rect 17773 13277 17785 13311
rect 17819 13277 17831 13311
rect 17773 13271 17831 13277
rect 3602 13240 3608 13252
rect 3563 13212 3608 13240
rect 3602 13200 3608 13212
rect 3660 13200 3666 13252
rect 4522 13200 4528 13252
rect 4580 13240 4586 13252
rect 4580 13212 6960 13240
rect 4580 13200 4586 13212
rect 6932 13184 6960 13212
rect 10695 13212 11284 13240
rect 6914 13132 6920 13184
rect 6972 13172 6978 13184
rect 7101 13175 7159 13181
rect 7101 13172 7113 13175
rect 6972 13144 7113 13172
rect 6972 13132 6978 13144
rect 7101 13141 7113 13144
rect 7147 13141 7159 13175
rect 7101 13135 7159 13141
rect 7837 13175 7895 13181
rect 7837 13141 7849 13175
rect 7883 13172 7895 13175
rect 9674 13172 9680 13184
rect 7883 13144 9680 13172
rect 7883 13141 7895 13144
rect 7837 13135 7895 13141
rect 9674 13132 9680 13144
rect 9732 13132 9738 13184
rect 10042 13132 10048 13184
rect 10100 13172 10106 13184
rect 10695 13172 10723 13212
rect 11146 13172 11152 13184
rect 10100 13144 10723 13172
rect 11107 13144 11152 13172
rect 10100 13132 10106 13144
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 11256 13172 11284 13212
rect 12710 13200 12716 13252
rect 12768 13240 12774 13252
rect 15289 13243 15347 13249
rect 15289 13240 15301 13243
rect 12768 13212 15301 13240
rect 12768 13200 12774 13212
rect 15289 13209 15301 13212
rect 15335 13209 15347 13243
rect 15289 13203 15347 13209
rect 15378 13200 15384 13252
rect 15436 13240 15442 13252
rect 17788 13240 17816 13271
rect 17954 13268 17960 13320
rect 18012 13308 18018 13320
rect 18322 13308 18328 13320
rect 18012 13280 18328 13308
rect 18012 13268 18018 13280
rect 18322 13268 18328 13280
rect 18380 13308 18386 13320
rect 18785 13311 18843 13317
rect 18785 13308 18797 13311
rect 18380 13280 18797 13308
rect 18380 13268 18386 13280
rect 18785 13277 18797 13280
rect 18831 13308 18843 13311
rect 19076 13308 19104 13416
rect 20898 13404 20904 13416
rect 20956 13404 20962 13456
rect 19426 13336 19432 13388
rect 19484 13336 19490 13388
rect 19702 13376 19708 13388
rect 19663 13348 19708 13376
rect 19702 13336 19708 13348
rect 19760 13336 19766 13388
rect 19444 13308 19472 13336
rect 19797 13311 19855 13317
rect 19797 13308 19809 13311
rect 18831 13280 19104 13308
rect 19352 13280 19809 13308
rect 18831 13277 18843 13280
rect 18785 13271 18843 13277
rect 19352 13240 19380 13280
rect 19797 13277 19809 13280
rect 19843 13277 19855 13311
rect 19797 13271 19855 13277
rect 19889 13311 19947 13317
rect 19889 13277 19901 13311
rect 19935 13277 19947 13311
rect 19889 13271 19947 13277
rect 15436 13212 17816 13240
rect 19260 13212 19380 13240
rect 15436 13200 15442 13212
rect 12250 13172 12256 13184
rect 11256 13144 12256 13172
rect 12250 13132 12256 13144
rect 12308 13132 12314 13184
rect 12986 13132 12992 13184
rect 13044 13172 13050 13184
rect 13357 13175 13415 13181
rect 13044 13144 13089 13172
rect 13044 13132 13050 13144
rect 13357 13141 13369 13175
rect 13403 13172 13415 13175
rect 13722 13172 13728 13184
rect 13403 13144 13728 13172
rect 13403 13141 13415 13144
rect 13357 13135 13415 13141
rect 13722 13132 13728 13144
rect 13780 13132 13786 13184
rect 13906 13172 13912 13184
rect 13867 13144 13912 13172
rect 13906 13132 13912 13144
rect 13964 13132 13970 13184
rect 14458 13132 14464 13184
rect 14516 13172 14522 13184
rect 14918 13172 14924 13184
rect 14516 13144 14924 13172
rect 14516 13132 14522 13144
rect 14918 13132 14924 13144
rect 14976 13132 14982 13184
rect 15470 13172 15476 13184
rect 15431 13144 15476 13172
rect 15470 13132 15476 13144
rect 15528 13132 15534 13184
rect 16390 13132 16396 13184
rect 16448 13172 16454 13184
rect 16485 13175 16543 13181
rect 16485 13172 16497 13175
rect 16448 13144 16497 13172
rect 16448 13132 16454 13144
rect 16485 13141 16497 13144
rect 16531 13172 16543 13175
rect 17862 13172 17868 13184
rect 16531 13144 17868 13172
rect 16531 13141 16543 13144
rect 16485 13135 16543 13141
rect 17862 13132 17868 13144
rect 17920 13132 17926 13184
rect 19260 13181 19288 13212
rect 19904 13184 19932 13271
rect 19245 13175 19303 13181
rect 19245 13141 19257 13175
rect 19291 13141 19303 13175
rect 19245 13135 19303 13141
rect 19334 13132 19340 13184
rect 19392 13172 19398 13184
rect 19392 13144 19437 13172
rect 19392 13132 19398 13144
rect 19886 13132 19892 13184
rect 19944 13132 19950 13184
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 1486 12928 1492 12980
rect 1544 12968 1550 12980
rect 1857 12971 1915 12977
rect 1857 12968 1869 12971
rect 1544 12940 1869 12968
rect 1544 12928 1550 12940
rect 1857 12937 1869 12940
rect 1903 12937 1915 12971
rect 4062 12968 4068 12980
rect 4023 12940 4068 12968
rect 1857 12931 1915 12937
rect 4062 12928 4068 12940
rect 4120 12928 4126 12980
rect 4246 12928 4252 12980
rect 4304 12968 4310 12980
rect 4304 12940 6040 12968
rect 4304 12928 4310 12940
rect 3970 12860 3976 12912
rect 4028 12900 4034 12912
rect 6012 12900 6040 12940
rect 6086 12928 6092 12980
rect 6144 12968 6150 12980
rect 6273 12971 6331 12977
rect 6273 12968 6285 12971
rect 6144 12940 6285 12968
rect 6144 12928 6150 12940
rect 6273 12937 6285 12940
rect 6319 12937 6331 12971
rect 7190 12968 7196 12980
rect 7151 12940 7196 12968
rect 6273 12931 6331 12937
rect 7190 12928 7196 12940
rect 7248 12928 7254 12980
rect 8478 12928 8484 12980
rect 8536 12968 8542 12980
rect 8938 12968 8944 12980
rect 8536 12940 8944 12968
rect 8536 12928 8542 12940
rect 8938 12928 8944 12940
rect 8996 12928 9002 12980
rect 9214 12968 9220 12980
rect 9175 12940 9220 12968
rect 9214 12928 9220 12940
rect 9272 12928 9278 12980
rect 10505 12971 10563 12977
rect 10505 12937 10517 12971
rect 10551 12968 10563 12971
rect 13998 12968 14004 12980
rect 10551 12940 14004 12968
rect 10551 12937 10563 12940
rect 10505 12931 10563 12937
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 14182 12968 14188 12980
rect 14143 12940 14188 12968
rect 14182 12928 14188 12940
rect 14240 12928 14246 12980
rect 15286 12968 15292 12980
rect 14568 12940 15292 12968
rect 6638 12900 6644 12912
rect 4028 12872 5764 12900
rect 6012 12872 6644 12900
rect 4028 12860 4034 12872
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12832 2559 12835
rect 2866 12832 2872 12844
rect 2547 12804 2872 12832
rect 2547 12801 2559 12804
rect 2501 12795 2559 12801
rect 2866 12792 2872 12804
rect 2924 12792 2930 12844
rect 3694 12832 3700 12844
rect 3655 12804 3700 12832
rect 3694 12792 3700 12804
rect 3752 12792 3758 12844
rect 4709 12835 4767 12841
rect 4709 12801 4721 12835
rect 4755 12832 4767 12835
rect 4798 12832 4804 12844
rect 4755 12804 4804 12832
rect 4755 12801 4767 12804
rect 4709 12795 4767 12801
rect 4798 12792 4804 12804
rect 4856 12792 4862 12844
rect 5626 12832 5632 12844
rect 5587 12804 5632 12832
rect 5626 12792 5632 12804
rect 5684 12792 5690 12844
rect 5736 12832 5764 12872
rect 6638 12860 6644 12872
rect 6696 12860 6702 12912
rect 8570 12860 8576 12912
rect 8628 12900 8634 12912
rect 8628 12872 11192 12900
rect 8628 12860 8634 12872
rect 9033 12835 9091 12841
rect 5736 12804 7696 12832
rect 3421 12767 3479 12773
rect 3421 12733 3433 12767
rect 3467 12764 3479 12767
rect 4246 12764 4252 12776
rect 3467 12736 4252 12764
rect 3467 12733 3479 12736
rect 3421 12727 3479 12733
rect 4246 12724 4252 12736
rect 4304 12724 4310 12776
rect 5442 12764 5448 12776
rect 5403 12736 5448 12764
rect 5442 12724 5448 12736
rect 5500 12724 5506 12776
rect 6089 12767 6147 12773
rect 6089 12733 6101 12767
rect 6135 12733 6147 12767
rect 7374 12764 7380 12776
rect 7335 12736 7380 12764
rect 6089 12727 6147 12733
rect 4433 12699 4491 12705
rect 4433 12696 4445 12699
rect 3068 12668 4445 12696
rect 1670 12588 1676 12640
rect 1728 12628 1734 12640
rect 2225 12631 2283 12637
rect 2225 12628 2237 12631
rect 1728 12600 2237 12628
rect 1728 12588 1734 12600
rect 2225 12597 2237 12600
rect 2271 12597 2283 12631
rect 2225 12591 2283 12597
rect 2317 12631 2375 12637
rect 2317 12597 2329 12631
rect 2363 12628 2375 12631
rect 2958 12628 2964 12640
rect 2363 12600 2964 12628
rect 2363 12597 2375 12600
rect 2317 12591 2375 12597
rect 2958 12588 2964 12600
rect 3016 12588 3022 12640
rect 3068 12637 3096 12668
rect 4433 12665 4445 12668
rect 4479 12665 4491 12699
rect 4433 12659 4491 12665
rect 5166 12656 5172 12708
rect 5224 12696 5230 12708
rect 6104 12696 6132 12727
rect 7374 12724 7380 12736
rect 7432 12724 7438 12776
rect 7561 12767 7619 12773
rect 7561 12733 7573 12767
rect 7607 12733 7619 12767
rect 7668 12764 7696 12804
rect 9033 12801 9045 12835
rect 9079 12832 9091 12835
rect 9769 12835 9827 12841
rect 9769 12832 9781 12835
rect 9079 12804 9781 12832
rect 9079 12801 9091 12804
rect 9033 12795 9091 12801
rect 9769 12801 9781 12804
rect 9815 12801 9827 12835
rect 9769 12795 9827 12801
rect 10318 12792 10324 12844
rect 10376 12792 10382 12844
rect 10502 12792 10508 12844
rect 10560 12832 10566 12844
rect 10686 12832 10692 12844
rect 10560 12804 10692 12832
rect 10560 12792 10566 12804
rect 10686 12792 10692 12804
rect 10744 12792 10750 12844
rect 10870 12792 10876 12844
rect 10928 12832 10934 12844
rect 11057 12835 11115 12841
rect 11057 12832 11069 12835
rect 10928 12804 11069 12832
rect 10928 12792 10934 12804
rect 11057 12801 11069 12804
rect 11103 12801 11115 12835
rect 11057 12795 11115 12801
rect 10336 12764 10364 12792
rect 7668 12736 10364 12764
rect 11164 12764 11192 12872
rect 11514 12860 11520 12912
rect 11572 12900 11578 12912
rect 11790 12900 11796 12912
rect 11572 12872 11796 12900
rect 11572 12860 11578 12872
rect 11790 12860 11796 12872
rect 11848 12860 11854 12912
rect 12526 12832 12532 12844
rect 11348 12804 11919 12832
rect 12487 12804 12532 12832
rect 11348 12764 11376 12804
rect 11164 12736 11376 12764
rect 11793 12767 11851 12773
rect 7561 12727 7619 12733
rect 11793 12733 11805 12767
rect 11839 12733 11851 12767
rect 11891 12764 11919 12804
rect 12526 12792 12532 12804
rect 12584 12792 12590 12844
rect 14568 12841 14596 12940
rect 15286 12928 15292 12940
rect 15344 12928 15350 12980
rect 15930 12928 15936 12980
rect 15988 12968 15994 12980
rect 16209 12971 16267 12977
rect 16209 12968 16221 12971
rect 15988 12940 16221 12968
rect 15988 12928 15994 12940
rect 16209 12937 16221 12940
rect 16255 12937 16267 12971
rect 16209 12931 16267 12937
rect 17862 12928 17868 12980
rect 17920 12968 17926 12980
rect 19429 12971 19487 12977
rect 17920 12940 19279 12968
rect 17920 12928 17926 12940
rect 14553 12835 14611 12841
rect 14553 12801 14565 12835
rect 14599 12801 14611 12835
rect 14553 12795 14611 12801
rect 16666 12792 16672 12844
rect 16724 12832 16730 12844
rect 16761 12835 16819 12841
rect 16761 12832 16773 12835
rect 16724 12804 16773 12832
rect 16724 12792 16730 12804
rect 16761 12801 16773 12804
rect 16807 12801 16819 12835
rect 16761 12795 16819 12801
rect 18056 12835 18114 12841
rect 18056 12801 18068 12835
rect 18102 12832 18114 12835
rect 18102 12804 18184 12832
rect 18102 12801 18114 12804
rect 18056 12795 18114 12801
rect 11891 12736 13851 12764
rect 11793 12727 11851 12733
rect 5224 12668 6132 12696
rect 5224 12656 5230 12668
rect 6822 12656 6828 12708
rect 6880 12696 6886 12708
rect 7190 12696 7196 12708
rect 6880 12668 7196 12696
rect 6880 12656 6886 12668
rect 7190 12656 7196 12668
rect 7248 12696 7254 12708
rect 7576 12696 7604 12727
rect 7248 12668 7604 12696
rect 7828 12699 7886 12705
rect 7248 12656 7254 12668
rect 7828 12665 7840 12699
rect 7874 12696 7886 12699
rect 8202 12696 8208 12708
rect 7874 12668 8208 12696
rect 7874 12665 7886 12668
rect 7828 12659 7886 12665
rect 8202 12656 8208 12668
rect 8260 12696 8266 12708
rect 9033 12699 9091 12705
rect 9033 12696 9045 12699
rect 8260 12668 9045 12696
rect 8260 12656 8266 12668
rect 9033 12665 9045 12668
rect 9079 12665 9091 12699
rect 9033 12659 9091 12665
rect 9677 12699 9735 12705
rect 9677 12665 9689 12699
rect 9723 12696 9735 12699
rect 10042 12696 10048 12708
rect 9723 12668 10048 12696
rect 9723 12665 9735 12668
rect 9677 12659 9735 12665
rect 10042 12656 10048 12668
rect 10100 12656 10106 12708
rect 10134 12656 10140 12708
rect 10192 12696 10198 12708
rect 11808 12696 11836 12727
rect 12066 12696 12072 12708
rect 10192 12668 11836 12696
rect 11891 12668 12072 12696
rect 10192 12656 10198 12668
rect 3053 12631 3111 12637
rect 3053 12597 3065 12631
rect 3099 12597 3111 12631
rect 3053 12591 3111 12597
rect 3234 12588 3240 12640
rect 3292 12628 3298 12640
rect 3513 12631 3571 12637
rect 3513 12628 3525 12631
rect 3292 12600 3525 12628
rect 3292 12588 3298 12600
rect 3513 12597 3525 12600
rect 3559 12597 3571 12631
rect 3513 12591 3571 12597
rect 4525 12631 4583 12637
rect 4525 12597 4537 12631
rect 4571 12628 4583 12631
rect 5077 12631 5135 12637
rect 5077 12628 5089 12631
rect 4571 12600 5089 12628
rect 4571 12597 4583 12600
rect 4525 12591 4583 12597
rect 5077 12597 5089 12600
rect 5123 12597 5135 12631
rect 5077 12591 5135 12597
rect 5537 12631 5595 12637
rect 5537 12597 5549 12631
rect 5583 12628 5595 12631
rect 6178 12628 6184 12640
rect 5583 12600 6184 12628
rect 5583 12597 5595 12600
rect 5537 12591 5595 12597
rect 6178 12588 6184 12600
rect 6236 12628 6242 12640
rect 8294 12628 8300 12640
rect 6236 12600 8300 12628
rect 6236 12588 6242 12600
rect 8294 12588 8300 12600
rect 8352 12588 8358 12640
rect 9585 12631 9643 12637
rect 9585 12597 9597 12631
rect 9631 12628 9643 12631
rect 10410 12628 10416 12640
rect 9631 12600 10416 12628
rect 9631 12597 9643 12600
rect 9585 12591 9643 12597
rect 10410 12588 10416 12600
rect 10468 12588 10474 12640
rect 10686 12588 10692 12640
rect 10744 12628 10750 12640
rect 10873 12631 10931 12637
rect 10873 12628 10885 12631
rect 10744 12600 10885 12628
rect 10744 12588 10750 12600
rect 10873 12597 10885 12600
rect 10919 12597 10931 12631
rect 10873 12591 10931 12597
rect 10965 12631 11023 12637
rect 10965 12597 10977 12631
rect 11011 12628 11023 12631
rect 11606 12628 11612 12640
rect 11011 12600 11612 12628
rect 11011 12597 11023 12600
rect 10965 12591 11023 12597
rect 11606 12588 11612 12600
rect 11664 12588 11670 12640
rect 11790 12588 11796 12640
rect 11848 12628 11854 12640
rect 11891 12628 11919 12668
rect 12066 12656 12072 12668
rect 12124 12656 12130 12708
rect 12796 12699 12854 12705
rect 12796 12665 12808 12699
rect 12842 12696 12854 12699
rect 12986 12696 12992 12708
rect 12842 12668 12992 12696
rect 12842 12665 12854 12668
rect 12796 12659 12854 12665
rect 12986 12656 12992 12668
rect 13044 12696 13050 12708
rect 13722 12696 13728 12708
rect 13044 12668 13728 12696
rect 13044 12656 13050 12668
rect 13722 12656 13728 12668
rect 13780 12656 13786 12708
rect 13823 12696 13851 12736
rect 13998 12724 14004 12776
rect 14056 12764 14062 12776
rect 14274 12764 14280 12776
rect 14056 12736 14280 12764
rect 14056 12724 14062 12736
rect 14274 12724 14280 12736
rect 14332 12724 14338 12776
rect 14369 12767 14427 12773
rect 14369 12733 14381 12767
rect 14415 12764 14427 12767
rect 14458 12764 14464 12776
rect 14415 12736 14464 12764
rect 14415 12733 14427 12736
rect 14369 12727 14427 12733
rect 14458 12724 14464 12736
rect 14516 12724 14522 12776
rect 15378 12764 15384 12776
rect 14752 12736 15384 12764
rect 14752 12696 14780 12736
rect 15378 12724 15384 12736
rect 15436 12724 15442 12776
rect 17218 12764 17224 12776
rect 15479 12736 16804 12764
rect 17179 12736 17224 12764
rect 13823 12668 14780 12696
rect 14820 12699 14878 12705
rect 14820 12665 14832 12699
rect 14866 12696 14878 12699
rect 15010 12696 15016 12708
rect 14866 12668 15016 12696
rect 14866 12665 14878 12668
rect 14820 12659 14878 12665
rect 15010 12656 15016 12668
rect 15068 12656 15074 12708
rect 11848 12600 11919 12628
rect 11977 12631 12035 12637
rect 11848 12588 11854 12600
rect 11977 12597 11989 12631
rect 12023 12628 12035 12631
rect 12434 12628 12440 12640
rect 12023 12600 12440 12628
rect 12023 12597 12035 12600
rect 11977 12591 12035 12597
rect 12434 12588 12440 12600
rect 12492 12588 12498 12640
rect 12710 12588 12716 12640
rect 12768 12628 12774 12640
rect 13909 12631 13967 12637
rect 13909 12628 13921 12631
rect 12768 12600 13921 12628
rect 12768 12588 12774 12600
rect 13909 12597 13921 12600
rect 13955 12628 13967 12631
rect 15479 12628 15507 12736
rect 16482 12656 16488 12708
rect 16540 12696 16546 12708
rect 16669 12699 16727 12705
rect 16669 12696 16681 12699
rect 16540 12668 16681 12696
rect 16540 12656 16546 12668
rect 16669 12665 16681 12668
rect 16715 12665 16727 12699
rect 16776 12696 16804 12736
rect 17218 12724 17224 12736
rect 17276 12724 17282 12776
rect 18156 12764 18184 12804
rect 19251 12764 19279 12940
rect 19429 12937 19441 12971
rect 19475 12968 19487 12971
rect 19518 12968 19524 12980
rect 19475 12940 19524 12968
rect 19475 12937 19487 12940
rect 19429 12931 19487 12937
rect 19518 12928 19524 12940
rect 19576 12928 19582 12980
rect 20898 12968 20904 12980
rect 20859 12940 20904 12968
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 19536 12832 19564 12928
rect 19536 12804 19656 12832
rect 19521 12767 19579 12773
rect 19521 12764 19533 12767
rect 18156 12736 18828 12764
rect 17497 12699 17555 12705
rect 16776 12668 17439 12696
rect 16669 12659 16727 12665
rect 15930 12628 15936 12640
rect 13955 12600 15507 12628
rect 15891 12600 15936 12628
rect 13955 12597 13967 12600
rect 13909 12591 13967 12597
rect 15930 12588 15936 12600
rect 15988 12588 15994 12640
rect 16577 12631 16635 12637
rect 16577 12597 16589 12631
rect 16623 12628 16635 12631
rect 17310 12628 17316 12640
rect 16623 12600 17316 12628
rect 16623 12597 16635 12600
rect 16577 12591 16635 12597
rect 17310 12588 17316 12600
rect 17368 12588 17374 12640
rect 17411 12628 17439 12668
rect 17497 12665 17509 12699
rect 17543 12696 17555 12699
rect 17954 12696 17960 12708
rect 17543 12668 17960 12696
rect 17543 12665 17555 12668
rect 17497 12659 17555 12665
rect 17954 12656 17960 12668
rect 18012 12656 18018 12708
rect 18046 12656 18052 12708
rect 18104 12696 18110 12708
rect 18156 12696 18184 12736
rect 18322 12705 18328 12708
rect 18104 12668 18184 12696
rect 18104 12656 18110 12668
rect 18316 12659 18328 12705
rect 18380 12696 18386 12708
rect 18800 12696 18828 12736
rect 19251 12736 19533 12764
rect 19251 12696 19279 12736
rect 19521 12733 19533 12736
rect 19567 12733 19579 12767
rect 19628 12764 19656 12804
rect 19777 12767 19835 12773
rect 19777 12764 19789 12767
rect 19628 12736 19789 12764
rect 19521 12727 19579 12733
rect 19777 12733 19789 12736
rect 19823 12733 19835 12767
rect 19777 12727 19835 12733
rect 18380 12668 18416 12696
rect 18800 12668 19279 12696
rect 18322 12656 18328 12659
rect 18380 12656 18386 12668
rect 20346 12628 20352 12640
rect 17411 12600 20352 12628
rect 20346 12588 20352 12600
rect 20404 12588 20410 12640
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 2314 12384 2320 12436
rect 2372 12424 2378 12436
rect 2372 12396 2452 12424
rect 2372 12384 2378 12396
rect 2130 12356 2136 12368
rect 1504 12328 2136 12356
rect 1504 12297 1532 12328
rect 2130 12316 2136 12328
rect 2188 12316 2194 12368
rect 1489 12291 1547 12297
rect 1489 12257 1501 12291
rect 1535 12257 1547 12291
rect 1489 12251 1547 12257
rect 1756 12291 1814 12297
rect 1756 12257 1768 12291
rect 1802 12288 1814 12291
rect 2314 12288 2320 12300
rect 1802 12260 2320 12288
rect 1802 12257 1814 12260
rect 1756 12251 1814 12257
rect 2314 12248 2320 12260
rect 2372 12248 2378 12300
rect 2424 12288 2452 12396
rect 2498 12384 2504 12436
rect 2556 12384 2562 12436
rect 2866 12424 2872 12436
rect 2827 12396 2872 12424
rect 2866 12384 2872 12396
rect 2924 12384 2930 12436
rect 3326 12424 3332 12436
rect 3287 12396 3332 12424
rect 3326 12384 3332 12396
rect 3384 12384 3390 12436
rect 4154 12384 4160 12436
rect 4212 12424 4218 12436
rect 4433 12427 4491 12433
rect 4433 12424 4445 12427
rect 4212 12396 4445 12424
rect 4212 12384 4218 12396
rect 4433 12393 4445 12396
rect 4479 12393 4491 12427
rect 4433 12387 4491 12393
rect 4525 12427 4583 12433
rect 4525 12393 4537 12427
rect 4571 12424 4583 12427
rect 5074 12424 5080 12436
rect 4571 12396 5080 12424
rect 4571 12393 4583 12396
rect 4525 12387 4583 12393
rect 5074 12384 5080 12396
rect 5132 12384 5138 12436
rect 7006 12384 7012 12436
rect 7064 12424 7070 12436
rect 7282 12424 7288 12436
rect 7064 12396 7288 12424
rect 7064 12384 7070 12396
rect 7282 12384 7288 12396
rect 7340 12384 7346 12436
rect 9674 12384 9680 12436
rect 9732 12424 9738 12436
rect 10137 12427 10195 12433
rect 10137 12424 10149 12427
rect 9732 12396 10149 12424
rect 9732 12384 9738 12396
rect 10137 12393 10149 12396
rect 10183 12393 10195 12427
rect 11790 12424 11796 12436
rect 10137 12387 10195 12393
rect 11072 12396 11652 12424
rect 11751 12396 11796 12424
rect 2516 12356 2544 12384
rect 2590 12356 2596 12368
rect 2516 12328 2596 12356
rect 2590 12316 2596 12328
rect 2648 12316 2654 12368
rect 7926 12316 7932 12368
rect 7984 12356 7990 12368
rect 11072 12356 11100 12396
rect 7984 12328 11100 12356
rect 11149 12359 11207 12365
rect 7984 12316 7990 12328
rect 11149 12325 11161 12359
rect 11195 12325 11207 12359
rect 11624 12356 11652 12396
rect 11790 12384 11796 12396
rect 11848 12384 11854 12436
rect 12161 12427 12219 12433
rect 12161 12393 12173 12427
rect 12207 12424 12219 12427
rect 12989 12427 13047 12433
rect 12207 12396 12940 12424
rect 12207 12393 12219 12396
rect 12161 12387 12219 12393
rect 12802 12356 12808 12368
rect 11624 12328 12808 12356
rect 11149 12319 11207 12325
rect 2498 12288 2504 12300
rect 2424 12260 2504 12288
rect 2498 12248 2504 12260
rect 2556 12248 2562 12300
rect 3142 12288 3148 12300
rect 3103 12260 3148 12288
rect 3142 12248 3148 12260
rect 3200 12248 3206 12300
rect 5442 12248 5448 12300
rect 5500 12288 5506 12300
rect 5804 12291 5862 12297
rect 5804 12288 5816 12291
rect 5500 12260 5816 12288
rect 5500 12248 5506 12260
rect 5804 12257 5816 12260
rect 5850 12288 5862 12291
rect 7190 12288 7196 12300
rect 5850 12260 7052 12288
rect 7151 12260 7196 12288
rect 5850 12257 5862 12260
rect 5804 12251 5862 12257
rect 3694 12180 3700 12232
rect 3752 12220 3758 12232
rect 4617 12223 4675 12229
rect 4617 12220 4629 12223
rect 3752 12192 4629 12220
rect 3752 12180 3758 12192
rect 4617 12189 4629 12192
rect 4663 12189 4675 12223
rect 4617 12183 4675 12189
rect 5537 12223 5595 12229
rect 5537 12189 5549 12223
rect 5583 12189 5595 12223
rect 5537 12183 5595 12189
rect 4522 12112 4528 12164
rect 4580 12152 4586 12164
rect 4890 12152 4896 12164
rect 4580 12124 4896 12152
rect 4580 12112 4586 12124
rect 4890 12112 4896 12124
rect 4948 12112 4954 12164
rect 3602 12044 3608 12096
rect 3660 12084 3666 12096
rect 4065 12087 4123 12093
rect 4065 12084 4077 12087
rect 3660 12056 4077 12084
rect 3660 12044 3666 12056
rect 4065 12053 4077 12056
rect 4111 12053 4123 12087
rect 5552 12084 5580 12183
rect 6730 12084 6736 12096
rect 5552 12056 6736 12084
rect 4065 12047 4123 12053
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 6914 12084 6920 12096
rect 6875 12056 6920 12084
rect 6914 12044 6920 12056
rect 6972 12044 6978 12096
rect 7024 12084 7052 12260
rect 7190 12248 7196 12260
rect 7248 12248 7254 12300
rect 7460 12291 7518 12297
rect 7460 12288 7472 12291
rect 7300 12260 7472 12288
rect 7300 12220 7328 12260
rect 7460 12257 7472 12260
rect 7506 12288 7518 12291
rect 7834 12288 7840 12300
rect 7506 12260 7840 12288
rect 7506 12257 7518 12260
rect 7460 12251 7518 12257
rect 7834 12248 7840 12260
rect 7892 12248 7898 12300
rect 8018 12248 8024 12300
rect 8076 12288 8082 12300
rect 10045 12291 10103 12297
rect 10045 12288 10057 12291
rect 8076 12260 10057 12288
rect 8076 12248 8082 12260
rect 10045 12257 10057 12260
rect 10091 12257 10103 12291
rect 11054 12288 11060 12300
rect 11015 12260 11060 12288
rect 10045 12251 10103 12257
rect 11054 12248 11060 12260
rect 11112 12248 11118 12300
rect 10229 12223 10287 12229
rect 10229 12220 10241 12223
rect 7208 12192 7328 12220
rect 8588 12192 10241 12220
rect 7208 12164 7236 12192
rect 7190 12112 7196 12164
rect 7248 12112 7254 12164
rect 8588 12161 8616 12192
rect 10229 12189 10241 12192
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 11164 12164 11192 12319
rect 12802 12316 12808 12328
rect 12860 12316 12866 12368
rect 12912 12356 12940 12396
rect 12989 12393 13001 12427
rect 13035 12424 13047 12427
rect 13630 12424 13636 12436
rect 13035 12396 13636 12424
rect 13035 12393 13047 12396
rect 12989 12387 13047 12393
rect 13630 12384 13636 12396
rect 13688 12384 13694 12436
rect 15286 12384 15292 12436
rect 15344 12424 15350 12436
rect 16390 12424 16396 12436
rect 15344 12396 16396 12424
rect 15344 12384 15350 12396
rect 16390 12384 16396 12396
rect 16448 12384 16454 12436
rect 16942 12384 16948 12436
rect 17000 12424 17006 12436
rect 17037 12427 17095 12433
rect 17037 12424 17049 12427
rect 17000 12396 17049 12424
rect 17000 12384 17006 12396
rect 17037 12393 17049 12396
rect 17083 12393 17095 12427
rect 17037 12387 17095 12393
rect 17862 12384 17868 12436
rect 17920 12424 17926 12436
rect 18414 12424 18420 12436
rect 17920 12396 18420 12424
rect 17920 12384 17926 12396
rect 18414 12384 18420 12396
rect 18472 12384 18478 12436
rect 19150 12384 19156 12436
rect 19208 12424 19214 12436
rect 19429 12427 19487 12433
rect 19429 12424 19441 12427
rect 19208 12396 19441 12424
rect 19208 12384 19214 12396
rect 19429 12393 19441 12396
rect 19475 12424 19487 12427
rect 19794 12424 19800 12436
rect 19475 12396 19800 12424
rect 19475 12393 19487 12396
rect 19429 12387 19487 12393
rect 19794 12384 19800 12396
rect 19852 12384 19858 12436
rect 13906 12356 13912 12368
rect 12912 12328 13912 12356
rect 13906 12316 13912 12328
rect 13964 12316 13970 12368
rect 14553 12359 14611 12365
rect 14553 12325 14565 12359
rect 14599 12356 14611 12359
rect 19521 12359 19579 12365
rect 19521 12356 19533 12359
rect 14599 12328 19533 12356
rect 14599 12325 14611 12328
rect 14553 12319 14611 12325
rect 19521 12325 19533 12328
rect 19567 12325 19579 12359
rect 19521 12319 19579 12325
rect 12253 12291 12311 12297
rect 12253 12257 12265 12291
rect 12299 12288 12311 12291
rect 12618 12288 12624 12300
rect 12299 12260 12624 12288
rect 12299 12257 12311 12260
rect 12253 12251 12311 12257
rect 12618 12248 12624 12260
rect 12676 12248 12682 12300
rect 13354 12288 13360 12300
rect 13315 12260 13360 12288
rect 13354 12248 13360 12260
rect 13412 12248 13418 12300
rect 15286 12288 15292 12300
rect 15247 12260 15292 12288
rect 15286 12248 15292 12260
rect 15344 12248 15350 12300
rect 15545 12291 15603 12297
rect 15545 12288 15557 12291
rect 15396 12260 15557 12288
rect 11241 12223 11299 12229
rect 11241 12189 11253 12223
rect 11287 12189 11299 12223
rect 11241 12183 11299 12189
rect 11517 12223 11575 12229
rect 11517 12189 11529 12223
rect 11563 12220 11575 12223
rect 12437 12223 12495 12229
rect 11563 12192 12388 12220
rect 11563 12189 11575 12192
rect 11517 12183 11575 12189
rect 8573 12155 8631 12161
rect 8573 12121 8585 12155
rect 8619 12121 8631 12155
rect 8573 12115 8631 12121
rect 8588 12084 8616 12115
rect 8754 12112 8760 12164
rect 8812 12152 8818 12164
rect 10689 12155 10747 12161
rect 10689 12152 10701 12155
rect 8812 12124 10701 12152
rect 8812 12112 8818 12124
rect 10689 12121 10701 12124
rect 10735 12121 10747 12155
rect 10689 12115 10747 12121
rect 11146 12112 11152 12164
rect 11204 12112 11210 12164
rect 7024 12056 8616 12084
rect 8662 12044 8668 12096
rect 8720 12084 8726 12096
rect 9677 12087 9735 12093
rect 9677 12084 9689 12087
rect 8720 12056 9689 12084
rect 8720 12044 8726 12056
rect 9677 12053 9689 12056
rect 9723 12053 9735 12087
rect 9677 12047 9735 12053
rect 9766 12044 9772 12096
rect 9824 12084 9830 12096
rect 11256 12084 11284 12183
rect 11330 12112 11336 12164
rect 11388 12152 11394 12164
rect 11698 12152 11704 12164
rect 11388 12124 11704 12152
rect 11388 12112 11394 12124
rect 11698 12112 11704 12124
rect 11756 12112 11762 12164
rect 12360 12152 12388 12192
rect 12437 12189 12449 12223
rect 12483 12220 12495 12223
rect 13262 12220 13268 12232
rect 12483 12192 13268 12220
rect 12483 12189 12495 12192
rect 12437 12183 12495 12189
rect 13262 12180 13268 12192
rect 13320 12180 13326 12232
rect 13449 12223 13507 12229
rect 13449 12189 13461 12223
rect 13495 12220 13507 12223
rect 13538 12220 13544 12232
rect 13495 12192 13544 12220
rect 13495 12189 13507 12192
rect 13449 12183 13507 12189
rect 13538 12180 13544 12192
rect 13596 12180 13602 12232
rect 13633 12223 13691 12229
rect 13633 12189 13645 12223
rect 13679 12220 13691 12223
rect 14182 12220 14188 12232
rect 13679 12192 14188 12220
rect 13679 12189 13691 12192
rect 13633 12183 13691 12189
rect 14182 12180 14188 12192
rect 14240 12180 14246 12232
rect 14642 12220 14648 12232
rect 14603 12192 14648 12220
rect 14642 12180 14648 12192
rect 14700 12180 14706 12232
rect 14829 12223 14887 12229
rect 14829 12189 14841 12223
rect 14875 12220 14887 12223
rect 15010 12220 15016 12232
rect 14875 12192 15016 12220
rect 14875 12189 14887 12192
rect 14829 12183 14887 12189
rect 15010 12180 15016 12192
rect 15068 12180 15074 12232
rect 15396 12220 15424 12260
rect 15545 12257 15557 12260
rect 15591 12288 15603 12291
rect 15930 12288 15936 12300
rect 15591 12260 15936 12288
rect 15591 12257 15603 12260
rect 15545 12251 15603 12257
rect 15930 12248 15936 12260
rect 15988 12248 15994 12300
rect 16022 12248 16028 12300
rect 16080 12288 16086 12300
rect 16850 12288 16856 12300
rect 16080 12260 16344 12288
rect 16811 12260 16856 12288
rect 16080 12248 16086 12260
rect 15304 12192 15424 12220
rect 16316 12220 16344 12260
rect 16850 12248 16856 12260
rect 16908 12248 16914 12300
rect 17589 12291 17647 12297
rect 17589 12257 17601 12291
rect 17635 12257 17647 12291
rect 18046 12288 18052 12300
rect 18007 12260 18052 12288
rect 17589 12251 17647 12257
rect 17604 12220 17632 12251
rect 18046 12248 18052 12260
rect 18104 12248 18110 12300
rect 18138 12248 18144 12300
rect 18196 12248 18202 12300
rect 18316 12291 18374 12297
rect 18316 12257 18328 12291
rect 18362 12288 18374 12291
rect 19334 12288 19340 12300
rect 18362 12260 19340 12288
rect 18362 12257 18374 12260
rect 18316 12251 18374 12257
rect 19334 12248 19340 12260
rect 19392 12288 19398 12300
rect 20530 12288 20536 12300
rect 19392 12260 20536 12288
rect 19392 12248 19398 12260
rect 20530 12248 20536 12260
rect 20588 12248 20594 12300
rect 16316 12192 17632 12220
rect 17681 12223 17739 12229
rect 12360 12124 13676 12152
rect 13648 12096 13676 12124
rect 14734 12112 14740 12164
rect 14792 12152 14798 12164
rect 15304 12152 15332 12192
rect 17681 12189 17693 12223
rect 17727 12220 17739 12223
rect 17770 12220 17776 12232
rect 17727 12192 17776 12220
rect 17727 12189 17739 12192
rect 17681 12183 17739 12189
rect 17770 12180 17776 12192
rect 17828 12180 17834 12232
rect 17865 12223 17923 12229
rect 17865 12189 17877 12223
rect 17911 12220 17923 12223
rect 18156 12220 18184 12248
rect 17911 12192 18184 12220
rect 17911 12189 17923 12192
rect 17865 12183 17923 12189
rect 14792 12124 15332 12152
rect 14792 12112 14798 12124
rect 12894 12084 12900 12096
rect 9824 12056 11284 12084
rect 12855 12056 12900 12084
rect 9824 12044 9830 12056
rect 12894 12044 12900 12056
rect 12952 12084 12958 12096
rect 13354 12084 13360 12096
rect 12952 12056 13360 12084
rect 12952 12044 12958 12056
rect 13354 12044 13360 12056
rect 13412 12044 13418 12096
rect 13630 12044 13636 12096
rect 13688 12044 13694 12096
rect 14185 12087 14243 12093
rect 14185 12053 14197 12087
rect 14231 12084 14243 12087
rect 15562 12084 15568 12096
rect 14231 12056 15568 12084
rect 14231 12053 14243 12056
rect 14185 12047 14243 12053
rect 15562 12044 15568 12056
rect 15620 12044 15626 12096
rect 15930 12044 15936 12096
rect 15988 12084 15994 12096
rect 16669 12087 16727 12093
rect 16669 12084 16681 12087
rect 15988 12056 16681 12084
rect 15988 12044 15994 12056
rect 16669 12053 16681 12056
rect 16715 12053 16727 12087
rect 16669 12047 16727 12053
rect 17221 12087 17279 12093
rect 17221 12053 17233 12087
rect 17267 12084 17279 12087
rect 19058 12084 19064 12096
rect 17267 12056 19064 12084
rect 17267 12053 17279 12056
rect 17221 12047 17279 12053
rect 19058 12044 19064 12056
rect 19116 12044 19122 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 2958 11840 2964 11892
rect 3016 11880 3022 11892
rect 3237 11883 3295 11889
rect 3237 11880 3249 11883
rect 3016 11852 3249 11880
rect 3016 11840 3022 11852
rect 3237 11849 3249 11852
rect 3283 11849 3295 11883
rect 3237 11843 3295 11849
rect 3510 11840 3516 11892
rect 3568 11880 3574 11892
rect 4798 11880 4804 11892
rect 3568 11852 4804 11880
rect 3568 11840 3574 11852
rect 4798 11840 4804 11852
rect 4856 11840 4862 11892
rect 5350 11840 5356 11892
rect 5408 11880 5414 11892
rect 5721 11883 5779 11889
rect 5721 11880 5733 11883
rect 5408 11852 5733 11880
rect 5408 11840 5414 11852
rect 5721 11849 5733 11852
rect 5767 11849 5779 11883
rect 5721 11843 5779 11849
rect 7650 11840 7656 11892
rect 7708 11880 7714 11892
rect 7837 11883 7895 11889
rect 7837 11880 7849 11883
rect 7708 11852 7849 11880
rect 7708 11840 7714 11852
rect 7837 11849 7849 11852
rect 7883 11849 7895 11883
rect 8018 11880 8024 11892
rect 7979 11852 8024 11880
rect 7837 11843 7895 11849
rect 8018 11840 8024 11852
rect 8076 11840 8082 11892
rect 8294 11840 8300 11892
rect 8352 11880 8358 11892
rect 9030 11880 9036 11892
rect 8352 11852 9036 11880
rect 8352 11840 8358 11852
rect 9030 11840 9036 11852
rect 9088 11840 9094 11892
rect 9306 11840 9312 11892
rect 9364 11880 9370 11892
rect 11425 11883 11483 11889
rect 11425 11880 11437 11883
rect 9364 11852 11437 11880
rect 9364 11840 9370 11852
rect 11425 11849 11437 11852
rect 11471 11849 11483 11883
rect 13354 11880 13360 11892
rect 11425 11843 11483 11849
rect 12452 11852 13360 11880
rect 3694 11812 3700 11824
rect 2608 11784 3700 11812
rect 1581 11679 1639 11685
rect 1581 11645 1593 11679
rect 1627 11645 1639 11679
rect 1581 11639 1639 11645
rect 1848 11679 1906 11685
rect 1848 11645 1860 11679
rect 1894 11676 1906 11679
rect 2608 11676 2636 11784
rect 3694 11772 3700 11784
rect 3752 11772 3758 11824
rect 4982 11772 4988 11824
rect 5040 11812 5046 11824
rect 7190 11812 7196 11824
rect 5040 11784 7196 11812
rect 5040 11772 5046 11784
rect 7190 11772 7196 11784
rect 7248 11772 7254 11824
rect 7668 11812 7696 11840
rect 7484 11784 7696 11812
rect 7760 11784 9812 11812
rect 3789 11747 3847 11753
rect 3789 11713 3801 11747
rect 3835 11713 3847 11747
rect 4246 11744 4252 11756
rect 4207 11716 4252 11744
rect 3789 11707 3847 11713
rect 3602 11676 3608 11688
rect 1894 11648 2636 11676
rect 3563 11648 3608 11676
rect 1894 11645 1906 11648
rect 1848 11639 1906 11645
rect 1596 11608 1624 11639
rect 3602 11636 3608 11648
rect 3660 11636 3666 11688
rect 2130 11608 2136 11620
rect 1596 11580 2136 11608
rect 2130 11568 2136 11580
rect 2188 11568 2194 11620
rect 3804 11608 3832 11707
rect 4246 11704 4252 11716
rect 4304 11704 4310 11756
rect 5353 11747 5411 11753
rect 5353 11713 5365 11747
rect 5399 11744 5411 11747
rect 5442 11744 5448 11756
rect 5399 11716 5448 11744
rect 5399 11713 5411 11716
rect 5353 11707 5411 11713
rect 5442 11704 5448 11716
rect 5500 11704 5506 11756
rect 6365 11747 6423 11753
rect 6365 11713 6377 11747
rect 6411 11744 6423 11747
rect 6914 11744 6920 11756
rect 6411 11716 6920 11744
rect 6411 11713 6423 11716
rect 6365 11707 6423 11713
rect 6914 11704 6920 11716
rect 6972 11704 6978 11756
rect 7484 11753 7512 11784
rect 7469 11747 7527 11753
rect 7469 11713 7481 11747
rect 7515 11713 7527 11747
rect 7650 11744 7656 11756
rect 7563 11716 7656 11744
rect 7469 11707 7527 11713
rect 7650 11704 7656 11716
rect 7708 11744 7714 11756
rect 7760 11744 7788 11784
rect 7708 11716 7788 11744
rect 7708 11704 7714 11716
rect 7834 11704 7840 11756
rect 7892 11744 7898 11756
rect 8573 11747 8631 11753
rect 8573 11744 8585 11747
rect 7892 11716 8585 11744
rect 7892 11704 7898 11716
rect 8573 11713 8585 11716
rect 8619 11744 8631 11747
rect 8938 11744 8944 11756
rect 8619 11716 8944 11744
rect 8619 11713 8631 11716
rect 8573 11707 8631 11713
rect 6181 11679 6239 11685
rect 6181 11645 6193 11679
rect 6227 11676 6239 11679
rect 8662 11676 8668 11688
rect 6227 11648 8668 11676
rect 6227 11645 6239 11648
rect 6181 11639 6239 11645
rect 8662 11636 8668 11648
rect 8720 11636 8726 11688
rect 8772 11676 8800 11716
rect 8938 11704 8944 11716
rect 8996 11704 9002 11756
rect 9214 11704 9220 11756
rect 9272 11744 9278 11756
rect 9784 11753 9812 11784
rect 10962 11772 10968 11824
rect 11020 11812 11026 11824
rect 11333 11815 11391 11821
rect 11333 11812 11345 11815
rect 11020 11784 11345 11812
rect 11020 11772 11026 11784
rect 11333 11781 11345 11784
rect 11379 11812 11391 11815
rect 12452 11812 12480 11852
rect 13354 11840 13360 11852
rect 13412 11840 13418 11892
rect 15194 11880 15200 11892
rect 15155 11852 15200 11880
rect 15194 11840 15200 11852
rect 15252 11840 15258 11892
rect 16209 11883 16267 11889
rect 16209 11880 16221 11883
rect 15304 11852 16221 11880
rect 11379 11784 12480 11812
rect 14185 11815 14243 11821
rect 11379 11781 11391 11784
rect 11333 11775 11391 11781
rect 14185 11781 14197 11815
rect 14231 11812 14243 11815
rect 15013 11815 15071 11821
rect 14231 11784 14964 11812
rect 14231 11781 14243 11784
rect 14185 11775 14243 11781
rect 9585 11747 9643 11753
rect 9585 11744 9597 11747
rect 9272 11716 9597 11744
rect 9272 11704 9278 11716
rect 9585 11713 9597 11716
rect 9631 11713 9643 11747
rect 9585 11707 9643 11713
rect 9769 11747 9827 11753
rect 9769 11713 9781 11747
rect 9815 11713 9827 11747
rect 9769 11707 9827 11713
rect 9784 11676 9812 11707
rect 9858 11704 9864 11756
rect 9916 11744 9922 11756
rect 9953 11747 10011 11753
rect 9953 11744 9965 11747
rect 9916 11716 9965 11744
rect 9916 11704 9922 11716
rect 9953 11713 9965 11716
rect 9999 11713 10011 11747
rect 11977 11747 12035 11753
rect 11977 11744 11989 11747
rect 9953 11707 10011 11713
rect 10980 11716 11989 11744
rect 10980 11676 11008 11716
rect 11977 11713 11989 11716
rect 12023 11713 12035 11747
rect 14734 11744 14740 11756
rect 14695 11716 14740 11744
rect 11977 11707 12035 11713
rect 14734 11704 14740 11716
rect 14792 11704 14798 11756
rect 14936 11744 14964 11784
rect 15013 11781 15025 11815
rect 15059 11812 15071 11815
rect 15304 11812 15332 11852
rect 16209 11849 16221 11852
rect 16255 11849 16267 11883
rect 17586 11880 17592 11892
rect 17547 11852 17592 11880
rect 16209 11843 16267 11849
rect 17586 11840 17592 11852
rect 17644 11840 17650 11892
rect 17770 11840 17776 11892
rect 17828 11880 17834 11892
rect 19150 11880 19156 11892
rect 17828 11852 19156 11880
rect 17828 11840 17834 11852
rect 19150 11840 19156 11852
rect 19208 11880 19214 11892
rect 19610 11880 19616 11892
rect 19208 11852 19616 11880
rect 19208 11840 19214 11852
rect 19610 11840 19616 11852
rect 19668 11840 19674 11892
rect 20901 11883 20959 11889
rect 20901 11849 20913 11883
rect 20947 11880 20959 11883
rect 21450 11880 21456 11892
rect 20947 11852 21456 11880
rect 20947 11849 20959 11852
rect 20901 11843 20959 11849
rect 21450 11840 21456 11852
rect 21508 11840 21514 11892
rect 15059 11784 15332 11812
rect 19521 11815 19579 11821
rect 15059 11781 15071 11784
rect 15013 11775 15071 11781
rect 19521 11781 19533 11815
rect 19567 11812 19579 11815
rect 19794 11812 19800 11824
rect 19567 11784 19800 11812
rect 19567 11781 19579 11784
rect 19521 11775 19579 11781
rect 19794 11772 19800 11784
rect 19852 11772 19858 11824
rect 15657 11747 15715 11753
rect 15657 11744 15669 11747
rect 14936 11716 15669 11744
rect 15657 11713 15669 11716
rect 15703 11713 15715 11747
rect 15657 11707 15715 11713
rect 15841 11747 15899 11753
rect 15841 11713 15853 11747
rect 15887 11744 15899 11747
rect 15930 11744 15936 11756
rect 15887 11716 15936 11744
rect 15887 11713 15899 11716
rect 15841 11707 15899 11713
rect 15930 11704 15936 11716
rect 15988 11704 15994 11756
rect 16025 11747 16083 11753
rect 16025 11713 16037 11747
rect 16071 11744 16083 11747
rect 16758 11744 16764 11756
rect 16071 11716 16764 11744
rect 16071 11713 16083 11716
rect 16025 11707 16083 11713
rect 16758 11704 16764 11716
rect 16816 11704 16822 11756
rect 16850 11704 16856 11756
rect 16908 11744 16914 11756
rect 20257 11747 20315 11753
rect 20257 11744 20269 11747
rect 16908 11716 20269 11744
rect 16908 11704 16914 11716
rect 20257 11713 20269 11716
rect 20303 11713 20315 11747
rect 20257 11707 20315 11713
rect 11790 11676 11796 11688
rect 8772 11648 9352 11676
rect 9784 11648 11008 11676
rect 11751 11648 11796 11676
rect 6089 11611 6147 11617
rect 6089 11608 6101 11611
rect 2976 11580 3832 11608
rect 4724 11580 6101 11608
rect 2314 11500 2320 11552
rect 2372 11540 2378 11552
rect 2976 11549 3004 11580
rect 2961 11543 3019 11549
rect 2961 11540 2973 11543
rect 2372 11512 2973 11540
rect 2372 11500 2378 11512
rect 2961 11509 2973 11512
rect 3007 11509 3019 11543
rect 2961 11503 3019 11509
rect 3050 11500 3056 11552
rect 3108 11540 3114 11552
rect 4724 11549 4752 11580
rect 6089 11577 6101 11580
rect 6135 11577 6147 11611
rect 9214 11608 9220 11620
rect 6089 11571 6147 11577
rect 7024 11580 9220 11608
rect 3697 11543 3755 11549
rect 3697 11540 3709 11543
rect 3108 11512 3709 11540
rect 3108 11500 3114 11512
rect 3697 11509 3709 11512
rect 3743 11509 3755 11543
rect 3697 11503 3755 11509
rect 4709 11543 4767 11549
rect 4709 11509 4721 11543
rect 4755 11509 4767 11543
rect 5074 11540 5080 11552
rect 5035 11512 5080 11540
rect 4709 11503 4767 11509
rect 5074 11500 5080 11512
rect 5132 11500 5138 11552
rect 5169 11543 5227 11549
rect 5169 11509 5181 11543
rect 5215 11540 5227 11543
rect 6822 11540 6828 11552
rect 5215 11512 6828 11540
rect 5215 11509 5227 11512
rect 5169 11503 5227 11509
rect 6822 11500 6828 11512
rect 6880 11500 6886 11552
rect 7024 11549 7052 11580
rect 9214 11568 9220 11580
rect 9272 11568 9278 11620
rect 9324 11608 9352 11648
rect 11790 11636 11796 11648
rect 11848 11676 11854 11688
rect 12250 11676 12256 11688
rect 11848 11648 12256 11676
rect 11848 11636 11854 11648
rect 12250 11636 12256 11648
rect 12308 11636 12314 11688
rect 12437 11679 12495 11685
rect 12437 11645 12449 11679
rect 12483 11676 12495 11679
rect 12526 11676 12532 11688
rect 12483 11648 12532 11676
rect 12483 11645 12495 11648
rect 12437 11639 12495 11645
rect 12526 11636 12532 11648
rect 12584 11636 12590 11688
rect 15553 11676 15559 11688
rect 15611 11685 15617 11688
rect 12627 11648 15148 11676
rect 15523 11648 15559 11676
rect 10220 11611 10278 11617
rect 9324 11580 10180 11608
rect 7009 11543 7067 11549
rect 7009 11509 7021 11543
rect 7055 11509 7067 11543
rect 7009 11503 7067 11509
rect 7098 11500 7104 11552
rect 7156 11540 7162 11552
rect 7377 11543 7435 11549
rect 7377 11540 7389 11543
rect 7156 11512 7389 11540
rect 7156 11500 7162 11512
rect 7377 11509 7389 11512
rect 7423 11509 7435 11543
rect 8386 11540 8392 11552
rect 8347 11512 8392 11540
rect 7377 11503 7435 11509
rect 8386 11500 8392 11512
rect 8444 11500 8450 11552
rect 8478 11500 8484 11552
rect 8536 11540 8542 11552
rect 9122 11540 9128 11552
rect 8536 11512 8581 11540
rect 9083 11512 9128 11540
rect 8536 11500 8542 11512
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 9493 11543 9551 11549
rect 9493 11509 9505 11543
rect 9539 11540 9551 11543
rect 9582 11540 9588 11552
rect 9539 11512 9588 11540
rect 9539 11509 9551 11512
rect 9493 11503 9551 11509
rect 9582 11500 9588 11512
rect 9640 11500 9646 11552
rect 10152 11540 10180 11580
rect 10220 11577 10232 11611
rect 10266 11608 10278 11611
rect 11606 11608 11612 11620
rect 10266 11580 11612 11608
rect 10266 11577 10278 11580
rect 10220 11571 10278 11577
rect 11606 11568 11612 11580
rect 11664 11608 11670 11620
rect 12627 11608 12655 11648
rect 11664 11580 12655 11608
rect 12704 11611 12762 11617
rect 11664 11568 11670 11580
rect 12704 11577 12716 11611
rect 12750 11608 12762 11611
rect 12802 11608 12808 11620
rect 12750 11580 12808 11608
rect 12750 11577 12762 11580
rect 12704 11571 12762 11577
rect 12802 11568 12808 11580
rect 12860 11568 12866 11620
rect 14645 11611 14703 11617
rect 14645 11577 14657 11611
rect 14691 11608 14703 11611
rect 15013 11611 15071 11617
rect 15013 11608 15025 11611
rect 14691 11580 15025 11608
rect 14691 11577 14703 11580
rect 14645 11571 14703 11577
rect 15013 11577 15025 11580
rect 15059 11577 15071 11611
rect 15120 11608 15148 11648
rect 15553 11636 15559 11648
rect 15611 11639 15623 11685
rect 15611 11636 15617 11639
rect 15746 11636 15752 11688
rect 15804 11676 15810 11688
rect 15804 11648 16160 11676
rect 15804 11636 15810 11648
rect 16132 11608 16160 11648
rect 17126 11636 17132 11688
rect 17184 11676 17190 11688
rect 17405 11679 17463 11685
rect 17405 11676 17417 11679
rect 17184 11648 17417 11676
rect 17184 11636 17190 11648
rect 17405 11645 17417 11648
rect 17451 11645 17463 11679
rect 17405 11639 17463 11645
rect 17678 11636 17684 11688
rect 17736 11676 17742 11688
rect 20714 11676 20720 11688
rect 17736 11648 20116 11676
rect 20675 11648 20720 11676
rect 17736 11636 17742 11648
rect 19610 11608 19616 11620
rect 15120 11580 15516 11608
rect 16132 11580 19616 11608
rect 15013 11571 15071 11577
rect 15488 11552 15516 11580
rect 19610 11568 19616 11580
rect 19668 11568 19674 11620
rect 20088 11617 20116 11648
rect 20714 11636 20720 11648
rect 20772 11636 20778 11688
rect 20073 11611 20131 11617
rect 20073 11577 20085 11611
rect 20119 11608 20131 11611
rect 20530 11608 20536 11620
rect 20119 11580 20536 11608
rect 20119 11577 20131 11580
rect 20073 11571 20131 11577
rect 20530 11568 20536 11580
rect 20588 11568 20594 11620
rect 11790 11540 11796 11552
rect 10152 11512 11796 11540
rect 11790 11500 11796 11512
rect 11848 11500 11854 11552
rect 11885 11543 11943 11549
rect 11885 11509 11897 11543
rect 11931 11540 11943 11543
rect 12986 11540 12992 11552
rect 11931 11512 12992 11540
rect 11931 11509 11943 11512
rect 11885 11503 11943 11509
rect 12986 11500 12992 11512
rect 13044 11500 13050 11552
rect 13817 11543 13875 11549
rect 13817 11509 13829 11543
rect 13863 11540 13875 11543
rect 13906 11540 13912 11552
rect 13863 11512 13912 11540
rect 13863 11509 13875 11512
rect 13817 11503 13875 11509
rect 13906 11500 13912 11512
rect 13964 11500 13970 11552
rect 14553 11543 14611 11549
rect 14553 11509 14565 11543
rect 14599 11540 14611 11543
rect 15286 11540 15292 11552
rect 14599 11512 15292 11540
rect 14599 11509 14611 11512
rect 14553 11503 14611 11509
rect 15286 11500 15292 11512
rect 15344 11500 15350 11552
rect 15470 11500 15476 11552
rect 15528 11500 15534 11552
rect 15562 11500 15568 11552
rect 15620 11540 15626 11552
rect 16025 11543 16083 11549
rect 16025 11540 16037 11543
rect 15620 11512 16037 11540
rect 15620 11500 15626 11512
rect 16025 11509 16037 11512
rect 16071 11509 16083 11543
rect 16025 11503 16083 11509
rect 16390 11500 16396 11552
rect 16448 11540 16454 11552
rect 16577 11543 16635 11549
rect 16577 11540 16589 11543
rect 16448 11512 16589 11540
rect 16448 11500 16454 11512
rect 16577 11509 16589 11512
rect 16623 11509 16635 11543
rect 16577 11503 16635 11509
rect 16666 11500 16672 11552
rect 16724 11540 16730 11552
rect 16724 11512 16769 11540
rect 16724 11500 16730 11512
rect 16942 11500 16948 11552
rect 17000 11540 17006 11552
rect 19705 11543 19763 11549
rect 19705 11540 19717 11543
rect 17000 11512 19717 11540
rect 17000 11500 17006 11512
rect 19705 11509 19717 11512
rect 19751 11509 19763 11543
rect 19705 11503 19763 11509
rect 19794 11500 19800 11552
rect 19852 11540 19858 11552
rect 20165 11543 20223 11549
rect 20165 11540 20177 11543
rect 19852 11512 20177 11540
rect 19852 11500 19858 11512
rect 20165 11509 20177 11512
rect 20211 11540 20223 11543
rect 20714 11540 20720 11552
rect 20211 11512 20720 11540
rect 20211 11509 20223 11512
rect 20165 11503 20223 11509
rect 20714 11500 20720 11512
rect 20772 11500 20778 11552
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 1949 11339 2007 11345
rect 1949 11305 1961 11339
rect 1995 11336 2007 11339
rect 2774 11336 2780 11348
rect 1995 11308 2780 11336
rect 1995 11305 2007 11308
rect 1949 11299 2007 11305
rect 2774 11296 2780 11308
rect 2832 11296 2838 11348
rect 3694 11336 3700 11348
rect 3655 11308 3700 11336
rect 3694 11296 3700 11308
rect 3752 11296 3758 11348
rect 4433 11339 4491 11345
rect 4433 11305 4445 11339
rect 4479 11336 4491 11339
rect 5074 11336 5080 11348
rect 4479 11308 5080 11336
rect 4479 11305 4491 11308
rect 4433 11299 4491 11305
rect 5074 11296 5080 11308
rect 5132 11296 5138 11348
rect 6457 11339 6515 11345
rect 6457 11305 6469 11339
rect 6503 11336 6515 11339
rect 7374 11336 7380 11348
rect 6503 11308 7380 11336
rect 6503 11305 6515 11308
rect 6457 11299 6515 11305
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 7650 11296 7656 11348
rect 7708 11336 7714 11348
rect 8113 11339 8171 11345
rect 8113 11336 8125 11339
rect 7708 11308 8125 11336
rect 7708 11296 7714 11308
rect 8113 11305 8125 11308
rect 8159 11305 8171 11339
rect 8113 11299 8171 11305
rect 8389 11339 8447 11345
rect 8389 11305 8401 11339
rect 8435 11336 8447 11339
rect 8478 11336 8484 11348
rect 8435 11308 8484 11336
rect 8435 11305 8447 11308
rect 8389 11299 8447 11305
rect 8478 11296 8484 11308
rect 8536 11296 8542 11348
rect 9858 11296 9864 11348
rect 9916 11336 9922 11348
rect 10134 11336 10140 11348
rect 9916 11308 10140 11336
rect 9916 11296 9922 11308
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 11054 11296 11060 11348
rect 11112 11336 11118 11348
rect 12802 11336 12808 11348
rect 11112 11308 12808 11336
rect 11112 11296 11118 11308
rect 12802 11296 12808 11308
rect 12860 11296 12866 11348
rect 13725 11339 13783 11345
rect 13725 11305 13737 11339
rect 13771 11336 13783 11339
rect 13814 11336 13820 11348
rect 13771 11308 13820 11336
rect 13771 11305 13783 11308
rect 13725 11299 13783 11305
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 13998 11296 14004 11348
rect 14056 11336 14062 11348
rect 14093 11339 14151 11345
rect 14093 11336 14105 11339
rect 14056 11308 14105 11336
rect 14056 11296 14062 11308
rect 14093 11305 14105 11308
rect 14139 11305 14151 11339
rect 14093 11299 14151 11305
rect 14185 11339 14243 11345
rect 14185 11305 14197 11339
rect 14231 11336 14243 11339
rect 14645 11339 14703 11345
rect 14645 11336 14657 11339
rect 14231 11308 14657 11336
rect 14231 11305 14243 11308
rect 14185 11299 14243 11305
rect 14645 11305 14657 11308
rect 14691 11305 14703 11339
rect 15286 11336 15292 11348
rect 15247 11308 15292 11336
rect 14645 11299 14703 11305
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 15654 11336 15660 11348
rect 15615 11308 15660 11336
rect 15654 11296 15660 11308
rect 15712 11296 15718 11348
rect 16301 11339 16359 11345
rect 16301 11305 16313 11339
rect 16347 11336 16359 11339
rect 16390 11336 16396 11348
rect 16347 11308 16396 11336
rect 16347 11305 16359 11308
rect 16301 11299 16359 11305
rect 16390 11296 16396 11308
rect 16448 11296 16454 11348
rect 16574 11296 16580 11348
rect 16632 11336 16638 11348
rect 16669 11339 16727 11345
rect 16669 11336 16681 11339
rect 16632 11308 16681 11336
rect 16632 11296 16638 11308
rect 16669 11305 16681 11308
rect 16715 11305 16727 11339
rect 16669 11299 16727 11305
rect 17310 11296 17316 11348
rect 17368 11336 17374 11348
rect 17773 11339 17831 11345
rect 17773 11336 17785 11339
rect 17368 11308 17785 11336
rect 17368 11296 17374 11308
rect 17773 11305 17785 11308
rect 17819 11305 17831 11339
rect 18782 11336 18788 11348
rect 18743 11308 18788 11336
rect 17773 11299 17831 11305
rect 18782 11296 18788 11308
rect 18840 11296 18846 11348
rect 19334 11296 19340 11348
rect 19392 11336 19398 11348
rect 20533 11339 20591 11345
rect 20533 11336 20545 11339
rect 19392 11308 20545 11336
rect 19392 11296 19398 11308
rect 20533 11305 20545 11308
rect 20579 11305 20591 11339
rect 20533 11299 20591 11305
rect 20806 11296 20812 11348
rect 20864 11336 20870 11348
rect 20901 11339 20959 11345
rect 20901 11336 20913 11339
rect 20864 11308 20913 11336
rect 20864 11296 20870 11308
rect 20901 11305 20913 11308
rect 20947 11305 20959 11339
rect 20901 11299 20959 11305
rect 2406 11228 2412 11280
rect 2464 11268 2470 11280
rect 4893 11271 4951 11277
rect 4893 11268 4905 11271
rect 2464 11240 4905 11268
rect 2464 11228 2470 11240
rect 4893 11237 4905 11240
rect 4939 11237 4951 11271
rect 4893 11231 4951 11237
rect 6914 11228 6920 11280
rect 6972 11277 6978 11280
rect 6972 11271 7036 11277
rect 6972 11237 6990 11271
rect 7024 11237 7036 11271
rect 8754 11268 8760 11280
rect 8715 11240 8760 11268
rect 6972 11231 7036 11237
rect 6972 11228 6978 11231
rect 8754 11228 8760 11240
rect 8812 11228 8818 11280
rect 9030 11228 9036 11280
rect 9088 11268 9094 11280
rect 9582 11268 9588 11280
rect 9088 11240 9588 11268
rect 9088 11228 9094 11240
rect 9582 11228 9588 11240
rect 9640 11228 9646 11280
rect 11330 11268 11336 11280
rect 10152 11240 11336 11268
rect 10152 11212 10180 11240
rect 11330 11228 11336 11240
rect 11388 11228 11394 11280
rect 12253 11271 12311 11277
rect 12253 11268 12265 11271
rect 11992 11240 12265 11268
rect 1762 11200 1768 11212
rect 1723 11172 1768 11200
rect 1762 11160 1768 11172
rect 1820 11160 1826 11212
rect 2130 11160 2136 11212
rect 2188 11200 2194 11212
rect 2317 11203 2375 11209
rect 2317 11200 2329 11203
rect 2188 11172 2329 11200
rect 2188 11160 2194 11172
rect 2317 11169 2329 11172
rect 2363 11169 2375 11203
rect 2317 11163 2375 11169
rect 2584 11203 2642 11209
rect 2584 11169 2596 11203
rect 2630 11200 2642 11203
rect 3786 11200 3792 11212
rect 2630 11172 3792 11200
rect 2630 11169 2642 11172
rect 2584 11163 2642 11169
rect 3786 11160 3792 11172
rect 3844 11160 3850 11212
rect 4801 11203 4859 11209
rect 4801 11169 4813 11203
rect 4847 11200 4859 11203
rect 5626 11200 5632 11212
rect 4847 11172 5632 11200
rect 4847 11169 4859 11172
rect 4801 11163 4859 11169
rect 5626 11160 5632 11172
rect 5684 11160 5690 11212
rect 5810 11200 5816 11212
rect 5771 11172 5816 11200
rect 5810 11160 5816 11172
rect 5868 11160 5874 11212
rect 6641 11203 6699 11209
rect 6641 11169 6653 11203
rect 6687 11200 6699 11203
rect 8849 11203 8907 11209
rect 6687 11172 8156 11200
rect 6687 11169 6699 11172
rect 6641 11163 6699 11169
rect 4982 11132 4988 11144
rect 4943 11104 4988 11132
rect 4982 11092 4988 11104
rect 5040 11092 5046 11144
rect 5905 11135 5963 11141
rect 5905 11132 5917 11135
rect 5092 11104 5917 11132
rect 5092 11064 5120 11104
rect 5905 11101 5917 11104
rect 5951 11101 5963 11135
rect 5905 11095 5963 11101
rect 5997 11135 6055 11141
rect 5997 11101 6009 11135
rect 6043 11132 6055 11135
rect 6730 11132 6736 11144
rect 6043 11104 6592 11132
rect 6691 11104 6736 11132
rect 6043 11101 6055 11104
rect 5997 11095 6055 11101
rect 3252 11036 5120 11064
rect 5445 11067 5503 11073
rect 2590 10956 2596 11008
rect 2648 10996 2654 11008
rect 3252 10996 3280 11036
rect 5445 11033 5457 11067
rect 5491 11064 5503 11067
rect 6086 11064 6092 11076
rect 5491 11036 6092 11064
rect 5491 11033 5503 11036
rect 5445 11027 5503 11033
rect 6086 11024 6092 11036
rect 6144 11024 6150 11076
rect 6564 11064 6592 11104
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 8128 11064 8156 11172
rect 8849 11169 8861 11203
rect 8895 11200 8907 11203
rect 9674 11200 9680 11212
rect 8895 11172 9680 11200
rect 8895 11169 8907 11172
rect 8849 11163 8907 11169
rect 9674 11160 9680 11172
rect 9732 11200 9738 11212
rect 10134 11200 10140 11212
rect 9732 11172 10140 11200
rect 9732 11160 9738 11172
rect 10134 11160 10140 11172
rect 10192 11160 10198 11212
rect 10318 11160 10324 11212
rect 10376 11200 10382 11212
rect 10505 11203 10563 11209
rect 10505 11200 10517 11203
rect 10376 11172 10517 11200
rect 10376 11160 10382 11172
rect 10505 11169 10517 11172
rect 10551 11169 10563 11203
rect 10505 11163 10563 11169
rect 8202 11092 8208 11144
rect 8260 11132 8266 11144
rect 8941 11135 8999 11141
rect 8941 11132 8953 11135
rect 8260 11104 8953 11132
rect 8260 11092 8266 11104
rect 8941 11101 8953 11104
rect 8987 11101 8999 11135
rect 8941 11095 8999 11101
rect 10042 11092 10048 11144
rect 10100 11132 10106 11144
rect 10778 11132 10784 11144
rect 10100 11104 10784 11132
rect 10100 11092 10106 11104
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 11054 11092 11060 11144
rect 11112 11132 11118 11144
rect 11514 11132 11520 11144
rect 11112 11104 11520 11132
rect 11112 11092 11118 11104
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 11992 11064 12020 11240
rect 12253 11237 12265 11240
rect 12299 11268 12311 11271
rect 14550 11268 14556 11280
rect 12299 11240 14556 11268
rect 12299 11237 12311 11240
rect 12253 11231 12311 11237
rect 14550 11228 14556 11240
rect 14608 11228 14614 11280
rect 14737 11271 14795 11277
rect 14737 11237 14749 11271
rect 14783 11268 14795 11271
rect 19420 11271 19478 11277
rect 14783 11240 16712 11268
rect 14783 11237 14795 11240
rect 14737 11231 14795 11237
rect 13078 11200 13084 11212
rect 13039 11172 13084 11200
rect 13078 11160 13084 11172
rect 13136 11160 13142 11212
rect 13630 11160 13636 11212
rect 13688 11200 13694 11212
rect 15654 11200 15660 11212
rect 13688 11172 15660 11200
rect 13688 11160 13694 11172
rect 15654 11160 15660 11172
rect 15712 11160 15718 11212
rect 15749 11203 15807 11209
rect 15749 11169 15761 11203
rect 15795 11200 15807 11203
rect 16574 11200 16580 11212
rect 15795 11172 16580 11200
rect 15795 11169 15807 11172
rect 15749 11163 15807 11169
rect 16574 11160 16580 11172
rect 16632 11160 16638 11212
rect 16684 11200 16712 11240
rect 16960 11240 18736 11268
rect 16960 11200 16988 11240
rect 16684 11172 16988 11200
rect 17034 11160 17040 11212
rect 17092 11200 17098 11212
rect 17678 11200 17684 11212
rect 17092 11172 17540 11200
rect 17639 11172 17684 11200
rect 17092 11160 17098 11172
rect 12250 11092 12256 11144
rect 12308 11132 12314 11144
rect 12308 11104 12940 11132
rect 12308 11092 12314 11104
rect 6564 11036 6776 11064
rect 8128 11036 12020 11064
rect 2648 10968 3280 10996
rect 6748 10996 6776 11036
rect 12526 11024 12532 11076
rect 12584 11064 12590 11076
rect 12713 11067 12771 11073
rect 12713 11064 12725 11067
rect 12584 11036 12725 11064
rect 12584 11024 12590 11036
rect 12713 11033 12725 11036
rect 12759 11033 12771 11067
rect 12912 11064 12940 11104
rect 12986 11092 12992 11144
rect 13044 11132 13050 11144
rect 13173 11135 13231 11141
rect 13173 11132 13185 11135
rect 13044 11104 13185 11132
rect 13044 11092 13050 11104
rect 13173 11101 13185 11104
rect 13219 11101 13231 11135
rect 13354 11132 13360 11144
rect 13315 11104 13360 11132
rect 13173 11095 13231 11101
rect 13354 11092 13360 11104
rect 13412 11132 13418 11144
rect 14274 11132 14280 11144
rect 13412 11104 14136 11132
rect 14235 11104 14280 11132
rect 13412 11092 13418 11104
rect 13814 11064 13820 11076
rect 12912 11036 13820 11064
rect 12713 11027 12771 11033
rect 13814 11024 13820 11036
rect 13872 11024 13878 11076
rect 14108 11064 14136 11104
rect 14274 11092 14280 11104
rect 14332 11092 14338 11144
rect 14642 11132 14648 11144
rect 14603 11104 14648 11132
rect 14642 11092 14648 11104
rect 14700 11092 14706 11144
rect 15010 11092 15016 11144
rect 15068 11132 15074 11144
rect 15562 11132 15568 11144
rect 15068 11104 15568 11132
rect 15068 11092 15074 11104
rect 15562 11092 15568 11104
rect 15620 11132 15626 11144
rect 16764 11141 16770 11144
rect 15841 11135 15899 11141
rect 15841 11132 15853 11135
rect 15620 11104 15853 11132
rect 15620 11092 15626 11104
rect 15841 11101 15853 11104
rect 15887 11101 15899 11135
rect 15841 11095 15899 11101
rect 16761 11095 16770 11141
rect 16822 11132 16828 11144
rect 16945 11135 17003 11141
rect 16822 11104 16861 11132
rect 16764 11092 16770 11095
rect 16822 11092 16828 11104
rect 16945 11101 16957 11135
rect 16991 11132 17003 11135
rect 17402 11132 17408 11144
rect 16991 11104 17408 11132
rect 16991 11101 17003 11104
rect 16945 11095 17003 11101
rect 17402 11092 17408 11104
rect 17460 11092 17466 11144
rect 17512 11132 17540 11172
rect 17678 11160 17684 11172
rect 17736 11160 17742 11212
rect 17954 11160 17960 11212
rect 18012 11200 18018 11212
rect 18601 11203 18659 11209
rect 18601 11200 18613 11203
rect 18012 11172 18613 11200
rect 18012 11160 18018 11172
rect 18601 11169 18613 11172
rect 18647 11169 18659 11203
rect 18708 11200 18736 11240
rect 19420 11237 19432 11271
rect 19466 11268 19478 11271
rect 20622 11268 20628 11280
rect 19466 11240 20628 11268
rect 19466 11237 19478 11240
rect 19420 11231 19478 11237
rect 20622 11228 20628 11240
rect 20680 11228 20686 11280
rect 20162 11200 20168 11212
rect 18708 11172 20168 11200
rect 18601 11163 18659 11169
rect 20162 11160 20168 11172
rect 20220 11160 20226 11212
rect 17865 11135 17923 11141
rect 17865 11132 17877 11135
rect 17512 11104 17877 11132
rect 17865 11101 17877 11104
rect 17911 11132 17923 11135
rect 18782 11132 18788 11144
rect 17911 11104 18788 11132
rect 17911 11101 17923 11104
rect 17865 11095 17923 11101
rect 18782 11092 18788 11104
rect 18840 11092 18846 11144
rect 18874 11092 18880 11144
rect 18932 11132 18938 11144
rect 19153 11135 19211 11141
rect 19153 11132 19165 11135
rect 18932 11104 19165 11132
rect 18932 11092 18938 11104
rect 19153 11101 19165 11104
rect 19199 11101 19211 11135
rect 19153 11095 19211 11101
rect 16482 11064 16488 11076
rect 14108 11036 16488 11064
rect 16482 11024 16488 11036
rect 16540 11024 16546 11076
rect 21266 11064 21272 11076
rect 16960 11036 18552 11064
rect 7374 10996 7380 11008
rect 6748 10968 7380 10996
rect 2648 10956 2654 10968
rect 7374 10956 7380 10968
rect 7432 10956 7438 11008
rect 8294 10956 8300 11008
rect 8352 10996 8358 11008
rect 8478 10996 8484 11008
rect 8352 10968 8484 10996
rect 8352 10956 8358 10968
rect 8478 10956 8484 10968
rect 8536 10956 8542 11008
rect 10502 10956 10508 11008
rect 10560 10996 10566 11008
rect 11974 10996 11980 11008
rect 10560 10968 11980 10996
rect 10560 10956 10566 10968
rect 11974 10956 11980 10968
rect 12032 10956 12038 11008
rect 13906 10956 13912 11008
rect 13964 10996 13970 11008
rect 16960 10996 16988 11036
rect 18524 11008 18552 11036
rect 20088 11036 21272 11064
rect 17310 10996 17316 11008
rect 13964 10968 16988 10996
rect 17271 10968 17316 10996
rect 13964 10956 13970 10968
rect 17310 10956 17316 10968
rect 17368 10956 17374 11008
rect 18506 10956 18512 11008
rect 18564 10956 18570 11008
rect 18782 10956 18788 11008
rect 18840 10996 18846 11008
rect 20088 10996 20116 11036
rect 21266 11024 21272 11036
rect 21324 11024 21330 11076
rect 18840 10968 20116 10996
rect 18840 10956 18846 10968
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 1670 10792 1676 10804
rect 1631 10764 1676 10792
rect 1670 10752 1676 10764
rect 1728 10752 1734 10804
rect 2958 10752 2964 10804
rect 3016 10792 3022 10804
rect 4801 10795 4859 10801
rect 4801 10792 4813 10795
rect 3016 10764 4813 10792
rect 3016 10752 3022 10764
rect 4801 10761 4813 10764
rect 4847 10761 4859 10795
rect 4801 10755 4859 10761
rect 5994 10752 6000 10804
rect 6052 10792 6058 10804
rect 6546 10792 6552 10804
rect 6052 10764 6552 10792
rect 6052 10752 6058 10764
rect 6546 10752 6552 10764
rect 6604 10752 6610 10804
rect 6822 10752 6828 10804
rect 6880 10792 6886 10804
rect 11517 10795 11575 10801
rect 11517 10792 11529 10795
rect 6880 10764 11529 10792
rect 6880 10752 6886 10764
rect 11517 10761 11529 10764
rect 11563 10761 11575 10795
rect 11517 10755 11575 10761
rect 13170 10752 13176 10804
rect 13228 10792 13234 10804
rect 13909 10795 13967 10801
rect 13228 10764 13860 10792
rect 13228 10752 13234 10764
rect 3786 10684 3792 10736
rect 3844 10724 3850 10736
rect 5350 10724 5356 10736
rect 3844 10696 5356 10724
rect 3844 10684 3850 10696
rect 2314 10656 2320 10668
rect 2275 10628 2320 10656
rect 2314 10616 2320 10628
rect 2372 10616 2378 10668
rect 3418 10616 3424 10668
rect 3476 10656 3482 10668
rect 4264 10665 4292 10696
rect 5350 10684 5356 10696
rect 5408 10724 5414 10736
rect 9766 10724 9772 10736
rect 5408 10696 9772 10724
rect 5408 10684 5414 10696
rect 9766 10684 9772 10696
rect 9824 10684 9830 10736
rect 11241 10727 11299 10733
rect 11241 10693 11253 10727
rect 11287 10724 11299 10727
rect 11606 10724 11612 10736
rect 11287 10696 11612 10724
rect 11287 10693 11299 10696
rect 11241 10687 11299 10693
rect 11606 10684 11612 10696
rect 11664 10684 11670 10736
rect 13832 10724 13860 10764
rect 13909 10761 13921 10795
rect 13955 10792 13967 10795
rect 13955 10764 16160 10792
rect 13955 10761 13967 10764
rect 13909 10755 13967 10761
rect 14001 10727 14059 10733
rect 14001 10724 14013 10727
rect 13832 10696 14013 10724
rect 14001 10693 14013 10696
rect 14047 10693 14059 10727
rect 14001 10687 14059 10693
rect 14093 10727 14151 10733
rect 14093 10693 14105 10727
rect 14139 10724 14151 10727
rect 15194 10724 15200 10736
rect 14139 10696 15200 10724
rect 14139 10693 14151 10696
rect 14093 10687 14151 10693
rect 15194 10684 15200 10696
rect 15252 10684 15258 10736
rect 16132 10724 16160 10764
rect 16574 10752 16580 10804
rect 16632 10792 16638 10804
rect 16853 10795 16911 10801
rect 16853 10792 16865 10795
rect 16632 10764 16865 10792
rect 16632 10752 16638 10764
rect 16853 10761 16865 10764
rect 16899 10761 16911 10795
rect 16853 10755 16911 10761
rect 20622 10752 20628 10804
rect 20680 10792 20686 10804
rect 20901 10795 20959 10801
rect 20901 10792 20913 10795
rect 20680 10764 20913 10792
rect 20680 10752 20686 10764
rect 20901 10761 20913 10764
rect 20947 10761 20959 10795
rect 20901 10755 20959 10761
rect 17218 10724 17224 10736
rect 16132 10696 17224 10724
rect 17218 10684 17224 10696
rect 17276 10684 17282 10736
rect 4065 10659 4123 10665
rect 4065 10656 4077 10659
rect 3476 10628 4077 10656
rect 3476 10616 3482 10628
rect 4065 10625 4077 10628
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 4249 10659 4307 10665
rect 4249 10625 4261 10659
rect 4295 10625 4307 10659
rect 5442 10656 5448 10668
rect 5403 10628 5448 10656
rect 4249 10619 4307 10625
rect 5442 10616 5448 10628
rect 5500 10616 5506 10668
rect 5626 10616 5632 10668
rect 5684 10656 5690 10668
rect 5905 10659 5963 10665
rect 5905 10656 5917 10659
rect 5684 10628 5917 10656
rect 5684 10616 5690 10628
rect 5905 10625 5917 10628
rect 5951 10625 5963 10659
rect 5905 10619 5963 10625
rect 5994 10616 6000 10668
rect 6052 10656 6058 10668
rect 7466 10656 7472 10668
rect 6052 10628 7328 10656
rect 7427 10628 7472 10656
rect 6052 10616 6058 10628
rect 1486 10548 1492 10600
rect 1544 10588 1550 10600
rect 1544 10560 3556 10588
rect 1544 10548 1550 10560
rect 2314 10480 2320 10532
rect 2372 10520 2378 10532
rect 2590 10520 2596 10532
rect 2372 10492 2596 10520
rect 2372 10480 2378 10492
rect 2590 10480 2596 10492
rect 2648 10480 2654 10532
rect 3528 10529 3556 10560
rect 4890 10548 4896 10600
rect 4948 10588 4954 10600
rect 7193 10591 7251 10597
rect 7193 10588 7205 10591
rect 4948 10560 7205 10588
rect 4948 10548 4954 10560
rect 7193 10557 7205 10560
rect 7239 10557 7251 10591
rect 7300 10588 7328 10628
rect 7466 10616 7472 10628
rect 7524 10656 7530 10668
rect 8202 10656 8208 10668
rect 7524 10628 8208 10656
rect 7524 10616 7530 10628
rect 8202 10616 8208 10628
rect 8260 10656 8266 10668
rect 8389 10659 8447 10665
rect 8389 10656 8401 10659
rect 8260 10628 8401 10656
rect 8260 10616 8266 10628
rect 8389 10625 8401 10628
rect 8435 10656 8447 10659
rect 9401 10659 9459 10665
rect 9401 10656 9413 10659
rect 8435 10628 9413 10656
rect 8435 10625 8447 10628
rect 8389 10619 8447 10625
rect 9401 10625 9413 10628
rect 9447 10625 9459 10659
rect 9401 10619 9459 10625
rect 11790 10616 11796 10668
rect 11848 10656 11854 10668
rect 12069 10659 12127 10665
rect 12069 10656 12081 10659
rect 11848 10628 12081 10656
rect 11848 10616 11854 10628
rect 12069 10625 12081 10628
rect 12115 10625 12127 10659
rect 12069 10619 12127 10625
rect 13722 10616 13728 10668
rect 13780 10656 13786 10668
rect 14274 10656 14280 10668
rect 13780 10628 14280 10656
rect 13780 10616 13786 10628
rect 14274 10616 14280 10628
rect 14332 10656 14338 10668
rect 14645 10659 14703 10665
rect 14645 10656 14657 10659
rect 14332 10628 14657 10656
rect 14332 10616 14338 10628
rect 14645 10625 14657 10628
rect 14691 10625 14703 10659
rect 17402 10656 17408 10668
rect 17363 10628 17408 10656
rect 14645 10619 14703 10625
rect 17402 10616 17408 10628
rect 17460 10616 17466 10668
rect 17862 10616 17868 10668
rect 17920 10616 17926 10668
rect 18506 10616 18512 10668
rect 18564 10656 18570 10668
rect 18601 10659 18659 10665
rect 18601 10656 18613 10659
rect 18564 10628 18613 10656
rect 18564 10616 18570 10628
rect 18601 10625 18613 10628
rect 18647 10625 18659 10659
rect 18601 10619 18659 10625
rect 8110 10588 8116 10600
rect 7300 10560 8116 10588
rect 7193 10551 7251 10557
rect 8110 10548 8116 10560
rect 8168 10548 8174 10600
rect 8297 10591 8355 10597
rect 8297 10557 8309 10591
rect 8343 10588 8355 10591
rect 9122 10588 9128 10600
rect 8343 10560 9128 10588
rect 8343 10557 8355 10560
rect 8297 10551 8355 10557
rect 9122 10548 9128 10560
rect 9180 10548 9186 10600
rect 9217 10591 9275 10597
rect 9217 10557 9229 10591
rect 9263 10588 9275 10591
rect 9306 10588 9312 10600
rect 9263 10560 9312 10588
rect 9263 10557 9275 10560
rect 9217 10551 9275 10557
rect 9306 10548 9312 10560
rect 9364 10548 9370 10600
rect 9674 10548 9680 10600
rect 9732 10588 9738 10600
rect 9861 10591 9919 10597
rect 9861 10588 9873 10591
rect 9732 10560 9873 10588
rect 9732 10548 9738 10560
rect 9861 10557 9873 10560
rect 9907 10557 9919 10591
rect 12250 10588 12256 10600
rect 9861 10551 9919 10557
rect 10060 10560 12256 10588
rect 3513 10523 3571 10529
rect 3513 10489 3525 10523
rect 3559 10520 3571 10523
rect 5261 10523 5319 10529
rect 3559 10492 4016 10520
rect 3559 10489 3571 10492
rect 3513 10483 3571 10489
rect 3988 10464 4016 10492
rect 5261 10489 5273 10523
rect 5307 10520 5319 10523
rect 6730 10520 6736 10532
rect 5307 10492 6736 10520
rect 5307 10489 5319 10492
rect 5261 10483 5319 10489
rect 6730 10480 6736 10492
rect 6788 10480 6794 10532
rect 7285 10523 7343 10529
rect 7285 10489 7297 10523
rect 7331 10520 7343 10523
rect 10060 10520 10088 10560
rect 12250 10548 12256 10560
rect 12308 10548 12314 10600
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 12704 10591 12762 10597
rect 12492 10560 12537 10588
rect 12492 10548 12498 10560
rect 12704 10557 12716 10591
rect 12750 10588 12762 10591
rect 12986 10588 12992 10600
rect 12750 10560 12992 10588
rect 12750 10557 12762 10560
rect 12704 10551 12762 10557
rect 12986 10548 12992 10560
rect 13044 10548 13050 10600
rect 13170 10548 13176 10600
rect 13228 10588 13234 10600
rect 13909 10591 13967 10597
rect 13909 10588 13921 10591
rect 13228 10560 13921 10588
rect 13228 10548 13234 10560
rect 13909 10557 13921 10560
rect 13955 10557 13967 10591
rect 13909 10551 13967 10557
rect 14001 10591 14059 10597
rect 14001 10557 14013 10591
rect 14047 10588 14059 10591
rect 14461 10591 14519 10597
rect 14461 10588 14473 10591
rect 14047 10560 14473 10588
rect 14047 10557 14059 10560
rect 14001 10551 14059 10557
rect 14461 10557 14473 10560
rect 14507 10588 14519 10591
rect 15010 10588 15016 10600
rect 14507 10560 15016 10588
rect 14507 10557 14519 10560
rect 14461 10551 14519 10557
rect 15010 10548 15016 10560
rect 15068 10548 15074 10600
rect 15197 10591 15255 10597
rect 15197 10557 15209 10591
rect 15243 10588 15255 10591
rect 15286 10588 15292 10600
rect 15243 10560 15292 10588
rect 15243 10557 15255 10560
rect 15197 10551 15255 10557
rect 15286 10548 15292 10560
rect 15344 10548 15350 10600
rect 15464 10591 15522 10597
rect 15464 10557 15476 10591
rect 15510 10588 15522 10591
rect 15930 10588 15936 10600
rect 15510 10560 15936 10588
rect 15510 10557 15522 10560
rect 15464 10551 15522 10557
rect 15930 10548 15936 10560
rect 15988 10548 15994 10600
rect 16574 10548 16580 10600
rect 16632 10588 16638 10600
rect 16850 10588 16856 10600
rect 16632 10560 16856 10588
rect 16632 10548 16638 10560
rect 16850 10548 16856 10560
rect 16908 10548 16914 10600
rect 17313 10591 17371 10597
rect 17313 10557 17325 10591
rect 17359 10588 17371 10591
rect 17880 10588 17908 10616
rect 18322 10588 18328 10600
rect 17359 10560 18328 10588
rect 17359 10557 17371 10560
rect 17313 10551 17371 10557
rect 18322 10548 18328 10560
rect 18380 10548 18386 10600
rect 18417 10591 18475 10597
rect 18417 10557 18429 10591
rect 18463 10588 18475 10591
rect 18690 10588 18696 10600
rect 18463 10560 18696 10588
rect 18463 10557 18475 10560
rect 18417 10551 18475 10557
rect 18690 10548 18696 10560
rect 18748 10548 18754 10600
rect 18874 10548 18880 10600
rect 18932 10588 18938 10600
rect 19521 10591 19579 10597
rect 19521 10588 19533 10591
rect 18932 10560 19533 10588
rect 18932 10548 18938 10560
rect 19521 10557 19533 10560
rect 19567 10557 19579 10591
rect 19521 10551 19579 10557
rect 7331 10492 10088 10520
rect 10128 10523 10186 10529
rect 7331 10489 7343 10492
rect 7285 10483 7343 10489
rect 10128 10489 10140 10523
rect 10174 10520 10186 10523
rect 10962 10520 10968 10532
rect 10174 10492 10968 10520
rect 10174 10489 10186 10492
rect 10128 10483 10186 10489
rect 10962 10480 10968 10492
rect 11020 10480 11026 10532
rect 11790 10480 11796 10532
rect 11848 10520 11854 10532
rect 12158 10520 12164 10532
rect 11848 10492 12164 10520
rect 11848 10480 11854 10492
rect 12158 10480 12164 10492
rect 12216 10480 12222 10532
rect 13354 10480 13360 10532
rect 13412 10520 13418 10532
rect 13722 10520 13728 10532
rect 13412 10492 13728 10520
rect 13412 10480 13418 10492
rect 13722 10480 13728 10492
rect 13780 10480 13786 10532
rect 17862 10520 17868 10532
rect 13832 10492 17868 10520
rect 1762 10412 1768 10464
rect 1820 10452 1826 10464
rect 2041 10455 2099 10461
rect 2041 10452 2053 10455
rect 1820 10424 2053 10452
rect 1820 10412 1826 10424
rect 2041 10421 2053 10424
rect 2087 10421 2099 10455
rect 2041 10415 2099 10421
rect 2130 10412 2136 10464
rect 2188 10452 2194 10464
rect 3602 10452 3608 10464
rect 2188 10424 2233 10452
rect 3563 10424 3608 10452
rect 2188 10412 2194 10424
rect 3602 10412 3608 10424
rect 3660 10412 3666 10464
rect 3970 10452 3976 10464
rect 3931 10424 3976 10452
rect 3970 10412 3976 10424
rect 4028 10412 4034 10464
rect 5166 10452 5172 10464
rect 5127 10424 5172 10452
rect 5166 10412 5172 10424
rect 5224 10412 5230 10464
rect 6178 10412 6184 10464
rect 6236 10452 6242 10464
rect 6825 10455 6883 10461
rect 6825 10452 6837 10455
rect 6236 10424 6837 10452
rect 6236 10412 6242 10424
rect 6825 10421 6837 10424
rect 6871 10421 6883 10455
rect 6825 10415 6883 10421
rect 7374 10412 7380 10464
rect 7432 10452 7438 10464
rect 7837 10455 7895 10461
rect 7837 10452 7849 10455
rect 7432 10424 7849 10452
rect 7432 10412 7438 10424
rect 7837 10421 7849 10424
rect 7883 10421 7895 10455
rect 7837 10415 7895 10421
rect 8205 10455 8263 10461
rect 8205 10421 8217 10455
rect 8251 10452 8263 10455
rect 8662 10452 8668 10464
rect 8251 10424 8668 10452
rect 8251 10421 8263 10424
rect 8205 10415 8263 10421
rect 8662 10412 8668 10424
rect 8720 10412 8726 10464
rect 8846 10452 8852 10464
rect 8807 10424 8852 10452
rect 8846 10412 8852 10424
rect 8904 10412 8910 10464
rect 9214 10412 9220 10464
rect 9272 10452 9278 10464
rect 9309 10455 9367 10461
rect 9309 10452 9321 10455
rect 9272 10424 9321 10452
rect 9272 10412 9278 10424
rect 9309 10421 9321 10424
rect 9355 10421 9367 10455
rect 9309 10415 9367 10421
rect 9582 10412 9588 10464
rect 9640 10452 9646 10464
rect 11885 10455 11943 10461
rect 11885 10452 11897 10455
rect 9640 10424 11897 10452
rect 9640 10412 9646 10424
rect 11885 10421 11897 10424
rect 11931 10421 11943 10455
rect 11885 10415 11943 10421
rect 11977 10455 12035 10461
rect 11977 10421 11989 10455
rect 12023 10452 12035 10455
rect 12710 10452 12716 10464
rect 12023 10424 12716 10452
rect 12023 10421 12035 10424
rect 11977 10415 12035 10421
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 12986 10412 12992 10464
rect 13044 10452 13050 10464
rect 13832 10461 13860 10492
rect 17862 10480 17868 10492
rect 17920 10480 17926 10532
rect 19788 10523 19846 10529
rect 19788 10489 19800 10523
rect 19834 10520 19846 10523
rect 20438 10520 20444 10532
rect 19834 10492 20444 10520
rect 19834 10489 19846 10492
rect 19788 10483 19846 10489
rect 20438 10480 20444 10492
rect 20496 10480 20502 10532
rect 13817 10455 13875 10461
rect 13817 10452 13829 10455
rect 13044 10424 13829 10452
rect 13044 10412 13050 10424
rect 13817 10421 13829 10424
rect 13863 10421 13875 10455
rect 13817 10415 13875 10421
rect 14182 10412 14188 10464
rect 14240 10452 14246 10464
rect 14553 10455 14611 10461
rect 14553 10452 14565 10455
rect 14240 10424 14565 10452
rect 14240 10412 14246 10424
rect 14553 10421 14565 10424
rect 14599 10421 14611 10455
rect 14553 10415 14611 10421
rect 15194 10412 15200 10464
rect 15252 10452 15258 10464
rect 16482 10452 16488 10464
rect 15252 10424 16488 10452
rect 15252 10412 15258 10424
rect 16482 10412 16488 10424
rect 16540 10412 16546 10464
rect 16577 10455 16635 10461
rect 16577 10421 16589 10455
rect 16623 10452 16635 10455
rect 16850 10452 16856 10464
rect 16623 10424 16856 10452
rect 16623 10421 16635 10424
rect 16577 10415 16635 10421
rect 16850 10412 16856 10424
rect 16908 10412 16914 10464
rect 17218 10452 17224 10464
rect 17179 10424 17224 10452
rect 17218 10412 17224 10424
rect 17276 10412 17282 10464
rect 17678 10412 17684 10464
rect 17736 10452 17742 10464
rect 18049 10455 18107 10461
rect 18049 10452 18061 10455
rect 17736 10424 18061 10452
rect 17736 10412 17742 10424
rect 18049 10421 18061 10424
rect 18095 10421 18107 10455
rect 18049 10415 18107 10421
rect 18509 10455 18567 10461
rect 18509 10421 18521 10455
rect 18555 10452 18567 10455
rect 18966 10452 18972 10464
rect 18555 10424 18972 10452
rect 18555 10421 18567 10424
rect 18509 10415 18567 10421
rect 18966 10412 18972 10424
rect 19024 10412 19030 10464
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 1762 10248 1768 10260
rect 1723 10220 1768 10248
rect 1762 10208 1768 10220
rect 1820 10208 1826 10260
rect 1854 10208 1860 10260
rect 1912 10248 1918 10260
rect 2225 10251 2283 10257
rect 2225 10248 2237 10251
rect 1912 10220 2237 10248
rect 1912 10208 1918 10220
rect 2225 10217 2237 10220
rect 2271 10217 2283 10251
rect 2225 10211 2283 10217
rect 2961 10251 3019 10257
rect 2961 10217 2973 10251
rect 3007 10248 3019 10251
rect 3050 10248 3056 10260
rect 3007 10220 3056 10248
rect 3007 10217 3019 10220
rect 2961 10211 3019 10217
rect 3050 10208 3056 10220
rect 3108 10208 3114 10260
rect 3329 10251 3387 10257
rect 3329 10217 3341 10251
rect 3375 10248 3387 10251
rect 3602 10248 3608 10260
rect 3375 10220 3608 10248
rect 3375 10217 3387 10220
rect 3329 10211 3387 10217
rect 3602 10208 3608 10220
rect 3660 10208 3666 10260
rect 5166 10208 5172 10260
rect 5224 10248 5230 10260
rect 5721 10251 5779 10257
rect 5721 10248 5733 10251
rect 5224 10220 5733 10248
rect 5224 10208 5230 10220
rect 5721 10217 5733 10220
rect 5767 10217 5779 10251
rect 5994 10248 6000 10260
rect 5721 10211 5779 10217
rect 5920 10220 6000 10248
rect 3421 10183 3479 10189
rect 3421 10149 3433 10183
rect 3467 10180 3479 10183
rect 3510 10180 3516 10192
rect 3467 10152 3516 10180
rect 3467 10149 3479 10152
rect 3421 10143 3479 10149
rect 3510 10140 3516 10152
rect 3568 10140 3574 10192
rect 5920 10180 5948 10220
rect 5994 10208 6000 10220
rect 6052 10208 6058 10260
rect 6178 10248 6184 10260
rect 6139 10220 6184 10248
rect 6178 10208 6184 10220
rect 6236 10208 6242 10260
rect 6288 10220 7779 10248
rect 6086 10180 6092 10192
rect 4264 10152 5948 10180
rect 6047 10152 6092 10180
rect 2133 10115 2191 10121
rect 2133 10081 2145 10115
rect 2179 10112 2191 10115
rect 2866 10112 2872 10124
rect 2179 10084 2872 10112
rect 2179 10081 2191 10084
rect 2133 10075 2191 10081
rect 2866 10072 2872 10084
rect 2924 10072 2930 10124
rect 3878 10072 3884 10124
rect 3936 10112 3942 10124
rect 4264 10112 4292 10152
rect 6086 10140 6092 10152
rect 6144 10140 6150 10192
rect 3936 10084 4292 10112
rect 4332 10115 4390 10121
rect 3936 10072 3942 10084
rect 4332 10081 4344 10115
rect 4378 10112 4390 10115
rect 5074 10112 5080 10124
rect 4378 10084 5080 10112
rect 4378 10081 4390 10084
rect 4332 10075 4390 10081
rect 5074 10072 5080 10084
rect 5132 10112 5138 10124
rect 6288 10112 6316 10220
rect 6638 10140 6644 10192
rect 6696 10180 6702 10192
rect 7098 10180 7104 10192
rect 6696 10152 7104 10180
rect 6696 10140 6702 10152
rect 7098 10140 7104 10152
rect 7156 10140 7162 10192
rect 7650 10189 7656 10192
rect 7644 10180 7656 10189
rect 7611 10152 7656 10180
rect 7644 10143 7656 10152
rect 7650 10140 7656 10143
rect 7708 10140 7714 10192
rect 7751 10180 7779 10220
rect 8202 10208 8208 10260
rect 8260 10248 8266 10260
rect 8757 10251 8815 10257
rect 8757 10248 8769 10251
rect 8260 10220 8769 10248
rect 8260 10208 8266 10220
rect 8757 10217 8769 10220
rect 8803 10217 8815 10251
rect 8757 10211 8815 10217
rect 10962 10208 10968 10260
rect 11020 10248 11026 10260
rect 11057 10251 11115 10257
rect 11057 10248 11069 10251
rect 11020 10220 11069 10248
rect 11020 10208 11026 10220
rect 11057 10217 11069 10220
rect 11103 10217 11115 10251
rect 11057 10211 11115 10217
rect 11146 10208 11152 10260
rect 11204 10248 11210 10260
rect 12345 10251 12403 10257
rect 12345 10248 12357 10251
rect 11204 10220 12357 10248
rect 11204 10208 11210 10220
rect 12345 10217 12357 10220
rect 12391 10217 12403 10251
rect 12345 10211 12403 10217
rect 12802 10208 12808 10260
rect 12860 10248 12866 10260
rect 16669 10251 16727 10257
rect 16669 10248 16681 10251
rect 12860 10220 16681 10248
rect 12860 10208 12866 10220
rect 16669 10217 16681 10220
rect 16715 10217 16727 10251
rect 17678 10248 17684 10260
rect 17639 10220 17684 10248
rect 16669 10211 16727 10217
rect 17678 10208 17684 10220
rect 17736 10208 17742 10260
rect 18601 10251 18659 10257
rect 18601 10217 18613 10251
rect 18647 10217 18659 10251
rect 18601 10211 18659 10217
rect 7751 10152 11836 10180
rect 7282 10112 7288 10124
rect 5132 10084 6316 10112
rect 7243 10084 7288 10112
rect 5132 10072 5138 10084
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 7377 10115 7435 10121
rect 7377 10081 7389 10115
rect 7423 10112 7435 10115
rect 8202 10112 8208 10124
rect 7423 10084 8208 10112
rect 7423 10081 7435 10084
rect 7377 10075 7435 10081
rect 8202 10072 8208 10084
rect 8260 10112 8266 10124
rect 9674 10112 9680 10124
rect 8260 10084 9680 10112
rect 8260 10072 8266 10084
rect 9674 10072 9680 10084
rect 9732 10072 9738 10124
rect 9944 10115 10002 10121
rect 9944 10081 9956 10115
rect 9990 10112 10002 10115
rect 10502 10112 10508 10124
rect 9990 10084 10508 10112
rect 9990 10081 10002 10084
rect 9944 10075 10002 10081
rect 10502 10072 10508 10084
rect 10560 10072 10566 10124
rect 10778 10072 10784 10124
rect 10836 10112 10842 10124
rect 11701 10115 11759 10121
rect 11701 10112 11713 10115
rect 10836 10084 11713 10112
rect 10836 10072 10842 10084
rect 11701 10081 11713 10084
rect 11747 10081 11759 10115
rect 11808 10112 11836 10152
rect 11974 10140 11980 10192
rect 12032 10180 12038 10192
rect 12713 10183 12771 10189
rect 12713 10180 12725 10183
rect 12032 10152 12725 10180
rect 12032 10140 12038 10152
rect 12713 10149 12725 10152
rect 12759 10180 12771 10183
rect 13630 10180 13636 10192
rect 12759 10152 13636 10180
rect 12759 10149 12771 10152
rect 12713 10143 12771 10149
rect 13630 10140 13636 10152
rect 13688 10140 13694 10192
rect 13817 10183 13875 10189
rect 13817 10149 13829 10183
rect 13863 10180 13875 10183
rect 15194 10180 15200 10192
rect 13863 10152 15200 10180
rect 13863 10149 13875 10152
rect 13817 10143 13875 10149
rect 15194 10140 15200 10152
rect 15252 10140 15258 10192
rect 18616 10180 18644 10211
rect 19794 10208 19800 10260
rect 19852 10248 19858 10260
rect 20070 10248 20076 10260
rect 19852 10220 20076 10248
rect 19852 10208 19858 10220
rect 20070 10208 20076 10220
rect 20128 10208 20134 10260
rect 20349 10251 20407 10257
rect 20349 10217 20361 10251
rect 20395 10248 20407 10251
rect 20438 10248 20444 10260
rect 20395 10220 20444 10248
rect 20395 10217 20407 10220
rect 20349 10211 20407 10217
rect 20438 10208 20444 10220
rect 20496 10208 20502 10260
rect 22462 10180 22468 10192
rect 15580 10152 15792 10180
rect 13725 10115 13783 10121
rect 11808 10084 13032 10112
rect 11701 10075 11759 10081
rect 2409 10047 2467 10053
rect 2409 10013 2421 10047
rect 2455 10044 2467 10047
rect 3602 10044 3608 10056
rect 2455 10016 2636 10044
rect 3563 10016 3608 10044
rect 2455 10013 2467 10016
rect 2409 10007 2467 10013
rect 2608 9908 2636 10016
rect 3602 10004 3608 10016
rect 3660 10004 3666 10056
rect 4062 10044 4068 10056
rect 4023 10016 4068 10044
rect 4062 10004 4068 10016
rect 4120 10004 4126 10056
rect 6178 10004 6184 10056
rect 6236 10044 6242 10056
rect 6273 10047 6331 10053
rect 6273 10044 6285 10047
rect 6236 10016 6285 10044
rect 6236 10004 6242 10016
rect 6273 10013 6285 10016
rect 6319 10013 6331 10047
rect 6273 10007 6331 10013
rect 11054 10004 11060 10056
rect 11112 10044 11118 10056
rect 11793 10047 11851 10053
rect 11793 10044 11805 10047
rect 11112 10016 11805 10044
rect 11112 10004 11118 10016
rect 11793 10013 11805 10016
rect 11839 10013 11851 10047
rect 11974 10044 11980 10056
rect 11935 10016 11980 10044
rect 11793 10007 11851 10013
rect 11974 10004 11980 10016
rect 12032 10004 12038 10056
rect 12802 10044 12808 10056
rect 12763 10016 12808 10044
rect 12802 10004 12808 10016
rect 12860 10004 12866 10056
rect 13004 10053 13032 10084
rect 13725 10081 13737 10115
rect 13771 10112 13783 10115
rect 14550 10112 14556 10124
rect 13771 10084 14320 10112
rect 14511 10084 14556 10112
rect 13771 10081 13783 10084
rect 13725 10075 13783 10081
rect 12989 10047 13047 10053
rect 12989 10013 13001 10047
rect 13035 10013 13047 10047
rect 12989 10007 13047 10013
rect 13909 10047 13967 10053
rect 13909 10013 13921 10047
rect 13955 10013 13967 10047
rect 13909 10007 13967 10013
rect 2774 9908 2780 9920
rect 2608 9880 2780 9908
rect 2774 9868 2780 9880
rect 2832 9908 2838 9920
rect 3620 9908 3648 10004
rect 5350 9936 5356 9988
rect 5408 9976 5414 9988
rect 5445 9979 5503 9985
rect 5445 9976 5457 9979
rect 5408 9948 5457 9976
rect 5408 9936 5414 9948
rect 5445 9945 5457 9948
rect 5491 9945 5503 9979
rect 7282 9976 7288 9988
rect 5445 9939 5503 9945
rect 5552 9948 7288 9976
rect 2832 9880 3648 9908
rect 2832 9868 2838 9880
rect 3970 9868 3976 9920
rect 4028 9908 4034 9920
rect 5552 9908 5580 9948
rect 7282 9936 7288 9948
rect 7340 9936 7346 9988
rect 8662 9936 8668 9988
rect 8720 9976 8726 9988
rect 9674 9976 9680 9988
rect 8720 9948 9680 9976
rect 8720 9936 8726 9948
rect 9674 9936 9680 9948
rect 9732 9936 9738 9988
rect 11698 9936 11704 9988
rect 11756 9976 11762 9988
rect 12158 9976 12164 9988
rect 11756 9948 12164 9976
rect 11756 9936 11762 9948
rect 12158 9936 12164 9948
rect 12216 9976 12222 9988
rect 13924 9976 13952 10007
rect 12216 9948 13952 9976
rect 12216 9936 12222 9948
rect 4028 9880 5580 9908
rect 4028 9868 4034 9880
rect 6914 9868 6920 9920
rect 6972 9908 6978 9920
rect 7101 9911 7159 9917
rect 7101 9908 7113 9911
rect 6972 9880 7113 9908
rect 6972 9868 6978 9880
rect 7101 9877 7113 9880
rect 7147 9877 7159 9911
rect 7101 9871 7159 9877
rect 7190 9868 7196 9920
rect 7248 9908 7254 9920
rect 10870 9908 10876 9920
rect 7248 9880 10876 9908
rect 7248 9868 7254 9880
rect 10870 9868 10876 9880
rect 10928 9868 10934 9920
rect 11054 9868 11060 9920
rect 11112 9908 11118 9920
rect 11333 9911 11391 9917
rect 11333 9908 11345 9911
rect 11112 9880 11345 9908
rect 11112 9868 11118 9880
rect 11333 9877 11345 9880
rect 11379 9877 11391 9911
rect 13354 9908 13360 9920
rect 13315 9880 13360 9908
rect 11333 9871 11391 9877
rect 13354 9868 13360 9880
rect 13412 9868 13418 9920
rect 14292 9908 14320 10084
rect 14550 10072 14556 10084
rect 14608 10072 14614 10124
rect 15013 10115 15071 10121
rect 15013 10081 15025 10115
rect 15059 10081 15071 10115
rect 15013 10075 15071 10081
rect 14458 10044 14464 10056
rect 14384 10016 14464 10044
rect 14384 9985 14412 10016
rect 14458 10004 14464 10016
rect 14516 10044 14522 10056
rect 15028 10044 15056 10075
rect 15286 10072 15292 10124
rect 15344 10112 15350 10124
rect 15580 10112 15608 10152
rect 15344 10084 15608 10112
rect 15657 10115 15715 10121
rect 15344 10072 15350 10084
rect 15657 10081 15669 10115
rect 15703 10081 15715 10115
rect 15764 10112 15792 10152
rect 17696 10152 18552 10180
rect 18616 10152 22468 10180
rect 17696 10124 17724 10152
rect 17678 10112 17684 10124
rect 15764 10084 17684 10112
rect 15657 10075 15715 10081
rect 14516 10016 15056 10044
rect 14516 10004 14522 10016
rect 15562 10004 15568 10056
rect 15620 10044 15626 10056
rect 15672 10044 15700 10075
rect 17678 10072 17684 10084
rect 17736 10072 17742 10124
rect 17773 10115 17831 10121
rect 17773 10081 17785 10115
rect 17819 10112 17831 10115
rect 17954 10112 17960 10124
rect 17819 10084 17960 10112
rect 17819 10081 17831 10084
rect 17773 10075 17831 10081
rect 17954 10072 17960 10084
rect 18012 10072 18018 10124
rect 18414 10112 18420 10124
rect 18375 10084 18420 10112
rect 18414 10072 18420 10084
rect 18472 10072 18478 10124
rect 18524 10112 18552 10152
rect 22462 10140 22468 10152
rect 22520 10140 22526 10192
rect 18874 10112 18880 10124
rect 18524 10084 18880 10112
rect 18874 10072 18880 10084
rect 18932 10112 18938 10124
rect 18969 10115 19027 10121
rect 18969 10112 18981 10115
rect 18932 10084 18981 10112
rect 18932 10072 18938 10084
rect 18969 10081 18981 10084
rect 19015 10081 19027 10115
rect 18969 10075 19027 10081
rect 19236 10115 19294 10121
rect 19236 10081 19248 10115
rect 19282 10112 19294 10115
rect 19518 10112 19524 10124
rect 19282 10084 19524 10112
rect 19282 10081 19294 10084
rect 19236 10075 19294 10081
rect 19518 10072 19524 10084
rect 19576 10072 19582 10124
rect 15620 10016 15700 10044
rect 15749 10047 15807 10053
rect 15620 10004 15626 10016
rect 15749 10013 15761 10047
rect 15795 10044 15807 10047
rect 15838 10044 15844 10056
rect 15795 10016 15844 10044
rect 15795 10013 15807 10016
rect 15749 10007 15807 10013
rect 15838 10004 15844 10016
rect 15896 10004 15902 10056
rect 15933 10047 15991 10053
rect 15933 10013 15945 10047
rect 15979 10044 15991 10047
rect 16022 10044 16028 10056
rect 15979 10016 16028 10044
rect 15979 10013 15991 10016
rect 15933 10007 15991 10013
rect 16022 10004 16028 10016
rect 16080 10004 16086 10056
rect 16758 10044 16764 10056
rect 16719 10016 16764 10044
rect 16758 10004 16764 10016
rect 16816 10004 16822 10056
rect 16850 10004 16856 10056
rect 16908 10044 16914 10056
rect 17862 10044 17868 10056
rect 16908 10016 16953 10044
rect 17823 10016 17868 10044
rect 16908 10004 16914 10016
rect 17862 10004 17868 10016
rect 17920 10004 17926 10056
rect 18322 10004 18328 10056
rect 18380 10044 18386 10056
rect 18690 10044 18696 10056
rect 18380 10016 18696 10044
rect 18380 10004 18386 10016
rect 18690 10004 18696 10016
rect 18748 10004 18754 10056
rect 14369 9979 14427 9985
rect 14369 9945 14381 9979
rect 14415 9945 14427 9979
rect 15289 9979 15347 9985
rect 14369 9939 14427 9945
rect 14476 9948 15240 9976
rect 14476 9908 14504 9948
rect 14292 9880 14504 9908
rect 14550 9868 14556 9920
rect 14608 9908 14614 9920
rect 14829 9911 14887 9917
rect 14829 9908 14841 9911
rect 14608 9880 14841 9908
rect 14608 9868 14614 9880
rect 14829 9877 14841 9880
rect 14875 9877 14887 9911
rect 15212 9908 15240 9948
rect 15289 9945 15301 9979
rect 15335 9976 15347 9979
rect 16114 9976 16120 9988
rect 15335 9948 16120 9976
rect 15335 9945 15347 9948
rect 15289 9939 15347 9945
rect 16114 9936 16120 9948
rect 16172 9936 16178 9988
rect 16224 9948 17439 9976
rect 16224 9908 16252 9948
rect 15212 9880 16252 9908
rect 16301 9911 16359 9917
rect 14829 9871 14887 9877
rect 16301 9877 16313 9911
rect 16347 9908 16359 9911
rect 16758 9908 16764 9920
rect 16347 9880 16764 9908
rect 16347 9877 16359 9880
rect 16301 9871 16359 9877
rect 16758 9868 16764 9880
rect 16816 9868 16822 9920
rect 17034 9868 17040 9920
rect 17092 9908 17098 9920
rect 17313 9911 17371 9917
rect 17313 9908 17325 9911
rect 17092 9880 17325 9908
rect 17092 9868 17098 9880
rect 17313 9877 17325 9880
rect 17359 9877 17371 9911
rect 17411 9908 17439 9948
rect 19334 9908 19340 9920
rect 17411 9880 19340 9908
rect 17313 9871 17371 9877
rect 19334 9868 19340 9880
rect 19392 9868 19398 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 1857 9707 1915 9713
rect 1857 9673 1869 9707
rect 1903 9704 1915 9707
rect 2130 9704 2136 9716
rect 1903 9676 2136 9704
rect 1903 9673 1915 9676
rect 1857 9667 1915 9673
rect 2130 9664 2136 9676
rect 2188 9664 2194 9716
rect 2866 9704 2872 9716
rect 2827 9676 2872 9704
rect 2866 9664 2872 9676
rect 2924 9664 2930 9716
rect 7190 9664 7196 9716
rect 7248 9704 7254 9716
rect 8294 9704 8300 9716
rect 7248 9676 8300 9704
rect 7248 9664 7254 9676
rect 8294 9664 8300 9676
rect 8352 9704 8358 9716
rect 13170 9704 13176 9716
rect 8352 9676 10364 9704
rect 8352 9664 8358 9676
rect 5350 9596 5356 9648
rect 5408 9636 5414 9648
rect 5408 9608 6868 9636
rect 5408 9596 5414 9608
rect 2038 9528 2044 9580
rect 2096 9568 2102 9580
rect 2317 9571 2375 9577
rect 2317 9568 2329 9571
rect 2096 9540 2329 9568
rect 2096 9528 2102 9540
rect 2317 9537 2329 9540
rect 2363 9537 2375 9571
rect 2317 9531 2375 9537
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 2774 9568 2780 9580
rect 2547 9540 2780 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 2774 9528 2780 9540
rect 2832 9528 2838 9580
rect 3513 9571 3571 9577
rect 3513 9537 3525 9571
rect 3559 9568 3571 9571
rect 3786 9568 3792 9580
rect 3559 9540 3792 9568
rect 3559 9537 3571 9540
rect 3513 9531 3571 9537
rect 3786 9528 3792 9540
rect 3844 9528 3850 9580
rect 5810 9528 5816 9580
rect 5868 9568 5874 9580
rect 5905 9571 5963 9577
rect 5905 9568 5917 9571
rect 5868 9540 5917 9568
rect 5868 9528 5874 9540
rect 5905 9537 5917 9540
rect 5951 9537 5963 9571
rect 6840 9568 6868 9608
rect 10336 9568 10364 9676
rect 12268 9676 13176 9704
rect 10502 9636 10508 9648
rect 10463 9608 10508 9636
rect 10502 9596 10508 9608
rect 10560 9596 10566 9648
rect 12268 9636 12296 9676
rect 13170 9664 13176 9676
rect 13228 9664 13234 9716
rect 14182 9664 14188 9716
rect 14240 9704 14246 9716
rect 15286 9704 15292 9716
rect 14240 9676 15292 9704
rect 14240 9664 14246 9676
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 15562 9664 15568 9716
rect 15620 9664 15626 9716
rect 15838 9664 15844 9716
rect 15896 9704 15902 9716
rect 16301 9707 16359 9713
rect 16301 9704 16313 9707
rect 15896 9676 16313 9704
rect 15896 9664 15902 9676
rect 16301 9673 16313 9676
rect 16347 9673 16359 9707
rect 16301 9667 16359 9673
rect 10612 9608 12296 9636
rect 15580 9636 15608 9664
rect 16206 9636 16212 9648
rect 15580 9608 16212 9636
rect 10612 9568 10640 9608
rect 16206 9596 16212 9608
rect 16264 9596 16270 9648
rect 19242 9596 19248 9648
rect 19300 9636 19306 9648
rect 20901 9639 20959 9645
rect 20901 9636 20913 9639
rect 19300 9608 20913 9636
rect 19300 9596 19306 9608
rect 20901 9605 20913 9608
rect 20947 9605 20959 9639
rect 20901 9599 20959 9605
rect 6840 9540 6960 9568
rect 10336 9540 10640 9568
rect 5905 9531 5963 9537
rect 2222 9500 2228 9512
rect 2183 9472 2228 9500
rect 2222 9460 2228 9472
rect 2280 9460 2286 9512
rect 3694 9460 3700 9512
rect 3752 9500 3758 9512
rect 4062 9500 4068 9512
rect 3752 9472 4068 9500
rect 3752 9460 3758 9472
rect 4062 9460 4068 9472
rect 4120 9500 4126 9512
rect 4249 9503 4307 9509
rect 4249 9500 4261 9503
rect 4120 9472 4261 9500
rect 4120 9460 4126 9472
rect 4249 9469 4261 9472
rect 4295 9469 4307 9503
rect 4249 9463 4307 9469
rect 4516 9503 4574 9509
rect 4516 9469 4528 9503
rect 4562 9500 4574 9503
rect 6178 9500 6184 9512
rect 4562 9472 6184 9500
rect 4562 9469 4574 9472
rect 4516 9463 4574 9469
rect 6178 9460 6184 9472
rect 6236 9460 6242 9512
rect 6822 9500 6828 9512
rect 6783 9472 6828 9500
rect 6822 9460 6828 9472
rect 6880 9460 6886 9512
rect 1397 9435 1455 9441
rect 1397 9401 1409 9435
rect 1443 9432 1455 9435
rect 3237 9435 3295 9441
rect 3237 9432 3249 9435
rect 1443 9404 3249 9432
rect 1443 9401 1455 9404
rect 1397 9395 1455 9401
rect 3237 9401 3249 9404
rect 3283 9401 3295 9435
rect 6932 9432 6960 9540
rect 11054 9528 11060 9580
rect 11112 9568 11118 9580
rect 11241 9571 11299 9577
rect 11241 9568 11253 9571
rect 11112 9540 11253 9568
rect 11112 9528 11118 9540
rect 11241 9537 11253 9540
rect 11287 9537 11299 9571
rect 11241 9531 11299 9537
rect 11333 9571 11391 9577
rect 11333 9537 11345 9571
rect 11379 9537 11391 9571
rect 14645 9571 14703 9577
rect 14645 9568 14657 9571
rect 11333 9531 11391 9537
rect 13740 9540 14657 9568
rect 7092 9503 7150 9509
rect 7092 9469 7104 9503
rect 7138 9500 7150 9503
rect 7466 9500 7472 9512
rect 7138 9472 7472 9500
rect 7138 9469 7150 9472
rect 7092 9463 7150 9469
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 8202 9460 8208 9512
rect 8260 9500 8266 9512
rect 9125 9503 9183 9509
rect 9125 9500 9137 9503
rect 8260 9472 9137 9500
rect 8260 9460 8266 9472
rect 9125 9469 9137 9472
rect 9171 9469 9183 9503
rect 9125 9463 9183 9469
rect 10502 9460 10508 9512
rect 10560 9500 10566 9512
rect 10870 9500 10876 9512
rect 10560 9472 10876 9500
rect 10560 9460 10566 9472
rect 10870 9460 10876 9472
rect 10928 9500 10934 9512
rect 11348 9500 11376 9531
rect 12434 9500 12440 9512
rect 10928 9472 11376 9500
rect 12347 9472 12440 9500
rect 10928 9460 10934 9472
rect 12434 9460 12440 9472
rect 12492 9460 12498 9512
rect 12704 9503 12762 9509
rect 12704 9469 12716 9503
rect 12750 9500 12762 9503
rect 12986 9500 12992 9512
rect 12750 9472 12992 9500
rect 12750 9469 12762 9472
rect 12704 9463 12762 9469
rect 12986 9460 12992 9472
rect 13044 9460 13050 9512
rect 9392 9435 9450 9441
rect 6932 9404 9352 9432
rect 3237 9395 3295 9401
rect 3326 9364 3332 9376
rect 3287 9336 3332 9364
rect 3326 9324 3332 9336
rect 3384 9324 3390 9376
rect 4062 9324 4068 9376
rect 4120 9364 4126 9376
rect 5350 9364 5356 9376
rect 4120 9336 5356 9364
rect 4120 9324 4126 9336
rect 5350 9324 5356 9336
rect 5408 9324 5414 9376
rect 5442 9324 5448 9376
rect 5500 9364 5506 9376
rect 5629 9367 5687 9373
rect 5629 9364 5641 9367
rect 5500 9336 5641 9364
rect 5500 9324 5506 9336
rect 5629 9333 5641 9336
rect 5675 9333 5687 9367
rect 5629 9327 5687 9333
rect 6178 9324 6184 9376
rect 6236 9364 6242 9376
rect 8205 9367 8263 9373
rect 8205 9364 8217 9367
rect 6236 9336 8217 9364
rect 6236 9324 6242 9336
rect 8205 9333 8217 9336
rect 8251 9333 8263 9367
rect 9324 9364 9352 9404
rect 9392 9401 9404 9435
rect 9438 9432 9450 9435
rect 9582 9432 9588 9444
rect 9438 9404 9588 9432
rect 9438 9401 9450 9404
rect 9392 9395 9450 9401
rect 9582 9392 9588 9404
rect 9640 9392 9646 9444
rect 10226 9392 10232 9444
rect 10284 9432 10290 9444
rect 10284 9404 10824 9432
rect 10284 9392 10290 9404
rect 10502 9364 10508 9376
rect 9324 9336 10508 9364
rect 8205 9327 8263 9333
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 10796 9373 10824 9404
rect 11698 9392 11704 9444
rect 11756 9432 11762 9444
rect 11793 9435 11851 9441
rect 11793 9432 11805 9435
rect 11756 9404 11805 9432
rect 11756 9392 11762 9404
rect 11793 9401 11805 9404
rect 11839 9401 11851 9435
rect 12452 9432 12480 9460
rect 13170 9432 13176 9444
rect 12452 9404 13176 9432
rect 11793 9395 11851 9401
rect 13170 9392 13176 9404
rect 13228 9432 13234 9444
rect 13740 9432 13768 9540
rect 14645 9537 14657 9540
rect 14691 9537 14703 9571
rect 16758 9568 16764 9580
rect 16719 9540 16764 9568
rect 14645 9531 14703 9537
rect 14660 9500 14688 9531
rect 16758 9528 16764 9540
rect 16816 9528 16822 9580
rect 16853 9571 16911 9577
rect 16853 9537 16865 9571
rect 16899 9537 16911 9571
rect 20346 9568 20352 9580
rect 20307 9540 20352 9568
rect 16853 9531 16911 9537
rect 15194 9500 15200 9512
rect 14660 9472 15200 9500
rect 15194 9460 15200 9472
rect 15252 9460 15258 9512
rect 16868 9500 16896 9531
rect 20346 9528 20352 9540
rect 20404 9528 20410 9580
rect 17402 9500 17408 9512
rect 15580 9472 16896 9500
rect 17363 9472 17408 9500
rect 15580 9444 15608 9472
rect 17402 9460 17408 9472
rect 17460 9460 17466 9512
rect 17678 9460 17684 9512
rect 17736 9500 17742 9512
rect 18049 9503 18107 9509
rect 18049 9500 18061 9503
rect 17736 9472 18061 9500
rect 17736 9460 17742 9472
rect 18049 9469 18061 9472
rect 18095 9469 18107 9503
rect 18049 9463 18107 9469
rect 18138 9460 18144 9512
rect 18196 9500 18202 9512
rect 19426 9500 19432 9512
rect 18196 9472 19432 9500
rect 18196 9460 18202 9472
rect 19426 9460 19432 9472
rect 19484 9460 19490 9512
rect 20714 9500 20720 9512
rect 20675 9472 20720 9500
rect 20714 9460 20720 9472
rect 20772 9460 20778 9512
rect 13228 9404 13768 9432
rect 14912 9435 14970 9441
rect 13228 9392 13234 9404
rect 14912 9401 14924 9435
rect 14958 9432 14970 9435
rect 15562 9432 15568 9444
rect 14958 9404 15568 9432
rect 14958 9401 14970 9404
rect 14912 9395 14970 9401
rect 15562 9392 15568 9404
rect 15620 9392 15626 9444
rect 17218 9432 17224 9444
rect 15672 9404 17224 9432
rect 10781 9367 10839 9373
rect 10781 9333 10793 9367
rect 10827 9333 10839 9367
rect 11146 9364 11152 9376
rect 11107 9336 11152 9364
rect 10781 9327 10839 9333
rect 11146 9324 11152 9336
rect 11204 9324 11210 9376
rect 13814 9364 13820 9376
rect 13775 9336 13820 9364
rect 13814 9324 13820 9336
rect 13872 9324 13878 9376
rect 14182 9364 14188 9376
rect 14143 9336 14188 9364
rect 14182 9324 14188 9336
rect 14240 9324 14246 9376
rect 14458 9324 14464 9376
rect 14516 9364 14522 9376
rect 15672 9364 15700 9404
rect 17218 9392 17224 9404
rect 17276 9392 17282 9444
rect 18316 9435 18374 9441
rect 18316 9401 18328 9435
rect 18362 9432 18374 9435
rect 18506 9432 18512 9444
rect 18362 9404 18512 9432
rect 18362 9401 18374 9404
rect 18316 9395 18374 9401
rect 18506 9392 18512 9404
rect 18564 9392 18570 9444
rect 16022 9364 16028 9376
rect 14516 9336 15700 9364
rect 15983 9336 16028 9364
rect 14516 9324 14522 9336
rect 16022 9324 16028 9336
rect 16080 9324 16086 9376
rect 16666 9364 16672 9376
rect 16627 9336 16672 9364
rect 16666 9324 16672 9336
rect 16724 9324 16730 9376
rect 17589 9367 17647 9373
rect 17589 9333 17601 9367
rect 17635 9364 17647 9367
rect 17862 9364 17868 9376
rect 17635 9336 17868 9364
rect 17635 9333 17647 9336
rect 17589 9327 17647 9333
rect 17862 9324 17868 9336
rect 17920 9324 17926 9376
rect 19429 9367 19487 9373
rect 19429 9333 19441 9367
rect 19475 9364 19487 9367
rect 19518 9364 19524 9376
rect 19475 9336 19524 9364
rect 19475 9333 19487 9336
rect 19429 9327 19487 9333
rect 19518 9324 19524 9336
rect 19576 9324 19582 9376
rect 19702 9364 19708 9376
rect 19663 9336 19708 9364
rect 19702 9324 19708 9336
rect 19760 9324 19766 9376
rect 20070 9364 20076 9376
rect 20031 9336 20076 9364
rect 20070 9324 20076 9336
rect 20128 9324 20134 9376
rect 20162 9324 20168 9376
rect 20220 9364 20226 9376
rect 20220 9336 20265 9364
rect 20220 9324 20226 9336
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 3697 9163 3755 9169
rect 3697 9129 3709 9163
rect 3743 9160 3755 9163
rect 5074 9160 5080 9172
rect 3743 9132 5080 9160
rect 3743 9129 3755 9132
rect 3697 9123 3755 9129
rect 5074 9120 5080 9132
rect 5132 9120 5138 9172
rect 5353 9163 5411 9169
rect 5353 9129 5365 9163
rect 5399 9160 5411 9163
rect 5718 9160 5724 9172
rect 5399 9132 5724 9160
rect 5399 9129 5411 9132
rect 5353 9123 5411 9129
rect 5718 9120 5724 9132
rect 5776 9120 5782 9172
rect 5905 9163 5963 9169
rect 5905 9129 5917 9163
rect 5951 9129 5963 9163
rect 6362 9160 6368 9172
rect 6323 9132 6368 9160
rect 5905 9123 5963 9129
rect 4890 9052 4896 9104
rect 4948 9092 4954 9104
rect 4948 9064 5580 9092
rect 4948 9052 4954 9064
rect 2590 9033 2596 9036
rect 2584 9024 2596 9033
rect 2551 8996 2596 9024
rect 2584 8987 2596 8996
rect 2590 8984 2596 8987
rect 2648 8984 2654 9036
rect 5166 8984 5172 9036
rect 5224 9024 5230 9036
rect 5261 9027 5319 9033
rect 5261 9024 5273 9027
rect 5224 8996 5273 9024
rect 5224 8984 5230 8996
rect 5261 8993 5273 8996
rect 5307 8993 5319 9027
rect 5261 8987 5319 8993
rect 1578 8916 1584 8968
rect 1636 8956 1642 8968
rect 2317 8959 2375 8965
rect 2317 8956 2329 8959
rect 1636 8928 2329 8956
rect 1636 8916 1642 8928
rect 2317 8925 2329 8928
rect 2363 8925 2375 8959
rect 2317 8919 2375 8925
rect 4338 8916 4344 8968
rect 4396 8956 4402 8968
rect 5074 8956 5080 8968
rect 4396 8928 5080 8956
rect 4396 8916 4402 8928
rect 5074 8916 5080 8928
rect 5132 8916 5138 8968
rect 5552 8965 5580 9064
rect 5810 9052 5816 9104
rect 5868 9092 5874 9104
rect 5920 9092 5948 9123
rect 6362 9120 6368 9132
rect 6420 9120 6426 9172
rect 6730 9120 6736 9172
rect 6788 9160 6794 9172
rect 6917 9163 6975 9169
rect 6917 9160 6929 9163
rect 6788 9132 6929 9160
rect 6788 9120 6794 9132
rect 6917 9129 6929 9132
rect 6963 9129 6975 9163
rect 6917 9123 6975 9129
rect 7285 9163 7343 9169
rect 7285 9129 7297 9163
rect 7331 9160 7343 9163
rect 7374 9160 7380 9172
rect 7331 9132 7380 9160
rect 7331 9129 7343 9132
rect 7285 9123 7343 9129
rect 7374 9120 7380 9132
rect 7432 9120 7438 9172
rect 8297 9163 8355 9169
rect 8297 9129 8309 9163
rect 8343 9160 8355 9163
rect 8938 9160 8944 9172
rect 8343 9132 8944 9160
rect 8343 9129 8355 9132
rect 8297 9123 8355 9129
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 10137 9163 10195 9169
rect 10137 9129 10149 9163
rect 10183 9160 10195 9163
rect 10226 9160 10232 9172
rect 10183 9132 10232 9160
rect 10183 9129 10195 9132
rect 10137 9123 10195 9129
rect 10226 9120 10232 9132
rect 10284 9120 10290 9172
rect 10781 9163 10839 9169
rect 10781 9129 10793 9163
rect 10827 9160 10839 9163
rect 11146 9160 11152 9172
rect 10827 9132 11152 9160
rect 10827 9129 10839 9132
rect 10781 9123 10839 9129
rect 11146 9120 11152 9132
rect 11204 9120 11210 9172
rect 11609 9163 11667 9169
rect 11609 9129 11621 9163
rect 11655 9160 11667 9163
rect 11698 9160 11704 9172
rect 11655 9132 11704 9160
rect 11655 9129 11667 9132
rect 11609 9123 11667 9129
rect 11698 9120 11704 9132
rect 11756 9120 11762 9172
rect 12161 9163 12219 9169
rect 12161 9129 12173 9163
rect 12207 9160 12219 9163
rect 13354 9160 13360 9172
rect 12207 9132 13360 9160
rect 12207 9129 12219 9132
rect 12161 9123 12219 9129
rect 13354 9120 13360 9132
rect 13412 9120 13418 9172
rect 14550 9120 14556 9172
rect 14608 9160 14614 9172
rect 14608 9132 16620 9160
rect 14608 9120 14614 9132
rect 5868 9064 5948 9092
rect 5868 9052 5874 9064
rect 6178 9052 6184 9104
rect 6236 9092 6242 9104
rect 8846 9092 8852 9104
rect 6236 9064 6684 9092
rect 6236 9052 6242 9064
rect 5626 8984 5632 9036
rect 5684 9024 5690 9036
rect 6273 9027 6331 9033
rect 6273 9024 6285 9027
rect 5684 8996 6285 9024
rect 5684 8984 5690 8996
rect 6273 8993 6285 8996
rect 6319 9024 6331 9027
rect 6362 9024 6368 9036
rect 6319 8996 6368 9024
rect 6319 8993 6331 8996
rect 6273 8987 6331 8993
rect 6362 8984 6368 8996
rect 6420 8984 6426 9036
rect 5537 8959 5595 8965
rect 5537 8925 5549 8959
rect 5583 8956 5595 8959
rect 6546 8956 6552 8968
rect 5583 8928 6552 8956
rect 5583 8925 5595 8928
rect 5537 8919 5595 8925
rect 6546 8916 6552 8928
rect 6604 8916 6610 8968
rect 6656 8956 6684 9064
rect 7392 9064 8852 9092
rect 7392 9033 7420 9064
rect 8846 9052 8852 9064
rect 8904 9052 8910 9104
rect 9582 9052 9588 9104
rect 9640 9092 9646 9104
rect 11422 9092 11428 9104
rect 9640 9064 11428 9092
rect 9640 9052 9646 9064
rect 11422 9052 11428 9064
rect 11480 9052 11486 9104
rect 13624 9095 13682 9101
rect 13624 9061 13636 9095
rect 13670 9092 13682 9095
rect 16022 9092 16028 9104
rect 13670 9064 16028 9092
rect 13670 9061 13682 9064
rect 13624 9055 13682 9061
rect 16022 9052 16028 9064
rect 16080 9052 16086 9104
rect 16592 9092 16620 9132
rect 16666 9120 16672 9172
rect 16724 9160 16730 9172
rect 16945 9163 17003 9169
rect 16945 9160 16957 9163
rect 16724 9132 16957 9160
rect 16724 9120 16730 9132
rect 16945 9129 16957 9132
rect 16991 9129 17003 9163
rect 16945 9123 17003 9129
rect 17313 9163 17371 9169
rect 17313 9129 17325 9163
rect 17359 9160 17371 9163
rect 17773 9163 17831 9169
rect 17773 9160 17785 9163
rect 17359 9132 17785 9160
rect 17359 9129 17371 9132
rect 17313 9123 17371 9129
rect 17773 9129 17785 9132
rect 17819 9129 17831 9163
rect 17954 9160 17960 9172
rect 17915 9132 17960 9160
rect 17773 9123 17831 9129
rect 17954 9120 17960 9132
rect 18012 9120 18018 9172
rect 18325 9163 18383 9169
rect 18325 9129 18337 9163
rect 18371 9160 18383 9163
rect 19702 9160 19708 9172
rect 18371 9132 19708 9160
rect 18371 9129 18383 9132
rect 18325 9123 18383 9129
rect 19702 9120 19708 9132
rect 19760 9120 19766 9172
rect 21174 9160 21180 9172
rect 20180 9132 21180 9160
rect 17862 9092 17868 9104
rect 16592 9064 17868 9092
rect 17862 9052 17868 9064
rect 17920 9052 17926 9104
rect 18417 9095 18475 9101
rect 18417 9061 18429 9095
rect 18463 9092 18475 9095
rect 18874 9092 18880 9104
rect 18463 9064 18880 9092
rect 18463 9061 18475 9064
rect 18417 9055 18475 9061
rect 18874 9052 18880 9064
rect 18932 9052 18938 9104
rect 19337 9095 19395 9101
rect 19337 9061 19349 9095
rect 19383 9092 19395 9095
rect 20180 9092 20208 9132
rect 21174 9120 21180 9132
rect 21232 9120 21238 9172
rect 19383 9064 20208 9092
rect 20257 9095 20315 9101
rect 19383 9061 19395 9064
rect 19337 9055 19395 9061
rect 20257 9061 20269 9095
rect 20303 9092 20315 9095
rect 20714 9092 20720 9104
rect 20303 9064 20720 9092
rect 20303 9061 20315 9064
rect 20257 9055 20315 9061
rect 20714 9052 20720 9064
rect 20772 9052 20778 9104
rect 7377 9027 7435 9033
rect 7377 8993 7389 9027
rect 7423 8993 7435 9027
rect 7377 8987 7435 8993
rect 8389 9027 8447 9033
rect 8389 8993 8401 9027
rect 8435 8993 8447 9027
rect 8389 8987 8447 8993
rect 7469 8959 7527 8965
rect 7469 8956 7481 8959
rect 6656 8928 7481 8956
rect 7469 8925 7481 8928
rect 7515 8925 7527 8959
rect 7469 8919 7527 8925
rect 4893 8891 4951 8897
rect 4893 8857 4905 8891
rect 4939 8888 4951 8891
rect 6730 8888 6736 8900
rect 4939 8860 6736 8888
rect 4939 8857 4951 8860
rect 4893 8851 4951 8857
rect 6730 8848 6736 8860
rect 6788 8848 6794 8900
rect 8404 8888 8432 8987
rect 9122 8984 9128 9036
rect 9180 9024 9186 9036
rect 10778 9024 10784 9036
rect 9180 8996 10784 9024
rect 9180 8984 9186 8996
rect 10778 8984 10784 8996
rect 10836 8984 10842 9036
rect 11149 9027 11207 9033
rect 11149 8993 11161 9027
rect 11195 9024 11207 9027
rect 11609 9027 11667 9033
rect 11609 9024 11621 9027
rect 11195 8996 11621 9024
rect 11195 8993 11207 8996
rect 11149 8987 11207 8993
rect 11609 8993 11621 8996
rect 11655 8993 11667 9027
rect 11609 8987 11667 8993
rect 11698 8984 11704 9036
rect 11756 9024 11762 9036
rect 12253 9027 12311 9033
rect 12253 9024 12265 9027
rect 11756 8996 12265 9024
rect 11756 8984 11762 8996
rect 12253 8993 12265 8996
rect 12299 8993 12311 9027
rect 13262 9024 13268 9036
rect 12253 8987 12311 8993
rect 13096 8996 13268 9024
rect 8573 8959 8631 8965
rect 8573 8925 8585 8959
rect 8619 8956 8631 8959
rect 8846 8956 8852 8968
rect 8619 8928 8852 8956
rect 8619 8925 8631 8928
rect 8573 8919 8631 8925
rect 8846 8916 8852 8928
rect 8904 8916 8910 8968
rect 10226 8956 10232 8968
rect 10187 8928 10232 8956
rect 10226 8916 10232 8928
rect 10284 8916 10290 8968
rect 10413 8959 10471 8965
rect 10413 8925 10425 8959
rect 10459 8956 10471 8959
rect 10962 8956 10968 8968
rect 10459 8928 10968 8956
rect 10459 8925 10471 8928
rect 10413 8919 10471 8925
rect 10962 8916 10968 8928
rect 11020 8916 11026 8968
rect 11238 8956 11244 8968
rect 11199 8928 11244 8956
rect 11238 8916 11244 8928
rect 11296 8916 11302 8968
rect 11422 8956 11428 8968
rect 11335 8928 11428 8956
rect 11422 8916 11428 8928
rect 11480 8956 11486 8968
rect 11974 8956 11980 8968
rect 11480 8928 11980 8956
rect 11480 8916 11486 8928
rect 11974 8916 11980 8928
rect 12032 8916 12038 8968
rect 12342 8956 12348 8968
rect 12303 8928 12348 8956
rect 12342 8916 12348 8928
rect 12400 8916 12406 8968
rect 12250 8888 12256 8900
rect 8404 8860 12256 8888
rect 12250 8848 12256 8860
rect 12308 8848 12314 8900
rect 12434 8848 12440 8900
rect 12492 8888 12498 8900
rect 13096 8888 13124 8996
rect 13262 8984 13268 8996
rect 13320 9024 13326 9036
rect 15378 9024 15384 9036
rect 13320 8996 15384 9024
rect 13320 8984 13326 8996
rect 15378 8984 15384 8996
rect 15436 8984 15442 9036
rect 15556 9027 15614 9033
rect 15556 8993 15568 9027
rect 15602 9024 15614 9027
rect 16666 9024 16672 9036
rect 15602 8996 16672 9024
rect 15602 8993 15614 8996
rect 15556 8987 15614 8993
rect 16666 8984 16672 8996
rect 16724 8984 16730 9036
rect 17405 9027 17463 9033
rect 17405 8993 17417 9027
rect 17451 9024 17463 9027
rect 19702 9024 19708 9036
rect 17451 8996 19708 9024
rect 17451 8993 17463 8996
rect 17405 8987 17463 8993
rect 19702 8984 19708 8996
rect 19760 8984 19766 9036
rect 19978 9024 19984 9036
rect 19939 8996 19984 9024
rect 19978 8984 19984 8996
rect 20036 8984 20042 9036
rect 13357 8959 13415 8965
rect 13357 8956 13369 8959
rect 13280 8928 13369 8956
rect 13280 8900 13308 8928
rect 13357 8925 13369 8928
rect 13403 8925 13415 8959
rect 13357 8919 13415 8925
rect 15194 8916 15200 8968
rect 15252 8956 15258 8968
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 15252 8928 15301 8956
rect 15252 8916 15258 8928
rect 15289 8925 15301 8928
rect 15335 8925 15347 8959
rect 16684 8956 16712 8984
rect 16850 8956 16856 8968
rect 16684 8928 16856 8956
rect 15289 8919 15347 8925
rect 16850 8916 16856 8928
rect 16908 8956 16914 8968
rect 17497 8959 17555 8965
rect 17497 8956 17509 8959
rect 16908 8928 17509 8956
rect 16908 8916 16914 8928
rect 17497 8925 17509 8928
rect 17543 8925 17555 8959
rect 18598 8956 18604 8968
rect 18559 8928 18604 8956
rect 17497 8919 17555 8925
rect 18598 8916 18604 8928
rect 18656 8916 18662 8968
rect 19242 8916 19248 8968
rect 19300 8956 19306 8968
rect 19429 8959 19487 8965
rect 19429 8956 19441 8959
rect 19300 8928 19441 8956
rect 19300 8916 19306 8928
rect 19429 8925 19441 8928
rect 19475 8925 19487 8959
rect 19610 8956 19616 8968
rect 19523 8928 19616 8956
rect 19429 8919 19487 8925
rect 19610 8916 19616 8928
rect 19668 8956 19674 8968
rect 20346 8956 20352 8968
rect 19668 8928 20352 8956
rect 19668 8916 19674 8928
rect 20346 8916 20352 8928
rect 20404 8916 20410 8968
rect 12492 8860 13124 8888
rect 12492 8848 12498 8860
rect 13262 8848 13268 8900
rect 13320 8848 13326 8900
rect 17773 8891 17831 8897
rect 17773 8857 17785 8891
rect 17819 8888 17831 8891
rect 18782 8888 18788 8900
rect 17819 8860 18788 8888
rect 17819 8857 17831 8860
rect 17773 8851 17831 8857
rect 18782 8848 18788 8860
rect 18840 8848 18846 8900
rect 18966 8888 18972 8900
rect 18927 8860 18972 8888
rect 18966 8848 18972 8860
rect 19024 8848 19030 8900
rect 7374 8780 7380 8832
rect 7432 8820 7438 8832
rect 7929 8823 7987 8829
rect 7929 8820 7941 8823
rect 7432 8792 7941 8820
rect 7432 8780 7438 8792
rect 7929 8789 7941 8792
rect 7975 8789 7987 8823
rect 7929 8783 7987 8789
rect 8018 8780 8024 8832
rect 8076 8820 8082 8832
rect 8386 8820 8392 8832
rect 8076 8792 8392 8820
rect 8076 8780 8082 8792
rect 8386 8780 8392 8792
rect 8444 8820 8450 8832
rect 8662 8820 8668 8832
rect 8444 8792 8668 8820
rect 8444 8780 8450 8792
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 9769 8823 9827 8829
rect 9769 8789 9781 8823
rect 9815 8820 9827 8823
rect 11146 8820 11152 8832
rect 9815 8792 11152 8820
rect 9815 8789 9827 8792
rect 9769 8783 9827 8789
rect 11146 8780 11152 8792
rect 11204 8780 11210 8832
rect 11793 8823 11851 8829
rect 11793 8789 11805 8823
rect 11839 8820 11851 8823
rect 13354 8820 13360 8832
rect 11839 8792 13360 8820
rect 11839 8789 11851 8792
rect 11793 8783 11851 8789
rect 13354 8780 13360 8792
rect 13412 8780 13418 8832
rect 14274 8780 14280 8832
rect 14332 8820 14338 8832
rect 14642 8820 14648 8832
rect 14332 8792 14648 8820
rect 14332 8780 14338 8792
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 14737 8823 14795 8829
rect 14737 8789 14749 8823
rect 14783 8820 14795 8823
rect 15194 8820 15200 8832
rect 14783 8792 15200 8820
rect 14783 8789 14795 8792
rect 14737 8783 14795 8789
rect 15194 8780 15200 8792
rect 15252 8820 15258 8832
rect 15470 8820 15476 8832
rect 15252 8792 15476 8820
rect 15252 8780 15258 8792
rect 15470 8780 15476 8792
rect 15528 8780 15534 8832
rect 15562 8780 15568 8832
rect 15620 8820 15626 8832
rect 16669 8823 16727 8829
rect 16669 8820 16681 8823
rect 15620 8792 16681 8820
rect 15620 8780 15626 8792
rect 16669 8789 16681 8792
rect 16715 8789 16727 8823
rect 16669 8783 16727 8789
rect 16758 8780 16764 8832
rect 16816 8820 16822 8832
rect 19978 8820 19984 8832
rect 16816 8792 19984 8820
rect 16816 8780 16822 8792
rect 19978 8780 19984 8792
rect 20036 8780 20042 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 3694 8576 3700 8628
rect 3752 8616 3758 8628
rect 6365 8619 6423 8625
rect 6365 8616 6377 8619
rect 3752 8588 6377 8616
rect 3752 8576 3758 8588
rect 6365 8585 6377 8588
rect 6411 8585 6423 8619
rect 6365 8579 6423 8585
rect 2590 8508 2596 8560
rect 2648 8548 2654 8560
rect 2777 8551 2835 8557
rect 2777 8548 2789 8551
rect 2648 8520 2789 8548
rect 2648 8508 2654 8520
rect 2777 8517 2789 8520
rect 2823 8517 2835 8551
rect 5077 8551 5135 8557
rect 5077 8548 5089 8551
rect 2777 8511 2835 8517
rect 4724 8520 5089 8548
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 1486 8412 1492 8424
rect 1443 8384 1492 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 1486 8372 1492 8384
rect 1544 8372 1550 8424
rect 3694 8412 3700 8424
rect 3655 8384 3700 8412
rect 3694 8372 3700 8384
rect 3752 8372 3758 8424
rect 4724 8412 4752 8520
rect 5077 8517 5089 8520
rect 5123 8548 5135 8551
rect 6380 8548 6408 8579
rect 9582 8576 9588 8628
rect 9640 8616 9646 8628
rect 9677 8619 9735 8625
rect 9677 8616 9689 8619
rect 9640 8588 9689 8616
rect 9640 8576 9646 8588
rect 9677 8585 9689 8588
rect 9723 8585 9735 8619
rect 9677 8579 9735 8585
rect 10226 8576 10232 8628
rect 10284 8616 10290 8628
rect 11149 8619 11207 8625
rect 11149 8616 11161 8619
rect 10284 8588 11161 8616
rect 10284 8576 10290 8588
rect 11149 8585 11161 8588
rect 11195 8585 11207 8619
rect 11149 8579 11207 8585
rect 13170 8576 13176 8628
rect 13228 8616 13234 8628
rect 13814 8616 13820 8628
rect 13228 8588 13820 8616
rect 13228 8576 13234 8588
rect 13814 8576 13820 8588
rect 13872 8576 13878 8628
rect 15105 8619 15163 8625
rect 15105 8585 15117 8619
rect 15151 8616 15163 8619
rect 15654 8616 15660 8628
rect 15151 8588 15660 8616
rect 15151 8585 15163 8588
rect 15105 8579 15163 8585
rect 15654 8576 15660 8588
rect 15712 8576 15718 8628
rect 16482 8576 16488 8628
rect 16540 8616 16546 8628
rect 17954 8616 17960 8628
rect 16540 8588 17960 8616
rect 16540 8576 16546 8588
rect 17954 8576 17960 8588
rect 18012 8576 18018 8628
rect 18049 8619 18107 8625
rect 18049 8585 18061 8619
rect 18095 8616 18107 8619
rect 18598 8616 18604 8628
rect 18095 8588 18604 8616
rect 18095 8585 18107 8588
rect 18049 8579 18107 8585
rect 18598 8576 18604 8588
rect 18656 8576 18662 8628
rect 18874 8576 18880 8628
rect 18932 8616 18938 8628
rect 19061 8619 19119 8625
rect 19061 8616 19073 8619
rect 18932 8588 19073 8616
rect 18932 8576 18938 8588
rect 19061 8585 19073 8588
rect 19107 8585 19119 8619
rect 19061 8579 19119 8585
rect 19426 8576 19432 8628
rect 19484 8616 19490 8628
rect 19484 8588 19564 8616
rect 19484 8576 19490 8588
rect 6822 8548 6828 8560
rect 5123 8520 5948 8548
rect 6380 8520 6828 8548
rect 5123 8517 5135 8520
rect 5077 8511 5135 8517
rect 5920 8489 5948 8520
rect 6822 8508 6828 8520
rect 6880 8508 6886 8560
rect 7006 8508 7012 8560
rect 7064 8548 7070 8560
rect 7064 8520 7328 8548
rect 7064 8508 7070 8520
rect 7300 8492 7328 8520
rect 9858 8508 9864 8560
rect 9916 8548 9922 8560
rect 10045 8551 10103 8557
rect 10045 8548 10057 8551
rect 9916 8520 10057 8548
rect 9916 8508 9922 8520
rect 10045 8517 10057 8520
rect 10091 8517 10103 8551
rect 10045 8511 10103 8517
rect 10137 8551 10195 8557
rect 10137 8517 10149 8551
rect 10183 8548 10195 8551
rect 11054 8548 11060 8560
rect 10183 8520 11060 8548
rect 10183 8517 10195 8520
rect 10137 8511 10195 8517
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8449 5963 8483
rect 7282 8480 7288 8492
rect 5905 8443 5963 8449
rect 6012 8452 7144 8480
rect 7243 8452 7288 8480
rect 3896 8384 4752 8412
rect 1664 8347 1722 8353
rect 1664 8313 1676 8347
rect 1710 8344 1722 8347
rect 2130 8344 2136 8356
rect 1710 8316 2136 8344
rect 1710 8313 1722 8316
rect 1664 8307 1722 8313
rect 2130 8304 2136 8316
rect 2188 8344 2194 8356
rect 3896 8344 3924 8384
rect 5166 8372 5172 8424
rect 5224 8412 5230 8424
rect 6012 8412 6040 8452
rect 5224 8384 6040 8412
rect 6549 8415 6607 8421
rect 5224 8372 5230 8384
rect 6549 8381 6561 8415
rect 6595 8412 6607 8415
rect 6914 8412 6920 8424
rect 6595 8384 6920 8412
rect 6595 8381 6607 8384
rect 6549 8375 6607 8381
rect 6914 8372 6920 8384
rect 6972 8372 6978 8424
rect 3970 8353 3976 8356
rect 2188 8316 3924 8344
rect 2188 8304 2194 8316
rect 3964 8307 3976 8353
rect 4028 8344 4034 8356
rect 5813 8347 5871 8353
rect 4028 8316 4064 8344
rect 4172 8316 5396 8344
rect 3970 8304 3976 8307
rect 4028 8304 4034 8316
rect 3878 8236 3884 8288
rect 3936 8276 3942 8288
rect 4172 8276 4200 8316
rect 5368 8285 5396 8316
rect 5813 8313 5825 8347
rect 5859 8344 5871 8347
rect 7006 8344 7012 8356
rect 5859 8316 7012 8344
rect 5859 8313 5871 8316
rect 5813 8307 5871 8313
rect 7006 8304 7012 8316
rect 7064 8304 7070 8356
rect 7116 8344 7144 8452
rect 7282 8440 7288 8452
rect 7340 8440 7346 8492
rect 7466 8480 7472 8492
rect 7427 8452 7472 8480
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 7193 8415 7251 8421
rect 7193 8381 7205 8415
rect 7239 8412 7251 8415
rect 8018 8412 8024 8424
rect 7239 8384 8024 8412
rect 7239 8381 7251 8384
rect 7193 8375 7251 8381
rect 8018 8372 8024 8384
rect 8076 8372 8082 8424
rect 8202 8372 8208 8424
rect 8260 8412 8266 8424
rect 8297 8415 8355 8421
rect 8297 8412 8309 8415
rect 8260 8384 8309 8412
rect 8260 8372 8266 8384
rect 8297 8381 8309 8384
rect 8343 8381 8355 8415
rect 9858 8412 9864 8424
rect 8297 8375 8355 8381
rect 8404 8384 9864 8412
rect 8404 8344 8432 8384
rect 9858 8372 9864 8384
rect 9916 8372 9922 8424
rect 7116 8316 8432 8344
rect 8564 8347 8622 8353
rect 8564 8313 8576 8347
rect 8610 8344 8622 8347
rect 8754 8344 8760 8356
rect 8610 8316 8760 8344
rect 8610 8313 8622 8316
rect 8564 8307 8622 8313
rect 8754 8304 8760 8316
rect 8812 8304 8818 8356
rect 9122 8304 9128 8356
rect 9180 8344 9186 8356
rect 10060 8344 10088 8511
rect 11054 8508 11060 8520
rect 11112 8508 11118 8560
rect 11606 8508 11612 8560
rect 11664 8548 11670 8560
rect 12342 8548 12348 8560
rect 11664 8520 12348 8548
rect 11664 8508 11670 8520
rect 12342 8508 12348 8520
rect 12400 8508 12406 8560
rect 14093 8551 14151 8557
rect 14093 8517 14105 8551
rect 14139 8548 14151 8551
rect 14139 8520 16896 8548
rect 14139 8517 14151 8520
rect 14093 8511 14151 8517
rect 10689 8483 10747 8489
rect 10689 8449 10701 8483
rect 10735 8449 10747 8483
rect 10689 8443 10747 8449
rect 10318 8372 10324 8424
rect 10376 8412 10382 8424
rect 10704 8412 10732 8443
rect 10870 8440 10876 8492
rect 10928 8480 10934 8492
rect 11701 8483 11759 8489
rect 11701 8480 11713 8483
rect 10928 8452 11713 8480
rect 10928 8440 10934 8452
rect 11701 8449 11713 8452
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 13998 8440 14004 8492
rect 14056 8480 14062 8492
rect 14274 8480 14280 8492
rect 14056 8452 14280 8480
rect 14056 8440 14062 8452
rect 14274 8440 14280 8452
rect 14332 8480 14338 8492
rect 14553 8483 14611 8489
rect 14553 8480 14565 8483
rect 14332 8452 14565 8480
rect 14332 8440 14338 8452
rect 14553 8449 14565 8452
rect 14599 8449 14611 8483
rect 14553 8443 14611 8449
rect 14642 8440 14648 8492
rect 14700 8480 14706 8492
rect 14737 8483 14795 8489
rect 14737 8480 14749 8483
rect 14700 8452 14749 8480
rect 14700 8440 14706 8452
rect 14737 8449 14749 8452
rect 14783 8480 14795 8483
rect 15378 8480 15384 8492
rect 14783 8452 15384 8480
rect 14783 8449 14795 8452
rect 14737 8443 14795 8449
rect 15378 8440 15384 8452
rect 15436 8440 15442 8492
rect 15562 8440 15568 8492
rect 15620 8480 15626 8492
rect 15657 8483 15715 8489
rect 15657 8480 15669 8483
rect 15620 8452 15669 8480
rect 15620 8440 15626 8452
rect 15657 8449 15669 8452
rect 15703 8449 15715 8483
rect 15657 8443 15715 8449
rect 15746 8440 15752 8492
rect 15804 8480 15810 8492
rect 16577 8483 16635 8489
rect 16577 8480 16589 8483
rect 15804 8452 16589 8480
rect 15804 8440 15810 8452
rect 16577 8449 16589 8452
rect 16623 8449 16635 8483
rect 16758 8480 16764 8492
rect 16719 8452 16764 8480
rect 16577 8443 16635 8449
rect 16758 8440 16764 8452
rect 16816 8440 16822 8492
rect 16868 8480 16896 8520
rect 17126 8508 17132 8560
rect 17184 8548 17190 8560
rect 17313 8551 17371 8557
rect 17313 8548 17325 8551
rect 17184 8520 17325 8548
rect 17184 8508 17190 8520
rect 17313 8517 17325 8520
rect 17359 8517 17371 8551
rect 17678 8548 17684 8560
rect 17639 8520 17684 8548
rect 17313 8511 17371 8517
rect 17678 8508 17684 8520
rect 17736 8508 17742 8560
rect 18230 8480 18236 8492
rect 16868 8452 18236 8480
rect 18230 8440 18236 8452
rect 18288 8440 18294 8492
rect 18693 8483 18751 8489
rect 18693 8449 18705 8483
rect 18739 8480 18751 8483
rect 19334 8480 19340 8492
rect 18739 8452 19340 8480
rect 18739 8449 18751 8452
rect 18693 8443 18751 8449
rect 19334 8440 19340 8452
rect 19392 8440 19398 8492
rect 19536 8489 19564 8588
rect 20073 8551 20131 8557
rect 20073 8517 20085 8551
rect 20119 8548 20131 8551
rect 20254 8548 20260 8560
rect 20119 8520 20260 8548
rect 20119 8517 20131 8520
rect 20073 8511 20131 8517
rect 20254 8508 20260 8520
rect 20312 8508 20318 8560
rect 19521 8483 19579 8489
rect 19521 8449 19533 8483
rect 19567 8449 19579 8483
rect 19521 8443 19579 8449
rect 19610 8440 19616 8492
rect 19668 8480 19674 8492
rect 20625 8483 20683 8489
rect 19668 8452 19713 8480
rect 19668 8440 19674 8452
rect 20625 8449 20637 8483
rect 20671 8449 20683 8483
rect 20625 8443 20683 8449
rect 10376 8384 10732 8412
rect 10376 8372 10382 8384
rect 10778 8372 10784 8424
rect 10836 8412 10842 8424
rect 11517 8415 11575 8421
rect 11517 8412 11529 8415
rect 10836 8384 11529 8412
rect 10836 8372 10842 8384
rect 11517 8381 11529 8384
rect 11563 8381 11575 8415
rect 11517 8375 11575 8381
rect 12066 8372 12072 8424
rect 12124 8412 12130 8424
rect 12437 8415 12495 8421
rect 12124 8384 12388 8412
rect 12124 8372 12130 8384
rect 10505 8347 10563 8353
rect 10505 8344 10517 8347
rect 9180 8316 10517 8344
rect 9180 8304 9186 8316
rect 10505 8313 10517 8316
rect 10551 8313 10563 8347
rect 10505 8307 10563 8313
rect 10597 8347 10655 8353
rect 10597 8313 10609 8347
rect 10643 8344 10655 8347
rect 12360 8344 12388 8384
rect 12437 8381 12449 8415
rect 12483 8412 12495 8415
rect 13262 8412 13268 8424
rect 12483 8384 13268 8412
rect 12483 8381 12495 8384
rect 12437 8375 12495 8381
rect 13262 8372 13268 8384
rect 13320 8372 13326 8424
rect 14182 8372 14188 8424
rect 14240 8412 14246 8424
rect 16485 8415 16543 8421
rect 16485 8412 16497 8415
rect 14240 8384 16497 8412
rect 14240 8372 14246 8384
rect 16485 8381 16497 8384
rect 16531 8381 16543 8415
rect 16485 8375 16543 8381
rect 17129 8415 17187 8421
rect 17129 8381 17141 8415
rect 17175 8381 17187 8415
rect 17862 8412 17868 8424
rect 17823 8384 17868 8412
rect 17129 8375 17187 8381
rect 12704 8347 12762 8353
rect 12704 8344 12716 8347
rect 10643 8316 12296 8344
rect 12360 8316 12716 8344
rect 10643 8313 10655 8316
rect 10597 8307 10655 8313
rect 3936 8248 4200 8276
rect 5353 8279 5411 8285
rect 3936 8236 3942 8248
rect 5353 8245 5365 8279
rect 5399 8245 5411 8279
rect 5718 8276 5724 8288
rect 5679 8248 5724 8276
rect 5353 8239 5411 8245
rect 5718 8236 5724 8248
rect 5776 8236 5782 8288
rect 6822 8276 6828 8288
rect 6783 8248 6828 8276
rect 6822 8236 6828 8248
rect 6880 8236 6886 8288
rect 9306 8236 9312 8288
rect 9364 8276 9370 8288
rect 9490 8276 9496 8288
rect 9364 8248 9496 8276
rect 9364 8236 9370 8248
rect 9490 8236 9496 8248
rect 9548 8236 9554 8288
rect 9858 8236 9864 8288
rect 9916 8276 9922 8288
rect 11609 8279 11667 8285
rect 11609 8276 11621 8279
rect 9916 8248 11621 8276
rect 9916 8236 9922 8248
rect 11609 8245 11621 8248
rect 11655 8245 11667 8279
rect 12268 8276 12296 8316
rect 12704 8313 12716 8316
rect 12750 8344 12762 8347
rect 15194 8344 15200 8356
rect 12750 8316 15200 8344
rect 12750 8313 12762 8316
rect 12704 8307 12762 8313
rect 15194 8304 15200 8316
rect 15252 8304 15258 8356
rect 15473 8347 15531 8353
rect 15473 8313 15485 8347
rect 15519 8344 15531 8347
rect 15519 8316 16160 8344
rect 15519 8313 15531 8316
rect 15473 8307 15531 8313
rect 12434 8276 12440 8288
rect 12268 8248 12440 8276
rect 11609 8239 11667 8245
rect 12434 8236 12440 8248
rect 12492 8236 12498 8288
rect 12986 8236 12992 8288
rect 13044 8276 13050 8288
rect 13817 8279 13875 8285
rect 13817 8276 13829 8279
rect 13044 8248 13829 8276
rect 13044 8236 13050 8248
rect 13817 8245 13829 8248
rect 13863 8245 13875 8279
rect 13817 8239 13875 8245
rect 13906 8236 13912 8288
rect 13964 8276 13970 8288
rect 14461 8279 14519 8285
rect 14461 8276 14473 8279
rect 13964 8248 14473 8276
rect 13964 8236 13970 8248
rect 14461 8245 14473 8248
rect 14507 8276 14519 8279
rect 15010 8276 15016 8288
rect 14507 8248 15016 8276
rect 14507 8245 14519 8248
rect 14461 8239 14519 8245
rect 15010 8236 15016 8248
rect 15068 8236 15074 8288
rect 15562 8276 15568 8288
rect 15523 8248 15568 8276
rect 15562 8236 15568 8248
rect 15620 8236 15626 8288
rect 16132 8285 16160 8316
rect 16298 8304 16304 8356
rect 16356 8344 16362 8356
rect 17144 8344 17172 8375
rect 17862 8372 17868 8384
rect 17920 8372 17926 8424
rect 19426 8412 19432 8424
rect 19387 8384 19432 8412
rect 19426 8372 19432 8384
rect 19484 8372 19490 8424
rect 19794 8372 19800 8424
rect 19852 8412 19858 8424
rect 20530 8412 20536 8424
rect 19852 8384 20536 8412
rect 19852 8372 19858 8384
rect 20530 8372 20536 8384
rect 20588 8412 20594 8424
rect 20640 8412 20668 8443
rect 20588 8384 20668 8412
rect 20588 8372 20594 8384
rect 16356 8316 17172 8344
rect 16356 8304 16362 8316
rect 17770 8304 17776 8356
rect 17828 8344 17834 8356
rect 18509 8347 18567 8353
rect 18509 8344 18521 8347
rect 17828 8316 18521 8344
rect 17828 8304 17834 8316
rect 18509 8313 18521 8316
rect 18555 8313 18567 8347
rect 18509 8307 18567 8313
rect 19702 8304 19708 8356
rect 19760 8344 19766 8356
rect 20438 8344 20444 8356
rect 19760 8316 20444 8344
rect 19760 8304 19766 8316
rect 20438 8304 20444 8316
rect 20496 8304 20502 8356
rect 16117 8279 16175 8285
rect 16117 8245 16129 8279
rect 16163 8245 16175 8279
rect 16117 8239 16175 8245
rect 17586 8236 17592 8288
rect 17644 8276 17650 8288
rect 18230 8276 18236 8288
rect 17644 8248 18236 8276
rect 17644 8236 17650 8248
rect 18230 8236 18236 8248
rect 18288 8236 18294 8288
rect 18414 8276 18420 8288
rect 18375 8248 18420 8276
rect 18414 8236 18420 8248
rect 18472 8236 18478 8288
rect 19978 8236 19984 8288
rect 20036 8276 20042 8288
rect 20533 8279 20591 8285
rect 20533 8276 20545 8279
rect 20036 8248 20545 8276
rect 20036 8236 20042 8248
rect 20533 8245 20545 8248
rect 20579 8276 20591 8279
rect 21358 8276 21364 8288
rect 20579 8248 21364 8276
rect 20579 8245 20591 8248
rect 20533 8239 20591 8245
rect 21358 8236 21364 8248
rect 21416 8236 21422 8288
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 2961 8075 3019 8081
rect 2961 8041 2973 8075
rect 3007 8072 3019 8075
rect 3050 8072 3056 8084
rect 3007 8044 3056 8072
rect 3007 8041 3019 8044
rect 2961 8035 3019 8041
rect 3050 8032 3056 8044
rect 3108 8072 3114 8084
rect 3326 8072 3332 8084
rect 3108 8044 3332 8072
rect 3108 8032 3114 8044
rect 3326 8032 3332 8044
rect 3384 8032 3390 8084
rect 5718 8032 5724 8084
rect 5776 8072 5782 8084
rect 5997 8075 6055 8081
rect 5997 8072 6009 8075
rect 5776 8044 6009 8072
rect 5776 8032 5782 8044
rect 5997 8041 6009 8044
rect 6043 8041 6055 8075
rect 5997 8035 6055 8041
rect 6365 8075 6423 8081
rect 6365 8041 6377 8075
rect 6411 8072 6423 8075
rect 6822 8072 6828 8084
rect 6411 8044 6828 8072
rect 6411 8041 6423 8044
rect 6365 8035 6423 8041
rect 6822 8032 6828 8044
rect 6880 8032 6886 8084
rect 7006 8072 7012 8084
rect 6967 8044 7012 8072
rect 7006 8032 7012 8044
rect 7064 8032 7070 8084
rect 7374 8072 7380 8084
rect 7335 8044 7380 8072
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 8573 8075 8631 8081
rect 8573 8041 8585 8075
rect 8619 8072 8631 8075
rect 8662 8072 8668 8084
rect 8619 8044 8668 8072
rect 8619 8041 8631 8044
rect 8573 8035 8631 8041
rect 8662 8032 8668 8044
rect 8720 8032 8726 8084
rect 9033 8075 9091 8081
rect 9033 8041 9045 8075
rect 9079 8072 9091 8075
rect 9677 8075 9735 8081
rect 9677 8072 9689 8075
rect 9079 8044 9689 8072
rect 9079 8041 9091 8044
rect 9033 8035 9091 8041
rect 9677 8041 9689 8044
rect 9723 8041 9735 8075
rect 9677 8035 9735 8041
rect 10045 8075 10103 8081
rect 10045 8041 10057 8075
rect 10091 8072 10103 8075
rect 10410 8072 10416 8084
rect 10091 8044 10416 8072
rect 10091 8041 10103 8044
rect 10045 8035 10103 8041
rect 10410 8032 10416 8044
rect 10468 8032 10474 8084
rect 10689 8075 10747 8081
rect 10689 8041 10701 8075
rect 10735 8072 10747 8075
rect 10778 8072 10784 8084
rect 10735 8044 10784 8072
rect 10735 8041 10747 8044
rect 10689 8035 10747 8041
rect 10778 8032 10784 8044
rect 10836 8032 10842 8084
rect 11054 8032 11060 8084
rect 11112 8072 11118 8084
rect 11149 8075 11207 8081
rect 11149 8072 11161 8075
rect 11112 8044 11161 8072
rect 11112 8032 11118 8044
rect 11149 8041 11161 8044
rect 11195 8041 11207 8075
rect 11698 8072 11704 8084
rect 11659 8044 11704 8072
rect 11149 8035 11207 8041
rect 11698 8032 11704 8044
rect 11756 8032 11762 8084
rect 12161 8075 12219 8081
rect 12161 8041 12173 8075
rect 12207 8072 12219 8075
rect 12713 8075 12771 8081
rect 12713 8072 12725 8075
rect 12207 8044 12725 8072
rect 12207 8041 12219 8044
rect 12161 8035 12219 8041
rect 12713 8041 12725 8044
rect 12759 8041 12771 8075
rect 12713 8035 12771 8041
rect 13538 8032 13544 8084
rect 13596 8072 13602 8084
rect 15289 8075 15347 8081
rect 13596 8044 14688 8072
rect 13596 8032 13602 8044
rect 3970 8004 3976 8016
rect 3620 7976 3976 8004
rect 1670 7896 1676 7948
rect 1728 7936 1734 7948
rect 1857 7939 1915 7945
rect 1857 7936 1869 7939
rect 1728 7908 1869 7936
rect 1728 7896 1734 7908
rect 1857 7905 1869 7908
rect 1903 7936 1915 7939
rect 2406 7936 2412 7948
rect 1903 7908 2412 7936
rect 1903 7905 1915 7908
rect 1857 7899 1915 7905
rect 2406 7896 2412 7908
rect 2464 7896 2470 7948
rect 2869 7939 2927 7945
rect 2869 7905 2881 7939
rect 2915 7936 2927 7939
rect 3513 7939 3571 7945
rect 3513 7936 3525 7939
rect 2915 7908 3525 7936
rect 2915 7905 2927 7908
rect 2869 7899 2927 7905
rect 3513 7905 3525 7908
rect 3559 7905 3571 7939
rect 3513 7899 3571 7905
rect 1949 7871 2007 7877
rect 1949 7837 1961 7871
rect 1995 7837 2007 7871
rect 1949 7831 2007 7837
rect 2133 7871 2191 7877
rect 2133 7837 2145 7871
rect 2179 7868 2191 7871
rect 3145 7871 3203 7877
rect 3145 7868 3157 7871
rect 2179 7840 3157 7868
rect 2179 7837 2191 7840
rect 2133 7831 2191 7837
rect 3145 7837 3157 7840
rect 3191 7868 3203 7871
rect 3620 7868 3648 7976
rect 3970 7964 3976 7976
rect 4028 8004 4034 8016
rect 4028 7976 5764 8004
rect 4028 7964 4034 7976
rect 3694 7896 3700 7948
rect 3752 7936 3758 7948
rect 4341 7939 4399 7945
rect 4341 7936 4353 7939
rect 3752 7908 4353 7936
rect 3752 7896 3758 7908
rect 4341 7905 4353 7908
rect 4387 7905 4399 7939
rect 4341 7899 4399 7905
rect 4608 7939 4666 7945
rect 4608 7905 4620 7939
rect 4654 7936 4666 7939
rect 4890 7936 4896 7948
rect 4654 7908 4896 7936
rect 4654 7905 4666 7908
rect 4608 7899 4666 7905
rect 4890 7896 4896 7908
rect 4948 7896 4954 7948
rect 3191 7840 3648 7868
rect 5736 7868 5764 7976
rect 5902 7964 5908 8016
rect 5960 8004 5966 8016
rect 6457 8007 6515 8013
rect 6457 8004 6469 8007
rect 5960 7976 6469 8004
rect 5960 7964 5966 7976
rect 6457 7973 6469 7976
rect 6503 7973 6515 8007
rect 6457 7967 6515 7973
rect 6730 7964 6736 8016
rect 6788 8004 6794 8016
rect 7469 8007 7527 8013
rect 7469 8004 7481 8007
rect 6788 7976 7481 8004
rect 6788 7964 6794 7976
rect 7469 7973 7481 7976
rect 7515 7973 7527 8007
rect 7469 7967 7527 7973
rect 8754 7964 8760 8016
rect 8812 8004 8818 8016
rect 12069 8007 12127 8013
rect 8812 7976 9720 8004
rect 8812 7964 8818 7976
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 8389 7939 8447 7945
rect 8389 7936 8401 7939
rect 6972 7908 8401 7936
rect 6972 7896 6978 7908
rect 8389 7905 8401 7908
rect 8435 7905 8447 7939
rect 8389 7899 8447 7905
rect 8941 7939 8999 7945
rect 8941 7905 8953 7939
rect 8987 7936 8999 7939
rect 9490 7936 9496 7948
rect 8987 7908 9496 7936
rect 8987 7905 8999 7908
rect 8941 7899 8999 7905
rect 9490 7896 9496 7908
rect 9548 7896 9554 7948
rect 6641 7871 6699 7877
rect 6641 7868 6653 7871
rect 5736 7840 6653 7868
rect 3191 7837 3203 7840
rect 3145 7831 3203 7837
rect 1964 7800 1992 7831
rect 4154 7800 4160 7812
rect 1964 7772 4160 7800
rect 4154 7760 4160 7772
rect 4212 7760 4218 7812
rect 5736 7809 5764 7840
rect 6641 7837 6653 7840
rect 6687 7868 6699 7871
rect 7561 7871 7619 7877
rect 7561 7868 7573 7871
rect 6687 7840 7573 7868
rect 6687 7837 6699 7840
rect 6641 7831 6699 7837
rect 7561 7837 7573 7840
rect 7607 7837 7619 7871
rect 7561 7831 7619 7837
rect 7650 7828 7656 7880
rect 7708 7868 7714 7880
rect 8110 7868 8116 7880
rect 7708 7840 8116 7868
rect 7708 7828 7714 7840
rect 8110 7828 8116 7840
rect 8168 7828 8174 7880
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7868 9275 7871
rect 9582 7868 9588 7880
rect 9263 7840 9588 7868
rect 9263 7837 9275 7840
rect 9217 7831 9275 7837
rect 9582 7828 9588 7840
rect 9640 7828 9646 7880
rect 9692 7868 9720 7976
rect 12069 7973 12081 8007
rect 12115 8004 12127 8007
rect 12526 8004 12532 8016
rect 12115 7976 12532 8004
rect 12115 7973 12127 7976
rect 12069 7967 12127 7973
rect 12526 7964 12532 7976
rect 12584 7964 12590 8016
rect 13906 8004 13912 8016
rect 12627 7976 13912 8004
rect 10137 7939 10195 7945
rect 10137 7905 10149 7939
rect 10183 7936 10195 7939
rect 10962 7936 10968 7948
rect 10183 7908 10968 7936
rect 10183 7905 10195 7908
rect 10137 7899 10195 7905
rect 10962 7896 10968 7908
rect 11020 7896 11026 7948
rect 11057 7939 11115 7945
rect 11057 7905 11069 7939
rect 11103 7936 11115 7939
rect 11606 7936 11612 7948
rect 11103 7908 11612 7936
rect 11103 7905 11115 7908
rect 11057 7899 11115 7905
rect 11606 7896 11612 7908
rect 11664 7896 11670 7948
rect 12627 7936 12655 7976
rect 13906 7964 13912 7976
rect 13964 7964 13970 8016
rect 14185 8007 14243 8013
rect 14185 7973 14197 8007
rect 14231 8004 14243 8007
rect 14458 8004 14464 8016
rect 14231 7976 14464 8004
rect 14231 7973 14243 7976
rect 14185 7967 14243 7973
rect 14458 7964 14464 7976
rect 14516 7964 14522 8016
rect 14660 8004 14688 8044
rect 15289 8041 15301 8075
rect 15335 8072 15347 8075
rect 15562 8072 15568 8084
rect 15335 8044 15568 8072
rect 15335 8041 15347 8044
rect 15289 8035 15347 8041
rect 15562 8032 15568 8044
rect 15620 8032 15626 8084
rect 17770 8072 17776 8084
rect 17144 8044 17776 8072
rect 15749 8007 15807 8013
rect 15749 8004 15761 8007
rect 14660 7976 15761 8004
rect 15749 7973 15761 7976
rect 15795 7973 15807 8007
rect 17144 8004 17172 8044
rect 17770 8032 17776 8044
rect 17828 8032 17834 8084
rect 17862 8032 17868 8084
rect 17920 8072 17926 8084
rect 18693 8075 18751 8081
rect 18693 8072 18705 8075
rect 17920 8044 18705 8072
rect 17920 8032 17926 8044
rect 18693 8041 18705 8044
rect 18739 8041 18751 8075
rect 18693 8035 18751 8041
rect 18966 8032 18972 8084
rect 19024 8072 19030 8084
rect 19153 8075 19211 8081
rect 19153 8072 19165 8075
rect 19024 8044 19165 8072
rect 19024 8032 19030 8044
rect 19153 8041 19165 8044
rect 19199 8041 19211 8075
rect 19153 8035 19211 8041
rect 19705 8075 19763 8081
rect 19705 8041 19717 8075
rect 19751 8072 19763 8075
rect 20162 8072 20168 8084
rect 19751 8044 20168 8072
rect 19751 8041 19763 8044
rect 19705 8035 19763 8041
rect 20162 8032 20168 8044
rect 20220 8032 20226 8084
rect 20901 8075 20959 8081
rect 20901 8041 20913 8075
rect 20947 8072 20959 8075
rect 20990 8072 20996 8084
rect 20947 8044 20996 8072
rect 20947 8041 20959 8044
rect 20901 8035 20959 8041
rect 20990 8032 20996 8044
rect 21048 8032 21054 8084
rect 17282 8007 17340 8013
rect 17282 8004 17294 8007
rect 17144 7976 17294 8004
rect 15749 7967 15807 7973
rect 17282 7973 17294 7976
rect 17328 7973 17340 8007
rect 17282 7967 17340 7973
rect 12084 7908 12655 7936
rect 13081 7939 13139 7945
rect 10318 7868 10324 7880
rect 9692 7840 10324 7868
rect 10318 7828 10324 7840
rect 10376 7828 10382 7880
rect 11333 7871 11391 7877
rect 11333 7837 11345 7871
rect 11379 7868 11391 7871
rect 11974 7868 11980 7880
rect 11379 7840 11980 7868
rect 11379 7837 11391 7840
rect 11333 7831 11391 7837
rect 11974 7828 11980 7840
rect 12032 7828 12038 7880
rect 5721 7803 5779 7809
rect 5721 7769 5733 7803
rect 5767 7769 5779 7803
rect 5721 7763 5779 7769
rect 5828 7772 8340 7800
rect 1489 7735 1547 7741
rect 1489 7701 1501 7735
rect 1535 7732 1547 7735
rect 1946 7732 1952 7744
rect 1535 7704 1952 7732
rect 1535 7701 1547 7704
rect 1489 7695 1547 7701
rect 1946 7692 1952 7704
rect 2004 7692 2010 7744
rect 2406 7692 2412 7744
rect 2464 7732 2470 7744
rect 2501 7735 2559 7741
rect 2501 7732 2513 7735
rect 2464 7704 2513 7732
rect 2464 7692 2470 7704
rect 2501 7701 2513 7704
rect 2547 7701 2559 7735
rect 2501 7695 2559 7701
rect 4062 7692 4068 7744
rect 4120 7732 4126 7744
rect 5828 7732 5856 7772
rect 4120 7704 5856 7732
rect 4120 7692 4126 7704
rect 5902 7692 5908 7744
rect 5960 7732 5966 7744
rect 6362 7732 6368 7744
rect 5960 7704 6368 7732
rect 5960 7692 5966 7704
rect 6362 7692 6368 7704
rect 6420 7692 6426 7744
rect 7374 7692 7380 7744
rect 7432 7732 7438 7744
rect 8202 7732 8208 7744
rect 7432 7704 8208 7732
rect 7432 7692 7438 7704
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 8312 7732 8340 7772
rect 10410 7760 10416 7812
rect 10468 7800 10474 7812
rect 11054 7800 11060 7812
rect 10468 7772 11060 7800
rect 10468 7760 10474 7772
rect 11054 7760 11060 7772
rect 11112 7760 11118 7812
rect 9858 7732 9864 7744
rect 8312 7704 9864 7732
rect 9858 7692 9864 7704
rect 9916 7692 9922 7744
rect 10962 7692 10968 7744
rect 11020 7732 11026 7744
rect 12084 7732 12112 7908
rect 13081 7905 13093 7939
rect 13127 7936 13139 7939
rect 13998 7936 14004 7948
rect 13127 7908 14004 7936
rect 13127 7905 13139 7908
rect 13081 7899 13139 7905
rect 13998 7896 14004 7908
rect 14056 7896 14062 7948
rect 14093 7939 14151 7945
rect 14093 7905 14105 7939
rect 14139 7936 14151 7939
rect 14139 7908 14688 7936
rect 14139 7905 14151 7908
rect 14093 7899 14151 7905
rect 12158 7828 12164 7880
rect 12216 7868 12222 7880
rect 12253 7871 12311 7877
rect 12253 7868 12265 7871
rect 12216 7840 12265 7868
rect 12216 7828 12222 7840
rect 12253 7837 12265 7840
rect 12299 7837 12311 7871
rect 12253 7831 12311 7837
rect 12434 7828 12440 7880
rect 12492 7868 12498 7880
rect 13173 7871 13231 7877
rect 13173 7868 13185 7871
rect 12492 7840 13185 7868
rect 12492 7828 12498 7840
rect 13173 7837 13185 7840
rect 13219 7837 13231 7871
rect 13173 7831 13231 7837
rect 13357 7871 13415 7877
rect 13357 7837 13369 7871
rect 13403 7868 13415 7871
rect 13722 7868 13728 7880
rect 13403 7840 13728 7868
rect 13403 7837 13415 7840
rect 13357 7831 13415 7837
rect 13722 7828 13728 7840
rect 13780 7828 13786 7880
rect 14277 7871 14335 7877
rect 14277 7837 14289 7871
rect 14323 7837 14335 7871
rect 14277 7831 14335 7837
rect 12710 7760 12716 7812
rect 12768 7800 12774 7812
rect 14292 7800 14320 7831
rect 12768 7772 14320 7800
rect 14660 7800 14688 7908
rect 15194 7896 15200 7948
rect 15252 7936 15258 7948
rect 15657 7939 15715 7945
rect 15657 7936 15669 7939
rect 15252 7908 15669 7936
rect 15252 7896 15258 7908
rect 15657 7905 15669 7908
rect 15703 7905 15715 7939
rect 15657 7899 15715 7905
rect 16390 7896 16396 7948
rect 16448 7936 16454 7948
rect 16485 7939 16543 7945
rect 16485 7936 16497 7939
rect 16448 7908 16497 7936
rect 16448 7896 16454 7908
rect 16485 7905 16497 7908
rect 16531 7905 16543 7939
rect 16485 7899 16543 7905
rect 16666 7896 16672 7948
rect 16724 7936 16730 7948
rect 17037 7939 17095 7945
rect 17037 7936 17049 7939
rect 16724 7908 17049 7936
rect 16724 7896 16730 7908
rect 17037 7905 17049 7908
rect 17083 7936 17095 7939
rect 17678 7936 17684 7948
rect 17083 7908 17684 7936
rect 17083 7905 17095 7908
rect 17037 7899 17095 7905
rect 17678 7896 17684 7908
rect 17736 7896 17742 7948
rect 17770 7896 17776 7948
rect 17828 7936 17834 7948
rect 19058 7936 19064 7948
rect 17828 7908 18644 7936
rect 19019 7908 19064 7936
rect 17828 7896 17834 7908
rect 14737 7871 14795 7877
rect 14737 7837 14749 7871
rect 14783 7868 14795 7871
rect 15562 7868 15568 7880
rect 14783 7840 15568 7868
rect 14783 7837 14795 7840
rect 14737 7831 14795 7837
rect 15562 7828 15568 7840
rect 15620 7828 15626 7880
rect 15933 7871 15991 7877
rect 15933 7837 15945 7871
rect 15979 7868 15991 7871
rect 16758 7868 16764 7880
rect 15979 7840 16764 7868
rect 15979 7837 15991 7840
rect 15933 7831 15991 7837
rect 16758 7828 16764 7840
rect 16816 7828 16822 7880
rect 18616 7868 18644 7908
rect 19058 7896 19064 7908
rect 19116 7896 19122 7948
rect 19702 7896 19708 7948
rect 19760 7936 19766 7948
rect 20073 7939 20131 7945
rect 20073 7936 20085 7939
rect 19760 7908 20085 7936
rect 19760 7896 19766 7908
rect 20073 7905 20085 7908
rect 20119 7905 20131 7939
rect 20073 7899 20131 7905
rect 19245 7871 19303 7877
rect 19245 7868 19257 7871
rect 18616 7840 19257 7868
rect 19245 7837 19257 7840
rect 19291 7868 19303 7871
rect 19334 7868 19340 7880
rect 19291 7840 19340 7868
rect 19291 7837 19303 7840
rect 19245 7831 19303 7837
rect 19334 7828 19340 7840
rect 19392 7868 19398 7880
rect 19794 7868 19800 7880
rect 19392 7840 19800 7868
rect 19392 7828 19398 7840
rect 19794 7828 19800 7840
rect 19852 7828 19858 7880
rect 19886 7828 19892 7880
rect 19944 7868 19950 7880
rect 20165 7871 20223 7877
rect 20165 7868 20177 7871
rect 19944 7840 20177 7868
rect 19944 7828 19950 7840
rect 20165 7837 20177 7840
rect 20211 7837 20223 7871
rect 20165 7831 20223 7837
rect 20257 7871 20315 7877
rect 20257 7837 20269 7871
rect 20303 7837 20315 7871
rect 20257 7831 20315 7837
rect 15654 7800 15660 7812
rect 14660 7772 15660 7800
rect 12768 7760 12774 7772
rect 15654 7760 15660 7772
rect 15712 7760 15718 7812
rect 16942 7800 16948 7812
rect 15764 7772 16948 7800
rect 11020 7704 12112 7732
rect 11020 7692 11026 7704
rect 12986 7692 12992 7744
rect 13044 7732 13050 7744
rect 13538 7732 13544 7744
rect 13044 7704 13544 7732
rect 13044 7692 13050 7704
rect 13538 7692 13544 7704
rect 13596 7692 13602 7744
rect 13722 7732 13728 7744
rect 13683 7704 13728 7732
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 13998 7692 14004 7744
rect 14056 7732 14062 7744
rect 15764 7732 15792 7772
rect 16942 7760 16948 7772
rect 17000 7760 17006 7812
rect 18230 7760 18236 7812
rect 18288 7760 18294 7812
rect 18417 7803 18475 7809
rect 18417 7769 18429 7803
rect 18463 7800 18475 7803
rect 18506 7800 18512 7812
rect 18463 7772 18512 7800
rect 18463 7769 18475 7772
rect 18417 7763 18475 7769
rect 18506 7760 18512 7772
rect 18564 7760 18570 7812
rect 18782 7760 18788 7812
rect 18840 7800 18846 7812
rect 20272 7800 20300 7831
rect 18840 7772 20300 7800
rect 18840 7760 18846 7772
rect 14056 7704 15792 7732
rect 14056 7692 14062 7704
rect 16298 7692 16304 7744
rect 16356 7732 16362 7744
rect 16574 7732 16580 7744
rect 16356 7704 16580 7732
rect 16356 7692 16362 7704
rect 16574 7692 16580 7704
rect 16632 7692 16638 7744
rect 16669 7735 16727 7741
rect 16669 7701 16681 7735
rect 16715 7732 16727 7735
rect 17678 7732 17684 7744
rect 16715 7704 17684 7732
rect 16715 7701 16727 7704
rect 16669 7695 16727 7701
rect 17678 7692 17684 7704
rect 17736 7692 17742 7744
rect 18248 7732 18276 7760
rect 19426 7732 19432 7744
rect 18248 7704 19432 7732
rect 19426 7692 19432 7704
rect 19484 7692 19490 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 4154 7528 4160 7540
rect 4115 7500 4160 7528
rect 4154 7488 4160 7500
rect 4212 7488 4218 7540
rect 4246 7488 4252 7540
rect 4304 7528 4310 7540
rect 6641 7531 6699 7537
rect 4304 7500 6408 7528
rect 4304 7488 4310 7500
rect 3881 7463 3939 7469
rect 3881 7429 3893 7463
rect 3927 7460 3939 7463
rect 3927 7432 4844 7460
rect 3927 7429 3939 7432
rect 3881 7423 3939 7429
rect 1946 7392 1952 7404
rect 1907 7364 1952 7392
rect 1946 7352 1952 7364
rect 2004 7352 2010 7404
rect 2130 7392 2136 7404
rect 2091 7364 2136 7392
rect 2130 7352 2136 7364
rect 2188 7352 2194 7404
rect 4816 7401 4844 7432
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7392 4859 7395
rect 4890 7392 4896 7404
rect 4847 7364 4896 7392
rect 4847 7361 4859 7364
rect 4801 7355 4859 7361
rect 4890 7352 4896 7364
rect 4948 7352 4954 7404
rect 5258 7352 5264 7404
rect 5316 7392 5322 7404
rect 6273 7395 6331 7401
rect 6273 7392 6285 7395
rect 5316 7364 6285 7392
rect 5316 7352 5322 7364
rect 6273 7361 6285 7364
rect 6319 7361 6331 7395
rect 6380 7392 6408 7500
rect 6641 7497 6653 7531
rect 6687 7528 6699 7531
rect 10042 7528 10048 7540
rect 6687 7500 10048 7528
rect 6687 7497 6699 7500
rect 6641 7491 6699 7497
rect 10042 7488 10048 7500
rect 10100 7528 10106 7540
rect 10962 7528 10968 7540
rect 10100 7500 10968 7528
rect 10100 7488 10106 7500
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 12434 7488 12440 7540
rect 12492 7528 12498 7540
rect 13265 7531 13323 7537
rect 12492 7500 12537 7528
rect 12492 7488 12498 7500
rect 13265 7497 13277 7531
rect 13311 7528 13323 7531
rect 13354 7528 13360 7540
rect 13311 7500 13360 7528
rect 13311 7497 13323 7500
rect 13265 7491 13323 7497
rect 13354 7488 13360 7500
rect 13412 7488 13418 7540
rect 13449 7531 13507 7537
rect 13449 7497 13461 7531
rect 13495 7497 13507 7531
rect 13449 7491 13507 7497
rect 8754 7460 8760 7472
rect 8715 7432 8760 7460
rect 8754 7420 8760 7432
rect 8812 7420 8818 7472
rect 9490 7460 9496 7472
rect 9451 7432 9496 7460
rect 9490 7420 9496 7432
rect 9548 7420 9554 7472
rect 11238 7460 11244 7472
rect 9968 7432 11244 7460
rect 7282 7392 7288 7404
rect 6380 7364 7288 7392
rect 6273 7355 6331 7361
rect 7282 7352 7288 7364
rect 7340 7392 7346 7404
rect 9398 7392 9404 7404
rect 7340 7364 7512 7392
rect 9359 7364 9404 7392
rect 7340 7352 7346 7364
rect 1857 7327 1915 7333
rect 1857 7293 1869 7327
rect 1903 7324 1915 7327
rect 2406 7324 2412 7336
rect 1903 7296 2412 7324
rect 1903 7293 1915 7296
rect 1857 7287 1915 7293
rect 2406 7284 2412 7296
rect 2464 7284 2470 7336
rect 2501 7327 2559 7333
rect 2501 7293 2513 7327
rect 2547 7324 2559 7327
rect 3694 7324 3700 7336
rect 2547 7296 3700 7324
rect 2547 7293 2559 7296
rect 2501 7287 2559 7293
rect 1578 7216 1584 7268
rect 1636 7256 1642 7268
rect 2516 7256 2544 7287
rect 3694 7284 3700 7296
rect 3752 7284 3758 7336
rect 7374 7324 7380 7336
rect 7335 7296 7380 7324
rect 7374 7284 7380 7296
rect 7432 7284 7438 7336
rect 7484 7324 7512 7364
rect 9398 7352 9404 7364
rect 9456 7392 9462 7404
rect 9968 7401 9996 7432
rect 11238 7420 11244 7432
rect 11296 7420 11302 7472
rect 13170 7460 13176 7472
rect 12176 7432 13176 7460
rect 9953 7395 10011 7401
rect 9953 7392 9965 7395
rect 9456 7364 9965 7392
rect 9456 7352 9462 7364
rect 9953 7361 9965 7364
rect 9999 7361 10011 7395
rect 9953 7355 10011 7361
rect 10137 7395 10195 7401
rect 10137 7361 10149 7395
rect 10183 7392 10195 7395
rect 10318 7392 10324 7404
rect 10183 7364 10324 7392
rect 10183 7361 10195 7364
rect 10137 7355 10195 7361
rect 10318 7352 10324 7364
rect 10376 7352 10382 7404
rect 10686 7392 10692 7404
rect 10428 7364 10692 7392
rect 9861 7327 9919 7333
rect 7484 7296 8524 7324
rect 1636 7228 2544 7256
rect 2768 7259 2826 7265
rect 1636 7216 1642 7228
rect 2768 7225 2780 7259
rect 2814 7256 2826 7259
rect 2866 7256 2872 7268
rect 2814 7228 2872 7256
rect 2814 7225 2826 7228
rect 2768 7219 2826 7225
rect 2866 7216 2872 7228
rect 2924 7216 2930 7268
rect 4525 7259 4583 7265
rect 4525 7225 4537 7259
rect 4571 7256 4583 7259
rect 4706 7256 4712 7268
rect 4571 7228 4712 7256
rect 4571 7225 4583 7228
rect 4525 7219 4583 7225
rect 4706 7216 4712 7228
rect 4764 7216 4770 7268
rect 6089 7259 6147 7265
rect 6089 7225 6101 7259
rect 6135 7256 6147 7259
rect 6270 7256 6276 7268
rect 6135 7228 6276 7256
rect 6135 7225 6147 7228
rect 6089 7219 6147 7225
rect 6270 7216 6276 7228
rect 6328 7216 6334 7268
rect 7466 7216 7472 7268
rect 7524 7256 7530 7268
rect 7622 7259 7680 7265
rect 7622 7256 7634 7259
rect 7524 7228 7634 7256
rect 7524 7216 7530 7228
rect 7622 7225 7634 7228
rect 7668 7225 7680 7259
rect 7622 7219 7680 7225
rect 1486 7188 1492 7200
rect 1447 7160 1492 7188
rect 1486 7148 1492 7160
rect 1544 7148 1550 7200
rect 4246 7148 4252 7200
rect 4304 7188 4310 7200
rect 4617 7191 4675 7197
rect 4617 7188 4629 7191
rect 4304 7160 4629 7188
rect 4304 7148 4310 7160
rect 4617 7157 4629 7160
rect 4663 7188 4675 7191
rect 5350 7188 5356 7200
rect 4663 7160 5356 7188
rect 4663 7157 4675 7160
rect 4617 7151 4675 7157
rect 5350 7148 5356 7160
rect 5408 7148 5414 7200
rect 5718 7188 5724 7200
rect 5679 7160 5724 7188
rect 5718 7148 5724 7160
rect 5776 7148 5782 7200
rect 6181 7191 6239 7197
rect 6181 7157 6193 7191
rect 6227 7188 6239 7191
rect 6641 7191 6699 7197
rect 6641 7188 6653 7191
rect 6227 7160 6653 7188
rect 6227 7157 6239 7160
rect 6181 7151 6239 7157
rect 6641 7157 6653 7160
rect 6687 7157 6699 7191
rect 8496 7188 8524 7296
rect 9861 7293 9873 7327
rect 9907 7324 9919 7327
rect 10428 7324 10456 7364
rect 10686 7352 10692 7364
rect 10744 7352 10750 7404
rect 10778 7352 10784 7404
rect 10836 7392 10842 7404
rect 11149 7395 11207 7401
rect 11149 7392 11161 7395
rect 10836 7364 11161 7392
rect 10836 7352 10842 7364
rect 11149 7361 11161 7364
rect 11195 7392 11207 7395
rect 12176 7392 12204 7432
rect 13170 7420 13176 7432
rect 13228 7420 13234 7472
rect 11195 7364 12204 7392
rect 11195 7361 11207 7364
rect 11149 7355 11207 7361
rect 12342 7352 12348 7404
rect 12400 7392 12406 7404
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 12400 7364 13001 7392
rect 12400 7352 12406 7364
rect 12989 7361 13001 7364
rect 13035 7361 13047 7395
rect 12989 7355 13047 7361
rect 13262 7352 13268 7404
rect 13320 7392 13326 7404
rect 13464 7392 13492 7491
rect 13538 7488 13544 7540
rect 13596 7528 13602 7540
rect 14185 7531 14243 7537
rect 14185 7528 14197 7531
rect 13596 7500 14197 7528
rect 13596 7488 13602 7500
rect 14185 7497 14197 7500
rect 14231 7497 14243 7531
rect 14366 7528 14372 7540
rect 14327 7500 14372 7528
rect 14185 7491 14243 7497
rect 14366 7488 14372 7500
rect 14424 7488 14430 7540
rect 14458 7488 14464 7540
rect 14516 7528 14522 7540
rect 17402 7528 17408 7540
rect 14516 7500 17408 7528
rect 14516 7488 14522 7500
rect 17402 7488 17408 7500
rect 17460 7488 17466 7540
rect 20530 7488 20536 7540
rect 20588 7528 20594 7540
rect 20717 7531 20775 7537
rect 20717 7528 20729 7531
rect 20588 7500 20729 7528
rect 20588 7488 20594 7500
rect 20717 7497 20729 7500
rect 20763 7497 20775 7531
rect 20717 7491 20775 7497
rect 13630 7420 13636 7472
rect 13688 7460 13694 7472
rect 13725 7463 13783 7469
rect 13725 7460 13737 7463
rect 13688 7432 13737 7460
rect 13688 7420 13694 7432
rect 13725 7429 13737 7432
rect 13771 7429 13783 7463
rect 13725 7423 13783 7429
rect 14001 7463 14059 7469
rect 14001 7429 14013 7463
rect 14047 7460 14059 7463
rect 15746 7460 15752 7472
rect 14047 7432 15752 7460
rect 14047 7429 14059 7432
rect 14001 7423 14059 7429
rect 15746 7420 15752 7432
rect 15804 7420 15810 7472
rect 18966 7460 18972 7472
rect 16500 7432 18972 7460
rect 14550 7392 14556 7404
rect 13320 7364 13492 7392
rect 13648 7364 14556 7392
rect 13320 7352 13326 7364
rect 9907 7296 10456 7324
rect 9907 7293 9919 7296
rect 9861 7287 9919 7293
rect 10502 7284 10508 7336
rect 10560 7324 10566 7336
rect 10965 7327 11023 7333
rect 10965 7324 10977 7327
rect 10560 7296 10977 7324
rect 10560 7284 10566 7296
rect 10965 7293 10977 7296
rect 11011 7293 11023 7327
rect 10965 7287 11023 7293
rect 11793 7327 11851 7333
rect 11793 7293 11805 7327
rect 11839 7324 11851 7327
rect 11974 7324 11980 7336
rect 11839 7296 11980 7324
rect 11839 7293 11851 7296
rect 11793 7287 11851 7293
rect 11974 7284 11980 7296
rect 12032 7284 12038 7336
rect 12805 7327 12863 7333
rect 12805 7293 12817 7327
rect 12851 7324 12863 7327
rect 13170 7324 13176 7336
rect 12851 7296 13176 7324
rect 12851 7293 12863 7296
rect 12805 7287 12863 7293
rect 13170 7284 13176 7296
rect 13228 7284 13234 7336
rect 13648 7333 13676 7364
rect 14550 7352 14556 7364
rect 14608 7352 14614 7404
rect 15013 7395 15071 7401
rect 15013 7361 15025 7395
rect 15059 7392 15071 7395
rect 15930 7392 15936 7404
rect 15059 7364 15936 7392
rect 15059 7361 15071 7364
rect 15013 7355 15071 7361
rect 15930 7352 15936 7364
rect 15988 7392 15994 7404
rect 16025 7395 16083 7401
rect 16025 7392 16037 7395
rect 15988 7364 16037 7392
rect 15988 7352 15994 7364
rect 16025 7361 16037 7364
rect 16071 7392 16083 7395
rect 16298 7392 16304 7404
rect 16071 7364 16304 7392
rect 16071 7361 16083 7364
rect 16025 7355 16083 7361
rect 16298 7352 16304 7364
rect 16356 7352 16362 7404
rect 13633 7327 13691 7333
rect 13633 7293 13645 7327
rect 13679 7293 13691 7327
rect 13633 7287 13691 7293
rect 13817 7327 13875 7333
rect 13817 7293 13829 7327
rect 13863 7293 13875 7327
rect 13817 7287 13875 7293
rect 8849 7259 8907 7265
rect 8849 7225 8861 7259
rect 8895 7256 8907 7259
rect 10873 7259 10931 7265
rect 10873 7256 10885 7259
rect 8895 7228 10885 7256
rect 8895 7225 8907 7228
rect 8849 7219 8907 7225
rect 10873 7225 10885 7228
rect 10919 7225 10931 7259
rect 10873 7219 10931 7225
rect 11238 7216 11244 7268
rect 11296 7256 11302 7268
rect 12897 7259 12955 7265
rect 11296 7228 12848 7256
rect 11296 7216 11302 7228
rect 9950 7188 9956 7200
rect 8496 7160 9956 7188
rect 6641 7151 6699 7157
rect 9950 7148 9956 7160
rect 10008 7148 10014 7200
rect 10502 7188 10508 7200
rect 10463 7160 10508 7188
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 10962 7148 10968 7200
rect 11020 7188 11026 7200
rect 11790 7188 11796 7200
rect 11020 7160 11796 7188
rect 11020 7148 11026 7160
rect 11790 7148 11796 7160
rect 11848 7148 11854 7200
rect 11977 7191 12035 7197
rect 11977 7157 11989 7191
rect 12023 7188 12035 7191
rect 12526 7188 12532 7200
rect 12023 7160 12532 7188
rect 12023 7157 12035 7160
rect 11977 7151 12035 7157
rect 12526 7148 12532 7160
rect 12584 7148 12590 7200
rect 12820 7188 12848 7228
rect 12897 7225 12909 7259
rect 12943 7256 12955 7259
rect 13265 7259 13323 7265
rect 13265 7256 13277 7259
rect 12943 7228 13277 7256
rect 12943 7225 12955 7228
rect 12897 7219 12955 7225
rect 13265 7225 13277 7228
rect 13311 7225 13323 7259
rect 13265 7219 13323 7225
rect 13725 7259 13783 7265
rect 13725 7225 13737 7259
rect 13771 7256 13783 7259
rect 13832 7256 13860 7287
rect 14090 7284 14096 7336
rect 14148 7324 14154 7336
rect 14185 7327 14243 7333
rect 14185 7324 14197 7327
rect 14148 7296 14197 7324
rect 14148 7284 14154 7296
rect 14185 7293 14197 7296
rect 14231 7293 14243 7327
rect 14185 7287 14243 7293
rect 14277 7327 14335 7333
rect 14277 7293 14289 7327
rect 14323 7324 14335 7327
rect 14829 7327 14887 7333
rect 14829 7324 14841 7327
rect 14323 7296 14841 7324
rect 14323 7293 14335 7296
rect 14277 7287 14335 7293
rect 14829 7293 14841 7296
rect 14875 7293 14887 7327
rect 14829 7287 14887 7293
rect 15286 7284 15292 7336
rect 15344 7324 15350 7336
rect 16209 7327 16267 7333
rect 16209 7324 16221 7327
rect 15344 7296 16221 7324
rect 15344 7284 15350 7296
rect 16209 7293 16221 7296
rect 16255 7293 16267 7327
rect 16209 7287 16267 7293
rect 13771 7228 13860 7256
rect 13771 7225 13783 7228
rect 13725 7219 13783 7225
rect 13906 7216 13912 7268
rect 13964 7256 13970 7268
rect 13964 7228 14780 7256
rect 13964 7216 13970 7228
rect 14090 7188 14096 7200
rect 12820 7160 14096 7188
rect 14090 7148 14096 7160
rect 14148 7148 14154 7200
rect 14185 7191 14243 7197
rect 14185 7157 14197 7191
rect 14231 7188 14243 7191
rect 14550 7188 14556 7200
rect 14231 7160 14556 7188
rect 14231 7157 14243 7160
rect 14185 7151 14243 7157
rect 14550 7148 14556 7160
rect 14608 7148 14614 7200
rect 14752 7197 14780 7228
rect 15470 7216 15476 7268
rect 15528 7256 15534 7268
rect 15841 7259 15899 7265
rect 15841 7256 15853 7259
rect 15528 7228 15853 7256
rect 15528 7216 15534 7228
rect 15841 7225 15853 7228
rect 15887 7225 15899 7259
rect 16500 7256 16528 7432
rect 18966 7420 18972 7432
rect 19024 7420 19030 7472
rect 17586 7392 17592 7404
rect 17499 7364 17592 7392
rect 17586 7352 17592 7364
rect 17644 7392 17650 7404
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 17644 7364 18613 7392
rect 17644 7352 17650 7364
rect 18601 7361 18613 7364
rect 18647 7392 18659 7395
rect 18690 7392 18696 7404
rect 18647 7364 18696 7392
rect 18647 7361 18659 7364
rect 18601 7355 18659 7361
rect 18690 7352 18696 7364
rect 18748 7352 18754 7404
rect 16850 7284 16856 7336
rect 16908 7324 16914 7336
rect 17313 7327 17371 7333
rect 17313 7324 17325 7327
rect 16908 7296 17325 7324
rect 16908 7284 16914 7296
rect 17313 7293 17325 7296
rect 17359 7293 17371 7327
rect 17313 7287 17371 7293
rect 17770 7284 17776 7336
rect 17828 7324 17834 7336
rect 18506 7324 18512 7336
rect 17828 7296 18512 7324
rect 17828 7284 17834 7296
rect 18506 7284 18512 7296
rect 18564 7284 18570 7336
rect 19242 7284 19248 7336
rect 19300 7324 19306 7336
rect 19337 7327 19395 7333
rect 19337 7324 19349 7327
rect 19300 7296 19349 7324
rect 19300 7284 19306 7296
rect 19337 7293 19349 7296
rect 19383 7293 19395 7327
rect 19337 7287 19395 7293
rect 19426 7284 19432 7336
rect 19484 7324 19490 7336
rect 19593 7327 19651 7333
rect 19593 7324 19605 7327
rect 19484 7296 19605 7324
rect 19484 7284 19490 7296
rect 19593 7293 19605 7296
rect 19639 7293 19651 7327
rect 19593 7287 19651 7293
rect 17405 7259 17463 7265
rect 17405 7256 17417 7259
rect 15841 7219 15899 7225
rect 16224 7228 16528 7256
rect 16776 7228 17417 7256
rect 14737 7191 14795 7197
rect 14737 7157 14749 7191
rect 14783 7188 14795 7191
rect 15010 7188 15016 7200
rect 14783 7160 15016 7188
rect 14783 7157 14795 7160
rect 14737 7151 14795 7157
rect 15010 7148 15016 7160
rect 15068 7148 15074 7200
rect 15378 7188 15384 7200
rect 15339 7160 15384 7188
rect 15378 7148 15384 7160
rect 15436 7148 15442 7200
rect 15749 7191 15807 7197
rect 15749 7157 15761 7191
rect 15795 7188 15807 7191
rect 16224 7188 16252 7228
rect 16776 7200 16804 7228
rect 17405 7225 17417 7228
rect 17451 7225 17463 7259
rect 17405 7219 17463 7225
rect 18417 7259 18475 7265
rect 18417 7225 18429 7259
rect 18463 7256 18475 7259
rect 19058 7256 19064 7268
rect 18463 7228 19064 7256
rect 18463 7225 18475 7228
rect 18417 7219 18475 7225
rect 19058 7216 19064 7228
rect 19116 7216 19122 7268
rect 15795 7160 16252 7188
rect 15795 7157 15807 7160
rect 15749 7151 15807 7157
rect 16298 7148 16304 7200
rect 16356 7188 16362 7200
rect 16393 7191 16451 7197
rect 16393 7188 16405 7191
rect 16356 7160 16405 7188
rect 16356 7148 16362 7160
rect 16393 7157 16405 7160
rect 16439 7157 16451 7191
rect 16758 7188 16764 7200
rect 16719 7160 16764 7188
rect 16393 7151 16451 7157
rect 16758 7148 16764 7160
rect 16816 7148 16822 7200
rect 16942 7188 16948 7200
rect 16903 7160 16948 7188
rect 16942 7148 16948 7160
rect 17000 7148 17006 7200
rect 17954 7148 17960 7200
rect 18012 7188 18018 7200
rect 18049 7191 18107 7197
rect 18049 7188 18061 7191
rect 18012 7160 18061 7188
rect 18012 7148 18018 7160
rect 18049 7157 18061 7160
rect 18095 7157 18107 7191
rect 18049 7151 18107 7157
rect 18322 7148 18328 7200
rect 18380 7188 18386 7200
rect 18509 7191 18567 7197
rect 18509 7188 18521 7191
rect 18380 7160 18521 7188
rect 18380 7148 18386 7160
rect 18509 7157 18521 7160
rect 18555 7157 18567 7191
rect 18509 7151 18567 7157
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 4890 6984 4896 6996
rect 4851 6956 4896 6984
rect 4890 6944 4896 6956
rect 4948 6944 4954 6996
rect 5902 6984 5908 6996
rect 5863 6956 5908 6984
rect 5902 6944 5908 6956
rect 5960 6944 5966 6996
rect 6086 6944 6092 6996
rect 6144 6984 6150 6996
rect 9398 6984 9404 6996
rect 6144 6956 9404 6984
rect 6144 6944 6150 6956
rect 9398 6944 9404 6956
rect 9456 6944 9462 6996
rect 9968 6956 10180 6984
rect 2406 6916 2412 6928
rect 2367 6888 2412 6916
rect 2406 6876 2412 6888
rect 2464 6876 2470 6928
rect 3970 6876 3976 6928
rect 4028 6916 4034 6928
rect 9968 6916 9996 6956
rect 4028 6888 9996 6916
rect 10152 6916 10180 6956
rect 11698 6944 11704 6996
rect 11756 6984 11762 6996
rect 12342 6984 12348 6996
rect 11756 6956 12348 6984
rect 11756 6944 11762 6956
rect 12342 6944 12348 6956
rect 12400 6944 12406 6996
rect 12526 6944 12532 6996
rect 12584 6984 12590 6996
rect 12584 6956 14320 6984
rect 12584 6944 12590 6956
rect 10870 6916 10876 6928
rect 10152 6888 10876 6916
rect 4028 6876 4034 6888
rect 10870 6876 10876 6888
rect 10928 6876 10934 6928
rect 12434 6916 12440 6928
rect 11348 6888 12440 6916
rect 3053 6851 3111 6857
rect 3053 6848 3065 6851
rect 2056 6820 3065 6848
rect 2056 6721 2084 6820
rect 3053 6817 3065 6820
rect 3099 6817 3111 6851
rect 7282 6848 7288 6860
rect 7243 6820 7288 6848
rect 3053 6811 3111 6817
rect 7282 6808 7288 6820
rect 7340 6808 7346 6860
rect 8294 6848 8300 6860
rect 8255 6820 8300 6848
rect 8294 6808 8300 6820
rect 8352 6808 8358 6860
rect 8386 6808 8392 6860
rect 8444 6848 8450 6860
rect 8444 6820 8489 6848
rect 8444 6808 8450 6820
rect 8662 6808 8668 6860
rect 8720 6848 8726 6860
rect 10042 6848 10048 6860
rect 8720 6820 9904 6848
rect 10003 6820 10048 6848
rect 8720 6808 8726 6820
rect 2501 6783 2559 6789
rect 2501 6749 2513 6783
rect 2547 6749 2559 6783
rect 2501 6743 2559 6749
rect 2685 6783 2743 6789
rect 2685 6749 2697 6783
rect 2731 6780 2743 6783
rect 2866 6780 2872 6792
rect 2731 6752 2872 6780
rect 2731 6749 2743 6752
rect 2685 6743 2743 6749
rect 2041 6715 2099 6721
rect 2041 6681 2053 6715
rect 2087 6681 2099 6715
rect 2516 6712 2544 6743
rect 2866 6740 2872 6752
rect 2924 6740 2930 6792
rect 3142 6740 3148 6792
rect 3200 6780 3206 6792
rect 3237 6783 3295 6789
rect 3237 6780 3249 6783
rect 3200 6752 3249 6780
rect 3200 6740 3206 6752
rect 3237 6749 3249 6752
rect 3283 6749 3295 6783
rect 3237 6743 3295 6749
rect 4433 6783 4491 6789
rect 4433 6749 4445 6783
rect 4479 6780 4491 6783
rect 4614 6780 4620 6792
rect 4479 6752 4620 6780
rect 4479 6749 4491 6752
rect 4433 6743 4491 6749
rect 4614 6740 4620 6752
rect 4672 6780 4678 6792
rect 4985 6783 5043 6789
rect 4985 6780 4997 6783
rect 4672 6752 4997 6780
rect 4672 6740 4678 6752
rect 4985 6749 4997 6752
rect 5031 6749 5043 6783
rect 4985 6743 5043 6749
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6780 5135 6783
rect 5258 6780 5264 6792
rect 5123 6752 5264 6780
rect 5123 6749 5135 6752
rect 5077 6743 5135 6749
rect 3510 6712 3516 6724
rect 2516 6684 3516 6712
rect 2041 6675 2099 6681
rect 3510 6672 3516 6684
rect 3568 6672 3574 6724
rect 4890 6672 4896 6724
rect 4948 6712 4954 6724
rect 5092 6712 5120 6743
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 5997 6783 6055 6789
rect 5997 6749 6009 6783
rect 6043 6780 6055 6783
rect 6086 6780 6092 6792
rect 6043 6752 6092 6780
rect 6043 6749 6055 6752
rect 5997 6743 6055 6749
rect 6086 6740 6092 6752
rect 6144 6740 6150 6792
rect 6181 6783 6239 6789
rect 6181 6749 6193 6783
rect 6227 6749 6239 6783
rect 6181 6743 6239 6749
rect 6196 6712 6224 6743
rect 6546 6740 6552 6792
rect 6604 6780 6610 6792
rect 7377 6783 7435 6789
rect 7377 6780 7389 6783
rect 6604 6752 7389 6780
rect 6604 6740 6610 6752
rect 7377 6749 7389 6752
rect 7423 6749 7435 6783
rect 7377 6743 7435 6749
rect 7561 6783 7619 6789
rect 7561 6749 7573 6783
rect 7607 6780 7619 6783
rect 7650 6780 7656 6792
rect 7607 6752 7656 6780
rect 7607 6749 7619 6752
rect 7561 6743 7619 6749
rect 7650 6740 7656 6752
rect 7708 6780 7714 6792
rect 8481 6783 8539 6789
rect 8481 6780 8493 6783
rect 7708 6752 8493 6780
rect 7708 6740 7714 6752
rect 8481 6749 8493 6752
rect 8527 6749 8539 6783
rect 8481 6743 8539 6749
rect 8754 6740 8760 6792
rect 8812 6780 8818 6792
rect 9766 6780 9772 6792
rect 8812 6752 9772 6780
rect 8812 6740 8818 6752
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 9876 6780 9904 6820
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 10137 6851 10195 6857
rect 10137 6817 10149 6851
rect 10183 6848 10195 6851
rect 10318 6848 10324 6860
rect 10183 6820 10324 6848
rect 10183 6817 10195 6820
rect 10137 6811 10195 6817
rect 10152 6780 10180 6811
rect 10318 6808 10324 6820
rect 10376 6808 10382 6860
rect 11348 6857 11376 6888
rect 12434 6876 12440 6888
rect 12492 6876 12498 6928
rect 13354 6916 13360 6928
rect 13315 6888 13360 6916
rect 13354 6876 13360 6888
rect 13412 6876 13418 6928
rect 13449 6919 13507 6925
rect 13449 6885 13461 6919
rect 13495 6916 13507 6919
rect 13722 6916 13728 6928
rect 13495 6888 13728 6916
rect 13495 6885 13507 6888
rect 13449 6879 13507 6885
rect 13722 6876 13728 6888
rect 13780 6876 13786 6928
rect 11333 6851 11391 6857
rect 11333 6817 11345 6851
rect 11379 6817 11391 6851
rect 11333 6811 11391 6817
rect 11600 6851 11658 6857
rect 11600 6817 11612 6851
rect 11646 6848 11658 6851
rect 12452 6848 12480 6876
rect 13262 6848 13268 6860
rect 11646 6820 12388 6848
rect 12452 6820 13268 6848
rect 11646 6817 11658 6820
rect 11600 6811 11658 6817
rect 9876 6752 10180 6780
rect 10229 6783 10287 6789
rect 10229 6749 10241 6783
rect 10275 6749 10287 6783
rect 10229 6743 10287 6749
rect 10873 6783 10931 6789
rect 10873 6749 10885 6783
rect 10919 6749 10931 6783
rect 12360 6780 12388 6820
rect 13262 6808 13268 6820
rect 13320 6808 13326 6860
rect 14292 6848 14320 6956
rect 14366 6944 14372 6996
rect 14424 6984 14430 6996
rect 14645 6987 14703 6993
rect 14645 6984 14657 6987
rect 14424 6956 14657 6984
rect 14424 6944 14430 6956
rect 14645 6953 14657 6956
rect 14691 6953 14703 6987
rect 14645 6947 14703 6953
rect 17586 6944 17592 6996
rect 17644 6984 17650 6996
rect 17957 6987 18015 6993
rect 17957 6984 17969 6987
rect 17644 6956 17969 6984
rect 17644 6944 17650 6956
rect 17957 6953 17969 6956
rect 18003 6953 18015 6987
rect 17957 6947 18015 6953
rect 19426 6944 19432 6996
rect 19484 6984 19490 6996
rect 20533 6987 20591 6993
rect 20533 6984 20545 6987
rect 19484 6956 20545 6984
rect 19484 6944 19490 6956
rect 20533 6953 20545 6956
rect 20579 6953 20591 6987
rect 20533 6947 20591 6953
rect 14553 6919 14611 6925
rect 14553 6885 14565 6919
rect 14599 6916 14611 6919
rect 15378 6916 15384 6928
rect 14599 6888 15384 6916
rect 14599 6885 14611 6888
rect 14553 6879 14611 6885
rect 15378 6876 15384 6888
rect 15436 6876 15442 6928
rect 15838 6876 15844 6928
rect 15896 6916 15902 6928
rect 19978 6916 19984 6928
rect 15896 6888 19984 6916
rect 15896 6876 15902 6888
rect 19978 6876 19984 6888
rect 20036 6876 20042 6928
rect 14366 6848 14372 6860
rect 14292 6820 14372 6848
rect 14366 6808 14372 6820
rect 14424 6808 14430 6860
rect 15194 6808 15200 6860
rect 15252 6848 15258 6860
rect 15749 6851 15807 6857
rect 15749 6848 15761 6851
rect 15252 6820 15761 6848
rect 15252 6808 15258 6820
rect 15749 6817 15761 6820
rect 15795 6817 15807 6851
rect 16482 6848 16488 6860
rect 15749 6811 15807 6817
rect 16040 6820 16488 6848
rect 13078 6780 13084 6792
rect 12360 6752 13084 6780
rect 10873 6743 10931 6749
rect 4948 6684 6224 6712
rect 4948 6672 4954 6684
rect 6196 6656 6224 6684
rect 9677 6715 9735 6721
rect 9677 6681 9689 6715
rect 9723 6712 9735 6715
rect 9858 6712 9864 6724
rect 9723 6684 9864 6712
rect 9723 6681 9735 6684
rect 9677 6675 9735 6681
rect 9858 6672 9864 6684
rect 9916 6672 9922 6724
rect 4525 6647 4583 6653
rect 4525 6613 4537 6647
rect 4571 6644 4583 6647
rect 5074 6644 5080 6656
rect 4571 6616 5080 6644
rect 4571 6613 4583 6616
rect 4525 6607 4583 6613
rect 5074 6604 5080 6616
rect 5132 6604 5138 6656
rect 5537 6647 5595 6653
rect 5537 6613 5549 6647
rect 5583 6644 5595 6647
rect 6086 6644 6092 6656
rect 5583 6616 6092 6644
rect 5583 6613 5595 6616
rect 5537 6607 5595 6613
rect 6086 6604 6092 6616
rect 6144 6604 6150 6656
rect 6178 6604 6184 6656
rect 6236 6604 6242 6656
rect 6730 6604 6736 6656
rect 6788 6644 6794 6656
rect 6917 6647 6975 6653
rect 6917 6644 6929 6647
rect 6788 6616 6929 6644
rect 6788 6604 6794 6616
rect 6917 6613 6929 6616
rect 6963 6613 6975 6647
rect 6917 6607 6975 6613
rect 7929 6647 7987 6653
rect 7929 6613 7941 6647
rect 7975 6644 7987 6647
rect 8294 6644 8300 6656
rect 7975 6616 8300 6644
rect 7975 6613 7987 6616
rect 7929 6607 7987 6613
rect 8294 6604 8300 6616
rect 8352 6604 8358 6656
rect 8754 6604 8760 6656
rect 8812 6644 8818 6656
rect 9306 6644 9312 6656
rect 8812 6616 9312 6644
rect 8812 6604 8818 6616
rect 9306 6604 9312 6616
rect 9364 6644 9370 6656
rect 10244 6644 10272 6743
rect 9364 6616 10272 6644
rect 10888 6644 10916 6743
rect 13078 6740 13084 6752
rect 13136 6740 13142 6792
rect 13587 6783 13645 6789
rect 13587 6749 13599 6783
rect 13633 6780 13645 6783
rect 13814 6780 13820 6792
rect 13633 6752 13820 6780
rect 13633 6749 13645 6752
rect 13587 6743 13645 6749
rect 13814 6740 13820 6752
rect 13872 6740 13878 6792
rect 14826 6780 14832 6792
rect 14787 6752 14832 6780
rect 14826 6740 14832 6752
rect 14884 6740 14890 6792
rect 16040 6789 16068 6820
rect 16482 6808 16488 6820
rect 16540 6848 16546 6860
rect 16833 6851 16891 6857
rect 16833 6848 16845 6851
rect 16540 6820 16845 6848
rect 16540 6808 16546 6820
rect 16833 6817 16845 6820
rect 16879 6817 16891 6851
rect 18506 6848 18512 6860
rect 18467 6820 18512 6848
rect 16833 6811 16891 6817
rect 18506 6808 18512 6820
rect 18564 6808 18570 6860
rect 19242 6848 19248 6860
rect 19168 6820 19248 6848
rect 15841 6783 15899 6789
rect 15841 6749 15853 6783
rect 15887 6749 15899 6783
rect 15841 6743 15899 6749
rect 16025 6783 16083 6789
rect 16025 6749 16037 6783
rect 16071 6749 16083 6783
rect 16574 6780 16580 6792
rect 16535 6752 16580 6780
rect 16025 6743 16083 6749
rect 12710 6712 12716 6724
rect 12671 6684 12716 6712
rect 12710 6672 12716 6684
rect 12768 6672 12774 6724
rect 12250 6644 12256 6656
rect 10888 6616 12256 6644
rect 9364 6604 9370 6616
rect 12250 6604 12256 6616
rect 12308 6604 12314 6656
rect 12989 6647 13047 6653
rect 12989 6613 13001 6647
rect 13035 6644 13047 6647
rect 13262 6644 13268 6656
rect 13035 6616 13268 6644
rect 13035 6613 13047 6616
rect 12989 6607 13047 6613
rect 13262 6604 13268 6616
rect 13320 6604 13326 6656
rect 14185 6647 14243 6653
rect 14185 6613 14197 6647
rect 14231 6644 14243 6647
rect 14918 6644 14924 6656
rect 14231 6616 14924 6644
rect 14231 6613 14243 6616
rect 14185 6607 14243 6613
rect 14918 6604 14924 6616
rect 14976 6604 14982 6656
rect 15378 6644 15384 6656
rect 15339 6616 15384 6644
rect 15378 6604 15384 6616
rect 15436 6604 15442 6656
rect 15856 6644 15884 6743
rect 16574 6740 16580 6752
rect 16632 6740 16638 6792
rect 18966 6740 18972 6792
rect 19024 6780 19030 6792
rect 19168 6789 19196 6820
rect 19242 6808 19248 6820
rect 19300 6808 19306 6860
rect 19420 6851 19478 6857
rect 19420 6817 19432 6851
rect 19466 6848 19478 6851
rect 20346 6848 20352 6860
rect 19466 6820 20352 6848
rect 19466 6817 19478 6820
rect 19420 6811 19478 6817
rect 20346 6808 20352 6820
rect 20404 6808 20410 6860
rect 19153 6783 19211 6789
rect 19153 6780 19165 6783
rect 19024 6752 19165 6780
rect 19024 6740 19030 6752
rect 19153 6749 19165 6752
rect 19199 6749 19211 6783
rect 19153 6743 19211 6749
rect 17586 6672 17592 6724
rect 17644 6712 17650 6724
rect 18874 6712 18880 6724
rect 17644 6684 18880 6712
rect 17644 6672 17650 6684
rect 18874 6672 18880 6684
rect 18932 6672 18938 6724
rect 20438 6672 20444 6724
rect 20496 6712 20502 6724
rect 21266 6712 21272 6724
rect 20496 6684 21272 6712
rect 20496 6672 20502 6684
rect 21266 6672 21272 6684
rect 21324 6672 21330 6724
rect 16850 6644 16856 6656
rect 15856 6616 16856 6644
rect 16850 6604 16856 6616
rect 16908 6604 16914 6656
rect 18693 6647 18751 6653
rect 18693 6613 18705 6647
rect 18739 6644 18751 6647
rect 19150 6644 19156 6656
rect 18739 6616 19156 6644
rect 18739 6613 18751 6616
rect 18693 6607 18751 6613
rect 19150 6604 19156 6616
rect 19208 6604 19214 6656
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 2866 6440 2872 6452
rect 2827 6412 2872 6440
rect 2866 6400 2872 6412
rect 2924 6400 2930 6452
rect 3510 6440 3516 6452
rect 3471 6412 3516 6440
rect 3510 6400 3516 6412
rect 3568 6400 3574 6452
rect 6178 6400 6184 6452
rect 6236 6440 6242 6452
rect 6236 6412 8616 6440
rect 6236 6400 6242 6412
rect 4614 6332 4620 6384
rect 4672 6372 4678 6384
rect 4672 6344 5212 6372
rect 4672 6332 4678 6344
rect 3142 6264 3148 6316
rect 3200 6304 3206 6316
rect 4065 6307 4123 6313
rect 4065 6304 4077 6307
rect 3200 6276 4077 6304
rect 3200 6264 3206 6276
rect 4065 6273 4077 6276
rect 4111 6273 4123 6307
rect 5074 6304 5080 6316
rect 5035 6276 5080 6304
rect 4065 6267 4123 6273
rect 5074 6264 5080 6276
rect 5132 6264 5138 6316
rect 5184 6313 5212 6344
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6273 5227 6307
rect 6086 6304 6092 6316
rect 6047 6276 6092 6304
rect 5169 6267 5227 6273
rect 6086 6264 6092 6276
rect 6144 6264 6150 6316
rect 6178 6264 6184 6316
rect 6236 6304 6242 6316
rect 6236 6276 6281 6304
rect 6236 6264 6242 6276
rect 7098 6264 7104 6316
rect 7156 6304 7162 6316
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 7156 6276 7389 6304
rect 7156 6264 7162 6276
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 7377 6267 7435 6273
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6304 7619 6307
rect 7650 6304 7656 6316
rect 7607 6276 7656 6304
rect 7607 6273 7619 6276
rect 7561 6267 7619 6273
rect 7650 6264 7656 6276
rect 7708 6264 7714 6316
rect 8588 6313 8616 6412
rect 9398 6400 9404 6452
rect 9456 6440 9462 6452
rect 10689 6443 10747 6449
rect 9456 6412 10640 6440
rect 9456 6400 9462 6412
rect 10612 6372 10640 6412
rect 10689 6409 10701 6443
rect 10735 6440 10747 6443
rect 12618 6440 12624 6452
rect 10735 6412 12624 6440
rect 10735 6409 10747 6412
rect 10689 6403 10747 6409
rect 12618 6400 12624 6412
rect 12676 6400 12682 6452
rect 13078 6400 13084 6452
rect 13136 6440 13142 6452
rect 13446 6440 13452 6452
rect 13136 6412 13452 6440
rect 13136 6400 13142 6412
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 14185 6443 14243 6449
rect 14185 6409 14197 6443
rect 14231 6440 14243 6443
rect 15194 6440 15200 6452
rect 14231 6412 15200 6440
rect 14231 6409 14243 6412
rect 14185 6403 14243 6409
rect 15194 6400 15200 6412
rect 15252 6400 15258 6452
rect 15378 6400 15384 6452
rect 15436 6440 15442 6452
rect 15436 6412 16436 6440
rect 15436 6400 15442 6412
rect 11790 6372 11796 6384
rect 10612 6344 11796 6372
rect 11790 6332 11796 6344
rect 11848 6332 11854 6384
rect 13998 6332 14004 6384
rect 14056 6372 14062 6384
rect 14642 6372 14648 6384
rect 14056 6344 14648 6372
rect 14056 6332 14062 6344
rect 14642 6332 14648 6344
rect 14700 6332 14706 6384
rect 16408 6372 16436 6412
rect 16482 6400 16488 6452
rect 16540 6440 16546 6452
rect 16577 6443 16635 6449
rect 16577 6440 16589 6443
rect 16540 6412 16589 6440
rect 16540 6400 16546 6412
rect 16577 6409 16589 6412
rect 16623 6409 16635 6443
rect 16850 6440 16856 6452
rect 16811 6412 16856 6440
rect 16577 6403 16635 6409
rect 16850 6400 16856 6412
rect 16908 6400 16914 6452
rect 17218 6400 17224 6452
rect 17276 6440 17282 6452
rect 19150 6440 19156 6452
rect 17276 6412 19156 6440
rect 17276 6400 17282 6412
rect 19150 6400 19156 6412
rect 19208 6400 19214 6452
rect 20346 6440 20352 6452
rect 20307 6412 20352 6440
rect 20346 6400 20352 6412
rect 20404 6400 20410 6452
rect 16408 6344 19012 6372
rect 8573 6307 8631 6313
rect 8573 6273 8585 6307
rect 8619 6304 8631 6307
rect 8849 6307 8907 6313
rect 8849 6304 8861 6307
rect 8619 6276 8861 6304
rect 8619 6273 8631 6276
rect 8573 6267 8631 6273
rect 8849 6273 8861 6276
rect 8895 6273 8907 6307
rect 8849 6267 8907 6273
rect 10134 6264 10140 6316
rect 10192 6304 10198 6316
rect 11149 6307 11207 6313
rect 11149 6304 11161 6307
rect 10192 6276 11161 6304
rect 10192 6264 10198 6276
rect 11149 6273 11161 6276
rect 11195 6273 11207 6307
rect 11149 6267 11207 6273
rect 11333 6307 11391 6313
rect 11333 6273 11345 6307
rect 11379 6304 11391 6307
rect 11698 6304 11704 6316
rect 11379 6276 11704 6304
rect 11379 6273 11391 6276
rect 11333 6267 11391 6273
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 1489 6239 1547 6245
rect 1489 6205 1501 6239
rect 1535 6236 1547 6239
rect 1578 6236 1584 6248
rect 1535 6208 1584 6236
rect 1535 6205 1547 6208
rect 1489 6199 1547 6205
rect 1578 6196 1584 6208
rect 1636 6196 1642 6248
rect 4985 6239 5043 6245
rect 4985 6205 4997 6239
rect 5031 6236 5043 6239
rect 5718 6236 5724 6248
rect 5031 6208 5724 6236
rect 5031 6205 5043 6208
rect 4985 6199 5043 6205
rect 5718 6196 5724 6208
rect 5776 6196 5782 6248
rect 6638 6196 6644 6248
rect 6696 6236 6702 6248
rect 8481 6239 8539 6245
rect 8481 6236 8493 6239
rect 6696 6208 8493 6236
rect 6696 6196 6702 6208
rect 8481 6205 8493 6208
rect 8527 6236 8539 6239
rect 8662 6236 8668 6248
rect 8527 6208 8668 6236
rect 8527 6205 8539 6208
rect 8481 6199 8539 6205
rect 8662 6196 8668 6208
rect 8720 6196 8726 6248
rect 9033 6239 9091 6245
rect 9033 6205 9045 6239
rect 9079 6236 9091 6239
rect 9122 6236 9128 6248
rect 9079 6208 9128 6236
rect 9079 6205 9091 6208
rect 9033 6199 9091 6205
rect 9122 6196 9128 6208
rect 9180 6196 9186 6248
rect 11808 6245 11836 6332
rect 11974 6264 11980 6316
rect 12032 6304 12038 6316
rect 12032 6276 12572 6304
rect 12032 6264 12038 6276
rect 11793 6239 11851 6245
rect 9232 6208 11744 6236
rect 1756 6171 1814 6177
rect 1756 6137 1768 6171
rect 1802 6168 1814 6171
rect 2314 6168 2320 6180
rect 1802 6140 2320 6168
rect 1802 6137 1814 6140
rect 1756 6131 1814 6137
rect 2314 6128 2320 6140
rect 2372 6128 2378 6180
rect 3881 6171 3939 6177
rect 3881 6137 3893 6171
rect 3927 6168 3939 6171
rect 5997 6171 6055 6177
rect 3927 6140 5672 6168
rect 3927 6137 3939 6140
rect 3881 6131 3939 6137
rect 5644 6109 5672 6140
rect 5997 6137 6009 6171
rect 6043 6168 6055 6171
rect 8389 6171 8447 6177
rect 6043 6140 8064 6168
rect 6043 6137 6055 6140
rect 5997 6131 6055 6137
rect 3973 6103 4031 6109
rect 3973 6069 3985 6103
rect 4019 6100 4031 6103
rect 4617 6103 4675 6109
rect 4617 6100 4629 6103
rect 4019 6072 4629 6100
rect 4019 6069 4031 6072
rect 3973 6063 4031 6069
rect 4617 6069 4629 6072
rect 4663 6069 4675 6103
rect 4617 6063 4675 6069
rect 5629 6103 5687 6109
rect 5629 6069 5641 6103
rect 5675 6069 5687 6103
rect 5629 6063 5687 6069
rect 6638 6060 6644 6112
rect 6696 6100 6702 6112
rect 6917 6103 6975 6109
rect 6917 6100 6929 6103
rect 6696 6072 6929 6100
rect 6696 6060 6702 6072
rect 6917 6069 6929 6072
rect 6963 6069 6975 6103
rect 7282 6100 7288 6112
rect 7243 6072 7288 6100
rect 6917 6063 6975 6069
rect 7282 6060 7288 6072
rect 7340 6060 7346 6112
rect 8036 6109 8064 6140
rect 8389 6137 8401 6171
rect 8435 6168 8447 6171
rect 9232 6168 9260 6208
rect 8435 6140 9260 6168
rect 9300 6171 9358 6177
rect 8435 6137 8447 6140
rect 8389 6131 8447 6137
rect 9300 6137 9312 6171
rect 9346 6168 9358 6171
rect 10870 6168 10876 6180
rect 9346 6140 10876 6168
rect 9346 6137 9358 6140
rect 9300 6131 9358 6137
rect 10870 6128 10876 6140
rect 10928 6128 10934 6180
rect 11716 6168 11744 6208
rect 11793 6205 11805 6239
rect 11839 6205 11851 6239
rect 12434 6236 12440 6248
rect 12395 6208 12440 6236
rect 11793 6199 11851 6205
rect 12434 6196 12440 6208
rect 12492 6196 12498 6248
rect 12342 6168 12348 6180
rect 11716 6140 12348 6168
rect 12342 6128 12348 6140
rect 12400 6128 12406 6180
rect 12544 6168 12572 6276
rect 14274 6264 14280 6316
rect 14332 6264 14338 6316
rect 14829 6307 14887 6313
rect 14829 6273 14841 6307
rect 14875 6304 14887 6307
rect 15194 6304 15200 6316
rect 14875 6276 15056 6304
rect 15155 6276 15200 6304
rect 14875 6273 14887 6276
rect 14829 6267 14887 6273
rect 12710 6245 12716 6248
rect 12704 6236 12716 6245
rect 12671 6208 12716 6236
rect 12704 6199 12716 6208
rect 12710 6196 12716 6199
rect 12768 6196 12774 6248
rect 12986 6196 12992 6248
rect 13044 6236 13050 6248
rect 14292 6236 14320 6264
rect 13044 6208 14320 6236
rect 13044 6196 13050 6208
rect 13630 6168 13636 6180
rect 12544 6140 13636 6168
rect 13630 6128 13636 6140
rect 13688 6128 13694 6180
rect 14274 6128 14280 6180
rect 14332 6168 14338 6180
rect 14645 6171 14703 6177
rect 14645 6168 14657 6171
rect 14332 6140 14657 6168
rect 14332 6128 14338 6140
rect 14645 6137 14657 6140
rect 14691 6137 14703 6171
rect 14645 6131 14703 6137
rect 14826 6128 14832 6180
rect 14884 6128 14890 6180
rect 15028 6168 15056 6276
rect 15194 6264 15200 6276
rect 15252 6264 15258 6316
rect 16482 6264 16488 6316
rect 16540 6304 16546 6316
rect 17405 6307 17463 6313
rect 17405 6304 17417 6307
rect 16540 6276 17417 6304
rect 16540 6264 16546 6276
rect 17405 6273 17417 6276
rect 17451 6273 17463 6307
rect 18984 6304 19012 6344
rect 20901 6307 20959 6313
rect 18984 6276 19104 6304
rect 17405 6267 17463 6273
rect 15212 6236 15240 6264
rect 16574 6236 16580 6248
rect 15212 6208 16580 6236
rect 16574 6196 16580 6208
rect 16632 6196 16638 6248
rect 16666 6196 16672 6248
rect 16724 6236 16730 6248
rect 17313 6239 17371 6245
rect 17313 6236 17325 6239
rect 16724 6208 17325 6236
rect 16724 6196 16730 6208
rect 17313 6205 17325 6208
rect 17359 6205 17371 6239
rect 17313 6199 17371 6205
rect 17586 6196 17592 6248
rect 17644 6236 17650 6248
rect 18417 6239 18475 6245
rect 18417 6236 18429 6239
rect 17644 6208 18429 6236
rect 17644 6196 17650 6208
rect 18417 6205 18429 6208
rect 18463 6205 18475 6239
rect 18966 6236 18972 6248
rect 18879 6208 18972 6236
rect 18417 6199 18475 6205
rect 18966 6196 18972 6208
rect 19024 6196 19030 6248
rect 19076 6236 19104 6276
rect 20901 6273 20913 6307
rect 20947 6304 20959 6307
rect 21082 6304 21088 6316
rect 20947 6276 21088 6304
rect 20947 6273 20959 6276
rect 20901 6267 20959 6273
rect 21082 6264 21088 6276
rect 21140 6264 21146 6316
rect 20625 6239 20683 6245
rect 20625 6236 20637 6239
rect 19076 6208 20637 6236
rect 20625 6205 20637 6208
rect 20671 6205 20683 6239
rect 20625 6199 20683 6205
rect 15464 6171 15522 6177
rect 15028 6140 15332 6168
rect 8021 6103 8079 6109
rect 8021 6069 8033 6103
rect 8067 6069 8079 6103
rect 8021 6063 8079 6069
rect 8849 6103 8907 6109
rect 8849 6069 8861 6103
rect 8895 6100 8907 6103
rect 9398 6100 9404 6112
rect 8895 6072 9404 6100
rect 8895 6069 8907 6072
rect 8849 6063 8907 6069
rect 9398 6060 9404 6072
rect 9456 6060 9462 6112
rect 9766 6060 9772 6112
rect 9824 6100 9830 6112
rect 10413 6103 10471 6109
rect 10413 6100 10425 6103
rect 9824 6072 10425 6100
rect 9824 6060 9830 6072
rect 10413 6069 10425 6072
rect 10459 6069 10471 6103
rect 10413 6063 10471 6069
rect 10962 6060 10968 6112
rect 11020 6100 11026 6112
rect 11057 6103 11115 6109
rect 11057 6100 11069 6103
rect 11020 6072 11069 6100
rect 11020 6060 11026 6072
rect 11057 6069 11069 6072
rect 11103 6069 11115 6103
rect 11057 6063 11115 6069
rect 11977 6103 12035 6109
rect 11977 6069 11989 6103
rect 12023 6100 12035 6103
rect 13078 6100 13084 6112
rect 12023 6072 13084 6100
rect 12023 6069 12035 6072
rect 11977 6063 12035 6069
rect 13078 6060 13084 6072
rect 13136 6060 13142 6112
rect 13814 6100 13820 6112
rect 13775 6072 13820 6100
rect 13814 6060 13820 6072
rect 13872 6060 13878 6112
rect 14550 6100 14556 6112
rect 14511 6072 14556 6100
rect 14550 6060 14556 6072
rect 14608 6060 14614 6112
rect 14844 6100 14872 6128
rect 15194 6100 15200 6112
rect 14844 6072 15200 6100
rect 15194 6060 15200 6072
rect 15252 6060 15258 6112
rect 15304 6100 15332 6140
rect 15464 6137 15476 6171
rect 15510 6168 15522 6171
rect 16482 6168 16488 6180
rect 15510 6140 16488 6168
rect 15510 6137 15522 6140
rect 15464 6131 15522 6137
rect 15479 6100 15507 6131
rect 16482 6128 16488 6140
rect 16540 6128 16546 6180
rect 16592 6168 16620 6196
rect 18984 6168 19012 6196
rect 16592 6140 19012 6168
rect 19236 6171 19294 6177
rect 19236 6137 19248 6171
rect 19282 6168 19294 6171
rect 19334 6168 19340 6180
rect 19282 6140 19340 6168
rect 19282 6137 19294 6140
rect 19236 6131 19294 6137
rect 19334 6128 19340 6140
rect 19392 6128 19398 6180
rect 15304 6072 15507 6100
rect 16666 6060 16672 6112
rect 16724 6100 16730 6112
rect 17221 6103 17279 6109
rect 17221 6100 17233 6103
rect 16724 6072 17233 6100
rect 16724 6060 16730 6072
rect 17221 6069 17233 6072
rect 17267 6069 17279 6103
rect 17221 6063 17279 6069
rect 18601 6103 18659 6109
rect 18601 6069 18613 6103
rect 18647 6100 18659 6103
rect 20990 6100 20996 6112
rect 18647 6072 20996 6100
rect 18647 6069 18659 6072
rect 18601 6063 18659 6069
rect 20990 6060 20996 6072
rect 21048 6060 21054 6112
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 2314 5856 2320 5908
rect 2372 5896 2378 5908
rect 3142 5896 3148 5908
rect 2372 5868 3148 5896
rect 2372 5856 2378 5868
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 3694 5856 3700 5908
rect 3752 5896 3758 5908
rect 4614 5896 4620 5908
rect 3752 5868 4620 5896
rect 3752 5856 3758 5868
rect 4614 5856 4620 5868
rect 4672 5896 4678 5908
rect 5445 5899 5503 5905
rect 5445 5896 5457 5899
rect 4672 5868 5457 5896
rect 4672 5856 4678 5868
rect 5445 5865 5457 5868
rect 5491 5896 5503 5899
rect 6178 5896 6184 5908
rect 5491 5868 6184 5896
rect 5491 5865 5503 5868
rect 5445 5859 5503 5865
rect 6178 5856 6184 5868
rect 6236 5856 6242 5908
rect 6638 5896 6644 5908
rect 6599 5868 6644 5896
rect 6638 5856 6644 5868
rect 6696 5856 6702 5908
rect 6730 5856 6736 5908
rect 6788 5896 6794 5908
rect 6788 5868 6833 5896
rect 6788 5856 6794 5868
rect 7282 5856 7288 5908
rect 7340 5896 7346 5908
rect 8941 5899 8999 5905
rect 8941 5896 8953 5899
rect 7340 5868 8953 5896
rect 7340 5856 7346 5868
rect 8941 5865 8953 5868
rect 8987 5865 8999 5899
rect 8941 5859 8999 5865
rect 9306 5856 9312 5908
rect 9364 5896 9370 5908
rect 11514 5896 11520 5908
rect 9364 5868 11520 5896
rect 9364 5856 9370 5868
rect 11514 5856 11520 5868
rect 11572 5856 11578 5908
rect 11793 5899 11851 5905
rect 11793 5865 11805 5899
rect 11839 5896 11851 5899
rect 14458 5896 14464 5908
rect 11839 5868 14464 5896
rect 11839 5865 11851 5868
rect 11793 5859 11851 5865
rect 14458 5856 14464 5868
rect 14516 5856 14522 5908
rect 16482 5856 16488 5908
rect 16540 5896 16546 5908
rect 16669 5899 16727 5905
rect 16669 5896 16681 5899
rect 16540 5868 16681 5896
rect 16540 5856 16546 5868
rect 16669 5865 16681 5868
rect 16715 5865 16727 5899
rect 16669 5859 16727 5865
rect 16945 5899 17003 5905
rect 16945 5865 16957 5899
rect 16991 5896 17003 5899
rect 18417 5899 18475 5905
rect 18417 5896 18429 5899
rect 16991 5868 18429 5896
rect 16991 5865 17003 5868
rect 16945 5859 17003 5865
rect 18417 5865 18429 5868
rect 18463 5865 18475 5899
rect 18417 5859 18475 5865
rect 19153 5899 19211 5905
rect 19153 5865 19165 5899
rect 19199 5896 19211 5899
rect 20714 5896 20720 5908
rect 19199 5868 20720 5896
rect 19199 5865 19211 5868
rect 19153 5859 19211 5865
rect 20714 5856 20720 5868
rect 20772 5856 20778 5908
rect 2032 5831 2090 5837
rect 2032 5797 2044 5831
rect 2078 5828 2090 5831
rect 2682 5828 2688 5840
rect 2078 5800 2688 5828
rect 2078 5797 2090 5800
rect 2032 5791 2090 5797
rect 2682 5788 2688 5800
rect 2740 5788 2746 5840
rect 4062 5788 4068 5840
rect 4120 5828 4126 5840
rect 7190 5828 7196 5840
rect 4120 5800 7196 5828
rect 4120 5788 4126 5800
rect 7190 5788 7196 5800
rect 7248 5788 7254 5840
rect 7374 5828 7380 5840
rect 7287 5800 7380 5828
rect 1578 5720 1584 5772
rect 1636 5760 1642 5772
rect 1765 5763 1823 5769
rect 1765 5760 1777 5763
rect 1636 5732 1777 5760
rect 1636 5720 1642 5732
rect 1765 5729 1777 5732
rect 1811 5760 1823 5763
rect 4332 5763 4390 5769
rect 1811 5732 4108 5760
rect 1811 5729 1823 5732
rect 1765 5723 1823 5729
rect 4080 5704 4108 5732
rect 4332 5729 4344 5763
rect 4378 5760 4390 5763
rect 4890 5760 4896 5772
rect 4378 5732 4896 5760
rect 4378 5729 4390 5732
rect 4332 5723 4390 5729
rect 4890 5720 4896 5732
rect 4948 5720 4954 5772
rect 5810 5720 5816 5772
rect 5868 5760 5874 5772
rect 7006 5760 7012 5772
rect 5868 5732 7012 5760
rect 5868 5720 5874 5732
rect 7006 5720 7012 5732
rect 7064 5720 7070 5772
rect 7300 5769 7328 5800
rect 7374 5788 7380 5800
rect 7432 5828 7438 5840
rect 8478 5828 8484 5840
rect 7432 5800 8484 5828
rect 7432 5788 7438 5800
rect 8478 5788 8484 5800
rect 8536 5788 8542 5840
rect 10686 5788 10692 5840
rect 10744 5828 10750 5840
rect 11701 5831 11759 5837
rect 11701 5828 11713 5831
rect 10744 5800 11713 5828
rect 10744 5788 10750 5800
rect 11701 5797 11713 5800
rect 11747 5797 11759 5831
rect 11701 5791 11759 5797
rect 12612 5831 12670 5837
rect 12612 5797 12624 5831
rect 12658 5828 12670 5831
rect 13814 5828 13820 5840
rect 12658 5800 13820 5828
rect 12658 5797 12670 5800
rect 12612 5791 12670 5797
rect 13814 5788 13820 5800
rect 13872 5788 13878 5840
rect 14093 5831 14151 5837
rect 14093 5797 14105 5831
rect 14139 5828 14151 5831
rect 14139 5800 14320 5828
rect 14139 5797 14151 5800
rect 14093 5791 14151 5797
rect 7285 5763 7343 5769
rect 7285 5729 7297 5763
rect 7331 5729 7343 5763
rect 7285 5723 7343 5729
rect 7552 5763 7610 5769
rect 7552 5729 7564 5763
rect 7598 5760 7610 5763
rect 9766 5760 9772 5772
rect 7598 5732 9772 5760
rect 7598 5729 7610 5732
rect 7552 5723 7610 5729
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 9944 5763 10002 5769
rect 9944 5729 9956 5763
rect 9990 5760 10002 5763
rect 12345 5763 12403 5769
rect 9990 5732 10824 5760
rect 9990 5729 10002 5732
rect 9944 5723 10002 5729
rect 10796 5704 10824 5732
rect 12345 5729 12357 5763
rect 12391 5760 12403 5763
rect 12434 5760 12440 5772
rect 12391 5732 12440 5760
rect 12391 5729 12403 5732
rect 12345 5723 12403 5729
rect 12434 5720 12440 5732
rect 12492 5720 12498 5772
rect 14292 5760 14320 5800
rect 15194 5788 15200 5840
rect 15252 5828 15258 5840
rect 15534 5831 15592 5837
rect 15534 5828 15546 5831
rect 15252 5800 15546 5828
rect 15252 5788 15258 5800
rect 15534 5797 15546 5800
rect 15580 5797 15592 5831
rect 15534 5791 15592 5797
rect 17313 5831 17371 5837
rect 17313 5797 17325 5831
rect 17359 5828 17371 5831
rect 17954 5828 17960 5840
rect 17359 5800 17960 5828
rect 17359 5797 17371 5800
rect 17313 5791 17371 5797
rect 17954 5788 17960 5800
rect 18012 5788 18018 5840
rect 14458 5760 14464 5772
rect 14292 5732 14464 5760
rect 14458 5720 14464 5732
rect 14516 5760 14522 5772
rect 14553 5763 14611 5769
rect 14553 5760 14565 5763
rect 14516 5732 14565 5760
rect 14516 5720 14522 5732
rect 14553 5729 14565 5732
rect 14599 5729 14611 5763
rect 14553 5723 14611 5729
rect 14645 5763 14703 5769
rect 14645 5729 14657 5763
rect 14691 5760 14703 5763
rect 15010 5760 15016 5772
rect 14691 5732 15016 5760
rect 14691 5729 14703 5732
rect 14645 5723 14703 5729
rect 15010 5720 15016 5732
rect 15068 5720 15074 5772
rect 15289 5763 15347 5769
rect 15289 5729 15301 5763
rect 15335 5760 15347 5763
rect 15378 5760 15384 5772
rect 15335 5732 15384 5760
rect 15335 5729 15347 5732
rect 15289 5723 15347 5729
rect 15378 5720 15384 5732
rect 15436 5720 15442 5772
rect 16942 5720 16948 5772
rect 17000 5760 17006 5772
rect 17405 5763 17463 5769
rect 17405 5760 17417 5763
rect 17000 5732 17417 5760
rect 17000 5720 17006 5732
rect 17405 5729 17417 5732
rect 17451 5729 17463 5763
rect 17405 5723 17463 5729
rect 18046 5720 18052 5772
rect 18104 5760 18110 5772
rect 18325 5763 18383 5769
rect 18325 5760 18337 5763
rect 18104 5732 18337 5760
rect 18104 5720 18110 5732
rect 18325 5729 18337 5732
rect 18371 5729 18383 5763
rect 18325 5723 18383 5729
rect 18874 5720 18880 5772
rect 18932 5760 18938 5772
rect 18969 5763 19027 5769
rect 18969 5760 18981 5763
rect 18932 5732 18981 5760
rect 18932 5720 18938 5732
rect 18969 5729 18981 5732
rect 19015 5729 19027 5763
rect 19886 5760 19892 5772
rect 19847 5732 19892 5760
rect 18969 5723 19027 5729
rect 19886 5720 19892 5732
rect 19944 5720 19950 5772
rect 2774 5652 2780 5704
rect 2832 5692 2838 5704
rect 3421 5695 3479 5701
rect 3421 5692 3433 5695
rect 2832 5664 3433 5692
rect 2832 5652 2838 5664
rect 3421 5661 3433 5664
rect 3467 5661 3479 5695
rect 4062 5692 4068 5704
rect 4023 5664 4068 5692
rect 3421 5655 3479 5661
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 6822 5692 6828 5704
rect 6783 5664 6828 5692
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 8478 5652 8484 5704
rect 8536 5692 8542 5704
rect 9122 5692 9128 5704
rect 8536 5664 9128 5692
rect 8536 5652 8542 5664
rect 9122 5652 9128 5664
rect 9180 5692 9186 5704
rect 9677 5695 9735 5701
rect 9677 5692 9689 5695
rect 9180 5664 9689 5692
rect 9180 5652 9186 5664
rect 9677 5661 9689 5664
rect 9723 5661 9735 5695
rect 9677 5655 9735 5661
rect 10778 5652 10784 5704
rect 10836 5692 10842 5704
rect 11790 5692 11796 5704
rect 10836 5664 11796 5692
rect 10836 5652 10842 5664
rect 11790 5652 11796 5664
rect 11848 5692 11854 5704
rect 11885 5695 11943 5701
rect 11885 5692 11897 5695
rect 11848 5664 11897 5692
rect 11848 5652 11854 5664
rect 11885 5661 11897 5664
rect 11931 5661 11943 5695
rect 14737 5695 14795 5701
rect 14737 5692 14749 5695
rect 11885 5655 11943 5661
rect 13740 5664 14749 5692
rect 8665 5627 8723 5633
rect 6012 5596 7328 5624
rect 3418 5516 3424 5568
rect 3476 5556 3482 5568
rect 6012 5556 6040 5596
rect 3476 5528 6040 5556
rect 3476 5516 3482 5528
rect 6086 5516 6092 5568
rect 6144 5556 6150 5568
rect 6273 5559 6331 5565
rect 6273 5556 6285 5559
rect 6144 5528 6285 5556
rect 6144 5516 6150 5528
rect 6273 5525 6285 5528
rect 6319 5525 6331 5559
rect 7300 5556 7328 5596
rect 8665 5593 8677 5627
rect 8711 5624 8723 5627
rect 9398 5624 9404 5636
rect 8711 5596 9404 5624
rect 8711 5593 8723 5596
rect 8665 5587 8723 5593
rect 9398 5584 9404 5596
rect 9456 5584 9462 5636
rect 10962 5584 10968 5636
rect 11020 5624 11026 5636
rect 11333 5627 11391 5633
rect 11333 5624 11345 5627
rect 11020 5596 11345 5624
rect 11020 5584 11026 5596
rect 11333 5593 11345 5596
rect 11379 5593 11391 5627
rect 11333 5587 11391 5593
rect 13740 5568 13768 5664
rect 14737 5661 14749 5664
rect 14783 5661 14795 5695
rect 14737 5655 14795 5661
rect 17310 5652 17316 5704
rect 17368 5692 17374 5704
rect 17497 5695 17555 5701
rect 17497 5692 17509 5695
rect 17368 5664 17509 5692
rect 17368 5652 17374 5664
rect 17497 5661 17509 5664
rect 17543 5661 17555 5695
rect 17497 5655 17555 5661
rect 18601 5695 18659 5701
rect 18601 5661 18613 5695
rect 18647 5692 18659 5695
rect 19334 5692 19340 5704
rect 18647 5664 19340 5692
rect 18647 5661 18659 5664
rect 18601 5655 18659 5661
rect 19334 5652 19340 5664
rect 19392 5652 19398 5704
rect 19981 5695 20039 5701
rect 19981 5661 19993 5695
rect 20027 5661 20039 5695
rect 19981 5655 20039 5661
rect 20165 5695 20223 5701
rect 20165 5661 20177 5695
rect 20211 5692 20223 5695
rect 20346 5692 20352 5704
rect 20211 5664 20352 5692
rect 20211 5661 20223 5664
rect 20165 5655 20223 5661
rect 13814 5584 13820 5636
rect 13872 5624 13878 5636
rect 14185 5627 14243 5633
rect 14185 5624 14197 5627
rect 13872 5596 14197 5624
rect 13872 5584 13878 5596
rect 14185 5593 14197 5596
rect 14231 5593 14243 5627
rect 14185 5587 14243 5593
rect 17957 5627 18015 5633
rect 17957 5593 17969 5627
rect 18003 5624 18015 5627
rect 19996 5624 20024 5655
rect 20346 5652 20352 5664
rect 20404 5652 20410 5704
rect 18003 5596 20024 5624
rect 18003 5593 18015 5596
rect 17957 5587 18015 5593
rect 8202 5556 8208 5568
rect 7300 5528 8208 5556
rect 6273 5519 6331 5525
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 8938 5516 8944 5568
rect 8996 5556 9002 5568
rect 10778 5556 10784 5568
rect 8996 5528 10784 5556
rect 8996 5516 9002 5528
rect 10778 5516 10784 5528
rect 10836 5516 10842 5568
rect 10870 5516 10876 5568
rect 10928 5556 10934 5568
rect 11057 5559 11115 5565
rect 11057 5556 11069 5559
rect 10928 5528 11069 5556
rect 10928 5516 10934 5528
rect 11057 5525 11069 5528
rect 11103 5525 11115 5559
rect 11057 5519 11115 5525
rect 11974 5516 11980 5568
rect 12032 5556 12038 5568
rect 13538 5556 13544 5568
rect 12032 5528 13544 5556
rect 12032 5516 12038 5528
rect 13538 5516 13544 5528
rect 13596 5516 13602 5568
rect 13722 5556 13728 5568
rect 13683 5528 13728 5556
rect 13722 5516 13728 5528
rect 13780 5516 13786 5568
rect 14090 5516 14096 5568
rect 14148 5556 14154 5568
rect 18782 5556 18788 5568
rect 14148 5528 18788 5556
rect 14148 5516 14154 5528
rect 18782 5516 18788 5528
rect 18840 5516 18846 5568
rect 19150 5516 19156 5568
rect 19208 5556 19214 5568
rect 19521 5559 19579 5565
rect 19521 5556 19533 5559
rect 19208 5528 19533 5556
rect 19208 5516 19214 5528
rect 19521 5525 19533 5528
rect 19567 5525 19579 5559
rect 19521 5519 19579 5525
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 2041 5355 2099 5361
rect 2041 5321 2053 5355
rect 2087 5352 2099 5355
rect 2406 5352 2412 5364
rect 2087 5324 2412 5352
rect 2087 5321 2099 5324
rect 2041 5315 2099 5321
rect 2406 5312 2412 5324
rect 2464 5312 2470 5364
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 12342 5352 12348 5364
rect 4120 5324 12348 5352
rect 4120 5312 4126 5324
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 12437 5355 12495 5361
rect 12437 5321 12449 5355
rect 12483 5352 12495 5355
rect 13354 5352 13360 5364
rect 12483 5324 13360 5352
rect 12483 5321 12495 5324
rect 12437 5315 12495 5321
rect 13354 5312 13360 5324
rect 13412 5312 13418 5364
rect 14274 5352 14280 5364
rect 14235 5324 14280 5352
rect 14274 5312 14280 5324
rect 14332 5312 14338 5364
rect 14550 5312 14556 5364
rect 14608 5352 14614 5364
rect 15289 5355 15347 5361
rect 15289 5352 15301 5355
rect 14608 5324 15301 5352
rect 14608 5312 14614 5324
rect 15289 5321 15301 5324
rect 15335 5321 15347 5355
rect 15289 5315 15347 5321
rect 16945 5355 17003 5361
rect 16945 5321 16957 5355
rect 16991 5352 17003 5355
rect 17954 5352 17960 5364
rect 16991 5324 17960 5352
rect 16991 5321 17003 5324
rect 16945 5315 17003 5321
rect 17954 5312 17960 5324
rect 18012 5312 18018 5364
rect 18049 5355 18107 5361
rect 18049 5321 18061 5355
rect 18095 5352 18107 5355
rect 19245 5355 19303 5361
rect 19245 5352 19257 5355
rect 18095 5324 19257 5352
rect 18095 5321 18107 5324
rect 18049 5315 18107 5321
rect 19245 5321 19257 5324
rect 19291 5321 19303 5355
rect 19245 5315 19303 5321
rect 19334 5312 19340 5364
rect 19392 5352 19398 5364
rect 20254 5352 20260 5364
rect 19392 5324 20260 5352
rect 19392 5312 19398 5324
rect 20254 5312 20260 5324
rect 20312 5352 20318 5364
rect 20717 5355 20775 5361
rect 20717 5352 20729 5355
rect 20312 5324 20729 5352
rect 20312 5312 20318 5324
rect 20717 5321 20729 5324
rect 20763 5321 20775 5355
rect 20717 5315 20775 5321
rect 6825 5287 6883 5293
rect 6825 5253 6837 5287
rect 6871 5284 6883 5287
rect 9585 5287 9643 5293
rect 6871 5256 9536 5284
rect 6871 5253 6883 5256
rect 6825 5247 6883 5253
rect 2314 5176 2320 5228
rect 2372 5216 2378 5228
rect 2593 5219 2651 5225
rect 2593 5216 2605 5219
rect 2372 5188 2605 5216
rect 2372 5176 2378 5188
rect 2593 5185 2605 5188
rect 2639 5185 2651 5219
rect 3694 5216 3700 5228
rect 2593 5179 2651 5185
rect 2792 5188 3700 5216
rect 2682 5108 2688 5160
rect 2740 5148 2746 5160
rect 2792 5148 2820 5188
rect 3694 5176 3700 5188
rect 3752 5176 3758 5228
rect 7466 5216 7472 5228
rect 7427 5188 7472 5216
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 7650 5176 7656 5228
rect 7708 5216 7714 5228
rect 8757 5219 8815 5225
rect 8757 5216 8769 5219
rect 7708 5188 8769 5216
rect 7708 5176 7714 5188
rect 8757 5185 8769 5188
rect 8803 5216 8815 5219
rect 8938 5216 8944 5228
rect 8803 5188 8944 5216
rect 8803 5185 8815 5188
rect 8757 5179 8815 5185
rect 8938 5176 8944 5188
rect 8996 5176 9002 5228
rect 9508 5216 9536 5256
rect 9585 5253 9597 5287
rect 9631 5284 9643 5287
rect 11790 5284 11796 5296
rect 9631 5256 11796 5284
rect 9631 5253 9643 5256
rect 9585 5247 9643 5253
rect 11790 5244 11796 5256
rect 11848 5244 11854 5296
rect 12253 5287 12311 5293
rect 12253 5253 12265 5287
rect 12299 5284 12311 5287
rect 14090 5284 14096 5296
rect 12299 5256 14096 5284
rect 12299 5253 12311 5256
rect 12253 5247 12311 5253
rect 14090 5244 14096 5256
rect 14148 5244 14154 5296
rect 14182 5244 14188 5296
rect 14240 5284 14246 5296
rect 18874 5284 18880 5296
rect 14240 5256 18880 5284
rect 14240 5244 14246 5256
rect 18874 5244 18880 5256
rect 18932 5244 18938 5296
rect 9674 5216 9680 5228
rect 9508 5188 9680 5216
rect 9674 5176 9680 5188
rect 9732 5176 9738 5228
rect 9766 5176 9772 5228
rect 9824 5216 9830 5228
rect 10137 5219 10195 5225
rect 10137 5216 10149 5219
rect 9824 5188 10149 5216
rect 9824 5176 9830 5188
rect 10137 5185 10149 5188
rect 10183 5185 10195 5219
rect 10137 5179 10195 5185
rect 10870 5176 10876 5228
rect 10928 5216 10934 5228
rect 11054 5216 11060 5228
rect 10928 5188 11060 5216
rect 10928 5176 10934 5188
rect 11054 5176 11060 5188
rect 11112 5216 11118 5228
rect 11149 5219 11207 5225
rect 11149 5216 11161 5219
rect 11112 5188 11161 5216
rect 11112 5176 11118 5188
rect 11149 5185 11161 5188
rect 11195 5185 11207 5219
rect 11149 5179 11207 5185
rect 11885 5219 11943 5225
rect 11885 5185 11897 5219
rect 11931 5216 11943 5219
rect 11974 5216 11980 5228
rect 11931 5188 11980 5216
rect 11931 5185 11943 5188
rect 11885 5179 11943 5185
rect 11974 5176 11980 5188
rect 12032 5176 12038 5228
rect 12710 5176 12716 5228
rect 12768 5216 12774 5228
rect 12989 5219 13047 5225
rect 12989 5216 13001 5219
rect 12768 5188 13001 5216
rect 12768 5176 12774 5188
rect 12989 5185 13001 5188
rect 13035 5185 13047 5219
rect 13630 5216 13636 5228
rect 13591 5188 13636 5216
rect 12989 5179 13047 5185
rect 13630 5176 13636 5188
rect 13688 5176 13694 5228
rect 14921 5219 14979 5225
rect 14921 5185 14933 5219
rect 14967 5216 14979 5219
rect 15194 5216 15200 5228
rect 14967 5188 15200 5216
rect 14967 5185 14979 5188
rect 14921 5179 14979 5185
rect 15194 5176 15200 5188
rect 15252 5216 15258 5228
rect 15838 5216 15844 5228
rect 15252 5188 15844 5216
rect 15252 5176 15258 5188
rect 15838 5176 15844 5188
rect 15896 5176 15902 5228
rect 17310 5176 17316 5228
rect 17368 5216 17374 5228
rect 17497 5219 17555 5225
rect 17497 5216 17509 5219
rect 17368 5188 17509 5216
rect 17368 5176 17374 5188
rect 17497 5185 17509 5188
rect 17543 5185 17555 5219
rect 17497 5179 17555 5185
rect 18601 5219 18659 5225
rect 18601 5185 18613 5219
rect 18647 5185 18659 5219
rect 18601 5179 18659 5185
rect 2740 5120 2820 5148
rect 2740 5108 2746 5120
rect 4154 5108 4160 5160
rect 4212 5148 4218 5160
rect 4341 5151 4399 5157
rect 4341 5148 4353 5151
rect 4212 5120 4353 5148
rect 4212 5108 4218 5120
rect 4341 5117 4353 5120
rect 4387 5117 4399 5151
rect 4341 5111 4399 5117
rect 4608 5151 4666 5157
rect 4608 5117 4620 5151
rect 4654 5148 4666 5151
rect 5442 5148 5448 5160
rect 4654 5120 5448 5148
rect 4654 5117 4666 5120
rect 4608 5111 4666 5117
rect 4356 5080 4384 5111
rect 5442 5108 5448 5120
rect 5500 5108 5506 5160
rect 8202 5108 8208 5160
rect 8260 5148 8266 5160
rect 8481 5151 8539 5157
rect 8481 5148 8493 5151
rect 8260 5120 8493 5148
rect 8260 5108 8266 5120
rect 8481 5117 8493 5120
rect 8527 5148 8539 5151
rect 9306 5148 9312 5160
rect 8527 5120 9312 5148
rect 8527 5117 8539 5120
rect 8481 5111 8539 5117
rect 9306 5108 9312 5120
rect 9364 5108 9370 5160
rect 9398 5108 9404 5160
rect 9456 5148 9462 5160
rect 10962 5148 10968 5160
rect 9456 5120 10824 5148
rect 10923 5120 10968 5148
rect 9456 5108 9462 5120
rect 5810 5080 5816 5092
rect 4356 5052 5816 5080
rect 5810 5040 5816 5052
rect 5868 5040 5874 5092
rect 7006 5040 7012 5092
rect 7064 5080 7070 5092
rect 8573 5083 8631 5089
rect 7064 5052 8524 5080
rect 7064 5040 7070 5052
rect 2406 5012 2412 5024
rect 2367 4984 2412 5012
rect 2406 4972 2412 4984
rect 2464 4972 2470 5024
rect 2501 5015 2559 5021
rect 2501 4981 2513 5015
rect 2547 5012 2559 5015
rect 3053 5015 3111 5021
rect 3053 5012 3065 5015
rect 2547 4984 3065 5012
rect 2547 4981 2559 4984
rect 2501 4975 2559 4981
rect 3053 4981 3065 4984
rect 3099 4981 3111 5015
rect 3053 4975 3111 4981
rect 3234 4972 3240 5024
rect 3292 5012 3298 5024
rect 3421 5015 3479 5021
rect 3421 5012 3433 5015
rect 3292 4984 3433 5012
rect 3292 4972 3298 4984
rect 3421 4981 3433 4984
rect 3467 4981 3479 5015
rect 3421 4975 3479 4981
rect 3510 4972 3516 5024
rect 3568 5012 3574 5024
rect 5718 5012 5724 5024
rect 3568 4984 3613 5012
rect 5679 4984 5724 5012
rect 3568 4972 3574 4984
rect 5718 4972 5724 4984
rect 5776 4972 5782 5024
rect 7190 5012 7196 5024
rect 7151 4984 7196 5012
rect 7190 4972 7196 4984
rect 7248 4972 7254 5024
rect 7282 4972 7288 5024
rect 7340 5012 7346 5024
rect 8113 5015 8171 5021
rect 7340 4984 7385 5012
rect 7340 4972 7346 4984
rect 8113 4981 8125 5015
rect 8159 5012 8171 5015
rect 8386 5012 8392 5024
rect 8159 4984 8392 5012
rect 8159 4981 8171 4984
rect 8113 4975 8171 4981
rect 8386 4972 8392 4984
rect 8444 4972 8450 5024
rect 8496 5012 8524 5052
rect 8573 5049 8585 5083
rect 8619 5080 8631 5083
rect 10134 5080 10140 5092
rect 8619 5052 10140 5080
rect 8619 5049 8631 5052
rect 8573 5043 8631 5049
rect 10134 5040 10140 5052
rect 10192 5040 10198 5092
rect 9122 5012 9128 5024
rect 8496 4984 9128 5012
rect 9122 4972 9128 4984
rect 9180 4972 9186 5024
rect 9674 4972 9680 5024
rect 9732 5012 9738 5024
rect 9953 5015 10011 5021
rect 9953 5012 9965 5015
rect 9732 4984 9965 5012
rect 9732 4972 9738 4984
rect 9953 4981 9965 4984
rect 9999 4981 10011 5015
rect 9953 4975 10011 4981
rect 10045 5015 10103 5021
rect 10045 4981 10057 5015
rect 10091 5012 10103 5015
rect 10597 5015 10655 5021
rect 10597 5012 10609 5015
rect 10091 4984 10609 5012
rect 10091 4981 10103 4984
rect 10045 4975 10103 4981
rect 10597 4981 10609 4984
rect 10643 4981 10655 5015
rect 10796 5012 10824 5120
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 11609 5151 11667 5157
rect 11609 5117 11621 5151
rect 11655 5148 11667 5151
rect 12434 5148 12440 5160
rect 11655 5120 12440 5148
rect 11655 5117 11667 5120
rect 11609 5111 11667 5117
rect 12434 5108 12440 5120
rect 12492 5108 12498 5160
rect 13449 5151 13507 5157
rect 13449 5117 13461 5151
rect 13495 5148 13507 5151
rect 13998 5148 14004 5160
rect 13495 5120 14004 5148
rect 13495 5117 13507 5120
rect 13449 5111 13507 5117
rect 13998 5108 14004 5120
rect 14056 5108 14062 5160
rect 15470 5148 15476 5160
rect 14108 5120 15476 5148
rect 11057 5083 11115 5089
rect 11057 5049 11069 5083
rect 11103 5080 11115 5083
rect 13630 5080 13636 5092
rect 11103 5052 13636 5080
rect 11103 5049 11115 5052
rect 11057 5043 11115 5049
rect 13630 5040 13636 5052
rect 13688 5040 13694 5092
rect 12253 5015 12311 5021
rect 12253 5012 12265 5015
rect 10796 4984 12265 5012
rect 10597 4975 10655 4981
rect 12253 4981 12265 4984
rect 12299 4981 12311 5015
rect 12802 5012 12808 5024
rect 12763 4984 12808 5012
rect 12253 4975 12311 4981
rect 12802 4972 12808 4984
rect 12860 4972 12866 5024
rect 12897 5015 12955 5021
rect 12897 4981 12909 5015
rect 12943 5012 12955 5015
rect 14108 5012 14136 5120
rect 15470 5108 15476 5120
rect 15528 5108 15534 5160
rect 15562 5108 15568 5160
rect 15620 5148 15626 5160
rect 15657 5151 15715 5157
rect 15657 5148 15669 5151
rect 15620 5120 15669 5148
rect 15620 5108 15626 5120
rect 15657 5117 15669 5120
rect 15703 5117 15715 5151
rect 15657 5111 15715 5117
rect 16114 5108 16120 5160
rect 16172 5148 16178 5160
rect 16393 5151 16451 5157
rect 16393 5148 16405 5151
rect 16172 5120 16405 5148
rect 16172 5108 16178 5120
rect 16393 5117 16405 5120
rect 16439 5117 16451 5151
rect 16393 5111 16451 5117
rect 16574 5108 16580 5160
rect 16632 5148 16638 5160
rect 18616 5148 18644 5179
rect 18690 5148 18696 5160
rect 16632 5120 18092 5148
rect 18616 5120 18696 5148
rect 16632 5108 16638 5120
rect 14182 5040 14188 5092
rect 14240 5080 14246 5092
rect 14737 5083 14795 5089
rect 14737 5080 14749 5083
rect 14240 5052 14749 5080
rect 14240 5040 14246 5052
rect 14737 5049 14749 5052
rect 14783 5049 14795 5083
rect 14737 5043 14795 5049
rect 15286 5040 15292 5092
rect 15344 5080 15350 5092
rect 15749 5083 15807 5089
rect 15749 5080 15761 5083
rect 15344 5052 15761 5080
rect 15344 5040 15350 5052
rect 15749 5049 15761 5052
rect 15795 5049 15807 5083
rect 15749 5043 15807 5049
rect 17313 5083 17371 5089
rect 17313 5049 17325 5083
rect 17359 5080 17371 5083
rect 17954 5080 17960 5092
rect 17359 5052 17960 5080
rect 17359 5049 17371 5052
rect 17313 5043 17371 5049
rect 17954 5040 17960 5052
rect 18012 5040 18018 5092
rect 18064 5080 18092 5120
rect 18690 5108 18696 5120
rect 18748 5108 18754 5160
rect 19337 5151 19395 5157
rect 19337 5117 19349 5151
rect 19383 5117 19395 5151
rect 19337 5111 19395 5117
rect 18064 5052 18552 5080
rect 12943 4984 14136 5012
rect 12943 4981 12955 4984
rect 12897 4975 12955 4981
rect 14274 4972 14280 5024
rect 14332 5012 14338 5024
rect 14645 5015 14703 5021
rect 14645 5012 14657 5015
rect 14332 4984 14657 5012
rect 14332 4972 14338 4984
rect 14645 4981 14657 4984
rect 14691 5012 14703 5015
rect 15194 5012 15200 5024
rect 14691 4984 15200 5012
rect 14691 4981 14703 4984
rect 14645 4975 14703 4981
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 16577 5015 16635 5021
rect 16577 4981 16589 5015
rect 16623 5012 16635 5015
rect 16850 5012 16856 5024
rect 16623 4984 16856 5012
rect 16623 4981 16635 4984
rect 16577 4975 16635 4981
rect 16850 4972 16856 4984
rect 16908 4972 16914 5024
rect 17402 4972 17408 5024
rect 17460 5012 17466 5024
rect 17460 4984 17505 5012
rect 17460 4972 17466 4984
rect 17586 4972 17592 5024
rect 17644 5012 17650 5024
rect 18524 5021 18552 5052
rect 18966 5040 18972 5092
rect 19024 5080 19030 5092
rect 19352 5080 19380 5111
rect 19426 5108 19432 5160
rect 19484 5148 19490 5160
rect 19593 5151 19651 5157
rect 19593 5148 19605 5151
rect 19484 5120 19605 5148
rect 19484 5108 19490 5120
rect 19593 5117 19605 5120
rect 19639 5117 19651 5151
rect 19593 5111 19651 5117
rect 19024 5052 19380 5080
rect 19024 5040 19030 5052
rect 18417 5015 18475 5021
rect 18417 5012 18429 5015
rect 17644 4984 18429 5012
rect 17644 4972 17650 4984
rect 18417 4981 18429 4984
rect 18463 4981 18475 5015
rect 18417 4975 18475 4981
rect 18509 5015 18567 5021
rect 18509 4981 18521 5015
rect 18555 4981 18567 5015
rect 18509 4975 18567 4981
rect 19245 5015 19303 5021
rect 19245 4981 19257 5015
rect 19291 5012 19303 5015
rect 19794 5012 19800 5024
rect 19291 4984 19800 5012
rect 19291 4981 19303 4984
rect 19245 4975 19303 4981
rect 19794 4972 19800 4984
rect 19852 4972 19858 5024
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 2041 4811 2099 4817
rect 2041 4777 2053 4811
rect 2087 4808 2099 4811
rect 2406 4808 2412 4820
rect 2087 4780 2412 4808
rect 2087 4777 2099 4780
rect 2041 4771 2099 4777
rect 2406 4768 2412 4780
rect 2464 4768 2470 4820
rect 4985 4811 5043 4817
rect 4985 4777 4997 4811
rect 5031 4808 5043 4811
rect 5442 4808 5448 4820
rect 5031 4780 5448 4808
rect 5031 4777 5043 4780
rect 4985 4771 5043 4777
rect 5442 4768 5448 4780
rect 5500 4808 5506 4820
rect 5537 4811 5595 4817
rect 5537 4808 5549 4811
rect 5500 4780 5549 4808
rect 5500 4768 5506 4780
rect 5537 4777 5549 4780
rect 5583 4777 5595 4811
rect 5537 4771 5595 4777
rect 7466 4768 7472 4820
rect 7524 4808 7530 4820
rect 7653 4811 7711 4817
rect 7653 4808 7665 4811
rect 7524 4780 7665 4808
rect 7524 4768 7530 4780
rect 7653 4777 7665 4780
rect 7699 4777 7711 4811
rect 8386 4808 8392 4820
rect 8347 4780 8392 4808
rect 7653 4771 7711 4777
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 9217 4811 9275 4817
rect 9217 4777 9229 4811
rect 9263 4808 9275 4811
rect 9398 4808 9404 4820
rect 9263 4780 9404 4808
rect 9263 4777 9275 4780
rect 9217 4771 9275 4777
rect 9398 4768 9404 4780
rect 9456 4768 9462 4820
rect 9674 4808 9680 4820
rect 9635 4780 9680 4808
rect 9674 4768 9680 4780
rect 9732 4768 9738 4820
rect 10045 4811 10103 4817
rect 10045 4777 10057 4811
rect 10091 4808 10103 4811
rect 10502 4808 10508 4820
rect 10091 4780 10508 4808
rect 10091 4777 10103 4780
rect 10045 4771 10103 4777
rect 10502 4768 10508 4780
rect 10560 4768 10566 4820
rect 11517 4811 11575 4817
rect 11517 4777 11529 4811
rect 11563 4808 11575 4811
rect 13814 4808 13820 4820
rect 11563 4780 13820 4808
rect 11563 4777 11575 4780
rect 11517 4771 11575 4777
rect 13814 4768 13820 4780
rect 13872 4768 13878 4820
rect 14182 4808 14188 4820
rect 14143 4780 14188 4808
rect 14182 4768 14188 4780
rect 14240 4768 14246 4820
rect 15838 4768 15844 4820
rect 15896 4808 15902 4820
rect 16669 4811 16727 4817
rect 16669 4808 16681 4811
rect 15896 4780 16681 4808
rect 15896 4768 15902 4780
rect 16669 4777 16681 4780
rect 16715 4777 16727 4811
rect 16669 4771 16727 4777
rect 17310 4768 17316 4820
rect 17368 4808 17374 4820
rect 18785 4811 18843 4817
rect 18785 4808 18797 4811
rect 17368 4780 18797 4808
rect 17368 4768 17374 4780
rect 18785 4777 18797 4780
rect 18831 4808 18843 4811
rect 19426 4808 19432 4820
rect 18831 4780 19432 4808
rect 18831 4777 18843 4780
rect 18785 4771 18843 4777
rect 19426 4768 19432 4780
rect 19484 4768 19490 4820
rect 19613 4811 19671 4817
rect 19613 4777 19625 4811
rect 19659 4808 19671 4811
rect 19886 4808 19892 4820
rect 19659 4780 19892 4808
rect 19659 4777 19671 4780
rect 19613 4771 19671 4777
rect 19886 4768 19892 4780
rect 19944 4768 19950 4820
rect 5810 4700 5816 4752
rect 5868 4740 5874 4752
rect 5868 4712 6316 4740
rect 5868 4700 5874 4712
rect 2409 4675 2467 4681
rect 2409 4641 2421 4675
rect 2455 4672 2467 4675
rect 2774 4672 2780 4684
rect 2455 4644 2780 4672
rect 2455 4641 2467 4644
rect 2409 4635 2467 4641
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 2958 4632 2964 4684
rect 3016 4672 3022 4684
rect 6288 4681 6316 4712
rect 6822 4700 6828 4752
rect 6880 4740 6886 4752
rect 8294 4740 8300 4752
rect 6880 4712 7604 4740
rect 8255 4712 8300 4740
rect 6880 4700 6886 4712
rect 3513 4675 3571 4681
rect 3513 4672 3525 4675
rect 3016 4644 3525 4672
rect 3016 4632 3022 4644
rect 3513 4641 3525 4644
rect 3559 4641 3571 4675
rect 3513 4635 3571 4641
rect 5445 4675 5503 4681
rect 5445 4641 5457 4675
rect 5491 4672 5503 4675
rect 6273 4675 6331 4681
rect 5491 4644 6224 4672
rect 5491 4641 5503 4644
rect 5445 4635 5503 4641
rect 2314 4564 2320 4616
rect 2372 4604 2378 4616
rect 2501 4607 2559 4613
rect 2501 4604 2513 4607
rect 2372 4576 2513 4604
rect 2372 4564 2378 4576
rect 2501 4573 2513 4576
rect 2547 4573 2559 4607
rect 2682 4604 2688 4616
rect 2643 4576 2688 4604
rect 2501 4567 2559 4573
rect 2682 4564 2688 4576
rect 2740 4564 2746 4616
rect 2866 4604 2872 4616
rect 2827 4576 2872 4604
rect 2866 4564 2872 4576
rect 2924 4564 2930 4616
rect 3602 4604 3608 4616
rect 3563 4576 3608 4604
rect 3602 4564 3608 4576
rect 3660 4564 3666 4616
rect 3789 4607 3847 4613
rect 3789 4573 3801 4607
rect 3835 4604 3847 4607
rect 4246 4604 4252 4616
rect 3835 4576 4252 4604
rect 3835 4573 3847 4576
rect 3789 4567 3847 4573
rect 4246 4564 4252 4576
rect 4304 4564 4310 4616
rect 5718 4604 5724 4616
rect 5679 4576 5724 4604
rect 5718 4564 5724 4576
rect 5776 4564 5782 4616
rect 2406 4496 2412 4548
rect 2464 4536 2470 4548
rect 3145 4539 3203 4545
rect 3145 4536 3157 4539
rect 2464 4508 3157 4536
rect 2464 4496 2470 4508
rect 3145 4505 3157 4508
rect 3191 4505 3203 4539
rect 3145 4499 3203 4505
rect 5074 4468 5080 4480
rect 5035 4440 5080 4468
rect 5074 4428 5080 4440
rect 5132 4428 5138 4480
rect 6196 4468 6224 4644
rect 6273 4641 6285 4675
rect 6319 4641 6331 4675
rect 6273 4635 6331 4641
rect 6540 4675 6598 4681
rect 6540 4641 6552 4675
rect 6586 4672 6598 4675
rect 6914 4672 6920 4684
rect 6586 4644 6920 4672
rect 6586 4641 6598 4644
rect 6540 4635 6598 4641
rect 6914 4632 6920 4644
rect 6972 4632 6978 4684
rect 7576 4604 7604 4712
rect 8294 4700 8300 4712
rect 8352 4700 8358 4752
rect 10318 4740 10324 4752
rect 9048 4712 10324 4740
rect 9048 4681 9076 4712
rect 10318 4700 10324 4712
rect 10376 4700 10382 4752
rect 11054 4740 11060 4752
rect 10520 4712 11060 4740
rect 9033 4675 9091 4681
rect 9033 4641 9045 4675
rect 9079 4641 9091 4675
rect 9033 4635 9091 4641
rect 8481 4607 8539 4613
rect 8481 4604 8493 4607
rect 7576 4576 8493 4604
rect 8481 4573 8493 4576
rect 8527 4573 8539 4607
rect 8481 4567 8539 4573
rect 10137 4607 10195 4613
rect 10137 4573 10149 4607
rect 10183 4573 10195 4607
rect 10137 4567 10195 4573
rect 10321 4607 10379 4613
rect 10321 4573 10333 4607
rect 10367 4604 10379 4607
rect 10520 4604 10548 4712
rect 11054 4700 11060 4712
rect 11112 4700 11118 4752
rect 11698 4700 11704 4752
rect 11756 4740 11762 4752
rect 12621 4743 12679 4749
rect 11756 4712 12572 4740
rect 11756 4700 11762 4712
rect 10689 4675 10747 4681
rect 10689 4641 10701 4675
rect 10735 4641 10747 4675
rect 10689 4635 10747 4641
rect 10367 4576 10548 4604
rect 10597 4607 10655 4613
rect 10367 4573 10379 4576
rect 10321 4567 10379 4573
rect 10597 4573 10609 4607
rect 10643 4604 10655 4607
rect 10704 4604 10732 4635
rect 11146 4632 11152 4684
rect 11204 4672 11210 4684
rect 11425 4675 11483 4681
rect 11425 4672 11437 4675
rect 11204 4644 11437 4672
rect 11204 4632 11210 4644
rect 11425 4641 11437 4644
rect 11471 4641 11483 4675
rect 12434 4672 12440 4684
rect 11425 4635 11483 4641
rect 11532 4644 12440 4672
rect 11532 4604 11560 4644
rect 12434 4632 12440 4644
rect 12492 4632 12498 4684
rect 12544 4672 12572 4712
rect 12621 4709 12633 4743
rect 12667 4740 12679 4743
rect 12667 4712 12940 4740
rect 12667 4709 12679 4712
rect 12621 4703 12679 4709
rect 12912 4672 12940 4712
rect 13906 4700 13912 4752
rect 13964 4740 13970 4752
rect 14645 4743 14703 4749
rect 14645 4740 14657 4743
rect 13964 4712 14657 4740
rect 13964 4700 13970 4712
rect 14645 4709 14657 4712
rect 14691 4709 14703 4743
rect 15556 4743 15614 4749
rect 15556 4740 15568 4743
rect 14645 4703 14703 4709
rect 14844 4712 15568 4740
rect 13081 4675 13139 4681
rect 13081 4672 13093 4675
rect 12544 4644 12848 4672
rect 12912 4644 13093 4672
rect 11698 4604 11704 4616
rect 10643 4576 11560 4604
rect 11659 4576 11704 4604
rect 10643 4573 10655 4576
rect 10597 4567 10655 4573
rect 9582 4536 9588 4548
rect 7208 4508 9588 4536
rect 7208 4468 7236 4508
rect 9582 4496 9588 4508
rect 9640 4496 9646 4548
rect 10152 4536 10180 4567
rect 11698 4564 11704 4576
rect 11756 4564 11762 4616
rect 11974 4564 11980 4616
rect 12032 4604 12038 4616
rect 12161 4607 12219 4613
rect 12161 4604 12173 4607
rect 12032 4576 12173 4604
rect 12032 4564 12038 4576
rect 12161 4573 12173 4576
rect 12207 4604 12219 4607
rect 12342 4604 12348 4616
rect 12207 4576 12348 4604
rect 12207 4573 12219 4576
rect 12161 4567 12219 4573
rect 12342 4564 12348 4576
rect 12400 4604 12406 4616
rect 12820 4613 12848 4644
rect 13081 4641 13093 4644
rect 13127 4641 13139 4675
rect 13262 4672 13268 4684
rect 13223 4644 13268 4672
rect 13081 4635 13139 4641
rect 13262 4632 13268 4644
rect 13320 4632 13326 4684
rect 14274 4632 14280 4684
rect 14332 4672 14338 4684
rect 14553 4675 14611 4681
rect 14553 4672 14565 4675
rect 14332 4644 14565 4672
rect 14332 4632 14338 4644
rect 14553 4641 14565 4644
rect 14599 4641 14611 4675
rect 14553 4635 14611 4641
rect 14844 4613 14872 4712
rect 15556 4709 15568 4712
rect 15602 4740 15614 4743
rect 15930 4740 15936 4752
rect 15602 4712 15936 4740
rect 15602 4709 15614 4712
rect 15556 4703 15614 4709
rect 15930 4700 15936 4712
rect 15988 4740 15994 4752
rect 16482 4740 16488 4752
rect 15988 4712 16488 4740
rect 15988 4700 15994 4712
rect 16482 4700 16488 4712
rect 16540 4700 16546 4752
rect 16942 4700 16948 4752
rect 17000 4740 17006 4752
rect 17672 4743 17730 4749
rect 17000 4712 17540 4740
rect 17000 4700 17006 4712
rect 15289 4675 15347 4681
rect 15289 4641 15301 4675
rect 15335 4672 15347 4675
rect 15378 4672 15384 4684
rect 15335 4644 15384 4672
rect 15335 4641 15347 4644
rect 15289 4635 15347 4641
rect 15378 4632 15384 4644
rect 15436 4672 15442 4684
rect 17405 4675 17463 4681
rect 17405 4672 17417 4675
rect 15436 4644 17417 4672
rect 15436 4632 15442 4644
rect 17405 4641 17417 4644
rect 17451 4641 17463 4675
rect 17512 4672 17540 4712
rect 17672 4709 17684 4743
rect 17718 4740 17730 4743
rect 18690 4740 18696 4752
rect 17718 4712 18696 4740
rect 17718 4709 17730 4712
rect 17672 4703 17730 4709
rect 18690 4700 18696 4712
rect 18748 4700 18754 4752
rect 20254 4740 20260 4752
rect 20180 4712 20260 4740
rect 19061 4675 19119 4681
rect 19061 4672 19073 4675
rect 17512 4644 19073 4672
rect 17405 4635 17463 4641
rect 19061 4641 19073 4644
rect 19107 4641 19119 4675
rect 19981 4675 20039 4681
rect 19981 4672 19993 4675
rect 19061 4635 19119 4641
rect 19904 4644 19993 4672
rect 12713 4607 12771 4613
rect 12713 4604 12725 4607
rect 12400 4576 12725 4604
rect 12400 4564 12406 4576
rect 12713 4573 12725 4576
rect 12759 4573 12771 4607
rect 12713 4567 12771 4573
rect 12805 4607 12863 4613
rect 12805 4573 12817 4607
rect 12851 4604 12863 4607
rect 13541 4607 13599 4613
rect 12851 4576 13492 4604
rect 12851 4573 12863 4576
rect 12805 4567 12863 4573
rect 10962 4536 10968 4548
rect 10152 4508 10968 4536
rect 10962 4496 10968 4508
rect 11020 4496 11026 4548
rect 11057 4539 11115 4545
rect 11057 4505 11069 4539
rect 11103 4536 11115 4539
rect 12986 4536 12992 4548
rect 11103 4508 12992 4536
rect 11103 4505 11115 4508
rect 11057 4499 11115 4505
rect 12986 4496 12992 4508
rect 13044 4496 13050 4548
rect 13464 4536 13492 4576
rect 13541 4573 13553 4607
rect 13587 4604 13599 4607
rect 14829 4607 14887 4613
rect 13587 4576 14596 4604
rect 13587 4573 13599 4576
rect 13541 4567 13599 4573
rect 14568 4548 14596 4576
rect 14829 4573 14841 4607
rect 14875 4573 14887 4607
rect 14829 4567 14887 4573
rect 13814 4536 13820 4548
rect 13464 4508 13820 4536
rect 13814 4496 13820 4508
rect 13872 4496 13878 4548
rect 14550 4496 14556 4548
rect 14608 4496 14614 4548
rect 19058 4496 19064 4548
rect 19116 4536 19122 4548
rect 19334 4536 19340 4548
rect 19116 4508 19340 4536
rect 19116 4496 19122 4508
rect 19334 4496 19340 4508
rect 19392 4496 19398 4548
rect 19904 4536 19932 4644
rect 19981 4641 19993 4644
rect 20027 4641 20039 4675
rect 19981 4635 20039 4641
rect 20070 4604 20076 4616
rect 20031 4576 20076 4604
rect 20070 4564 20076 4576
rect 20128 4564 20134 4616
rect 20180 4613 20208 4712
rect 20254 4700 20260 4712
rect 20312 4700 20318 4752
rect 20165 4607 20223 4613
rect 20165 4573 20177 4607
rect 20211 4573 20223 4607
rect 20165 4567 20223 4573
rect 20254 4564 20260 4616
rect 20312 4604 20318 4616
rect 20901 4607 20959 4613
rect 20901 4604 20913 4607
rect 20312 4576 20913 4604
rect 20312 4564 20318 4576
rect 20901 4573 20913 4576
rect 20947 4573 20959 4607
rect 20901 4567 20959 4573
rect 19978 4536 19984 4548
rect 19904 4508 19984 4536
rect 19978 4496 19984 4508
rect 20036 4496 20042 4548
rect 7926 4468 7932 4480
rect 6196 4440 7236 4468
rect 7887 4440 7932 4468
rect 7926 4428 7932 4440
rect 7984 4428 7990 4480
rect 8294 4428 8300 4480
rect 8352 4468 8358 4480
rect 8846 4468 8852 4480
rect 8352 4440 8852 4468
rect 8352 4428 8358 4440
rect 8846 4428 8852 4440
rect 8904 4428 8910 4480
rect 9122 4428 9128 4480
rect 9180 4468 9186 4480
rect 10597 4471 10655 4477
rect 10597 4468 10609 4471
rect 9180 4440 10609 4468
rect 9180 4428 9186 4440
rect 10597 4437 10609 4440
rect 10643 4437 10655 4471
rect 10597 4431 10655 4437
rect 10873 4471 10931 4477
rect 10873 4437 10885 4471
rect 10919 4468 10931 4471
rect 11974 4468 11980 4480
rect 10919 4440 11980 4468
rect 10919 4437 10931 4440
rect 10873 4431 10931 4437
rect 11974 4428 11980 4440
rect 12032 4428 12038 4480
rect 12253 4471 12311 4477
rect 12253 4437 12265 4471
rect 12299 4468 12311 4471
rect 12894 4468 12900 4480
rect 12299 4440 12900 4468
rect 12299 4437 12311 4440
rect 12253 4431 12311 4437
rect 12894 4428 12900 4440
rect 12952 4428 12958 4480
rect 13081 4471 13139 4477
rect 13081 4437 13093 4471
rect 13127 4468 13139 4471
rect 15102 4468 15108 4480
rect 13127 4440 15108 4468
rect 13127 4437 13139 4440
rect 13081 4431 13139 4437
rect 15102 4428 15108 4440
rect 15160 4428 15166 4480
rect 19245 4471 19303 4477
rect 19245 4437 19257 4471
rect 19291 4468 19303 4471
rect 20438 4468 20444 4480
rect 19291 4440 20444 4468
rect 19291 4437 19303 4440
rect 19245 4431 19303 4437
rect 20438 4428 20444 4440
rect 20496 4428 20502 4480
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 3510 4224 3516 4276
rect 3568 4264 3574 4276
rect 4065 4267 4123 4273
rect 4065 4264 4077 4267
rect 3568 4236 4077 4264
rect 3568 4224 3574 4236
rect 4065 4233 4077 4236
rect 4111 4233 4123 4267
rect 4893 4267 4951 4273
rect 4893 4264 4905 4267
rect 4065 4227 4123 4233
rect 4448 4236 4905 4264
rect 4154 4156 4160 4208
rect 4212 4196 4218 4208
rect 4338 4196 4344 4208
rect 4212 4168 4344 4196
rect 4212 4156 4218 4168
rect 4338 4156 4344 4168
rect 4396 4156 4402 4208
rect 3418 4088 3424 4140
rect 3476 4128 3482 4140
rect 4448 4128 4476 4236
rect 4893 4233 4905 4236
rect 4939 4233 4951 4267
rect 4893 4227 4951 4233
rect 7009 4267 7067 4273
rect 7009 4233 7021 4267
rect 7055 4264 7067 4267
rect 7282 4264 7288 4276
rect 7055 4236 7288 4264
rect 7055 4233 7067 4236
rect 7009 4227 7067 4233
rect 7282 4224 7288 4236
rect 7340 4224 7346 4276
rect 10134 4264 10140 4276
rect 10095 4236 10140 4264
rect 10134 4224 10140 4236
rect 10192 4224 10198 4276
rect 10962 4224 10968 4276
rect 11020 4264 11026 4276
rect 13906 4264 13912 4276
rect 11020 4236 13912 4264
rect 11020 4224 11026 4236
rect 13906 4224 13912 4236
rect 13964 4224 13970 4276
rect 13998 4224 14004 4276
rect 14056 4264 14062 4276
rect 16206 4264 16212 4276
rect 14056 4236 16212 4264
rect 14056 4224 14062 4236
rect 16206 4224 16212 4236
rect 16264 4224 16270 4276
rect 17954 4224 17960 4276
rect 18012 4264 18018 4276
rect 18049 4267 18107 4273
rect 18049 4264 18061 4267
rect 18012 4236 18061 4264
rect 18012 4224 18018 4236
rect 18049 4233 18061 4236
rect 18095 4233 18107 4267
rect 18049 4227 18107 4233
rect 19426 4224 19432 4276
rect 19484 4224 19490 4276
rect 19610 4224 19616 4276
rect 19668 4264 19674 4276
rect 19705 4267 19763 4273
rect 19705 4264 19717 4267
rect 19668 4236 19717 4264
rect 19668 4224 19674 4236
rect 19705 4233 19717 4236
rect 19751 4233 19763 4267
rect 19705 4227 19763 4233
rect 19889 4267 19947 4273
rect 19889 4233 19901 4267
rect 19935 4264 19947 4267
rect 19978 4264 19984 4276
rect 19935 4236 19984 4264
rect 19935 4233 19947 4236
rect 19889 4227 19947 4233
rect 19978 4224 19984 4236
rect 20036 4224 20042 4276
rect 5718 4196 5724 4208
rect 5552 4168 5724 4196
rect 3476 4100 4476 4128
rect 4617 4131 4675 4137
rect 3476 4088 3482 4100
rect 4617 4097 4629 4131
rect 4663 4128 4675 4131
rect 4890 4128 4896 4140
rect 4663 4100 4896 4128
rect 4663 4097 4675 4100
rect 4617 4091 4675 4097
rect 4890 4088 4896 4100
rect 4948 4088 4954 4140
rect 5552 4137 5580 4168
rect 5718 4156 5724 4168
rect 5776 4156 5782 4208
rect 6914 4196 6920 4208
rect 6380 4168 6920 4196
rect 6380 4137 6408 4168
rect 6914 4156 6920 4168
rect 6972 4196 6978 4208
rect 11149 4199 11207 4205
rect 6972 4168 7604 4196
rect 6972 4156 6978 4168
rect 7576 4137 7604 4168
rect 11149 4165 11161 4199
rect 11195 4196 11207 4199
rect 11882 4196 11888 4208
rect 11195 4168 11888 4196
rect 11195 4165 11207 4168
rect 11149 4159 11207 4165
rect 11882 4156 11888 4168
rect 11940 4156 11946 4208
rect 13814 4196 13820 4208
rect 13775 4168 13820 4196
rect 13814 4156 13820 4168
rect 13872 4196 13878 4208
rect 15289 4199 15347 4205
rect 13872 4168 14688 4196
rect 13872 4156 13878 4168
rect 5537 4131 5595 4137
rect 5537 4097 5549 4131
rect 5583 4097 5595 4131
rect 6365 4131 6423 4137
rect 5537 4091 5595 4097
rect 5920 4100 6316 4128
rect 2041 4063 2099 4069
rect 2041 4029 2053 4063
rect 2087 4060 2099 4063
rect 2682 4060 2688 4072
rect 2087 4032 2688 4060
rect 2087 4029 2099 4032
rect 2041 4023 2099 4029
rect 2682 4020 2688 4032
rect 2740 4020 2746 4072
rect 4706 4020 4712 4072
rect 4764 4060 4770 4072
rect 5353 4063 5411 4069
rect 4764 4032 5120 4060
rect 4764 4020 4770 4032
rect 2308 3995 2366 4001
rect 2308 3961 2320 3995
rect 2354 3992 2366 3995
rect 2498 3992 2504 4004
rect 2354 3964 2504 3992
rect 2354 3961 2366 3964
rect 2308 3955 2366 3961
rect 2498 3952 2504 3964
rect 2556 3952 2562 4004
rect 3142 3952 3148 4004
rect 3200 3992 3206 4004
rect 3878 3992 3884 4004
rect 3200 3964 3884 3992
rect 3200 3952 3206 3964
rect 3878 3952 3884 3964
rect 3936 3952 3942 4004
rect 4154 3952 4160 4004
rect 4212 3992 4218 4004
rect 4433 3995 4491 4001
rect 4433 3992 4445 3995
rect 4212 3964 4445 3992
rect 4212 3952 4218 3964
rect 4433 3961 4445 3964
rect 4479 3992 4491 3995
rect 4982 3992 4988 4004
rect 4479 3964 4988 3992
rect 4479 3961 4491 3964
rect 4433 3955 4491 3961
rect 4982 3952 4988 3964
rect 5040 3952 5046 4004
rect 5092 3992 5120 4032
rect 5353 4029 5365 4063
rect 5399 4060 5411 4063
rect 5920 4060 5948 4100
rect 6086 4060 6092 4072
rect 5399 4032 5948 4060
rect 6047 4032 6092 4060
rect 5399 4029 5411 4032
rect 5353 4023 5411 4029
rect 6086 4020 6092 4032
rect 6144 4020 6150 4072
rect 6288 4060 6316 4100
rect 6365 4097 6377 4131
rect 6411 4097 6423 4131
rect 6365 4091 6423 4097
rect 7561 4131 7619 4137
rect 7561 4097 7573 4131
rect 7607 4097 7619 4131
rect 7561 4091 7619 4097
rect 10502 4088 10508 4140
rect 10560 4128 10566 4140
rect 10597 4131 10655 4137
rect 10597 4128 10609 4131
rect 10560 4100 10609 4128
rect 10560 4088 10566 4100
rect 10597 4097 10609 4100
rect 10643 4097 10655 4131
rect 10597 4091 10655 4097
rect 10689 4131 10747 4137
rect 10689 4097 10701 4131
rect 10735 4097 10747 4131
rect 11698 4128 11704 4140
rect 11659 4100 11704 4128
rect 10689 4091 10747 4097
rect 6638 4060 6644 4072
rect 6288 4032 6644 4060
rect 6638 4020 6644 4032
rect 6696 4020 6702 4072
rect 7469 4063 7527 4069
rect 7469 4029 7481 4063
rect 7515 4060 7527 4063
rect 7926 4060 7932 4072
rect 7515 4032 7932 4060
rect 7515 4029 7527 4032
rect 7469 4023 7527 4029
rect 7926 4020 7932 4032
rect 7984 4020 7990 4072
rect 8478 4060 8484 4072
rect 8439 4032 8484 4060
rect 8478 4020 8484 4032
rect 8536 4020 8542 4072
rect 8748 4063 8806 4069
rect 8748 4029 8760 4063
rect 8794 4060 8806 4063
rect 10134 4060 10140 4072
rect 8794 4032 10140 4060
rect 8794 4029 8806 4032
rect 8748 4023 8806 4029
rect 10134 4020 10140 4032
rect 10192 4060 10198 4072
rect 10704 4060 10732 4091
rect 11698 4088 11704 4100
rect 11756 4088 11762 4140
rect 11790 4088 11796 4140
rect 11848 4128 11854 4140
rect 11848 4100 12572 4128
rect 11848 4088 11854 4100
rect 10192 4032 10732 4060
rect 12437 4063 12495 4069
rect 10192 4020 10198 4032
rect 12437 4029 12449 4063
rect 12483 4029 12495 4063
rect 12544 4060 12572 4100
rect 14458 4088 14464 4140
rect 14516 4128 14522 4140
rect 14660 4137 14688 4168
rect 15289 4165 15301 4199
rect 15335 4165 15347 4199
rect 15289 4159 15347 4165
rect 14553 4131 14611 4137
rect 14553 4128 14565 4131
rect 14516 4100 14565 4128
rect 14516 4088 14522 4100
rect 14553 4097 14565 4100
rect 14599 4097 14611 4131
rect 14553 4091 14611 4097
rect 14645 4131 14703 4137
rect 14645 4097 14657 4131
rect 14691 4097 14703 4131
rect 14645 4091 14703 4097
rect 12544 4032 12839 4060
rect 12437 4023 12495 4029
rect 5258 3992 5264 4004
rect 5092 3964 5264 3992
rect 5258 3952 5264 3964
rect 5316 3952 5322 4004
rect 7190 3992 7196 4004
rect 5736 3964 7196 3992
rect 2406 3884 2412 3936
rect 2464 3924 2470 3936
rect 2866 3924 2872 3936
rect 2464 3896 2872 3924
rect 2464 3884 2470 3896
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 3421 3927 3479 3933
rect 3421 3893 3433 3927
rect 3467 3924 3479 3927
rect 3510 3924 3516 3936
rect 3467 3896 3516 3924
rect 3467 3893 3479 3896
rect 3421 3887 3479 3893
rect 3510 3884 3516 3896
rect 3568 3884 3574 3936
rect 3970 3884 3976 3936
rect 4028 3924 4034 3936
rect 5736 3933 5764 3964
rect 7190 3952 7196 3964
rect 7248 3952 7254 4004
rect 7650 3952 7656 4004
rect 7708 3992 7714 4004
rect 10042 3992 10048 4004
rect 7708 3964 10048 3992
rect 7708 3952 7714 3964
rect 10042 3952 10048 3964
rect 10100 3992 10106 4004
rect 10226 3992 10232 4004
rect 10100 3964 10232 3992
rect 10100 3952 10106 3964
rect 10226 3952 10232 3964
rect 10284 3952 10290 4004
rect 12452 3992 12480 4023
rect 12704 3995 12762 4001
rect 12452 3964 12664 3992
rect 12636 3936 12664 3964
rect 12704 3961 12716 3995
rect 12750 3961 12762 3995
rect 12811 3992 12839 4032
rect 13814 4020 13820 4072
rect 13872 4060 13878 4072
rect 14274 4060 14280 4072
rect 13872 4032 14280 4060
rect 13872 4020 13878 4032
rect 14274 4020 14280 4032
rect 14332 4020 14338 4072
rect 15304 4060 15332 4159
rect 16482 4156 16488 4208
rect 16540 4196 16546 4208
rect 18690 4196 18696 4208
rect 16540 4168 16896 4196
rect 16540 4156 16546 4168
rect 15838 4128 15844 4140
rect 15799 4100 15844 4128
rect 15838 4088 15844 4100
rect 15896 4088 15902 4140
rect 16868 4137 16896 4168
rect 18616 4168 18696 4196
rect 16853 4131 16911 4137
rect 16853 4097 16865 4131
rect 16899 4097 16911 4131
rect 16853 4091 16911 4097
rect 17770 4088 17776 4140
rect 17828 4128 17834 4140
rect 17954 4128 17960 4140
rect 17828 4100 17960 4128
rect 17828 4088 17834 4100
rect 17954 4088 17960 4100
rect 18012 4088 18018 4140
rect 18616 4137 18644 4168
rect 18690 4156 18696 4168
rect 18748 4156 18754 4208
rect 18601 4131 18659 4137
rect 18601 4097 18613 4131
rect 18647 4097 18659 4131
rect 19153 4131 19211 4137
rect 19153 4128 19165 4131
rect 18601 4091 18659 4097
rect 18708 4100 19165 4128
rect 16574 4060 16580 4072
rect 15304 4032 16580 4060
rect 16574 4020 16580 4032
rect 16632 4020 16638 4072
rect 16666 4020 16672 4072
rect 16724 4060 16730 4072
rect 16761 4063 16819 4069
rect 16761 4060 16773 4063
rect 16724 4032 16773 4060
rect 16724 4020 16730 4032
rect 16761 4029 16773 4032
rect 16807 4029 16819 4063
rect 17405 4063 17463 4069
rect 16761 4023 16819 4029
rect 16868 4032 17172 4060
rect 16868 3992 16896 4032
rect 12811 3964 16896 3992
rect 17144 3992 17172 4032
rect 17405 4029 17417 4063
rect 17451 4060 17463 4063
rect 18708 4060 18736 4100
rect 19153 4097 19165 4100
rect 19199 4097 19211 4131
rect 19444 4128 19472 4224
rect 20441 4131 20499 4137
rect 20441 4128 20453 4131
rect 19444 4100 20453 4128
rect 19153 4091 19211 4097
rect 20441 4097 20453 4100
rect 20487 4128 20499 4131
rect 20530 4128 20536 4140
rect 20487 4100 20536 4128
rect 20487 4097 20499 4100
rect 20441 4091 20499 4097
rect 20530 4088 20536 4100
rect 20588 4088 20594 4140
rect 17451 4032 18736 4060
rect 18969 4063 19027 4069
rect 17451 4029 17463 4032
rect 17405 4023 17463 4029
rect 18969 4029 18981 4063
rect 19015 4029 19027 4063
rect 20254 4060 20260 4072
rect 20215 4032 20260 4060
rect 18969 4023 19027 4029
rect 18984 3992 19012 4023
rect 20254 4020 20260 4032
rect 20312 4020 20318 4072
rect 17144 3964 19012 3992
rect 12704 3955 12762 3961
rect 4525 3927 4583 3933
rect 4525 3924 4537 3927
rect 4028 3896 4537 3924
rect 4028 3884 4034 3896
rect 4525 3893 4537 3896
rect 4571 3893 4583 3927
rect 4525 3887 4583 3893
rect 5721 3927 5779 3933
rect 5721 3893 5733 3927
rect 5767 3893 5779 3927
rect 5721 3887 5779 3893
rect 6181 3927 6239 3933
rect 6181 3893 6193 3927
rect 6227 3924 6239 3927
rect 6914 3924 6920 3936
rect 6227 3896 6920 3924
rect 6227 3893 6239 3896
rect 6181 3887 6239 3893
rect 6914 3884 6920 3896
rect 6972 3884 6978 3936
rect 7374 3924 7380 3936
rect 7335 3896 7380 3924
rect 7374 3884 7380 3896
rect 7432 3884 7438 3936
rect 8938 3884 8944 3936
rect 8996 3924 9002 3936
rect 9306 3924 9312 3936
rect 8996 3896 9312 3924
rect 8996 3884 9002 3896
rect 9306 3884 9312 3896
rect 9364 3924 9370 3936
rect 9861 3927 9919 3933
rect 9861 3924 9873 3927
rect 9364 3896 9873 3924
rect 9364 3884 9370 3896
rect 9861 3893 9873 3896
rect 9907 3893 9919 3927
rect 9861 3887 9919 3893
rect 10505 3927 10563 3933
rect 10505 3893 10517 3927
rect 10551 3924 10563 3927
rect 10594 3924 10600 3936
rect 10551 3896 10600 3924
rect 10551 3893 10563 3896
rect 10505 3887 10563 3893
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 11238 3884 11244 3936
rect 11296 3924 11302 3936
rect 11517 3927 11575 3933
rect 11517 3924 11529 3927
rect 11296 3896 11529 3924
rect 11296 3884 11302 3896
rect 11517 3893 11529 3896
rect 11563 3893 11575 3927
rect 11517 3887 11575 3893
rect 11609 3927 11667 3933
rect 11609 3893 11621 3927
rect 11655 3924 11667 3927
rect 12434 3924 12440 3936
rect 11655 3896 12440 3924
rect 11655 3893 11667 3896
rect 11609 3887 11667 3893
rect 12434 3884 12440 3896
rect 12492 3884 12498 3936
rect 12618 3884 12624 3936
rect 12676 3884 12682 3936
rect 12719 3924 12747 3955
rect 19610 3952 19616 4004
rect 19668 3992 19674 4004
rect 20349 3995 20407 4001
rect 20349 3992 20361 3995
rect 19668 3964 20361 3992
rect 19668 3952 19674 3964
rect 20349 3961 20361 3964
rect 20395 3961 20407 3995
rect 20349 3955 20407 3961
rect 13722 3924 13728 3936
rect 12719 3896 13728 3924
rect 13722 3884 13728 3896
rect 13780 3884 13786 3936
rect 14090 3924 14096 3936
rect 14051 3896 14096 3924
rect 14090 3884 14096 3896
rect 14148 3884 14154 3936
rect 14274 3884 14280 3936
rect 14332 3924 14338 3936
rect 14461 3927 14519 3933
rect 14461 3924 14473 3927
rect 14332 3896 14473 3924
rect 14332 3884 14338 3896
rect 14461 3893 14473 3896
rect 14507 3893 14519 3927
rect 14461 3887 14519 3893
rect 15378 3884 15384 3936
rect 15436 3924 15442 3936
rect 15657 3927 15715 3933
rect 15657 3924 15669 3927
rect 15436 3896 15669 3924
rect 15436 3884 15442 3896
rect 15657 3893 15669 3896
rect 15703 3893 15715 3927
rect 15657 3887 15715 3893
rect 15749 3927 15807 3933
rect 15749 3893 15761 3927
rect 15795 3924 15807 3927
rect 16301 3927 16359 3933
rect 16301 3924 16313 3927
rect 15795 3896 16313 3924
rect 15795 3893 15807 3896
rect 15749 3887 15807 3893
rect 16301 3893 16313 3896
rect 16347 3893 16359 3927
rect 16301 3887 16359 3893
rect 16574 3884 16580 3936
rect 16632 3924 16638 3936
rect 16669 3927 16727 3933
rect 16669 3924 16681 3927
rect 16632 3896 16681 3924
rect 16632 3884 16638 3896
rect 16669 3893 16681 3896
rect 16715 3893 16727 3927
rect 17586 3924 17592 3936
rect 17547 3896 17592 3924
rect 16669 3887 16727 3893
rect 17586 3884 17592 3896
rect 17644 3884 17650 3936
rect 17770 3884 17776 3936
rect 17828 3924 17834 3936
rect 18417 3927 18475 3933
rect 18417 3924 18429 3927
rect 17828 3896 18429 3924
rect 17828 3884 17834 3896
rect 18417 3893 18429 3896
rect 18463 3893 18475 3927
rect 18417 3887 18475 3893
rect 18509 3927 18567 3933
rect 18509 3893 18521 3927
rect 18555 3924 18567 3927
rect 18782 3924 18788 3936
rect 18555 3896 18788 3924
rect 18555 3893 18567 3896
rect 18509 3887 18567 3893
rect 18782 3884 18788 3896
rect 18840 3884 18846 3936
rect 19886 3884 19892 3936
rect 19944 3924 19950 3936
rect 20254 3924 20260 3936
rect 19944 3896 20260 3924
rect 19944 3884 19950 3896
rect 20254 3884 20260 3896
rect 20312 3884 20318 3936
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 1949 3723 2007 3729
rect 1949 3689 1961 3723
rect 1995 3689 2007 3723
rect 1949 3683 2007 3689
rect 2317 3723 2375 3729
rect 2317 3689 2329 3723
rect 2363 3720 2375 3723
rect 2406 3720 2412 3732
rect 2363 3692 2412 3720
rect 2363 3689 2375 3692
rect 2317 3683 2375 3689
rect 1964 3652 1992 3683
rect 2406 3680 2412 3692
rect 2464 3680 2470 3732
rect 2958 3720 2964 3732
rect 2919 3692 2964 3720
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 3418 3720 3424 3732
rect 3379 3692 3424 3720
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 3602 3680 3608 3732
rect 3660 3720 3666 3732
rect 4065 3723 4123 3729
rect 4065 3720 4077 3723
rect 3660 3692 4077 3720
rect 3660 3680 3666 3692
rect 4065 3689 4077 3692
rect 4111 3689 4123 3723
rect 4065 3683 4123 3689
rect 4433 3723 4491 3729
rect 4433 3689 4445 3723
rect 4479 3720 4491 3723
rect 5074 3720 5080 3732
rect 4479 3692 5080 3720
rect 4479 3689 4491 3692
rect 4433 3683 4491 3689
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 7006 3680 7012 3732
rect 7064 3720 7070 3732
rect 7101 3723 7159 3729
rect 7101 3720 7113 3723
rect 7064 3692 7113 3720
rect 7064 3680 7070 3692
rect 7101 3689 7113 3692
rect 7147 3689 7159 3723
rect 7374 3720 7380 3732
rect 7335 3692 7380 3720
rect 7101 3683 7159 3689
rect 7374 3680 7380 3692
rect 7432 3680 7438 3732
rect 7745 3723 7803 3729
rect 7745 3689 7757 3723
rect 7791 3720 7803 3723
rect 8573 3723 8631 3729
rect 8573 3720 8585 3723
rect 7791 3692 8585 3720
rect 7791 3689 7803 3692
rect 7745 3683 7803 3689
rect 8573 3689 8585 3692
rect 8619 3689 8631 3723
rect 11514 3720 11520 3732
rect 8573 3683 8631 3689
rect 9692 3692 10916 3720
rect 11475 3692 11520 3720
rect 3329 3655 3387 3661
rect 3329 3652 3341 3655
rect 1964 3624 3341 3652
rect 3329 3621 3341 3624
rect 3375 3621 3387 3655
rect 3329 3615 3387 3621
rect 4338 3612 4344 3664
rect 4396 3652 4402 3664
rect 4890 3652 4896 3664
rect 4396 3624 4896 3652
rect 4396 3612 4402 3624
rect 4890 3612 4896 3624
rect 4948 3612 4954 3664
rect 8205 3655 8263 3661
rect 8205 3621 8217 3655
rect 8251 3652 8263 3655
rect 9692 3652 9720 3692
rect 8251 3624 9720 3652
rect 8251 3621 8263 3624
rect 8205 3615 8263 3621
rect 9766 3612 9772 3664
rect 9824 3652 9830 3664
rect 9824 3624 10824 3652
rect 9824 3612 9830 3624
rect 2409 3587 2467 3593
rect 2409 3553 2421 3587
rect 2455 3584 2467 3587
rect 3050 3584 3056 3596
rect 2455 3556 3056 3584
rect 2455 3553 2467 3556
rect 2409 3547 2467 3553
rect 3050 3544 3056 3556
rect 3108 3544 3114 3596
rect 3789 3587 3847 3593
rect 3789 3584 3801 3587
rect 3344 3556 3801 3584
rect 2498 3476 2504 3528
rect 2556 3516 2562 3528
rect 2593 3519 2651 3525
rect 2593 3516 2605 3519
rect 2556 3488 2605 3516
rect 2556 3476 2562 3488
rect 2593 3485 2605 3488
rect 2639 3516 2651 3519
rect 3344 3516 3372 3556
rect 3789 3553 3801 3556
rect 3835 3553 3847 3587
rect 3789 3547 3847 3553
rect 4525 3587 4583 3593
rect 4525 3553 4537 3587
rect 4571 3584 4583 3587
rect 4706 3584 4712 3596
rect 4571 3556 4712 3584
rect 4571 3553 4583 3556
rect 4525 3547 4583 3553
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 5074 3544 5080 3596
rect 5132 3584 5138 3596
rect 5534 3584 5540 3596
rect 5132 3556 5540 3584
rect 5132 3544 5138 3556
rect 5534 3544 5540 3556
rect 5592 3544 5598 3596
rect 5721 3587 5779 3593
rect 5721 3553 5733 3587
rect 5767 3584 5779 3587
rect 5810 3584 5816 3596
rect 5767 3556 5816 3584
rect 5767 3553 5779 3556
rect 5721 3547 5779 3553
rect 5810 3544 5816 3556
rect 5868 3544 5874 3596
rect 5988 3587 6046 3593
rect 5988 3553 6000 3587
rect 6034 3584 6046 3587
rect 6822 3584 6828 3596
rect 6034 3556 6828 3584
rect 6034 3553 6046 3556
rect 5988 3547 6046 3553
rect 6822 3544 6828 3556
rect 6880 3584 6886 3596
rect 6880 3556 7972 3584
rect 6880 3544 6886 3556
rect 3510 3516 3516 3528
rect 2639 3488 3372 3516
rect 3471 3488 3516 3516
rect 2639 3485 2651 3488
rect 2593 3479 2651 3485
rect 3510 3476 3516 3488
rect 3568 3516 3574 3528
rect 7944 3525 7972 3556
rect 8754 3544 8760 3596
rect 8812 3584 8818 3596
rect 8941 3587 8999 3593
rect 8941 3584 8953 3587
rect 8812 3556 8953 3584
rect 8812 3544 8818 3556
rect 8941 3553 8953 3556
rect 8987 3553 8999 3587
rect 8941 3547 8999 3553
rect 9033 3587 9091 3593
rect 9033 3553 9045 3587
rect 9079 3584 9091 3587
rect 9398 3584 9404 3596
rect 9079 3556 9404 3584
rect 9079 3553 9091 3556
rect 9033 3547 9091 3553
rect 4617 3519 4675 3525
rect 4617 3516 4629 3519
rect 3568 3488 4629 3516
rect 3568 3476 3574 3488
rect 4617 3485 4629 3488
rect 4663 3485 4675 3519
rect 4617 3479 4675 3485
rect 7837 3519 7895 3525
rect 7837 3485 7849 3519
rect 7883 3485 7895 3519
rect 7837 3479 7895 3485
rect 7929 3519 7987 3525
rect 7929 3485 7941 3519
rect 7975 3516 7987 3519
rect 8202 3516 8208 3528
rect 7975 3488 8208 3516
rect 7975 3485 7987 3488
rect 7929 3479 7987 3485
rect 7852 3448 7880 3479
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 8386 3476 8392 3528
rect 8444 3516 8450 3528
rect 8481 3519 8539 3525
rect 8481 3516 8493 3519
rect 8444 3488 8493 3516
rect 8444 3476 8450 3488
rect 8481 3485 8493 3488
rect 8527 3516 8539 3519
rect 9048 3516 9076 3547
rect 9398 3544 9404 3556
rect 9456 3544 9462 3596
rect 10045 3587 10103 3593
rect 10045 3553 10057 3587
rect 10091 3584 10103 3587
rect 10226 3584 10232 3596
rect 10091 3556 10232 3584
rect 10091 3553 10103 3556
rect 10045 3547 10103 3553
rect 10226 3544 10232 3556
rect 10284 3544 10290 3596
rect 10796 3593 10824 3624
rect 10781 3587 10839 3593
rect 10781 3553 10793 3587
rect 10827 3553 10839 3587
rect 10888 3584 10916 3692
rect 11514 3680 11520 3692
rect 11572 3680 11578 3732
rect 11882 3720 11888 3732
rect 11843 3692 11888 3720
rect 11882 3680 11888 3692
rect 11940 3680 11946 3732
rect 11977 3723 12035 3729
rect 11977 3689 11989 3723
rect 12023 3720 12035 3723
rect 13998 3720 14004 3732
rect 12023 3692 13860 3720
rect 13911 3692 14004 3720
rect 12023 3689 12035 3692
rect 11977 3683 12035 3689
rect 11054 3652 11060 3664
rect 11015 3624 11060 3652
rect 11054 3612 11060 3624
rect 11112 3612 11118 3664
rect 12894 3652 12900 3664
rect 12855 3624 12900 3652
rect 12894 3612 12900 3624
rect 12952 3612 12958 3664
rect 13832 3652 13860 3692
rect 13998 3680 14004 3692
rect 14056 3720 14062 3732
rect 15194 3720 15200 3732
rect 14056 3692 15200 3720
rect 14056 3680 14062 3692
rect 15194 3680 15200 3692
rect 15252 3680 15258 3732
rect 15378 3720 15384 3732
rect 15339 3692 15384 3720
rect 15378 3680 15384 3692
rect 15436 3680 15442 3732
rect 15746 3680 15752 3732
rect 15804 3720 15810 3732
rect 16114 3720 16120 3732
rect 15804 3692 16120 3720
rect 15804 3680 15810 3692
rect 16114 3680 16120 3692
rect 16172 3680 16178 3732
rect 17310 3720 17316 3732
rect 17271 3692 17316 3720
rect 17310 3680 17316 3692
rect 17368 3680 17374 3732
rect 17402 3680 17408 3732
rect 17460 3720 17466 3732
rect 17865 3723 17923 3729
rect 17865 3720 17877 3723
rect 17460 3692 17877 3720
rect 17460 3680 17466 3692
rect 17865 3689 17877 3692
rect 17911 3689 17923 3723
rect 17865 3683 17923 3689
rect 18233 3723 18291 3729
rect 18233 3689 18245 3723
rect 18279 3720 18291 3723
rect 19058 3720 19064 3732
rect 18279 3692 19064 3720
rect 18279 3689 18291 3692
rect 18233 3683 18291 3689
rect 19058 3680 19064 3692
rect 19116 3680 19122 3732
rect 19613 3723 19671 3729
rect 19613 3689 19625 3723
rect 19659 3720 19671 3723
rect 20070 3720 20076 3732
rect 19659 3692 20076 3720
rect 19659 3689 19671 3692
rect 19613 3683 19671 3689
rect 20070 3680 20076 3692
rect 20128 3680 20134 3732
rect 14090 3652 14096 3664
rect 13832 3624 14096 3652
rect 14090 3612 14096 3624
rect 14148 3612 14154 3664
rect 15102 3612 15108 3664
rect 15160 3652 15166 3664
rect 16393 3655 16451 3661
rect 16393 3652 16405 3655
rect 15160 3624 16405 3652
rect 15160 3612 15166 3624
rect 16393 3621 16405 3624
rect 16439 3621 16451 3655
rect 16393 3615 16451 3621
rect 17221 3655 17279 3661
rect 17221 3621 17233 3655
rect 17267 3652 17279 3655
rect 17494 3652 17500 3664
rect 17267 3624 17500 3652
rect 17267 3621 17279 3624
rect 17221 3615 17279 3621
rect 17494 3612 17500 3624
rect 17552 3612 17558 3664
rect 17681 3655 17739 3661
rect 17681 3621 17693 3655
rect 17727 3652 17739 3655
rect 17954 3652 17960 3664
rect 17727 3624 17960 3652
rect 17727 3621 17739 3624
rect 17681 3615 17739 3621
rect 17954 3612 17960 3624
rect 18012 3612 18018 3664
rect 18156 3624 18359 3652
rect 11882 3584 11888 3596
rect 10888 3556 11888 3584
rect 10781 3547 10839 3553
rect 11882 3544 11888 3556
rect 11940 3544 11946 3596
rect 12986 3584 12992 3596
rect 12947 3556 12992 3584
rect 12986 3544 12992 3556
rect 13044 3544 13050 3596
rect 13538 3544 13544 3596
rect 13596 3584 13602 3596
rect 13909 3587 13967 3593
rect 13909 3584 13921 3587
rect 13596 3556 13921 3584
rect 13596 3544 13602 3556
rect 13909 3553 13921 3556
rect 13955 3553 13967 3587
rect 14550 3584 14556 3596
rect 14511 3556 14556 3584
rect 13909 3547 13967 3553
rect 14550 3544 14556 3556
rect 14608 3544 14614 3596
rect 15378 3544 15384 3596
rect 15436 3584 15442 3596
rect 15749 3587 15807 3593
rect 15749 3584 15761 3587
rect 15436 3556 15761 3584
rect 15436 3544 15442 3556
rect 15749 3553 15761 3556
rect 15795 3553 15807 3587
rect 15749 3547 15807 3553
rect 15841 3587 15899 3593
rect 15841 3553 15853 3587
rect 15887 3584 15899 3587
rect 15887 3556 16988 3584
rect 15887 3553 15899 3556
rect 15841 3547 15899 3553
rect 8527 3488 9076 3516
rect 9217 3519 9275 3525
rect 8527 3485 8539 3488
rect 8481 3479 8539 3485
rect 9217 3485 9229 3519
rect 9263 3516 9275 3519
rect 9306 3516 9312 3528
rect 9263 3488 9312 3516
rect 9263 3485 9275 3488
rect 9217 3479 9275 3485
rect 9306 3476 9312 3488
rect 9364 3516 9370 3528
rect 10137 3519 10195 3525
rect 9364 3488 9904 3516
rect 9364 3476 9370 3488
rect 9677 3451 9735 3457
rect 9677 3448 9689 3451
rect 7852 3420 9689 3448
rect 9677 3417 9689 3420
rect 9723 3417 9735 3451
rect 9677 3411 9735 3417
rect 3789 3383 3847 3389
rect 3789 3349 3801 3383
rect 3835 3380 3847 3383
rect 5718 3380 5724 3392
rect 3835 3352 5724 3380
rect 3835 3349 3847 3352
rect 3789 3343 3847 3349
rect 5718 3340 5724 3352
rect 5776 3340 5782 3392
rect 6638 3340 6644 3392
rect 6696 3380 6702 3392
rect 8205 3383 8263 3389
rect 8205 3380 8217 3383
rect 6696 3352 8217 3380
rect 6696 3340 6702 3352
rect 8205 3349 8217 3352
rect 8251 3349 8263 3383
rect 9876 3380 9904 3488
rect 10137 3485 10149 3519
rect 10183 3485 10195 3519
rect 10137 3479 10195 3485
rect 10152 3448 10180 3479
rect 10318 3476 10324 3528
rect 10376 3516 10382 3528
rect 10502 3516 10508 3528
rect 10376 3488 10421 3516
rect 10463 3488 10508 3516
rect 10376 3476 10382 3488
rect 10502 3476 10508 3488
rect 10560 3476 10566 3528
rect 11790 3476 11796 3528
rect 11848 3516 11854 3528
rect 12161 3519 12219 3525
rect 12161 3516 12173 3519
rect 11848 3488 12173 3516
rect 11848 3476 11854 3488
rect 12161 3485 12173 3488
rect 12207 3516 12219 3519
rect 13081 3519 13139 3525
rect 13081 3516 13093 3519
rect 12207 3488 13093 3516
rect 12207 3485 12219 3488
rect 12161 3479 12219 3485
rect 13081 3485 13093 3488
rect 13127 3485 13139 3519
rect 13081 3479 13139 3485
rect 13722 3476 13728 3528
rect 13780 3516 13786 3528
rect 14090 3516 14096 3528
rect 13780 3488 14096 3516
rect 13780 3476 13786 3488
rect 14090 3476 14096 3488
rect 14148 3476 14154 3528
rect 16025 3519 16083 3525
rect 16025 3485 16037 3519
rect 16071 3516 16083 3519
rect 16482 3516 16488 3528
rect 16071 3488 16488 3516
rect 16071 3485 16083 3488
rect 16025 3479 16083 3485
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 16960 3516 16988 3556
rect 17034 3544 17040 3596
rect 17092 3584 17098 3596
rect 18156 3584 18184 3624
rect 17092 3556 18184 3584
rect 18331 3584 18359 3624
rect 18506 3612 18512 3664
rect 18564 3652 18570 3664
rect 19153 3655 19211 3661
rect 19153 3652 19165 3655
rect 18564 3624 19165 3652
rect 18564 3612 18570 3624
rect 19153 3621 19165 3624
rect 19199 3621 19211 3655
rect 19153 3615 19211 3621
rect 19334 3612 19340 3664
rect 19392 3652 19398 3664
rect 20806 3652 20812 3664
rect 19392 3624 20812 3652
rect 19392 3612 19398 3624
rect 20806 3612 20812 3624
rect 20864 3612 20870 3664
rect 18877 3587 18935 3593
rect 18877 3584 18889 3587
rect 18331 3556 18889 3584
rect 17092 3544 17098 3556
rect 18877 3553 18889 3556
rect 18923 3553 18935 3587
rect 18877 3547 18935 3553
rect 19610 3544 19616 3596
rect 19668 3584 19674 3596
rect 19981 3587 20039 3593
rect 19981 3584 19993 3587
rect 19668 3556 19993 3584
rect 19668 3544 19674 3556
rect 19981 3553 19993 3556
rect 20027 3553 20039 3587
rect 19981 3547 20039 3553
rect 17310 3516 17316 3528
rect 16960 3488 17316 3516
rect 17310 3476 17316 3488
rect 17368 3476 17374 3528
rect 17494 3516 17500 3528
rect 17407 3488 17500 3516
rect 17494 3476 17500 3488
rect 17552 3516 17558 3528
rect 17681 3519 17739 3525
rect 17681 3516 17693 3519
rect 17552 3488 17693 3516
rect 17552 3476 17558 3488
rect 17681 3485 17693 3488
rect 17727 3485 17739 3519
rect 17681 3479 17739 3485
rect 17954 3476 17960 3528
rect 18012 3516 18018 3528
rect 18325 3519 18383 3525
rect 18325 3516 18337 3519
rect 18012 3488 18337 3516
rect 18012 3476 18018 3488
rect 18325 3485 18337 3488
rect 18371 3485 18383 3519
rect 18325 3479 18383 3485
rect 18509 3519 18567 3525
rect 18509 3485 18521 3519
rect 18555 3516 18567 3519
rect 18690 3516 18696 3528
rect 18555 3488 18696 3516
rect 18555 3485 18567 3488
rect 18509 3479 18567 3485
rect 18690 3476 18696 3488
rect 18748 3476 18754 3528
rect 19334 3476 19340 3528
rect 19392 3516 19398 3528
rect 19702 3516 19708 3528
rect 19392 3488 19708 3516
rect 19392 3476 19398 3488
rect 19702 3476 19708 3488
rect 19760 3476 19766 3528
rect 19794 3476 19800 3528
rect 19852 3516 19858 3528
rect 20073 3519 20131 3525
rect 20073 3516 20085 3519
rect 19852 3488 20085 3516
rect 19852 3476 19858 3488
rect 20073 3485 20085 3488
rect 20119 3485 20131 3519
rect 20073 3479 20131 3485
rect 20257 3519 20315 3525
rect 20257 3485 20269 3519
rect 20303 3516 20315 3519
rect 20530 3516 20536 3528
rect 20303 3488 20536 3516
rect 20303 3485 20315 3488
rect 20257 3479 20315 3485
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 10520 3448 10548 3476
rect 10152 3420 10548 3448
rect 10594 3408 10600 3460
rect 10652 3448 10658 3460
rect 11606 3448 11612 3460
rect 10652 3420 11612 3448
rect 10652 3408 10658 3420
rect 11606 3408 11612 3420
rect 11664 3408 11670 3460
rect 12526 3448 12532 3460
rect 12487 3420 12532 3448
rect 12526 3408 12532 3420
rect 12584 3408 12590 3460
rect 13541 3451 13599 3457
rect 13541 3417 13553 3451
rect 13587 3448 13599 3451
rect 14274 3448 14280 3460
rect 13587 3420 14280 3448
rect 13587 3417 13599 3420
rect 13541 3411 13599 3417
rect 14274 3408 14280 3420
rect 14332 3408 14338 3460
rect 14826 3408 14832 3460
rect 14884 3448 14890 3460
rect 14884 3420 17540 3448
rect 14884 3408 14890 3420
rect 10318 3380 10324 3392
rect 9876 3352 10324 3380
rect 8205 3343 8263 3349
rect 10318 3340 10324 3352
rect 10376 3340 10382 3392
rect 13998 3340 14004 3392
rect 14056 3380 14062 3392
rect 14737 3383 14795 3389
rect 14737 3380 14749 3383
rect 14056 3352 14749 3380
rect 14056 3340 14062 3352
rect 14737 3349 14749 3352
rect 14783 3349 14795 3383
rect 14737 3343 14795 3349
rect 16853 3383 16911 3389
rect 16853 3349 16865 3383
rect 16899 3380 16911 3383
rect 17402 3380 17408 3392
rect 16899 3352 17408 3380
rect 16899 3349 16911 3352
rect 16853 3343 16911 3349
rect 17402 3340 17408 3352
rect 17460 3340 17466 3392
rect 17512 3380 17540 3420
rect 17586 3408 17592 3460
rect 17644 3448 17650 3460
rect 17644 3420 20392 3448
rect 17644 3408 17650 3420
rect 19334 3380 19340 3392
rect 17512 3352 19340 3380
rect 19334 3340 19340 3352
rect 19392 3340 19398 3392
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 19702 3380 19708 3392
rect 19484 3352 19708 3380
rect 19484 3340 19490 3352
rect 19702 3340 19708 3352
rect 19760 3340 19766 3392
rect 20364 3380 20392 3420
rect 20438 3408 20444 3460
rect 20496 3448 20502 3460
rect 21634 3448 21640 3460
rect 20496 3420 21640 3448
rect 20496 3408 20502 3420
rect 21634 3408 21640 3420
rect 21692 3408 21698 3460
rect 21174 3380 21180 3392
rect 20364 3352 21180 3380
rect 21174 3340 21180 3352
rect 21232 3340 21238 3392
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 2038 3136 2044 3188
rect 2096 3176 2102 3188
rect 2133 3179 2191 3185
rect 2133 3176 2145 3179
rect 2096 3148 2145 3176
rect 2096 3136 2102 3148
rect 2133 3145 2145 3148
rect 2179 3145 2191 3179
rect 2133 3139 2191 3145
rect 2682 3136 2688 3188
rect 2740 3176 2746 3188
rect 2740 3148 3188 3176
rect 2740 3136 2746 3148
rect 2590 3000 2596 3052
rect 2648 3040 2654 3052
rect 2685 3043 2743 3049
rect 2685 3040 2697 3043
rect 2648 3012 2697 3040
rect 2648 3000 2654 3012
rect 2685 3009 2697 3012
rect 2731 3009 2743 3043
rect 2685 3003 2743 3009
rect 1486 2932 1492 2984
rect 1544 2972 1550 2984
rect 3160 2981 3188 3148
rect 3326 3136 3332 3188
rect 3384 3176 3390 3188
rect 3384 3148 4200 3176
rect 3384 3136 3390 3148
rect 4172 3040 4200 3148
rect 4246 3136 4252 3188
rect 4304 3176 4310 3188
rect 4525 3179 4583 3185
rect 4525 3176 4537 3179
rect 4304 3148 4537 3176
rect 4304 3136 4310 3148
rect 4525 3145 4537 3148
rect 4571 3176 4583 3179
rect 6086 3176 6092 3188
rect 4571 3148 4660 3176
rect 4571 3145 4583 3148
rect 4525 3139 4583 3145
rect 4632 3120 4660 3148
rect 4724 3148 6092 3176
rect 4614 3068 4620 3120
rect 4672 3068 4678 3120
rect 4724 3040 4752 3148
rect 6086 3136 6092 3148
rect 6144 3136 6150 3188
rect 6181 3179 6239 3185
rect 6181 3145 6193 3179
rect 6227 3176 6239 3179
rect 7466 3176 7472 3188
rect 6227 3148 7472 3176
rect 6227 3145 6239 3148
rect 6181 3139 6239 3145
rect 7466 3136 7472 3148
rect 7524 3136 7530 3188
rect 7558 3136 7564 3188
rect 7616 3176 7622 3188
rect 8202 3176 8208 3188
rect 7616 3148 8208 3176
rect 7616 3136 7622 3148
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 8754 3136 8760 3188
rect 8812 3176 8818 3188
rect 10134 3176 10140 3188
rect 8812 3148 9996 3176
rect 10095 3148 10140 3176
rect 8812 3136 8818 3148
rect 9968 3108 9996 3148
rect 10134 3136 10140 3148
rect 10192 3136 10198 3188
rect 10686 3176 10692 3188
rect 10428 3148 10692 3176
rect 10428 3108 10456 3148
rect 10686 3136 10692 3148
rect 10744 3136 10750 3188
rect 11790 3176 11796 3188
rect 11751 3148 11796 3176
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 12434 3136 12440 3188
rect 12492 3176 12498 3188
rect 12492 3148 12537 3176
rect 12492 3136 12498 3148
rect 13170 3136 13176 3188
rect 13228 3176 13234 3188
rect 14461 3179 14519 3185
rect 13228 3148 13952 3176
rect 13228 3136 13234 3148
rect 9968 3080 10456 3108
rect 11882 3068 11888 3120
rect 11940 3108 11946 3120
rect 13814 3108 13820 3120
rect 11940 3080 13820 3108
rect 11940 3068 11946 3080
rect 13814 3068 13820 3080
rect 13872 3068 13878 3120
rect 13924 3108 13952 3148
rect 14461 3145 14473 3179
rect 14507 3176 14519 3179
rect 14642 3176 14648 3188
rect 14507 3148 14648 3176
rect 14507 3145 14519 3148
rect 14461 3139 14519 3145
rect 14642 3136 14648 3148
rect 14700 3136 14706 3188
rect 15470 3176 15476 3188
rect 15431 3148 15476 3176
rect 15470 3136 15476 3148
rect 15528 3136 15534 3188
rect 18417 3179 18475 3185
rect 18417 3145 18429 3179
rect 18463 3176 18475 3179
rect 20622 3176 20628 3188
rect 18463 3148 20628 3176
rect 18463 3145 18475 3148
rect 18417 3139 18475 3145
rect 20622 3136 20628 3148
rect 20680 3136 20686 3188
rect 16945 3111 17003 3117
rect 13924 3080 14872 3108
rect 4172 3012 4752 3040
rect 5810 3000 5816 3052
rect 5868 3040 5874 3052
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 5868 3012 6837 3040
rect 5868 3000 5874 3012
rect 6825 3009 6837 3012
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 11606 3000 11612 3052
rect 11664 3040 11670 3052
rect 12158 3040 12164 3052
rect 11664 3012 12164 3040
rect 11664 3000 11670 3012
rect 12158 3000 12164 3012
rect 12216 3000 12222 3052
rect 12986 3040 12992 3052
rect 12947 3012 12992 3040
rect 12986 3000 12992 3012
rect 13044 3040 13050 3052
rect 14001 3043 14059 3049
rect 14001 3040 14013 3043
rect 13044 3012 14013 3040
rect 13044 3000 13050 3012
rect 14001 3009 14013 3012
rect 14047 3040 14059 3043
rect 14090 3040 14096 3052
rect 14047 3012 14096 3040
rect 14047 3009 14059 3012
rect 14001 3003 14059 3009
rect 14090 3000 14096 3012
rect 14148 3000 14154 3052
rect 2501 2975 2559 2981
rect 2501 2972 2513 2975
rect 1544 2944 2513 2972
rect 1544 2932 1550 2944
rect 2501 2941 2513 2944
rect 2547 2941 2559 2975
rect 2501 2935 2559 2941
rect 3145 2975 3203 2981
rect 3145 2941 3157 2975
rect 3191 2972 3203 2975
rect 4801 2975 4859 2981
rect 4801 2972 4813 2975
rect 3191 2944 4813 2972
rect 3191 2941 3203 2944
rect 3145 2935 3203 2941
rect 4801 2941 4813 2944
rect 4847 2972 4859 2975
rect 5828 2972 5856 3000
rect 8386 2972 8392 2984
rect 4847 2944 5856 2972
rect 7024 2944 8392 2972
rect 4847 2941 4859 2944
rect 4801 2935 4859 2941
rect 1026 2864 1032 2916
rect 1084 2904 1090 2916
rect 2222 2904 2228 2916
rect 1084 2876 2228 2904
rect 1084 2864 1090 2876
rect 2222 2864 2228 2876
rect 2280 2904 2286 2916
rect 3412 2907 3470 2913
rect 2280 2876 3372 2904
rect 2280 2864 2286 2876
rect 2593 2839 2651 2845
rect 2593 2805 2605 2839
rect 2639 2836 2651 2839
rect 3142 2836 3148 2848
rect 2639 2808 3148 2836
rect 2639 2805 2651 2808
rect 2593 2799 2651 2805
rect 3142 2796 3148 2808
rect 3200 2796 3206 2848
rect 3344 2836 3372 2876
rect 3412 2873 3424 2907
rect 3458 2904 3470 2907
rect 3510 2904 3516 2916
rect 3458 2876 3516 2904
rect 3458 2873 3470 2876
rect 3412 2867 3470 2873
rect 3510 2864 3516 2876
rect 3568 2864 3574 2916
rect 4154 2864 4160 2916
rect 4212 2904 4218 2916
rect 5046 2907 5104 2913
rect 5046 2904 5058 2907
rect 4212 2876 5058 2904
rect 4212 2864 4218 2876
rect 5046 2873 5058 2876
rect 5092 2873 5104 2907
rect 5046 2867 5104 2873
rect 5534 2864 5540 2916
rect 5592 2904 5598 2916
rect 5994 2904 6000 2916
rect 5592 2876 6000 2904
rect 5592 2864 5598 2876
rect 5994 2864 6000 2876
rect 6052 2864 6058 2916
rect 7024 2904 7052 2944
rect 8386 2932 8392 2944
rect 8444 2932 8450 2984
rect 8478 2932 8484 2984
rect 8536 2972 8542 2984
rect 8757 2975 8815 2981
rect 8757 2972 8769 2975
rect 8536 2944 8769 2972
rect 8536 2932 8542 2944
rect 8757 2941 8769 2944
rect 8803 2972 8815 2975
rect 10413 2975 10471 2981
rect 10413 2972 10425 2975
rect 8803 2944 10425 2972
rect 8803 2941 8815 2944
rect 8757 2935 8815 2941
rect 10413 2941 10425 2944
rect 10459 2941 10471 2975
rect 10413 2935 10471 2941
rect 10680 2975 10738 2981
rect 10680 2941 10692 2975
rect 10726 2972 10738 2975
rect 11698 2972 11704 2984
rect 10726 2944 11704 2972
rect 10726 2941 10738 2944
rect 10680 2935 10738 2941
rect 11698 2932 11704 2944
rect 11756 2932 11762 2984
rect 12894 2972 12900 2984
rect 12855 2944 12900 2972
rect 12894 2932 12900 2944
rect 12952 2932 12958 2984
rect 14734 2972 14740 2984
rect 13004 2944 14740 2972
rect 7098 2913 7104 2916
rect 6196 2876 7052 2904
rect 6196 2836 6224 2876
rect 7092 2867 7104 2913
rect 7156 2904 7162 2916
rect 7156 2876 7192 2904
rect 7098 2864 7104 2867
rect 7156 2864 7162 2876
rect 7466 2864 7472 2916
rect 7524 2904 7530 2916
rect 8662 2904 8668 2916
rect 7524 2876 8668 2904
rect 7524 2864 7530 2876
rect 8662 2864 8668 2876
rect 8720 2864 8726 2916
rect 9030 2913 9036 2916
rect 9024 2904 9036 2913
rect 8991 2876 9036 2904
rect 9024 2867 9036 2876
rect 9030 2864 9036 2867
rect 9088 2864 9094 2916
rect 10226 2864 10232 2916
rect 10284 2904 10290 2916
rect 12805 2907 12863 2913
rect 12805 2904 12817 2907
rect 10284 2876 12817 2904
rect 10284 2864 10290 2876
rect 12805 2873 12817 2876
rect 12851 2873 12863 2907
rect 12805 2867 12863 2873
rect 3344 2808 6224 2836
rect 6270 2796 6276 2848
rect 6328 2836 6334 2848
rect 8478 2836 8484 2848
rect 6328 2808 8484 2836
rect 6328 2796 6334 2808
rect 8478 2796 8484 2808
rect 8536 2796 8542 2848
rect 9398 2796 9404 2848
rect 9456 2836 9462 2848
rect 13004 2836 13032 2944
rect 14734 2932 14740 2944
rect 14792 2932 14798 2984
rect 14844 2981 14872 3080
rect 16945 3077 16957 3111
rect 16991 3108 17003 3111
rect 19518 3108 19524 3120
rect 16991 3080 19524 3108
rect 16991 3077 17003 3080
rect 16945 3071 17003 3077
rect 19518 3068 19524 3080
rect 19576 3068 19582 3120
rect 20530 3108 20536 3120
rect 19720 3080 20536 3108
rect 15102 3040 15108 3052
rect 15063 3012 15108 3040
rect 15102 3000 15108 3012
rect 15160 3000 15166 3052
rect 15286 3000 15292 3052
rect 15344 3040 15350 3052
rect 16114 3040 16120 3052
rect 15344 3012 15884 3040
rect 16075 3012 16120 3040
rect 15344 3000 15350 3012
rect 15856 2981 15884 3012
rect 16114 3000 16120 3012
rect 16172 3000 16178 3052
rect 17494 3040 17500 3052
rect 17455 3012 17500 3040
rect 17494 3000 17500 3012
rect 17552 3000 17558 3052
rect 17586 3000 17592 3052
rect 17644 3040 17650 3052
rect 18877 3043 18935 3049
rect 18877 3040 18889 3043
rect 17644 3012 18889 3040
rect 17644 3000 17650 3012
rect 18877 3009 18889 3012
rect 18923 3009 18935 3043
rect 18877 3003 18935 3009
rect 19061 3043 19119 3049
rect 19061 3009 19073 3043
rect 19107 3040 19119 3043
rect 19334 3040 19340 3052
rect 19107 3012 19340 3040
rect 19107 3009 19119 3012
rect 19061 3003 19119 3009
rect 19334 3000 19340 3012
rect 19392 3000 19398 3052
rect 19720 3040 19748 3080
rect 19886 3040 19892 3052
rect 19444 3012 19748 3040
rect 19847 3012 19892 3040
rect 14829 2975 14887 2981
rect 14829 2941 14841 2975
rect 14875 2941 14887 2975
rect 14829 2935 14887 2941
rect 15841 2975 15899 2981
rect 15841 2941 15853 2975
rect 15887 2941 15899 2975
rect 15841 2935 15899 2941
rect 17405 2975 17463 2981
rect 17405 2941 17417 2975
rect 17451 2972 17463 2975
rect 18322 2972 18328 2984
rect 17451 2944 18328 2972
rect 17451 2941 17463 2944
rect 17405 2935 17463 2941
rect 18322 2932 18328 2944
rect 18380 2932 18386 2984
rect 19242 2932 19248 2984
rect 19300 2972 19306 2984
rect 19444 2972 19472 3012
rect 19886 3000 19892 3012
rect 19944 3000 19950 3052
rect 19996 3049 20024 3080
rect 20530 3068 20536 3080
rect 20588 3068 20594 3120
rect 19981 3043 20039 3049
rect 19981 3009 19993 3043
rect 20027 3009 20039 3043
rect 19981 3003 20039 3009
rect 19794 2972 19800 2984
rect 19300 2944 19472 2972
rect 19755 2944 19800 2972
rect 19300 2932 19306 2944
rect 19794 2932 19800 2944
rect 19852 2932 19858 2984
rect 20254 2932 20260 2984
rect 20312 2972 20318 2984
rect 20533 2975 20591 2981
rect 20533 2972 20545 2975
rect 20312 2944 20545 2972
rect 20312 2932 20318 2944
rect 20533 2941 20545 2944
rect 20579 2941 20591 2975
rect 20533 2935 20591 2941
rect 14366 2864 14372 2916
rect 14424 2904 14430 2916
rect 14921 2907 14979 2913
rect 14921 2904 14933 2907
rect 14424 2876 14933 2904
rect 14424 2864 14430 2876
rect 14921 2873 14933 2876
rect 14967 2904 14979 2907
rect 15010 2904 15016 2916
rect 14967 2876 15016 2904
rect 14967 2873 14979 2876
rect 14921 2867 14979 2873
rect 15010 2864 15016 2876
rect 15068 2864 15074 2916
rect 15286 2864 15292 2916
rect 15344 2904 15350 2916
rect 15933 2907 15991 2913
rect 15933 2904 15945 2907
rect 15344 2876 15945 2904
rect 15344 2864 15350 2876
rect 15933 2873 15945 2876
rect 15979 2873 15991 2907
rect 16758 2904 16764 2916
rect 15933 2867 15991 2873
rect 16040 2876 16764 2904
rect 9456 2808 13032 2836
rect 13449 2839 13507 2845
rect 9456 2796 9462 2808
rect 13449 2805 13461 2839
rect 13495 2836 13507 2839
rect 13538 2836 13544 2848
rect 13495 2808 13544 2836
rect 13495 2805 13507 2808
rect 13449 2799 13507 2805
rect 13538 2796 13544 2808
rect 13596 2796 13602 2848
rect 13814 2836 13820 2848
rect 13775 2808 13820 2836
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 13906 2796 13912 2848
rect 13964 2836 13970 2848
rect 16040 2836 16068 2876
rect 16758 2864 16764 2876
rect 16816 2864 16822 2916
rect 17313 2907 17371 2913
rect 17313 2873 17325 2907
rect 17359 2904 17371 2907
rect 17862 2904 17868 2916
rect 17359 2876 17868 2904
rect 17359 2873 17371 2876
rect 17313 2867 17371 2873
rect 17862 2864 17868 2876
rect 17920 2864 17926 2916
rect 18506 2904 18512 2916
rect 18340 2876 18512 2904
rect 13964 2808 16068 2836
rect 13964 2796 13970 2808
rect 16298 2796 16304 2848
rect 16356 2836 16362 2848
rect 18340 2836 18368 2876
rect 18506 2864 18512 2876
rect 18564 2864 18570 2916
rect 18785 2907 18843 2913
rect 18785 2873 18797 2907
rect 18831 2904 18843 2907
rect 18831 2876 19472 2904
rect 18831 2873 18843 2876
rect 18785 2867 18843 2873
rect 19444 2845 19472 2876
rect 16356 2808 18368 2836
rect 19429 2839 19487 2845
rect 16356 2796 16362 2808
rect 19429 2805 19441 2839
rect 19475 2805 19487 2839
rect 19429 2799 19487 2805
rect 20717 2839 20775 2845
rect 20717 2805 20729 2839
rect 20763 2836 20775 2839
rect 22094 2836 22100 2848
rect 20763 2808 22100 2836
rect 20763 2805 20775 2808
rect 20717 2799 20775 2805
rect 22094 2796 22100 2808
rect 22152 2796 22158 2848
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 2222 2632 2228 2644
rect 2183 2604 2228 2632
rect 2222 2592 2228 2604
rect 2280 2592 2286 2644
rect 2774 2632 2780 2644
rect 2735 2604 2780 2632
rect 2774 2592 2780 2604
rect 2832 2632 2838 2644
rect 3329 2635 3387 2641
rect 3329 2632 3341 2635
rect 2832 2604 3341 2632
rect 2832 2592 2838 2604
rect 3329 2601 3341 2604
rect 3375 2601 3387 2635
rect 3329 2595 3387 2601
rect 4617 2635 4675 2641
rect 4617 2601 4629 2635
rect 4663 2632 4675 2635
rect 4706 2632 4712 2644
rect 4663 2604 4712 2632
rect 4663 2601 4675 2604
rect 4617 2595 4675 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 5077 2635 5135 2641
rect 5077 2601 5089 2635
rect 5123 2632 5135 2635
rect 5166 2632 5172 2644
rect 5123 2604 5172 2632
rect 5123 2601 5135 2604
rect 5077 2595 5135 2601
rect 1946 2524 1952 2576
rect 2004 2564 2010 2576
rect 2133 2567 2191 2573
rect 2133 2564 2145 2567
rect 2004 2536 2145 2564
rect 2004 2524 2010 2536
rect 2133 2533 2145 2536
rect 2179 2564 2191 2567
rect 3142 2564 3148 2576
rect 2179 2536 3148 2564
rect 2179 2533 2191 2536
rect 2133 2527 2191 2533
rect 3142 2524 3148 2536
rect 3200 2524 3206 2576
rect 3418 2564 3424 2576
rect 3379 2536 3424 2564
rect 3418 2524 3424 2536
rect 3476 2524 3482 2576
rect 4525 2567 4583 2573
rect 4525 2533 4537 2567
rect 4571 2564 4583 2567
rect 5092 2564 5120 2595
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 5813 2635 5871 2641
rect 5813 2601 5825 2635
rect 5859 2601 5871 2635
rect 5813 2595 5871 2601
rect 4571 2536 5120 2564
rect 5828 2564 5856 2595
rect 6086 2592 6092 2644
rect 6144 2632 6150 2644
rect 6181 2635 6239 2641
rect 6181 2632 6193 2635
rect 6144 2604 6193 2632
rect 6144 2592 6150 2604
rect 6181 2601 6193 2604
rect 6227 2601 6239 2635
rect 6914 2632 6920 2644
rect 6875 2604 6920 2632
rect 6181 2595 6239 2601
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 7377 2635 7435 2641
rect 7377 2601 7389 2635
rect 7423 2632 7435 2635
rect 7929 2635 7987 2641
rect 7929 2632 7941 2635
rect 7423 2604 7941 2632
rect 7423 2601 7435 2604
rect 7377 2595 7435 2601
rect 7929 2601 7941 2604
rect 7975 2601 7987 2635
rect 7929 2595 7987 2601
rect 9309 2635 9367 2641
rect 9309 2601 9321 2635
rect 9355 2601 9367 2635
rect 10226 2632 10232 2644
rect 10187 2604 10232 2632
rect 9309 2595 9367 2601
rect 7285 2567 7343 2573
rect 7285 2564 7297 2567
rect 5828 2536 7297 2564
rect 4571 2533 4583 2536
rect 4525 2527 4583 2533
rect 7285 2533 7297 2536
rect 7331 2533 7343 2567
rect 8294 2564 8300 2576
rect 8255 2536 8300 2564
rect 7285 2527 7343 2533
rect 8294 2524 8300 2536
rect 8352 2564 8358 2576
rect 9324 2564 9352 2595
rect 10226 2592 10232 2604
rect 10284 2592 10290 2644
rect 10321 2635 10379 2641
rect 10321 2601 10333 2635
rect 10367 2632 10379 2635
rect 10686 2632 10692 2644
rect 10367 2604 10692 2632
rect 10367 2601 10379 2604
rect 10321 2595 10379 2601
rect 10686 2592 10692 2604
rect 10744 2592 10750 2644
rect 10781 2635 10839 2641
rect 10781 2601 10793 2635
rect 10827 2632 10839 2635
rect 10962 2632 10968 2644
rect 10827 2604 10968 2632
rect 10827 2601 10839 2604
rect 10781 2595 10839 2601
rect 10962 2592 10968 2604
rect 11020 2592 11026 2644
rect 12253 2635 12311 2641
rect 12253 2601 12265 2635
rect 12299 2632 12311 2635
rect 12342 2632 12348 2644
rect 12299 2604 12348 2632
rect 12299 2601 12311 2604
rect 12253 2595 12311 2601
rect 12342 2592 12348 2604
rect 12400 2592 12406 2644
rect 12713 2635 12771 2641
rect 12713 2601 12725 2635
rect 12759 2632 12771 2635
rect 12802 2632 12808 2644
rect 12759 2604 12808 2632
rect 12759 2601 12771 2604
rect 12713 2595 12771 2601
rect 12802 2592 12808 2604
rect 12860 2592 12866 2644
rect 13173 2635 13231 2641
rect 13173 2601 13185 2635
rect 13219 2632 13231 2635
rect 13446 2632 13452 2644
rect 13219 2604 13452 2632
rect 13219 2601 13231 2604
rect 13173 2595 13231 2601
rect 13446 2592 13452 2604
rect 13504 2592 13510 2644
rect 13630 2592 13636 2644
rect 13688 2632 13694 2644
rect 13725 2635 13783 2641
rect 13725 2632 13737 2635
rect 13688 2604 13737 2632
rect 13688 2592 13694 2604
rect 13725 2601 13737 2604
rect 13771 2601 13783 2635
rect 13725 2595 13783 2601
rect 13906 2592 13912 2644
rect 13964 2632 13970 2644
rect 14093 2635 14151 2641
rect 14093 2632 14105 2635
rect 13964 2604 14105 2632
rect 13964 2592 13970 2604
rect 14093 2601 14105 2604
rect 14139 2601 14151 2635
rect 14093 2595 14151 2601
rect 14185 2635 14243 2641
rect 14185 2601 14197 2635
rect 14231 2632 14243 2635
rect 15194 2632 15200 2644
rect 14231 2604 15200 2632
rect 14231 2601 14243 2604
rect 14185 2595 14243 2601
rect 10502 2564 10508 2576
rect 8352 2536 9260 2564
rect 9324 2536 10508 2564
rect 8352 2524 8358 2536
rect 4985 2499 5043 2505
rect 4985 2465 4997 2499
rect 5031 2496 5043 2499
rect 8754 2496 8760 2508
rect 5031 2468 8760 2496
rect 5031 2465 5043 2468
rect 4985 2459 5043 2465
rect 8754 2456 8760 2468
rect 8812 2456 8818 2508
rect 9125 2499 9183 2505
rect 9125 2465 9137 2499
rect 9171 2465 9183 2499
rect 9232 2496 9260 2536
rect 10502 2524 10508 2536
rect 10560 2524 10566 2576
rect 11140 2567 11198 2573
rect 11140 2533 11152 2567
rect 11186 2564 11198 2567
rect 11790 2564 11796 2576
rect 11186 2536 11796 2564
rect 11186 2533 11198 2536
rect 11140 2527 11198 2533
rect 11790 2524 11796 2536
rect 11848 2524 11854 2576
rect 12986 2564 12992 2576
rect 12176 2536 12992 2564
rect 10226 2496 10232 2508
rect 9232 2468 10232 2496
rect 9125 2459 9183 2465
rect 2409 2431 2467 2437
rect 2409 2397 2421 2431
rect 2455 2397 2467 2431
rect 3510 2428 3516 2440
rect 3471 2400 3516 2428
rect 2409 2391 2467 2397
rect 2424 2360 2452 2391
rect 3510 2388 3516 2400
rect 3568 2388 3574 2440
rect 5261 2431 5319 2437
rect 5261 2397 5273 2431
rect 5307 2428 5319 2431
rect 5718 2428 5724 2440
rect 5307 2400 5724 2428
rect 5307 2397 5319 2400
rect 5261 2391 5319 2397
rect 5718 2388 5724 2400
rect 5776 2388 5782 2440
rect 6270 2428 6276 2440
rect 6231 2400 6276 2428
rect 6270 2388 6276 2400
rect 6328 2388 6334 2440
rect 6457 2431 6515 2437
rect 6457 2397 6469 2431
rect 6503 2428 6515 2431
rect 7098 2428 7104 2440
rect 6503 2400 7104 2428
rect 6503 2397 6515 2400
rect 6457 2391 6515 2397
rect 7098 2388 7104 2400
rect 7156 2388 7162 2440
rect 7558 2428 7564 2440
rect 7519 2400 7564 2428
rect 7558 2388 7564 2400
rect 7616 2388 7622 2440
rect 7837 2431 7895 2437
rect 7837 2397 7849 2431
rect 7883 2428 7895 2431
rect 8386 2428 8392 2440
rect 7883 2400 8392 2428
rect 7883 2397 7895 2400
rect 7837 2391 7895 2397
rect 8386 2388 8392 2400
rect 8444 2388 8450 2440
rect 8481 2431 8539 2437
rect 8481 2397 8493 2431
rect 8527 2397 8539 2431
rect 9140 2428 9168 2459
rect 10226 2456 10232 2468
rect 10284 2456 10290 2508
rect 12176 2496 12204 2536
rect 12986 2524 12992 2536
rect 13044 2524 13050 2576
rect 15120 2564 15148 2604
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 15473 2635 15531 2641
rect 15473 2601 15485 2635
rect 15519 2632 15531 2635
rect 15654 2632 15660 2644
rect 15519 2604 15660 2632
rect 15519 2601 15531 2604
rect 15473 2595 15531 2601
rect 15654 2592 15660 2604
rect 15712 2592 15718 2644
rect 15930 2632 15936 2644
rect 15891 2604 15936 2632
rect 15930 2592 15936 2604
rect 15988 2592 15994 2644
rect 16022 2592 16028 2644
rect 16080 2632 16086 2644
rect 16485 2635 16543 2641
rect 16485 2632 16497 2635
rect 16080 2604 16497 2632
rect 16080 2592 16086 2604
rect 16485 2601 16497 2604
rect 16531 2601 16543 2635
rect 16942 2632 16948 2644
rect 16903 2604 16948 2632
rect 16485 2595 16543 2601
rect 16942 2592 16948 2604
rect 17000 2592 17006 2644
rect 19058 2632 19064 2644
rect 19019 2604 19064 2632
rect 19058 2592 19064 2604
rect 19116 2592 19122 2644
rect 19518 2632 19524 2644
rect 19479 2604 19524 2632
rect 19518 2592 19524 2604
rect 19576 2592 19582 2644
rect 20073 2635 20131 2641
rect 20073 2601 20085 2635
rect 20119 2601 20131 2635
rect 20438 2632 20444 2644
rect 20399 2604 20444 2632
rect 20073 2595 20131 2601
rect 15746 2564 15752 2576
rect 15120 2536 15752 2564
rect 15746 2524 15752 2536
rect 15804 2524 15810 2576
rect 19429 2567 19487 2573
rect 19429 2533 19441 2567
rect 19475 2564 19487 2567
rect 20088 2564 20116 2595
rect 20438 2592 20444 2604
rect 20496 2592 20502 2644
rect 19475 2536 20116 2564
rect 19475 2533 19487 2536
rect 19429 2527 19487 2533
rect 20530 2524 20536 2576
rect 20588 2564 20594 2576
rect 20588 2536 20668 2564
rect 20588 2524 20594 2536
rect 10520 2468 12204 2496
rect 10134 2428 10140 2440
rect 9140 2400 10140 2428
rect 8481 2391 8539 2397
rect 3050 2360 3056 2372
rect 2424 2332 3056 2360
rect 3050 2320 3056 2332
rect 3108 2320 3114 2372
rect 3142 2320 3148 2372
rect 3200 2360 3206 2372
rect 7116 2360 7144 2388
rect 8496 2360 8524 2391
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 10520 2437 10548 2468
rect 12250 2456 12256 2508
rect 12308 2496 12314 2508
rect 13081 2499 13139 2505
rect 13081 2496 13093 2499
rect 12308 2468 13093 2496
rect 12308 2456 12314 2468
rect 13081 2465 13093 2468
rect 13127 2465 13139 2499
rect 13081 2459 13139 2465
rect 13814 2456 13820 2508
rect 13872 2496 13878 2508
rect 14829 2499 14887 2505
rect 14829 2496 14841 2499
rect 13872 2468 14841 2496
rect 13872 2456 13878 2468
rect 14829 2465 14841 2468
rect 14875 2465 14887 2499
rect 14829 2459 14887 2465
rect 15102 2456 15108 2508
rect 15160 2496 15166 2508
rect 15841 2499 15899 2505
rect 15841 2496 15853 2499
rect 15160 2468 15853 2496
rect 15160 2456 15166 2468
rect 15841 2465 15853 2468
rect 15887 2465 15899 2499
rect 15841 2459 15899 2465
rect 16853 2499 16911 2505
rect 16853 2465 16865 2499
rect 16899 2496 16911 2499
rect 17218 2496 17224 2508
rect 16899 2468 17224 2496
rect 16899 2465 16911 2468
rect 16853 2459 16911 2465
rect 17218 2456 17224 2468
rect 17276 2456 17282 2508
rect 17310 2456 17316 2508
rect 17368 2496 17374 2508
rect 17497 2499 17555 2505
rect 17497 2496 17509 2499
rect 17368 2468 17509 2496
rect 17368 2456 17374 2468
rect 17497 2465 17509 2468
rect 17543 2465 17555 2499
rect 17497 2459 17555 2465
rect 17770 2456 17776 2508
rect 17828 2496 17834 2508
rect 18509 2499 18567 2505
rect 18509 2496 18521 2499
rect 17828 2468 18521 2496
rect 17828 2456 17834 2468
rect 18509 2465 18521 2468
rect 18555 2465 18567 2499
rect 18509 2459 18567 2465
rect 10505 2431 10563 2437
rect 10505 2397 10517 2431
rect 10551 2397 10563 2431
rect 10505 2391 10563 2397
rect 10873 2431 10931 2437
rect 10873 2397 10885 2431
rect 10919 2397 10931 2431
rect 13354 2428 13360 2440
rect 13315 2400 13360 2428
rect 10873 2391 10931 2397
rect 9306 2360 9312 2372
rect 3200 2332 7052 2360
rect 7116 2332 9312 2360
rect 3200 2320 3206 2332
rect 1762 2292 1768 2304
rect 1723 2264 1768 2292
rect 1762 2252 1768 2264
rect 1820 2252 1826 2304
rect 2958 2292 2964 2304
rect 2919 2264 2964 2292
rect 2958 2252 2964 2264
rect 3016 2252 3022 2304
rect 7024 2292 7052 2332
rect 9306 2320 9312 2332
rect 9364 2320 9370 2372
rect 9861 2363 9919 2369
rect 9861 2329 9873 2363
rect 9907 2360 9919 2363
rect 10781 2363 10839 2369
rect 10781 2360 10793 2363
rect 9907 2332 10793 2360
rect 9907 2329 9919 2332
rect 9861 2323 9919 2329
rect 10781 2329 10793 2332
rect 10827 2329 10839 2363
rect 10781 2323 10839 2329
rect 7837 2295 7895 2301
rect 7837 2292 7849 2295
rect 7024 2264 7849 2292
rect 7837 2261 7849 2264
rect 7883 2261 7895 2295
rect 10888 2292 10916 2391
rect 13354 2388 13360 2400
rect 13412 2388 13418 2440
rect 13906 2388 13912 2440
rect 13964 2428 13970 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 13964 2400 14289 2428
rect 13964 2388 13970 2400
rect 14277 2397 14289 2400
rect 14323 2428 14335 2431
rect 15010 2428 15016 2440
rect 14323 2400 15016 2428
rect 14323 2397 14335 2400
rect 14277 2391 14335 2397
rect 15010 2388 15016 2400
rect 15068 2388 15074 2440
rect 16025 2431 16083 2437
rect 16025 2397 16037 2431
rect 16071 2428 16083 2431
rect 16114 2428 16120 2440
rect 16071 2400 16120 2428
rect 16071 2397 16083 2400
rect 16025 2391 16083 2397
rect 13372 2360 13400 2388
rect 16040 2360 16068 2391
rect 16114 2388 16120 2400
rect 16172 2428 16178 2440
rect 17037 2431 17095 2437
rect 17037 2428 17049 2431
rect 16172 2400 17049 2428
rect 16172 2388 16178 2400
rect 17037 2397 17049 2400
rect 17083 2397 17095 2431
rect 17037 2391 17095 2397
rect 17681 2431 17739 2437
rect 17681 2397 17693 2431
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 13372 2332 16068 2360
rect 16390 2320 16396 2372
rect 16448 2360 16454 2372
rect 17696 2360 17724 2391
rect 19334 2388 19340 2440
rect 19392 2428 19398 2440
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 19392 2400 19625 2428
rect 19392 2388 19398 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 19613 2391 19671 2397
rect 20346 2388 20352 2440
rect 20404 2428 20410 2440
rect 20640 2437 20668 2536
rect 20533 2431 20591 2437
rect 20533 2428 20545 2431
rect 20404 2400 20545 2428
rect 20404 2388 20410 2400
rect 20533 2397 20545 2400
rect 20579 2397 20591 2431
rect 20533 2391 20591 2397
rect 20625 2431 20683 2437
rect 20625 2397 20637 2431
rect 20671 2397 20683 2431
rect 20625 2391 20683 2397
rect 20254 2360 20260 2372
rect 16448 2332 17724 2360
rect 18616 2332 20260 2360
rect 16448 2320 16454 2332
rect 12618 2292 12624 2304
rect 10888 2264 12624 2292
rect 7837 2255 7895 2261
rect 12618 2252 12624 2264
rect 12676 2252 12682 2304
rect 14182 2252 14188 2304
rect 14240 2292 14246 2304
rect 14918 2292 14924 2304
rect 14240 2264 14924 2292
rect 14240 2252 14246 2264
rect 14918 2252 14924 2264
rect 14976 2252 14982 2304
rect 15013 2295 15071 2301
rect 15013 2261 15025 2295
rect 15059 2292 15071 2295
rect 18616 2292 18644 2332
rect 20254 2320 20260 2332
rect 20312 2320 20318 2372
rect 15059 2264 18644 2292
rect 18693 2295 18751 2301
rect 15059 2261 15071 2264
rect 15013 2255 15071 2261
rect 18693 2261 18705 2295
rect 18739 2292 18751 2295
rect 22554 2292 22560 2304
rect 18739 2264 22560 2292
rect 18739 2261 18751 2264
rect 18693 2255 18751 2261
rect 22554 2252 22560 2264
rect 22612 2252 22618 2304
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 2866 2048 2872 2100
rect 2924 2088 2930 2100
rect 3418 2088 3424 2100
rect 2924 2060 3424 2088
rect 2924 2048 2930 2060
rect 3418 2048 3424 2060
rect 3476 2088 3482 2100
rect 6270 2088 6276 2100
rect 3476 2060 6276 2088
rect 3476 2048 3482 2060
rect 6270 2048 6276 2060
rect 6328 2088 6334 2100
rect 20162 2088 20168 2100
rect 6328 2060 20168 2088
rect 6328 2048 6334 2060
rect 20162 2048 20168 2060
rect 20220 2048 20226 2100
rect 1762 1980 1768 2032
rect 1820 2020 1826 2032
rect 15102 2020 15108 2032
rect 1820 1992 15108 2020
rect 1820 1980 1826 1992
rect 15102 1980 15108 1992
rect 15160 1980 15166 2032
rect 16850 1980 16856 2032
rect 16908 2020 16914 2032
rect 18966 2020 18972 2032
rect 16908 1992 18972 2020
rect 16908 1980 16914 1992
rect 18966 1980 18972 1992
rect 19024 1980 19030 2032
rect 2958 1912 2964 1964
rect 3016 1952 3022 1964
rect 15286 1952 15292 1964
rect 3016 1924 15292 1952
rect 3016 1912 3022 1924
rect 15286 1912 15292 1924
rect 15344 1912 15350 1964
rect 8754 1844 8760 1896
rect 8812 1884 8818 1896
rect 15194 1884 15200 1896
rect 8812 1856 15200 1884
rect 8812 1844 8818 1856
rect 15194 1844 15200 1856
rect 15252 1844 15258 1896
rect 3050 1776 3056 1828
rect 3108 1816 3114 1828
rect 3510 1816 3516 1828
rect 3108 1788 3516 1816
rect 3108 1776 3114 1788
rect 3510 1776 3516 1788
rect 3568 1816 3574 1828
rect 3568 1788 5580 1816
rect 3568 1776 3574 1788
rect 5552 1748 5580 1788
rect 8386 1776 8392 1828
rect 8444 1816 8450 1828
rect 10594 1816 10600 1828
rect 8444 1788 10600 1816
rect 8444 1776 8450 1788
rect 10594 1776 10600 1788
rect 10652 1776 10658 1828
rect 12066 1748 12072 1760
rect 5552 1720 12072 1748
rect 12066 1708 12072 1720
rect 12124 1708 12130 1760
rect 1486 1640 1492 1692
rect 1544 1680 1550 1692
rect 8846 1680 8852 1692
rect 1544 1652 8852 1680
rect 1544 1640 1550 1652
rect 8846 1640 8852 1652
rect 8904 1640 8910 1692
rect 10502 1640 10508 1692
rect 10560 1680 10566 1692
rect 16666 1680 16672 1692
rect 10560 1652 16672 1680
rect 10560 1640 10566 1652
rect 16666 1640 16672 1652
rect 16724 1640 16730 1692
rect 2406 1572 2412 1624
rect 2464 1612 2470 1624
rect 8294 1612 8300 1624
rect 2464 1584 8300 1612
rect 2464 1572 2470 1584
rect 8294 1572 8300 1584
rect 8352 1572 8358 1624
rect 3234 1300 3240 1352
rect 3292 1340 3298 1352
rect 4982 1340 4988 1352
rect 3292 1312 4988 1340
rect 3292 1300 3298 1312
rect 4982 1300 4988 1312
rect 5040 1300 5046 1352
rect 16758 1300 16764 1352
rect 16816 1340 16822 1352
rect 17954 1340 17960 1352
rect 16816 1312 17960 1340
rect 16816 1300 16822 1312
rect 17954 1300 17960 1312
rect 18012 1300 18018 1352
rect 566 1232 572 1284
rect 624 1272 630 1284
rect 7650 1272 7656 1284
rect 624 1244 7656 1272
rect 624 1232 630 1244
rect 7650 1232 7656 1244
rect 7708 1232 7714 1284
rect 13078 1096 13084 1148
rect 13136 1136 13142 1148
rect 15378 1136 15384 1148
rect 13136 1108 15384 1136
rect 13136 1096 13142 1108
rect 15378 1096 15384 1108
rect 15436 1096 15442 1148
rect 19794 552 19800 604
rect 19852 592 19858 604
rect 20990 592 20996 604
rect 19852 564 20996 592
rect 19852 552 19858 564
rect 20990 552 20996 564
rect 21048 552 21054 604
<< via1 >>
rect 3056 22176 3108 22228
rect 3700 22176 3752 22228
rect 9680 20408 9732 20460
rect 10876 20408 10928 20460
rect 16672 20408 16724 20460
rect 7380 20340 7432 20392
rect 8208 20340 8260 20392
rect 10232 20340 10284 20392
rect 17776 20340 17828 20392
rect 3608 20272 3660 20324
rect 16304 20272 16356 20324
rect 3332 20204 3384 20256
rect 15384 20204 15436 20256
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 2872 20000 2924 20052
rect 3332 20000 3384 20052
rect 3608 20043 3660 20052
rect 3608 20009 3617 20043
rect 3617 20009 3651 20043
rect 3651 20009 3660 20043
rect 3608 20000 3660 20009
rect 1860 19864 1912 19916
rect 2136 19864 2188 19916
rect 3332 19864 3384 19916
rect 5724 20000 5776 20052
rect 9772 20043 9824 20052
rect 9772 20009 9781 20043
rect 9781 20009 9815 20043
rect 9815 20009 9824 20043
rect 9772 20000 9824 20009
rect 8024 19932 8076 19984
rect 5172 19864 5224 19916
rect 6920 19907 6972 19916
rect 6920 19873 6929 19907
rect 6929 19873 6963 19907
rect 6963 19873 6972 19907
rect 6920 19864 6972 19873
rect 7748 19864 7800 19916
rect 9864 19932 9916 19984
rect 9956 19932 10008 19984
rect 13268 20000 13320 20052
rect 14464 20000 14516 20052
rect 18972 20043 19024 20052
rect 18972 20009 18981 20043
rect 18981 20009 19015 20043
rect 19015 20009 19024 20043
rect 18972 20000 19024 20009
rect 19248 20000 19300 20052
rect 8852 19907 8904 19916
rect 8852 19873 8861 19907
rect 8861 19873 8895 19907
rect 8895 19873 8904 19907
rect 8852 19864 8904 19873
rect 9680 19864 9732 19916
rect 10508 19864 10560 19916
rect 11888 19907 11940 19916
rect 11888 19873 11897 19907
rect 11897 19873 11931 19907
rect 11931 19873 11940 19907
rect 11888 19864 11940 19873
rect 13452 19907 13504 19916
rect 13452 19873 13461 19907
rect 13461 19873 13495 19907
rect 13495 19873 13504 19907
rect 13452 19864 13504 19873
rect 14280 19864 14332 19916
rect 15200 19864 15252 19916
rect 17960 19932 18012 19984
rect 2780 19728 2832 19780
rect 8208 19796 8260 19848
rect 8944 19839 8996 19848
rect 8944 19805 8953 19839
rect 8953 19805 8987 19839
rect 8987 19805 8996 19839
rect 8944 19796 8996 19805
rect 9220 19796 9272 19848
rect 10416 19839 10468 19848
rect 10416 19805 10425 19839
rect 10425 19805 10459 19839
rect 10459 19805 10468 19839
rect 10416 19796 10468 19805
rect 10692 19796 10744 19848
rect 11704 19796 11756 19848
rect 12440 19796 12492 19848
rect 13544 19839 13596 19848
rect 13544 19805 13553 19839
rect 13553 19805 13587 19839
rect 13587 19805 13596 19839
rect 13544 19796 13596 19805
rect 13728 19839 13780 19848
rect 13728 19805 13737 19839
rect 13737 19805 13771 19839
rect 13771 19805 13780 19839
rect 13728 19796 13780 19805
rect 14372 19796 14424 19848
rect 14648 19839 14700 19848
rect 14648 19805 14657 19839
rect 14657 19805 14691 19839
rect 14691 19805 14700 19839
rect 14648 19796 14700 19805
rect 15384 19796 15436 19848
rect 17408 19864 17460 19916
rect 18880 19864 18932 19916
rect 20076 19864 20128 19916
rect 20996 19864 21048 19916
rect 17040 19839 17092 19848
rect 17040 19805 17049 19839
rect 17049 19805 17083 19839
rect 17083 19805 17092 19839
rect 17040 19796 17092 19805
rect 20444 19839 20496 19848
rect 20444 19805 20453 19839
rect 20453 19805 20487 19839
rect 20487 19805 20496 19839
rect 20444 19796 20496 19805
rect 14464 19728 14516 19780
rect 18972 19728 19024 19780
rect 4712 19660 4764 19712
rect 5356 19660 5408 19712
rect 8116 19660 8168 19712
rect 8300 19660 8352 19712
rect 10416 19660 10468 19712
rect 12900 19660 12952 19712
rect 14188 19660 14240 19712
rect 18788 19660 18840 19712
rect 19892 19703 19944 19712
rect 19892 19669 19901 19703
rect 19901 19669 19935 19703
rect 19935 19669 19944 19703
rect 19892 19660 19944 19669
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 3148 19456 3200 19508
rect 3332 19456 3384 19508
rect 8024 19456 8076 19508
rect 8300 19456 8352 19508
rect 12348 19456 12400 19508
rect 12440 19456 12492 19508
rect 1676 19252 1728 19304
rect 1124 19184 1176 19236
rect 2688 19252 2740 19304
rect 2872 19295 2924 19304
rect 2872 19261 2881 19295
rect 2881 19261 2915 19295
rect 2915 19261 2924 19295
rect 2872 19252 2924 19261
rect 3056 19252 3108 19304
rect 10232 19388 10284 19440
rect 13728 19456 13780 19508
rect 19340 19499 19392 19508
rect 19340 19465 19349 19499
rect 19349 19465 19383 19499
rect 19383 19465 19392 19499
rect 19340 19456 19392 19465
rect 3516 19252 3568 19304
rect 4712 19295 4764 19304
rect 4712 19261 4721 19295
rect 4721 19261 4755 19295
rect 4755 19261 4764 19295
rect 4712 19252 4764 19261
rect 2964 19116 3016 19168
rect 3884 19116 3936 19168
rect 3976 19116 4028 19168
rect 4712 19116 4764 19168
rect 5356 19252 5408 19304
rect 6460 19252 6512 19304
rect 6736 19184 6788 19236
rect 7656 19252 7708 19304
rect 7564 19184 7616 19236
rect 8116 19184 8168 19236
rect 10416 19252 10468 19304
rect 10784 19252 10836 19304
rect 11244 19252 11296 19304
rect 12348 19252 12400 19304
rect 9128 19184 9180 19236
rect 11428 19184 11480 19236
rect 11704 19184 11756 19236
rect 7288 19116 7340 19168
rect 8668 19116 8720 19168
rect 9220 19116 9272 19168
rect 10232 19116 10284 19168
rect 13084 19252 13136 19304
rect 14464 19295 14516 19304
rect 13176 19184 13228 19236
rect 14464 19261 14473 19295
rect 14473 19261 14507 19295
rect 14507 19261 14516 19295
rect 14464 19252 14516 19261
rect 15016 19252 15068 19304
rect 18880 19388 18932 19440
rect 16212 19320 16264 19372
rect 17132 19320 17184 19372
rect 20352 19363 20404 19372
rect 20352 19329 20361 19363
rect 20361 19329 20395 19363
rect 20395 19329 20404 19363
rect 20352 19320 20404 19329
rect 15936 19252 15988 19304
rect 16120 19295 16172 19304
rect 16120 19261 16129 19295
rect 16129 19261 16163 19295
rect 16163 19261 16172 19295
rect 16120 19252 16172 19261
rect 16580 19252 16632 19304
rect 12256 19116 12308 19168
rect 12992 19116 13044 19168
rect 15108 19159 15160 19168
rect 15108 19125 15117 19159
rect 15117 19125 15151 19159
rect 15151 19125 15160 19159
rect 15108 19116 15160 19125
rect 15476 19116 15528 19168
rect 18420 19295 18472 19304
rect 18420 19261 18429 19295
rect 18429 19261 18463 19295
rect 18463 19261 18472 19295
rect 18420 19252 18472 19261
rect 18512 19116 18564 19168
rect 18696 19116 18748 19168
rect 18880 19116 18932 19168
rect 20168 19252 20220 19304
rect 21272 19252 21324 19304
rect 19340 19184 19392 19236
rect 20628 19184 20680 19236
rect 19708 19159 19760 19168
rect 19708 19125 19717 19159
rect 19717 19125 19751 19159
rect 19751 19125 19760 19159
rect 19708 19116 19760 19125
rect 19892 19116 19944 19168
rect 20168 19159 20220 19168
rect 20168 19125 20177 19159
rect 20177 19125 20211 19159
rect 20211 19125 20220 19159
rect 20904 19159 20956 19168
rect 20168 19116 20220 19125
rect 20904 19125 20913 19159
rect 20913 19125 20947 19159
rect 20947 19125 20956 19159
rect 20904 19116 20956 19125
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 1768 18955 1820 18964
rect 1768 18921 1777 18955
rect 1777 18921 1811 18955
rect 1811 18921 1820 18955
rect 1768 18912 1820 18921
rect 2504 18912 2556 18964
rect 4068 18912 4120 18964
rect 4712 18955 4764 18964
rect 4712 18921 4721 18955
rect 4721 18921 4755 18955
rect 4755 18921 4764 18955
rect 4712 18912 4764 18921
rect 7288 18912 7340 18964
rect 7656 18912 7708 18964
rect 8208 18912 8260 18964
rect 8944 18912 8996 18964
rect 1860 18844 1912 18896
rect 10968 18912 11020 18964
rect 11428 18955 11480 18964
rect 11428 18921 11437 18955
rect 11437 18921 11471 18955
rect 11471 18921 11480 18955
rect 11428 18912 11480 18921
rect 12072 18912 12124 18964
rect 12440 18912 12492 18964
rect 16672 18955 16724 18964
rect 1584 18819 1636 18828
rect 1584 18785 1593 18819
rect 1593 18785 1627 18819
rect 1627 18785 1636 18819
rect 1584 18776 1636 18785
rect 2228 18776 2280 18828
rect 664 18708 716 18760
rect 2044 18640 2096 18692
rect 3056 18640 3108 18692
rect 3424 18776 3476 18828
rect 3516 18751 3568 18760
rect 3516 18717 3525 18751
rect 3525 18717 3559 18751
rect 3559 18717 3568 18751
rect 3516 18708 3568 18717
rect 4344 18776 4396 18828
rect 5264 18776 5316 18828
rect 6736 18819 6788 18828
rect 6736 18785 6745 18819
rect 6745 18785 6779 18819
rect 6779 18785 6788 18819
rect 6736 18776 6788 18785
rect 8300 18776 8352 18828
rect 5356 18751 5408 18760
rect 3424 18640 3476 18692
rect 3608 18640 3660 18692
rect 4344 18640 4396 18692
rect 5356 18717 5365 18751
rect 5365 18717 5399 18751
rect 5399 18717 5408 18751
rect 5356 18708 5408 18717
rect 6184 18751 6236 18760
rect 6184 18717 6193 18751
rect 6193 18717 6227 18751
rect 6227 18717 6236 18751
rect 6184 18708 6236 18717
rect 6460 18708 6512 18760
rect 11152 18844 11204 18896
rect 16672 18921 16681 18955
rect 16681 18921 16715 18955
rect 16715 18921 16724 18955
rect 16672 18912 16724 18921
rect 18604 18955 18656 18964
rect 8668 18776 8720 18828
rect 11704 18776 11756 18828
rect 13820 18887 13872 18896
rect 13820 18853 13843 18887
rect 13843 18853 13872 18887
rect 13820 18844 13872 18853
rect 14096 18844 14148 18896
rect 17776 18887 17828 18896
rect 17776 18853 17785 18887
rect 17785 18853 17819 18887
rect 17819 18853 17828 18887
rect 17776 18844 17828 18853
rect 17960 18844 18012 18896
rect 18604 18921 18613 18955
rect 18613 18921 18647 18955
rect 18647 18921 18656 18955
rect 18604 18912 18656 18921
rect 19432 18955 19484 18964
rect 19432 18921 19441 18955
rect 19441 18921 19475 18955
rect 19475 18921 19484 18955
rect 19432 18912 19484 18921
rect 19616 18844 19668 18896
rect 4160 18572 4212 18624
rect 6736 18640 6788 18692
rect 9128 18751 9180 18760
rect 9128 18717 9137 18751
rect 9137 18717 9171 18751
rect 9171 18717 9180 18751
rect 9128 18708 9180 18717
rect 12256 18751 12308 18760
rect 9496 18640 9548 18692
rect 9588 18640 9640 18692
rect 12256 18717 12265 18751
rect 12265 18717 12299 18751
rect 12299 18717 12308 18751
rect 12256 18708 12308 18717
rect 15292 18776 15344 18828
rect 15660 18819 15712 18828
rect 15660 18785 15669 18819
rect 15669 18785 15703 18819
rect 15703 18785 15712 18819
rect 15660 18776 15712 18785
rect 17868 18819 17920 18828
rect 12992 18708 13044 18760
rect 13360 18708 13412 18760
rect 15752 18751 15804 18760
rect 15752 18717 15761 18751
rect 15761 18717 15795 18751
rect 15795 18717 15804 18751
rect 15752 18708 15804 18717
rect 16212 18708 16264 18760
rect 16672 18708 16724 18760
rect 17868 18785 17877 18819
rect 17877 18785 17911 18819
rect 17911 18785 17920 18819
rect 17868 18776 17920 18785
rect 18604 18776 18656 18828
rect 19984 18776 20036 18828
rect 17592 18708 17644 18760
rect 18512 18708 18564 18760
rect 20352 18751 20404 18760
rect 20352 18717 20361 18751
rect 20361 18717 20395 18751
rect 20395 18717 20404 18751
rect 20352 18708 20404 18717
rect 13452 18640 13504 18692
rect 5356 18572 5408 18624
rect 9680 18572 9732 18624
rect 13176 18572 13228 18624
rect 21548 18640 21600 18692
rect 15016 18572 15068 18624
rect 16028 18572 16080 18624
rect 16304 18615 16356 18624
rect 16304 18581 16313 18615
rect 16313 18581 16347 18615
rect 16347 18581 16356 18615
rect 16304 18572 16356 18581
rect 17684 18572 17736 18624
rect 19800 18615 19852 18624
rect 19800 18581 19809 18615
rect 19809 18581 19843 18615
rect 19843 18581 19852 18615
rect 19800 18572 19852 18581
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 2780 18368 2832 18420
rect 3056 18368 3108 18420
rect 3424 18368 3476 18420
rect 3700 18368 3752 18420
rect 4988 18368 5040 18420
rect 5172 18411 5224 18420
rect 5172 18377 5181 18411
rect 5181 18377 5215 18411
rect 5215 18377 5224 18411
rect 5172 18368 5224 18377
rect 6184 18368 6236 18420
rect 8116 18368 8168 18420
rect 8668 18368 8720 18420
rect 8852 18368 8904 18420
rect 9036 18368 9088 18420
rect 9404 18368 9456 18420
rect 9496 18368 9548 18420
rect 9680 18368 9732 18420
rect 9956 18411 10008 18420
rect 9956 18377 9965 18411
rect 9965 18377 9999 18411
rect 9999 18377 10008 18411
rect 9956 18368 10008 18377
rect 10416 18368 10468 18420
rect 1768 18207 1820 18216
rect 1768 18173 1777 18207
rect 1777 18173 1811 18207
rect 1811 18173 1820 18207
rect 1768 18164 1820 18173
rect 2320 18207 2372 18216
rect 2320 18173 2329 18207
rect 2329 18173 2363 18207
rect 2363 18173 2372 18207
rect 2320 18164 2372 18173
rect 3056 18164 3108 18216
rect 3608 18232 3660 18284
rect 3884 18232 3936 18284
rect 4712 18275 4764 18284
rect 4712 18241 4721 18275
rect 4721 18241 4755 18275
rect 4755 18241 4764 18275
rect 4712 18232 4764 18241
rect 5540 18232 5592 18284
rect 4068 18164 4120 18216
rect 9772 18300 9824 18352
rect 8116 18232 8168 18284
rect 8300 18232 8352 18284
rect 9036 18232 9088 18284
rect 9128 18232 9180 18284
rect 9680 18232 9732 18284
rect 1492 18096 1544 18148
rect 3792 18096 3844 18148
rect 4528 18139 4580 18148
rect 4528 18105 4537 18139
rect 4537 18105 4571 18139
rect 4571 18105 4580 18139
rect 4528 18096 4580 18105
rect 4712 18096 4764 18148
rect 6276 18164 6328 18216
rect 13544 18368 13596 18420
rect 13728 18368 13780 18420
rect 15752 18368 15804 18420
rect 16948 18368 17000 18420
rect 18696 18368 18748 18420
rect 19248 18368 19300 18420
rect 19340 18368 19392 18420
rect 19616 18368 19668 18420
rect 22008 18368 22060 18420
rect 13268 18300 13320 18352
rect 13452 18300 13504 18352
rect 10968 18232 11020 18284
rect 11796 18164 11848 18216
rect 12256 18232 12308 18284
rect 13912 18232 13964 18284
rect 14096 18232 14148 18284
rect 12624 18164 12676 18216
rect 16764 18300 16816 18352
rect 17500 18300 17552 18352
rect 18236 18300 18288 18352
rect 14372 18275 14424 18284
rect 14372 18241 14381 18275
rect 14381 18241 14415 18275
rect 14415 18241 14424 18275
rect 14372 18232 14424 18241
rect 15568 18232 15620 18284
rect 16948 18232 17000 18284
rect 17316 18275 17368 18284
rect 17316 18241 17325 18275
rect 17325 18241 17359 18275
rect 17359 18241 17368 18275
rect 17316 18232 17368 18241
rect 20352 18300 20404 18352
rect 19524 18232 19576 18284
rect 3240 18028 3292 18080
rect 4160 18071 4212 18080
rect 4160 18037 4169 18071
rect 4169 18037 4203 18071
rect 4203 18037 4212 18071
rect 4160 18028 4212 18037
rect 4896 18028 4948 18080
rect 6460 18028 6512 18080
rect 12532 18096 12584 18148
rect 18604 18164 18656 18216
rect 19156 18164 19208 18216
rect 7472 18071 7524 18080
rect 7472 18037 7481 18071
rect 7481 18037 7515 18071
rect 7515 18037 7524 18071
rect 7472 18028 7524 18037
rect 7656 18028 7708 18080
rect 8208 18028 8260 18080
rect 9496 18028 9548 18080
rect 10416 18028 10468 18080
rect 12799 18028 12851 18080
rect 13084 18028 13136 18080
rect 16488 18096 16540 18148
rect 18696 18096 18748 18148
rect 19340 18096 19392 18148
rect 20720 18139 20772 18148
rect 20720 18105 20729 18139
rect 20729 18105 20763 18139
rect 20763 18105 20772 18139
rect 20720 18096 20772 18105
rect 14188 18071 14240 18080
rect 14188 18037 14197 18071
rect 14197 18037 14231 18071
rect 14231 18037 14240 18071
rect 14188 18028 14240 18037
rect 14280 18071 14332 18080
rect 14280 18037 14289 18071
rect 14289 18037 14323 18071
rect 14323 18037 14332 18071
rect 15200 18071 15252 18080
rect 14280 18028 14332 18037
rect 15200 18037 15209 18071
rect 15209 18037 15243 18071
rect 15243 18037 15252 18071
rect 15200 18028 15252 18037
rect 15476 18028 15528 18080
rect 17224 18071 17276 18080
rect 17224 18037 17233 18071
rect 17233 18037 17267 18071
rect 17267 18037 17276 18071
rect 17224 18028 17276 18037
rect 18052 18071 18104 18080
rect 18052 18037 18061 18071
rect 18061 18037 18095 18071
rect 18095 18037 18104 18071
rect 18052 18028 18104 18037
rect 18604 18028 18656 18080
rect 19432 18071 19484 18080
rect 19432 18037 19441 18071
rect 19441 18037 19475 18071
rect 19475 18037 19484 18071
rect 19432 18028 19484 18037
rect 19800 18071 19852 18080
rect 19800 18037 19809 18071
rect 19809 18037 19843 18071
rect 19843 18037 19852 18071
rect 19800 18028 19852 18037
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 1676 17867 1728 17876
rect 1676 17833 1685 17867
rect 1685 17833 1719 17867
rect 1719 17833 1728 17867
rect 1676 17824 1728 17833
rect 1952 17824 2004 17876
rect 3240 17824 3292 17876
rect 4252 17824 4304 17876
rect 4988 17824 5040 17876
rect 6828 17824 6880 17876
rect 7288 17867 7340 17876
rect 7288 17833 7297 17867
rect 7297 17833 7331 17867
rect 7331 17833 7340 17867
rect 7288 17824 7340 17833
rect 2320 17799 2372 17808
rect 2320 17765 2329 17799
rect 2329 17765 2363 17799
rect 2363 17765 2372 17799
rect 2320 17756 2372 17765
rect 4160 17756 4212 17808
rect 3056 17688 3108 17740
rect 3516 17688 3568 17740
rect 4804 17688 4856 17740
rect 5540 17688 5592 17740
rect 7472 17688 7524 17740
rect 7748 17824 7800 17876
rect 7840 17756 7892 17808
rect 12164 17824 12216 17876
rect 12808 17867 12860 17876
rect 12808 17833 12817 17867
rect 12817 17833 12851 17867
rect 12851 17833 12860 17867
rect 12808 17824 12860 17833
rect 13452 17824 13504 17876
rect 14188 17824 14240 17876
rect 15292 17867 15344 17876
rect 15292 17833 15301 17867
rect 15301 17833 15335 17867
rect 15335 17833 15344 17867
rect 15292 17824 15344 17833
rect 16580 17824 16632 17876
rect 16764 17867 16816 17876
rect 16764 17833 16773 17867
rect 16773 17833 16807 17867
rect 16807 17833 16816 17867
rect 16764 17824 16816 17833
rect 19800 17824 19852 17876
rect 10508 17756 10560 17808
rect 13084 17756 13136 17808
rect 13268 17799 13320 17808
rect 13268 17765 13277 17799
rect 13277 17765 13311 17799
rect 13311 17765 13320 17799
rect 13268 17756 13320 17765
rect 13544 17756 13596 17808
rect 15108 17756 15160 17808
rect 10048 17731 10100 17740
rect 2780 17620 2832 17672
rect 3608 17663 3660 17672
rect 3608 17629 3617 17663
rect 3617 17629 3651 17663
rect 3651 17629 3660 17663
rect 3608 17620 3660 17629
rect 4160 17620 4212 17672
rect 4620 17663 4672 17672
rect 4620 17629 4629 17663
rect 4629 17629 4663 17663
rect 4663 17629 4672 17663
rect 4620 17620 4672 17629
rect 5080 17663 5132 17672
rect 5080 17629 5089 17663
rect 5089 17629 5123 17663
rect 5123 17629 5132 17663
rect 5080 17620 5132 17629
rect 5172 17620 5224 17672
rect 10048 17697 10057 17731
rect 10057 17697 10091 17731
rect 10091 17697 10100 17731
rect 10048 17688 10100 17697
rect 10784 17688 10836 17740
rect 11704 17688 11756 17740
rect 4712 17552 4764 17604
rect 2872 17484 2924 17536
rect 5264 17484 5316 17536
rect 5448 17484 5500 17536
rect 7748 17663 7800 17672
rect 7748 17629 7757 17663
rect 7757 17629 7791 17663
rect 7791 17629 7800 17663
rect 7748 17620 7800 17629
rect 8944 17663 8996 17672
rect 8944 17629 8953 17663
rect 8953 17629 8987 17663
rect 8987 17629 8996 17663
rect 8944 17620 8996 17629
rect 9036 17663 9088 17672
rect 9036 17629 9045 17663
rect 9045 17629 9079 17663
rect 9079 17629 9088 17663
rect 9036 17620 9088 17629
rect 9220 17620 9272 17672
rect 9404 17620 9456 17672
rect 6644 17484 6696 17536
rect 7748 17484 7800 17536
rect 9128 17552 9180 17604
rect 12256 17620 12308 17672
rect 13912 17688 13964 17740
rect 15660 17731 15712 17740
rect 15660 17697 15669 17731
rect 15669 17697 15703 17731
rect 15703 17697 15712 17731
rect 15660 17688 15712 17697
rect 15936 17688 15988 17740
rect 13820 17620 13872 17672
rect 15016 17620 15068 17672
rect 16580 17688 16632 17740
rect 16764 17688 16816 17740
rect 17132 17688 17184 17740
rect 19616 17756 19668 17808
rect 19984 17756 20036 17808
rect 16856 17663 16908 17672
rect 16856 17629 16865 17663
rect 16865 17629 16899 17663
rect 16899 17629 16908 17663
rect 17776 17663 17828 17672
rect 16856 17620 16908 17629
rect 17776 17629 17785 17663
rect 17785 17629 17819 17663
rect 17819 17629 17828 17663
rect 17776 17620 17828 17629
rect 19708 17688 19760 17740
rect 19800 17688 19852 17740
rect 20168 17688 20220 17740
rect 18788 17663 18840 17672
rect 18788 17629 18797 17663
rect 18797 17629 18831 17663
rect 18831 17629 18840 17663
rect 18788 17620 18840 17629
rect 18972 17663 19024 17672
rect 18972 17629 18981 17663
rect 18981 17629 19015 17663
rect 19015 17629 19024 17663
rect 19984 17663 20036 17672
rect 18972 17620 19024 17629
rect 10508 17484 10560 17536
rect 12624 17484 12676 17536
rect 19340 17552 19392 17604
rect 19984 17629 19993 17663
rect 19993 17629 20027 17663
rect 20027 17629 20036 17663
rect 19984 17620 20036 17629
rect 20904 17484 20956 17536
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 3516 17280 3568 17332
rect 3608 17280 3660 17332
rect 5540 17323 5592 17332
rect 1952 17187 2004 17196
rect 1952 17153 1961 17187
rect 1961 17153 1995 17187
rect 1995 17153 2004 17187
rect 1952 17144 2004 17153
rect 2136 17187 2188 17196
rect 2136 17153 2145 17187
rect 2145 17153 2179 17187
rect 2179 17153 2188 17187
rect 2136 17144 2188 17153
rect 5540 17289 5549 17323
rect 5549 17289 5583 17323
rect 5583 17289 5592 17323
rect 5540 17280 5592 17289
rect 7840 17280 7892 17332
rect 8208 17280 8260 17332
rect 8944 17280 8996 17332
rect 9220 17280 9272 17332
rect 11152 17323 11204 17332
rect 11152 17289 11161 17323
rect 11161 17289 11195 17323
rect 11195 17289 11204 17323
rect 11152 17280 11204 17289
rect 14188 17280 14240 17332
rect 4160 17212 4212 17264
rect 5264 17212 5316 17264
rect 11428 17212 11480 17264
rect 11612 17212 11664 17264
rect 17316 17280 17368 17332
rect 17868 17280 17920 17332
rect 17960 17280 18012 17332
rect 20168 17280 20220 17332
rect 18420 17212 18472 17264
rect 1400 17076 1452 17128
rect 2504 17119 2556 17128
rect 2504 17085 2513 17119
rect 2513 17085 2547 17119
rect 2547 17085 2556 17119
rect 2504 17076 2556 17085
rect 6552 17144 6604 17196
rect 6920 17144 6972 17196
rect 2964 17008 3016 17060
rect 3148 17008 3200 17060
rect 7012 17076 7064 17128
rect 9128 17144 9180 17196
rect 10508 17144 10560 17196
rect 5172 17008 5224 17060
rect 6920 17008 6972 17060
rect 7748 17008 7800 17060
rect 2872 16940 2924 16992
rect 3332 16940 3384 16992
rect 4896 16940 4948 16992
rect 7104 16983 7156 16992
rect 7104 16949 7113 16983
rect 7113 16949 7147 16983
rect 7147 16949 7156 16983
rect 7104 16940 7156 16949
rect 9864 17076 9916 17128
rect 9956 17076 10008 17128
rect 12256 17144 12308 17196
rect 13820 17144 13872 17196
rect 14188 17144 14240 17196
rect 19340 17144 19392 17196
rect 20536 17187 20588 17196
rect 20536 17153 20545 17187
rect 20545 17153 20579 17187
rect 20579 17153 20588 17187
rect 20536 17144 20588 17153
rect 12532 17119 12584 17128
rect 12532 17085 12541 17119
rect 12541 17085 12575 17119
rect 12575 17085 12584 17119
rect 12532 17076 12584 17085
rect 13360 17076 13412 17128
rect 14280 17119 14332 17128
rect 14280 17085 14289 17119
rect 14289 17085 14323 17119
rect 14323 17085 14332 17119
rect 14280 17076 14332 17085
rect 14372 17076 14424 17128
rect 15016 17076 15068 17128
rect 16212 17119 16264 17128
rect 8852 17008 8904 17060
rect 9404 17008 9456 17060
rect 13452 17051 13504 17060
rect 8484 16940 8536 16992
rect 9496 16983 9548 16992
rect 9496 16949 9505 16983
rect 9505 16949 9539 16983
rect 9539 16949 9548 16983
rect 9496 16940 9548 16949
rect 9680 16940 9732 16992
rect 13452 17017 13461 17051
rect 13461 17017 13495 17051
rect 13495 17017 13504 17051
rect 13452 17008 13504 17017
rect 16212 17085 16221 17119
rect 16221 17085 16255 17119
rect 16255 17085 16264 17119
rect 16212 17076 16264 17085
rect 16856 17076 16908 17128
rect 16948 17076 17000 17128
rect 19248 17076 19300 17128
rect 20904 17187 20956 17196
rect 20904 17153 20913 17187
rect 20913 17153 20947 17187
rect 20947 17153 20956 17187
rect 20904 17144 20956 17153
rect 12440 16940 12492 16992
rect 15568 16940 15620 16992
rect 18328 17008 18380 17060
rect 17132 16940 17184 16992
rect 18052 16983 18104 16992
rect 18052 16949 18061 16983
rect 18061 16949 18095 16983
rect 18095 16949 18104 16983
rect 18052 16940 18104 16949
rect 18144 16940 18196 16992
rect 20812 17008 20864 17060
rect 18880 16940 18932 16992
rect 19248 16983 19300 16992
rect 19248 16949 19257 16983
rect 19257 16949 19291 16983
rect 19291 16949 19300 16983
rect 19248 16940 19300 16949
rect 19340 16983 19392 16992
rect 19340 16949 19349 16983
rect 19349 16949 19383 16983
rect 19383 16949 19392 16983
rect 19340 16940 19392 16949
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 1584 16779 1636 16788
rect 1584 16745 1593 16779
rect 1593 16745 1627 16779
rect 1627 16745 1636 16779
rect 1584 16736 1636 16745
rect 2320 16779 2372 16788
rect 204 16668 256 16720
rect 2320 16745 2329 16779
rect 2329 16745 2363 16779
rect 2363 16745 2372 16779
rect 2320 16736 2372 16745
rect 2412 16736 2464 16788
rect 2780 16736 2832 16788
rect 4252 16736 4304 16788
rect 5448 16779 5500 16788
rect 5448 16745 5457 16779
rect 5457 16745 5491 16779
rect 5491 16745 5500 16779
rect 5448 16736 5500 16745
rect 7104 16736 7156 16788
rect 7472 16779 7524 16788
rect 7472 16745 7481 16779
rect 7481 16745 7515 16779
rect 7515 16745 7524 16779
rect 7472 16736 7524 16745
rect 8576 16736 8628 16788
rect 9128 16736 9180 16788
rect 11704 16779 11756 16788
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 4712 16668 4764 16720
rect 7656 16668 7708 16720
rect 2412 16575 2464 16584
rect 2412 16541 2421 16575
rect 2421 16541 2455 16575
rect 2455 16541 2464 16575
rect 2412 16532 2464 16541
rect 3608 16575 3660 16584
rect 3332 16464 3384 16516
rect 3608 16541 3617 16575
rect 3617 16541 3651 16575
rect 3651 16541 3660 16575
rect 3608 16532 3660 16541
rect 4160 16600 4212 16652
rect 6736 16600 6788 16652
rect 9680 16668 9732 16720
rect 11704 16745 11713 16779
rect 11713 16745 11747 16779
rect 11747 16745 11756 16779
rect 11704 16736 11756 16745
rect 11888 16736 11940 16788
rect 11520 16668 11572 16720
rect 8208 16643 8260 16652
rect 4344 16532 4396 16584
rect 5264 16532 5316 16584
rect 5540 16464 5592 16516
rect 6460 16532 6512 16584
rect 7104 16575 7156 16584
rect 7104 16541 7113 16575
rect 7113 16541 7147 16575
rect 7147 16541 7156 16575
rect 7104 16532 7156 16541
rect 8208 16609 8231 16643
rect 8231 16609 8260 16643
rect 8208 16600 8260 16609
rect 8484 16600 8536 16652
rect 9128 16600 9180 16652
rect 10416 16600 10468 16652
rect 11152 16600 11204 16652
rect 12072 16600 12124 16652
rect 15016 16736 15068 16788
rect 16856 16736 16908 16788
rect 17408 16736 17460 16788
rect 14372 16668 14424 16720
rect 13268 16600 13320 16652
rect 13360 16600 13412 16652
rect 14188 16600 14240 16652
rect 15844 16668 15896 16720
rect 17132 16668 17184 16720
rect 12532 16575 12584 16584
rect 6184 16396 6236 16448
rect 6460 16439 6512 16448
rect 6460 16405 6469 16439
rect 6469 16405 6503 16439
rect 6503 16405 6512 16439
rect 6460 16396 6512 16405
rect 7564 16396 7616 16448
rect 12532 16541 12541 16575
rect 12541 16541 12575 16575
rect 12575 16541 12584 16575
rect 12532 16532 12584 16541
rect 12624 16575 12676 16584
rect 12624 16541 12633 16575
rect 12633 16541 12667 16575
rect 12667 16541 12676 16575
rect 12624 16532 12676 16541
rect 11428 16464 11480 16516
rect 12440 16464 12492 16516
rect 15568 16643 15620 16652
rect 15568 16609 15602 16643
rect 15602 16609 15620 16643
rect 17776 16736 17828 16788
rect 18236 16736 18288 16788
rect 18512 16736 18564 16788
rect 18788 16736 18840 16788
rect 19984 16779 20036 16788
rect 19984 16745 19993 16779
rect 19993 16745 20027 16779
rect 20027 16745 20036 16779
rect 19984 16736 20036 16745
rect 18052 16668 18104 16720
rect 15568 16600 15620 16609
rect 9680 16396 9732 16448
rect 11888 16396 11940 16448
rect 14924 16396 14976 16448
rect 17316 16532 17368 16584
rect 17776 16600 17828 16652
rect 18512 16643 18564 16652
rect 18512 16609 18521 16643
rect 18521 16609 18555 16643
rect 18555 16609 18564 16643
rect 18512 16600 18564 16609
rect 19064 16600 19116 16652
rect 21364 16668 21416 16720
rect 20904 16643 20956 16652
rect 18420 16532 18472 16584
rect 18788 16575 18840 16584
rect 18788 16541 18797 16575
rect 18797 16541 18831 16575
rect 18831 16541 18840 16575
rect 18788 16532 18840 16541
rect 19616 16575 19668 16584
rect 19616 16541 19625 16575
rect 19625 16541 19659 16575
rect 19659 16541 19668 16575
rect 19616 16532 19668 16541
rect 19708 16532 19760 16584
rect 20536 16575 20588 16584
rect 20536 16541 20545 16575
rect 20545 16541 20579 16575
rect 20579 16541 20588 16575
rect 20536 16532 20588 16541
rect 16580 16464 16632 16516
rect 17776 16464 17828 16516
rect 16212 16396 16264 16448
rect 16856 16396 16908 16448
rect 20904 16609 20913 16643
rect 20913 16609 20947 16643
rect 20947 16609 20956 16643
rect 20904 16600 20956 16609
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 1676 16235 1728 16244
rect 1676 16201 1685 16235
rect 1685 16201 1719 16235
rect 1719 16201 1728 16235
rect 1676 16192 1728 16201
rect 2504 16192 2556 16244
rect 4712 16235 4764 16244
rect 1676 15988 1728 16040
rect 2504 15963 2556 15972
rect 2504 15929 2513 15963
rect 2513 15929 2547 15963
rect 2547 15929 2556 15963
rect 2504 15920 2556 15929
rect 2780 16056 2832 16108
rect 4712 16201 4721 16235
rect 4721 16201 4755 16235
rect 4755 16201 4764 16235
rect 4712 16192 4764 16201
rect 6920 16192 6972 16244
rect 7012 16192 7064 16244
rect 7472 16192 7524 16244
rect 8116 16192 8168 16244
rect 8208 16192 8260 16244
rect 8944 16192 8996 16244
rect 6184 16124 6236 16176
rect 7104 16124 7156 16176
rect 11152 16192 11204 16244
rect 12624 16192 12676 16244
rect 12808 16192 12860 16244
rect 14464 16192 14516 16244
rect 14648 16192 14700 16244
rect 5264 16099 5316 16108
rect 5264 16065 5273 16099
rect 5273 16065 5307 16099
rect 5307 16065 5316 16099
rect 5264 16056 5316 16065
rect 6828 16056 6880 16108
rect 7012 16056 7064 16108
rect 3148 15988 3200 16040
rect 6460 15988 6512 16040
rect 7288 15988 7340 16040
rect 7564 15988 7616 16040
rect 7748 16031 7800 16040
rect 7748 15997 7782 16031
rect 7782 15997 7800 16031
rect 7748 15988 7800 15997
rect 9588 15988 9640 16040
rect 9680 15988 9732 16040
rect 15200 16192 15252 16244
rect 17132 16192 17184 16244
rect 18512 16192 18564 16244
rect 19616 16192 19668 16244
rect 12256 16056 12308 16108
rect 13360 16056 13412 16108
rect 13636 16056 13688 16108
rect 20904 16124 20956 16176
rect 21180 16124 21232 16176
rect 12440 15988 12492 16040
rect 3516 15920 3568 15972
rect 2412 15895 2464 15904
rect 2412 15861 2421 15895
rect 2421 15861 2455 15895
rect 2455 15861 2464 15895
rect 2412 15852 2464 15861
rect 2596 15852 2648 15904
rect 5540 15920 5592 15972
rect 14464 15988 14516 16040
rect 15844 16056 15896 16108
rect 17776 16056 17828 16108
rect 18788 16056 18840 16108
rect 20444 16099 20496 16108
rect 15384 15988 15436 16040
rect 16672 15988 16724 16040
rect 20444 16065 20453 16099
rect 20453 16065 20487 16099
rect 20487 16065 20496 16099
rect 20444 16056 20496 16065
rect 20628 15988 20680 16040
rect 10048 15920 10100 15972
rect 10876 15920 10928 15972
rect 13820 15963 13872 15972
rect 13820 15929 13829 15963
rect 13829 15929 13863 15963
rect 13863 15929 13872 15963
rect 13820 15920 13872 15929
rect 3700 15852 3752 15904
rect 6920 15852 6972 15904
rect 7104 15895 7156 15904
rect 7104 15861 7113 15895
rect 7113 15861 7147 15895
rect 7147 15861 7156 15895
rect 7104 15852 7156 15861
rect 12348 15852 12400 15904
rect 12532 15852 12584 15904
rect 12716 15852 12768 15904
rect 13176 15852 13228 15904
rect 13452 15895 13504 15904
rect 13452 15861 13461 15895
rect 13461 15861 13495 15895
rect 13495 15861 13504 15895
rect 13452 15852 13504 15861
rect 13544 15852 13596 15904
rect 14004 15920 14056 15972
rect 15844 15852 15896 15904
rect 16488 15852 16540 15904
rect 16672 15895 16724 15904
rect 16672 15861 16681 15895
rect 16681 15861 16715 15895
rect 16715 15861 16724 15895
rect 16672 15852 16724 15861
rect 19616 15852 19668 15904
rect 19984 15852 20036 15904
rect 20260 15895 20312 15904
rect 20260 15861 20269 15895
rect 20269 15861 20303 15895
rect 20303 15861 20312 15895
rect 20260 15852 20312 15861
rect 20352 15895 20404 15904
rect 20352 15861 20361 15895
rect 20361 15861 20395 15895
rect 20395 15861 20404 15895
rect 20352 15852 20404 15861
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 1492 15648 1544 15700
rect 2596 15648 2648 15700
rect 3332 15691 3384 15700
rect 3332 15657 3341 15691
rect 3341 15657 3375 15691
rect 3375 15657 3384 15691
rect 3332 15648 3384 15657
rect 4160 15648 4212 15700
rect 5080 15648 5132 15700
rect 6828 15648 6880 15700
rect 3700 15580 3752 15632
rect 4252 15580 4304 15632
rect 1584 15512 1636 15564
rect 2044 15512 2096 15564
rect 4896 15512 4948 15564
rect 2504 15444 2556 15496
rect 2780 15444 2832 15496
rect 3516 15487 3568 15496
rect 3516 15453 3525 15487
rect 3525 15453 3559 15487
rect 3559 15453 3568 15487
rect 3516 15444 3568 15453
rect 5448 15512 5500 15564
rect 6184 15512 6236 15564
rect 5540 15444 5592 15496
rect 3976 15376 4028 15428
rect 4068 15308 4120 15360
rect 6368 15308 6420 15360
rect 7748 15648 7800 15700
rect 8208 15648 8260 15700
rect 9680 15648 9732 15700
rect 10416 15648 10468 15700
rect 11888 15648 11940 15700
rect 7104 15580 7156 15632
rect 9036 15555 9088 15564
rect 7012 15444 7064 15496
rect 9036 15521 9045 15555
rect 9045 15521 9079 15555
rect 9079 15521 9088 15555
rect 9036 15512 9088 15521
rect 9680 15555 9732 15564
rect 9680 15521 9689 15555
rect 9689 15521 9723 15555
rect 9723 15521 9732 15555
rect 9680 15512 9732 15521
rect 10508 15512 10560 15564
rect 10968 15512 11020 15564
rect 12532 15648 12584 15700
rect 13636 15648 13688 15700
rect 15844 15648 15896 15700
rect 16672 15648 16724 15700
rect 12808 15580 12860 15632
rect 13084 15580 13136 15632
rect 14372 15580 14424 15632
rect 9220 15444 9272 15496
rect 11152 15444 11204 15496
rect 11888 15444 11940 15496
rect 12440 15512 12492 15564
rect 15016 15555 15068 15564
rect 15016 15521 15025 15555
rect 15025 15521 15059 15555
rect 15059 15521 15068 15555
rect 15016 15512 15068 15521
rect 16580 15580 16632 15632
rect 21364 15648 21416 15700
rect 17408 15580 17460 15632
rect 19708 15580 19760 15632
rect 19156 15555 19208 15564
rect 19156 15521 19165 15555
rect 19165 15521 19199 15555
rect 19199 15521 19208 15555
rect 19156 15512 19208 15521
rect 19432 15512 19484 15564
rect 12256 15444 12308 15496
rect 9496 15376 9548 15428
rect 10876 15376 10928 15428
rect 13544 15444 13596 15496
rect 14004 15376 14056 15428
rect 15568 15444 15620 15496
rect 16212 15376 16264 15428
rect 18788 15444 18840 15496
rect 20076 15487 20128 15496
rect 12440 15308 12492 15360
rect 12808 15351 12860 15360
rect 12808 15317 12817 15351
rect 12817 15317 12851 15351
rect 12851 15317 12860 15351
rect 12808 15308 12860 15317
rect 13820 15351 13872 15360
rect 13820 15317 13829 15351
rect 13829 15317 13863 15351
rect 13863 15317 13872 15351
rect 13820 15308 13872 15317
rect 14280 15308 14332 15360
rect 16764 15308 16816 15360
rect 20076 15453 20085 15487
rect 20085 15453 20119 15487
rect 20119 15453 20128 15487
rect 20076 15444 20128 15453
rect 17040 15308 17092 15360
rect 17960 15308 18012 15360
rect 18512 15308 18564 15360
rect 19340 15308 19392 15360
rect 19616 15351 19668 15360
rect 19616 15317 19625 15351
rect 19625 15317 19659 15351
rect 19659 15317 19668 15351
rect 19616 15308 19668 15317
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 3424 15147 3476 15156
rect 3424 15113 3433 15147
rect 3433 15113 3467 15147
rect 3467 15113 3476 15147
rect 3424 15104 3476 15113
rect 3976 15104 4028 15156
rect 5448 15104 5500 15156
rect 6368 15147 6420 15156
rect 6368 15113 6377 15147
rect 6377 15113 6411 15147
rect 6411 15113 6420 15147
rect 6368 15104 6420 15113
rect 7196 15104 7248 15156
rect 7472 15104 7524 15156
rect 7656 15147 7708 15156
rect 7656 15113 7665 15147
rect 7665 15113 7699 15147
rect 7699 15113 7708 15147
rect 7656 15104 7708 15113
rect 8576 15104 8628 15156
rect 8944 15104 8996 15156
rect 10324 15104 10376 15156
rect 12716 15104 12768 15156
rect 3148 15036 3200 15088
rect 5172 15079 5224 15088
rect 5172 15045 5181 15079
rect 5181 15045 5215 15079
rect 5215 15045 5224 15079
rect 5172 15036 5224 15045
rect 6184 15036 6236 15088
rect 6552 15036 6604 15088
rect 7564 15036 7616 15088
rect 13176 15036 13228 15088
rect 1676 15011 1728 15020
rect 1676 14977 1685 15011
rect 1685 14977 1719 15011
rect 1719 14977 1728 15011
rect 1676 14968 1728 14977
rect 2964 14968 3016 15020
rect 7472 15011 7524 15020
rect 7472 14977 7481 15011
rect 7481 14977 7515 15011
rect 7515 14977 7524 15011
rect 7472 14968 7524 14977
rect 8208 15011 8260 15020
rect 8208 14977 8217 15011
rect 8217 14977 8251 15011
rect 8251 14977 8260 15011
rect 8208 14968 8260 14977
rect 9312 14968 9364 15020
rect 9772 14968 9824 15020
rect 10968 14968 11020 15020
rect 12440 14968 12492 15020
rect 13268 14968 13320 15020
rect 14280 15104 14332 15156
rect 15384 15036 15436 15088
rect 1492 14943 1544 14952
rect 1492 14909 1501 14943
rect 1501 14909 1535 14943
rect 1535 14909 1544 14943
rect 1492 14900 1544 14909
rect 2872 14900 2924 14952
rect 3424 14900 3476 14952
rect 3516 14900 3568 14952
rect 7656 14900 7708 14952
rect 5448 14832 5500 14884
rect 6092 14832 6144 14884
rect 6920 14832 6972 14884
rect 7932 14832 7984 14884
rect 2044 14764 2096 14816
rect 2596 14807 2648 14816
rect 2596 14773 2605 14807
rect 2605 14773 2639 14807
rect 2639 14773 2648 14807
rect 2596 14764 2648 14773
rect 3884 14764 3936 14816
rect 4160 14764 4212 14816
rect 4620 14764 4672 14816
rect 6552 14764 6604 14816
rect 6828 14807 6880 14816
rect 6828 14773 6837 14807
rect 6837 14773 6871 14807
rect 6871 14773 6880 14807
rect 6828 14764 6880 14773
rect 8576 14764 8628 14816
rect 9220 14807 9272 14816
rect 9220 14773 9229 14807
rect 9229 14773 9263 14807
rect 9263 14773 9272 14807
rect 9220 14764 9272 14773
rect 9312 14807 9364 14816
rect 9312 14773 9321 14807
rect 9321 14773 9355 14807
rect 9355 14773 9364 14807
rect 9312 14764 9364 14773
rect 9772 14764 9824 14816
rect 10232 14807 10284 14816
rect 10232 14773 10241 14807
rect 10241 14773 10275 14807
rect 10275 14773 10284 14807
rect 10232 14764 10284 14773
rect 11152 14900 11204 14952
rect 11152 14764 11204 14816
rect 12532 14900 12584 14952
rect 11980 14764 12032 14816
rect 12256 14764 12308 14816
rect 12532 14764 12584 14816
rect 13728 14832 13780 14884
rect 13912 14900 13964 14952
rect 16856 15104 16908 15156
rect 16672 15036 16724 15088
rect 17224 15036 17276 15088
rect 18052 15036 18104 15088
rect 19432 15104 19484 15156
rect 20076 15147 20128 15156
rect 20076 15113 20085 15147
rect 20085 15113 20119 15147
rect 20119 15113 20128 15147
rect 20076 15104 20128 15113
rect 16764 14968 16816 15020
rect 17960 14968 18012 15020
rect 18512 15011 18564 15020
rect 18512 14977 18521 15011
rect 18521 14977 18555 15011
rect 18555 14977 18564 15011
rect 18512 14968 18564 14977
rect 15108 14832 15160 14884
rect 17408 14900 17460 14952
rect 19248 15036 19300 15088
rect 19340 14968 19392 15020
rect 16212 14832 16264 14884
rect 16856 14832 16908 14884
rect 19616 14832 19668 14884
rect 14280 14764 14332 14816
rect 15292 14764 15344 14816
rect 15752 14764 15804 14816
rect 17408 14764 17460 14816
rect 19064 14764 19116 14816
rect 19432 14807 19484 14816
rect 19432 14773 19441 14807
rect 19441 14773 19475 14807
rect 19475 14773 19484 14807
rect 19432 14764 19484 14773
rect 19892 14764 19944 14816
rect 20168 14764 20220 14816
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 1492 14560 1544 14612
rect 5356 14560 5408 14612
rect 6828 14560 6880 14612
rect 6920 14560 6972 14612
rect 7564 14560 7616 14612
rect 9128 14560 9180 14612
rect 10232 14560 10284 14612
rect 10324 14560 10376 14612
rect 3148 14492 3200 14544
rect 3516 14535 3568 14544
rect 3516 14501 3525 14535
rect 3525 14501 3559 14535
rect 3559 14501 3568 14535
rect 3516 14492 3568 14501
rect 4252 14492 4304 14544
rect 1492 14467 1544 14476
rect 1492 14433 1501 14467
rect 1501 14433 1535 14467
rect 1535 14433 1544 14467
rect 1492 14424 1544 14433
rect 3240 14467 3292 14476
rect 3240 14433 3249 14467
rect 3249 14433 3283 14467
rect 3283 14433 3292 14467
rect 3240 14424 3292 14433
rect 1768 14399 1820 14408
rect 1768 14365 1777 14399
rect 1777 14365 1811 14399
rect 1811 14365 1820 14399
rect 1768 14356 1820 14365
rect 2964 14356 3016 14408
rect 3516 14288 3568 14340
rect 2228 14263 2280 14272
rect 2228 14229 2237 14263
rect 2237 14229 2271 14263
rect 2271 14229 2280 14263
rect 2228 14220 2280 14229
rect 2596 14220 2648 14272
rect 4896 14424 4948 14476
rect 5540 14424 5592 14476
rect 5632 14424 5684 14476
rect 3976 14356 4028 14408
rect 6460 14424 6512 14476
rect 7840 14467 7892 14476
rect 7840 14433 7849 14467
rect 7849 14433 7883 14467
rect 7883 14433 7892 14467
rect 7840 14424 7892 14433
rect 8576 14492 8628 14544
rect 11980 14560 12032 14612
rect 12164 14603 12216 14612
rect 12164 14569 12173 14603
rect 12173 14569 12207 14603
rect 12207 14569 12216 14603
rect 12164 14560 12216 14569
rect 12716 14560 12768 14612
rect 13820 14560 13872 14612
rect 15292 14560 15344 14612
rect 17868 14560 17920 14612
rect 19156 14560 19208 14612
rect 19432 14560 19484 14612
rect 11336 14492 11388 14544
rect 7472 14399 7524 14408
rect 7472 14365 7481 14399
rect 7481 14365 7515 14399
rect 7515 14365 7524 14399
rect 8392 14399 8444 14408
rect 7472 14356 7524 14365
rect 8392 14365 8401 14399
rect 8401 14365 8435 14399
rect 8435 14365 8444 14399
rect 8392 14356 8444 14365
rect 4804 14220 4856 14272
rect 5540 14220 5592 14272
rect 6920 14263 6972 14272
rect 6920 14229 6929 14263
rect 6929 14229 6963 14263
rect 6963 14229 6972 14263
rect 6920 14220 6972 14229
rect 8668 14424 8720 14476
rect 10048 14467 10100 14476
rect 10048 14433 10057 14467
rect 10057 14433 10091 14467
rect 10091 14433 10100 14467
rect 10048 14424 10100 14433
rect 12992 14492 13044 14544
rect 12532 14467 12584 14476
rect 12532 14433 12541 14467
rect 12541 14433 12575 14467
rect 12575 14433 12584 14467
rect 12532 14424 12584 14433
rect 14924 14424 14976 14476
rect 15384 14424 15436 14476
rect 16948 14424 17000 14476
rect 20168 14467 20220 14476
rect 10232 14356 10284 14408
rect 10968 14356 11020 14408
rect 14004 14356 14056 14408
rect 15292 14399 15344 14408
rect 11704 14288 11756 14340
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 17040 14356 17092 14408
rect 19064 14399 19116 14408
rect 11612 14220 11664 14272
rect 12716 14220 12768 14272
rect 13728 14220 13780 14272
rect 15660 14220 15712 14272
rect 17040 14220 17092 14272
rect 19064 14365 19073 14399
rect 19073 14365 19107 14399
rect 19107 14365 19116 14399
rect 19064 14356 19116 14365
rect 20168 14433 20177 14467
rect 20177 14433 20211 14467
rect 20211 14433 20220 14467
rect 20168 14424 20220 14433
rect 19432 14356 19484 14408
rect 18788 14288 18840 14340
rect 19616 14331 19668 14340
rect 19616 14297 19625 14331
rect 19625 14297 19659 14331
rect 19659 14297 19668 14331
rect 20352 14399 20404 14408
rect 20352 14365 20361 14399
rect 20361 14365 20395 14399
rect 20395 14365 20404 14399
rect 20352 14356 20404 14365
rect 19616 14288 19668 14297
rect 17868 14220 17920 14272
rect 19248 14220 19300 14272
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 2872 14016 2924 14068
rect 3792 14016 3844 14068
rect 4068 14016 4120 14068
rect 4068 13880 4120 13932
rect 2412 13812 2464 13864
rect 2136 13744 2188 13796
rect 3976 13812 4028 13864
rect 4528 13855 4580 13864
rect 4528 13821 4537 13855
rect 4537 13821 4571 13855
rect 4571 13821 4580 13855
rect 4528 13812 4580 13821
rect 3608 13744 3660 13796
rect 4804 13855 4856 13864
rect 4804 13821 4838 13855
rect 4838 13821 4856 13855
rect 4804 13812 4856 13821
rect 6092 13812 6144 13864
rect 6276 13812 6328 13864
rect 9220 14016 9272 14068
rect 9864 13948 9916 14000
rect 14188 14016 14240 14068
rect 17960 14016 18012 14068
rect 19432 14059 19484 14068
rect 19432 14025 19441 14059
rect 19441 14025 19475 14059
rect 19475 14025 19484 14059
rect 19432 14016 19484 14025
rect 19708 14059 19760 14068
rect 19708 14025 19717 14059
rect 19717 14025 19751 14059
rect 19751 14025 19760 14059
rect 19708 14016 19760 14025
rect 8208 13880 8260 13932
rect 13544 13948 13596 14000
rect 6828 13855 6880 13864
rect 6828 13821 6837 13855
rect 6837 13821 6871 13855
rect 6871 13821 6880 13855
rect 6828 13812 6880 13821
rect 8392 13812 8444 13864
rect 9772 13812 9824 13864
rect 12440 13880 12492 13932
rect 12624 13880 12676 13932
rect 13268 13880 13320 13932
rect 10416 13855 10468 13864
rect 10416 13821 10425 13855
rect 10425 13821 10459 13855
rect 10459 13821 10468 13855
rect 10416 13812 10468 13821
rect 11152 13812 11204 13864
rect 12808 13855 12860 13864
rect 12808 13821 12817 13855
rect 12817 13821 12851 13855
rect 12851 13821 12860 13855
rect 12808 13812 12860 13821
rect 13452 13812 13504 13864
rect 13636 13812 13688 13864
rect 16580 13948 16632 14000
rect 14188 13880 14240 13932
rect 15292 13855 15344 13864
rect 15292 13821 15301 13855
rect 15301 13821 15335 13855
rect 15335 13821 15344 13855
rect 15292 13812 15344 13821
rect 17408 13880 17460 13932
rect 17868 13812 17920 13864
rect 1860 13719 1912 13728
rect 1860 13685 1869 13719
rect 1869 13685 1903 13719
rect 1903 13685 1912 13719
rect 1860 13676 1912 13685
rect 2504 13676 2556 13728
rect 3700 13676 3752 13728
rect 4252 13719 4304 13728
rect 4252 13685 4261 13719
rect 4261 13685 4295 13719
rect 4295 13685 4304 13719
rect 4252 13676 4304 13685
rect 5632 13676 5684 13728
rect 5816 13676 5868 13728
rect 7380 13744 7432 13796
rect 13084 13744 13136 13796
rect 8208 13719 8260 13728
rect 8208 13685 8217 13719
rect 8217 13685 8251 13719
rect 8251 13685 8260 13719
rect 8208 13676 8260 13685
rect 8300 13676 8352 13728
rect 8576 13676 8628 13728
rect 9128 13676 9180 13728
rect 9496 13676 9548 13728
rect 12348 13676 12400 13728
rect 12440 13676 12492 13728
rect 13360 13676 13412 13728
rect 13820 13719 13872 13728
rect 13820 13685 13829 13719
rect 13829 13685 13863 13719
rect 13863 13685 13872 13719
rect 13820 13676 13872 13685
rect 15752 13744 15804 13796
rect 16764 13744 16816 13796
rect 16948 13744 17000 13796
rect 17960 13744 18012 13796
rect 21088 13812 21140 13864
rect 18328 13787 18380 13796
rect 18328 13753 18362 13787
rect 18362 13753 18380 13787
rect 18328 13744 18380 13753
rect 16672 13719 16724 13728
rect 16672 13685 16681 13719
rect 16681 13685 16715 13719
rect 16715 13685 16724 13719
rect 16672 13676 16724 13685
rect 17224 13676 17276 13728
rect 19432 13744 19484 13796
rect 19616 13744 19668 13796
rect 18972 13676 19024 13728
rect 19892 13676 19944 13728
rect 20904 13719 20956 13728
rect 20904 13685 20913 13719
rect 20913 13685 20947 13719
rect 20947 13685 20956 13719
rect 20904 13676 20956 13685
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 3240 13472 3292 13524
rect 5540 13515 5592 13524
rect 5540 13481 5549 13515
rect 5549 13481 5583 13515
rect 5583 13481 5592 13515
rect 5540 13472 5592 13481
rect 5172 13404 5224 13456
rect 6920 13472 6972 13524
rect 7196 13472 7248 13524
rect 7748 13472 7800 13524
rect 8300 13515 8352 13524
rect 8300 13481 8309 13515
rect 8309 13481 8343 13515
rect 8343 13481 8352 13515
rect 8300 13472 8352 13481
rect 12440 13472 12492 13524
rect 13084 13472 13136 13524
rect 1952 13336 2004 13388
rect 2136 13336 2188 13388
rect 2872 13336 2924 13388
rect 4068 13336 4120 13388
rect 5816 13336 5868 13388
rect 7196 13336 7248 13388
rect 8392 13404 8444 13456
rect 10692 13404 10744 13456
rect 4804 13268 4856 13320
rect 5724 13268 5776 13320
rect 8484 13311 8536 13320
rect 8484 13277 8493 13311
rect 8493 13277 8527 13311
rect 8527 13277 8536 13311
rect 8484 13268 8536 13277
rect 9864 13336 9916 13388
rect 10968 13336 11020 13388
rect 12624 13404 12676 13456
rect 12348 13336 12400 13388
rect 12440 13336 12492 13388
rect 13728 13404 13780 13456
rect 14188 13404 14240 13456
rect 15016 13404 15068 13456
rect 17132 13472 17184 13524
rect 17960 13472 18012 13524
rect 18788 13472 18840 13524
rect 13452 13336 13504 13388
rect 13912 13336 13964 13388
rect 15108 13336 15160 13388
rect 15384 13336 15436 13388
rect 15568 13336 15620 13388
rect 15936 13379 15988 13388
rect 15936 13345 15945 13379
rect 15945 13345 15979 13379
rect 15979 13345 15988 13379
rect 18420 13404 18472 13456
rect 15936 13336 15988 13345
rect 16764 13379 16816 13388
rect 16764 13345 16773 13379
rect 16773 13345 16807 13379
rect 16807 13345 16816 13379
rect 16764 13336 16816 13345
rect 16948 13336 17000 13388
rect 18972 13336 19024 13388
rect 9220 13268 9272 13320
rect 13360 13268 13412 13320
rect 14648 13268 14700 13320
rect 15476 13268 15528 13320
rect 16028 13311 16080 13320
rect 16028 13277 16037 13311
rect 16037 13277 16071 13311
rect 16071 13277 16080 13311
rect 16028 13268 16080 13277
rect 3608 13243 3660 13252
rect 3608 13209 3617 13243
rect 3617 13209 3651 13243
rect 3651 13209 3660 13243
rect 3608 13200 3660 13209
rect 4528 13200 4580 13252
rect 6920 13132 6972 13184
rect 9680 13132 9732 13184
rect 10048 13132 10100 13184
rect 11152 13175 11204 13184
rect 11152 13141 11161 13175
rect 11161 13141 11195 13175
rect 11195 13141 11204 13175
rect 11152 13132 11204 13141
rect 12716 13200 12768 13252
rect 15384 13200 15436 13252
rect 17960 13311 18012 13320
rect 17960 13277 17969 13311
rect 17969 13277 18003 13311
rect 18003 13277 18012 13311
rect 17960 13268 18012 13277
rect 18328 13268 18380 13320
rect 20904 13404 20956 13456
rect 19432 13336 19484 13388
rect 19708 13379 19760 13388
rect 19708 13345 19717 13379
rect 19717 13345 19751 13379
rect 19751 13345 19760 13379
rect 19708 13336 19760 13345
rect 12256 13132 12308 13184
rect 12992 13175 13044 13184
rect 12992 13141 13001 13175
rect 13001 13141 13035 13175
rect 13035 13141 13044 13175
rect 12992 13132 13044 13141
rect 13728 13132 13780 13184
rect 13912 13175 13964 13184
rect 13912 13141 13921 13175
rect 13921 13141 13955 13175
rect 13955 13141 13964 13175
rect 13912 13132 13964 13141
rect 14464 13132 14516 13184
rect 14924 13132 14976 13184
rect 15476 13175 15528 13184
rect 15476 13141 15485 13175
rect 15485 13141 15519 13175
rect 15519 13141 15528 13175
rect 15476 13132 15528 13141
rect 16396 13132 16448 13184
rect 17868 13132 17920 13184
rect 19340 13175 19392 13184
rect 19340 13141 19349 13175
rect 19349 13141 19383 13175
rect 19383 13141 19392 13175
rect 19340 13132 19392 13141
rect 19892 13132 19944 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 1492 12928 1544 12980
rect 4068 12971 4120 12980
rect 4068 12937 4077 12971
rect 4077 12937 4111 12971
rect 4111 12937 4120 12971
rect 4068 12928 4120 12937
rect 4252 12928 4304 12980
rect 3976 12860 4028 12912
rect 6092 12928 6144 12980
rect 7196 12971 7248 12980
rect 7196 12937 7205 12971
rect 7205 12937 7239 12971
rect 7239 12937 7248 12971
rect 7196 12928 7248 12937
rect 8484 12928 8536 12980
rect 8944 12971 8996 12980
rect 8944 12937 8953 12971
rect 8953 12937 8987 12971
rect 8987 12937 8996 12971
rect 8944 12928 8996 12937
rect 9220 12971 9272 12980
rect 9220 12937 9229 12971
rect 9229 12937 9263 12971
rect 9263 12937 9272 12971
rect 9220 12928 9272 12937
rect 14004 12928 14056 12980
rect 14188 12971 14240 12980
rect 14188 12937 14197 12971
rect 14197 12937 14231 12971
rect 14231 12937 14240 12971
rect 14188 12928 14240 12937
rect 2872 12792 2924 12844
rect 3700 12835 3752 12844
rect 3700 12801 3709 12835
rect 3709 12801 3743 12835
rect 3743 12801 3752 12835
rect 3700 12792 3752 12801
rect 4804 12792 4856 12844
rect 5632 12835 5684 12844
rect 5632 12801 5641 12835
rect 5641 12801 5675 12835
rect 5675 12801 5684 12835
rect 5632 12792 5684 12801
rect 6644 12860 6696 12912
rect 8576 12860 8628 12912
rect 4252 12724 4304 12776
rect 5448 12767 5500 12776
rect 5448 12733 5457 12767
rect 5457 12733 5491 12767
rect 5491 12733 5500 12767
rect 5448 12724 5500 12733
rect 7380 12767 7432 12776
rect 1676 12588 1728 12640
rect 2964 12588 3016 12640
rect 5172 12656 5224 12708
rect 7380 12733 7389 12767
rect 7389 12733 7423 12767
rect 7423 12733 7432 12767
rect 7380 12724 7432 12733
rect 10324 12792 10376 12844
rect 10508 12792 10560 12844
rect 10692 12792 10744 12844
rect 10876 12792 10928 12844
rect 11520 12860 11572 12912
rect 11796 12860 11848 12912
rect 12532 12835 12584 12844
rect 12532 12801 12541 12835
rect 12541 12801 12575 12835
rect 12575 12801 12584 12835
rect 12532 12792 12584 12801
rect 15292 12928 15344 12980
rect 15936 12928 15988 12980
rect 17868 12928 17920 12980
rect 16672 12792 16724 12844
rect 6828 12656 6880 12708
rect 7196 12656 7248 12708
rect 8208 12656 8260 12708
rect 10048 12656 10100 12708
rect 10140 12656 10192 12708
rect 3240 12588 3292 12640
rect 6184 12588 6236 12640
rect 8300 12588 8352 12640
rect 10416 12588 10468 12640
rect 10692 12588 10744 12640
rect 11612 12588 11664 12640
rect 11796 12588 11848 12640
rect 12072 12656 12124 12708
rect 12992 12656 13044 12708
rect 13728 12656 13780 12708
rect 14004 12724 14056 12776
rect 14280 12724 14332 12776
rect 14464 12724 14516 12776
rect 15384 12724 15436 12776
rect 17224 12767 17276 12776
rect 15016 12656 15068 12708
rect 12440 12588 12492 12640
rect 12716 12588 12768 12640
rect 16488 12656 16540 12708
rect 17224 12733 17233 12767
rect 17233 12733 17267 12767
rect 17267 12733 17276 12767
rect 17224 12724 17276 12733
rect 19524 12928 19576 12980
rect 20904 12971 20956 12980
rect 20904 12937 20913 12971
rect 20913 12937 20947 12971
rect 20947 12937 20956 12971
rect 20904 12928 20956 12937
rect 15936 12631 15988 12640
rect 15936 12597 15945 12631
rect 15945 12597 15979 12631
rect 15979 12597 15988 12631
rect 15936 12588 15988 12597
rect 17316 12588 17368 12640
rect 17960 12656 18012 12708
rect 18052 12656 18104 12708
rect 18328 12699 18380 12708
rect 18328 12665 18362 12699
rect 18362 12665 18380 12699
rect 18328 12656 18380 12665
rect 20352 12588 20404 12640
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 2320 12384 2372 12436
rect 2136 12316 2188 12368
rect 2320 12248 2372 12300
rect 2504 12384 2556 12436
rect 2872 12427 2924 12436
rect 2872 12393 2881 12427
rect 2881 12393 2915 12427
rect 2915 12393 2924 12427
rect 2872 12384 2924 12393
rect 3332 12427 3384 12436
rect 3332 12393 3341 12427
rect 3341 12393 3375 12427
rect 3375 12393 3384 12427
rect 3332 12384 3384 12393
rect 4160 12384 4212 12436
rect 5080 12384 5132 12436
rect 7012 12384 7064 12436
rect 7288 12384 7340 12436
rect 9680 12384 9732 12436
rect 11796 12427 11848 12436
rect 2596 12316 2648 12368
rect 7932 12316 7984 12368
rect 11796 12393 11805 12427
rect 11805 12393 11839 12427
rect 11839 12393 11848 12427
rect 11796 12384 11848 12393
rect 2504 12248 2556 12300
rect 3148 12291 3200 12300
rect 3148 12257 3157 12291
rect 3157 12257 3191 12291
rect 3191 12257 3200 12291
rect 3148 12248 3200 12257
rect 5448 12248 5500 12300
rect 7196 12291 7248 12300
rect 3700 12180 3752 12232
rect 4528 12112 4580 12164
rect 4896 12112 4948 12164
rect 3608 12044 3660 12096
rect 6736 12044 6788 12096
rect 6920 12087 6972 12096
rect 6920 12053 6929 12087
rect 6929 12053 6963 12087
rect 6963 12053 6972 12087
rect 6920 12044 6972 12053
rect 7196 12257 7205 12291
rect 7205 12257 7239 12291
rect 7239 12257 7248 12291
rect 7196 12248 7248 12257
rect 7840 12248 7892 12300
rect 8024 12248 8076 12300
rect 11060 12291 11112 12300
rect 11060 12257 11069 12291
rect 11069 12257 11103 12291
rect 11103 12257 11112 12291
rect 11060 12248 11112 12257
rect 7196 12112 7248 12164
rect 12808 12316 12860 12368
rect 13636 12384 13688 12436
rect 15292 12384 15344 12436
rect 16396 12384 16448 12436
rect 16948 12384 17000 12436
rect 17868 12384 17920 12436
rect 18420 12384 18472 12436
rect 19156 12384 19208 12436
rect 19800 12384 19852 12436
rect 13912 12316 13964 12368
rect 12624 12248 12676 12300
rect 13360 12291 13412 12300
rect 13360 12257 13369 12291
rect 13369 12257 13403 12291
rect 13403 12257 13412 12291
rect 13360 12248 13412 12257
rect 15292 12291 15344 12300
rect 15292 12257 15301 12291
rect 15301 12257 15335 12291
rect 15335 12257 15344 12291
rect 15292 12248 15344 12257
rect 8760 12112 8812 12164
rect 11152 12112 11204 12164
rect 8668 12044 8720 12096
rect 9772 12044 9824 12096
rect 11336 12112 11388 12164
rect 11704 12112 11756 12164
rect 13268 12180 13320 12232
rect 13544 12180 13596 12232
rect 14188 12180 14240 12232
rect 14648 12223 14700 12232
rect 14648 12189 14657 12223
rect 14657 12189 14691 12223
rect 14691 12189 14700 12223
rect 14648 12180 14700 12189
rect 15016 12180 15068 12232
rect 15936 12248 15988 12300
rect 16028 12248 16080 12300
rect 16856 12291 16908 12300
rect 16856 12257 16865 12291
rect 16865 12257 16899 12291
rect 16899 12257 16908 12291
rect 16856 12248 16908 12257
rect 18052 12291 18104 12300
rect 18052 12257 18061 12291
rect 18061 12257 18095 12291
rect 18095 12257 18104 12291
rect 18052 12248 18104 12257
rect 18144 12248 18196 12300
rect 19340 12248 19392 12300
rect 20536 12248 20588 12300
rect 14740 12112 14792 12164
rect 17776 12180 17828 12232
rect 12900 12087 12952 12096
rect 12900 12053 12909 12087
rect 12909 12053 12943 12087
rect 12943 12053 12952 12087
rect 12900 12044 12952 12053
rect 13360 12044 13412 12096
rect 13636 12044 13688 12096
rect 15568 12044 15620 12096
rect 15936 12044 15988 12096
rect 19064 12044 19116 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 2964 11840 3016 11892
rect 3516 11840 3568 11892
rect 4804 11840 4856 11892
rect 5356 11840 5408 11892
rect 7656 11840 7708 11892
rect 8024 11883 8076 11892
rect 8024 11849 8033 11883
rect 8033 11849 8067 11883
rect 8067 11849 8076 11883
rect 8024 11840 8076 11849
rect 8300 11840 8352 11892
rect 9036 11840 9088 11892
rect 9312 11840 9364 11892
rect 3700 11772 3752 11824
rect 4988 11772 5040 11824
rect 7196 11772 7248 11824
rect 4252 11747 4304 11756
rect 3608 11679 3660 11688
rect 3608 11645 3617 11679
rect 3617 11645 3651 11679
rect 3651 11645 3660 11679
rect 3608 11636 3660 11645
rect 2136 11568 2188 11620
rect 4252 11713 4261 11747
rect 4261 11713 4295 11747
rect 4295 11713 4304 11747
rect 4252 11704 4304 11713
rect 5448 11704 5500 11756
rect 6920 11704 6972 11756
rect 7656 11747 7708 11756
rect 7656 11713 7665 11747
rect 7665 11713 7699 11747
rect 7699 11713 7708 11747
rect 7656 11704 7708 11713
rect 7840 11704 7892 11756
rect 8668 11636 8720 11688
rect 8944 11704 8996 11756
rect 9220 11704 9272 11756
rect 10968 11772 11020 11824
rect 13360 11840 13412 11892
rect 15200 11883 15252 11892
rect 15200 11849 15209 11883
rect 15209 11849 15243 11883
rect 15243 11849 15252 11883
rect 15200 11840 15252 11849
rect 9864 11704 9916 11756
rect 14740 11747 14792 11756
rect 14740 11713 14749 11747
rect 14749 11713 14783 11747
rect 14783 11713 14792 11747
rect 14740 11704 14792 11713
rect 17592 11883 17644 11892
rect 17592 11849 17601 11883
rect 17601 11849 17635 11883
rect 17635 11849 17644 11883
rect 17592 11840 17644 11849
rect 17776 11840 17828 11892
rect 19156 11840 19208 11892
rect 19616 11840 19668 11892
rect 21456 11840 21508 11892
rect 19800 11772 19852 11824
rect 15936 11704 15988 11756
rect 16764 11747 16816 11756
rect 16764 11713 16773 11747
rect 16773 11713 16807 11747
rect 16807 11713 16816 11747
rect 16764 11704 16816 11713
rect 16856 11704 16908 11756
rect 11796 11679 11848 11688
rect 2320 11500 2372 11552
rect 3056 11500 3108 11552
rect 5080 11543 5132 11552
rect 5080 11509 5089 11543
rect 5089 11509 5123 11543
rect 5123 11509 5132 11543
rect 5080 11500 5132 11509
rect 6828 11500 6880 11552
rect 9220 11568 9272 11620
rect 11796 11645 11805 11679
rect 11805 11645 11839 11679
rect 11839 11645 11848 11679
rect 11796 11636 11848 11645
rect 12256 11636 12308 11688
rect 12532 11636 12584 11688
rect 15559 11679 15611 11688
rect 7104 11500 7156 11552
rect 8392 11543 8444 11552
rect 8392 11509 8401 11543
rect 8401 11509 8435 11543
rect 8435 11509 8444 11543
rect 8392 11500 8444 11509
rect 8484 11543 8536 11552
rect 8484 11509 8493 11543
rect 8493 11509 8527 11543
rect 8527 11509 8536 11543
rect 9128 11543 9180 11552
rect 8484 11500 8536 11509
rect 9128 11509 9137 11543
rect 9137 11509 9171 11543
rect 9171 11509 9180 11543
rect 9128 11500 9180 11509
rect 9588 11500 9640 11552
rect 11612 11568 11664 11620
rect 12808 11568 12860 11620
rect 15559 11645 15577 11679
rect 15577 11645 15611 11679
rect 15559 11636 15611 11645
rect 15752 11636 15804 11688
rect 17132 11636 17184 11688
rect 17684 11636 17736 11688
rect 20720 11679 20772 11688
rect 19616 11568 19668 11620
rect 20720 11645 20729 11679
rect 20729 11645 20763 11679
rect 20763 11645 20772 11679
rect 20720 11636 20772 11645
rect 20536 11568 20588 11620
rect 11796 11500 11848 11552
rect 12992 11500 13044 11552
rect 13912 11500 13964 11552
rect 15292 11500 15344 11552
rect 15476 11500 15528 11552
rect 15568 11500 15620 11552
rect 16396 11500 16448 11552
rect 16672 11543 16724 11552
rect 16672 11509 16681 11543
rect 16681 11509 16715 11543
rect 16715 11509 16724 11543
rect 16672 11500 16724 11509
rect 16948 11500 17000 11552
rect 19800 11500 19852 11552
rect 20720 11500 20772 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 2780 11296 2832 11348
rect 3700 11339 3752 11348
rect 3700 11305 3709 11339
rect 3709 11305 3743 11339
rect 3743 11305 3752 11339
rect 3700 11296 3752 11305
rect 5080 11296 5132 11348
rect 7380 11296 7432 11348
rect 7656 11296 7708 11348
rect 8484 11296 8536 11348
rect 9864 11296 9916 11348
rect 10140 11296 10192 11348
rect 11060 11296 11112 11348
rect 12808 11296 12860 11348
rect 13820 11296 13872 11348
rect 14004 11296 14056 11348
rect 15292 11339 15344 11348
rect 15292 11305 15301 11339
rect 15301 11305 15335 11339
rect 15335 11305 15344 11339
rect 15292 11296 15344 11305
rect 15660 11339 15712 11348
rect 15660 11305 15669 11339
rect 15669 11305 15703 11339
rect 15703 11305 15712 11339
rect 15660 11296 15712 11305
rect 16396 11296 16448 11348
rect 16580 11296 16632 11348
rect 17316 11296 17368 11348
rect 18788 11339 18840 11348
rect 18788 11305 18797 11339
rect 18797 11305 18831 11339
rect 18831 11305 18840 11339
rect 18788 11296 18840 11305
rect 19340 11296 19392 11348
rect 20812 11296 20864 11348
rect 2412 11228 2464 11280
rect 6920 11228 6972 11280
rect 8760 11271 8812 11280
rect 8760 11237 8769 11271
rect 8769 11237 8803 11271
rect 8803 11237 8812 11271
rect 8760 11228 8812 11237
rect 9036 11228 9088 11280
rect 9588 11228 9640 11280
rect 11336 11228 11388 11280
rect 1768 11203 1820 11212
rect 1768 11169 1777 11203
rect 1777 11169 1811 11203
rect 1811 11169 1820 11203
rect 1768 11160 1820 11169
rect 2136 11160 2188 11212
rect 3792 11160 3844 11212
rect 5632 11160 5684 11212
rect 5816 11203 5868 11212
rect 5816 11169 5825 11203
rect 5825 11169 5859 11203
rect 5859 11169 5868 11203
rect 5816 11160 5868 11169
rect 4988 11135 5040 11144
rect 4988 11101 4997 11135
rect 4997 11101 5031 11135
rect 5031 11101 5040 11135
rect 4988 11092 5040 11101
rect 6736 11135 6788 11144
rect 2596 10956 2648 11008
rect 6092 11024 6144 11076
rect 6736 11101 6745 11135
rect 6745 11101 6779 11135
rect 6779 11101 6788 11135
rect 6736 11092 6788 11101
rect 9680 11160 9732 11212
rect 10140 11160 10192 11212
rect 10324 11160 10376 11212
rect 8208 11092 8260 11144
rect 10048 11092 10100 11144
rect 10784 11092 10836 11144
rect 11060 11092 11112 11144
rect 11520 11092 11572 11144
rect 14556 11228 14608 11280
rect 13084 11203 13136 11212
rect 13084 11169 13093 11203
rect 13093 11169 13127 11203
rect 13127 11169 13136 11203
rect 13084 11160 13136 11169
rect 13636 11160 13688 11212
rect 15660 11160 15712 11212
rect 16580 11160 16632 11212
rect 17040 11160 17092 11212
rect 17684 11203 17736 11212
rect 12256 11092 12308 11144
rect 12532 11024 12584 11076
rect 12992 11092 13044 11144
rect 13360 11135 13412 11144
rect 13360 11101 13369 11135
rect 13369 11101 13403 11135
rect 13403 11101 13412 11135
rect 14280 11135 14332 11144
rect 13360 11092 13412 11101
rect 13820 11024 13872 11076
rect 14280 11101 14289 11135
rect 14289 11101 14323 11135
rect 14323 11101 14332 11135
rect 14280 11092 14332 11101
rect 14648 11135 14700 11144
rect 14648 11101 14657 11135
rect 14657 11101 14691 11135
rect 14691 11101 14700 11135
rect 14648 11092 14700 11101
rect 15016 11092 15068 11144
rect 15568 11092 15620 11144
rect 16770 11135 16822 11144
rect 16770 11101 16773 11135
rect 16773 11101 16807 11135
rect 16807 11101 16822 11135
rect 16770 11092 16822 11101
rect 17408 11092 17460 11144
rect 17684 11169 17693 11203
rect 17693 11169 17727 11203
rect 17727 11169 17736 11203
rect 17684 11160 17736 11169
rect 17960 11160 18012 11212
rect 20628 11228 20680 11280
rect 20168 11160 20220 11212
rect 18788 11092 18840 11144
rect 18880 11092 18932 11144
rect 16488 11024 16540 11076
rect 7380 10956 7432 11008
rect 8300 10956 8352 11008
rect 8484 10956 8536 11008
rect 10508 10956 10560 11008
rect 11980 10956 12032 11008
rect 13912 10956 13964 11008
rect 17316 10999 17368 11008
rect 17316 10965 17325 10999
rect 17325 10965 17359 10999
rect 17359 10965 17368 10999
rect 17316 10956 17368 10965
rect 18512 10956 18564 11008
rect 18788 10956 18840 11008
rect 21272 11024 21324 11076
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 1676 10795 1728 10804
rect 1676 10761 1685 10795
rect 1685 10761 1719 10795
rect 1719 10761 1728 10795
rect 1676 10752 1728 10761
rect 2964 10752 3016 10804
rect 6000 10752 6052 10804
rect 6552 10752 6604 10804
rect 6828 10752 6880 10804
rect 13176 10752 13228 10804
rect 3792 10684 3844 10736
rect 2320 10659 2372 10668
rect 2320 10625 2329 10659
rect 2329 10625 2363 10659
rect 2363 10625 2372 10659
rect 2320 10616 2372 10625
rect 3424 10616 3476 10668
rect 5356 10684 5408 10736
rect 9772 10684 9824 10736
rect 11612 10684 11664 10736
rect 15200 10684 15252 10736
rect 16580 10752 16632 10804
rect 20628 10752 20680 10804
rect 17224 10684 17276 10736
rect 5448 10659 5500 10668
rect 5448 10625 5457 10659
rect 5457 10625 5491 10659
rect 5491 10625 5500 10659
rect 5448 10616 5500 10625
rect 5632 10616 5684 10668
rect 6000 10616 6052 10668
rect 7472 10659 7524 10668
rect 1492 10548 1544 10600
rect 2320 10480 2372 10532
rect 2596 10480 2648 10532
rect 4896 10548 4948 10600
rect 7472 10625 7481 10659
rect 7481 10625 7515 10659
rect 7515 10625 7524 10659
rect 7472 10616 7524 10625
rect 8208 10616 8260 10668
rect 11796 10616 11848 10668
rect 13728 10616 13780 10668
rect 14280 10616 14332 10668
rect 17408 10659 17460 10668
rect 17408 10625 17417 10659
rect 17417 10625 17451 10659
rect 17451 10625 17460 10659
rect 17408 10616 17460 10625
rect 17868 10616 17920 10668
rect 18512 10616 18564 10668
rect 8116 10548 8168 10600
rect 9128 10548 9180 10600
rect 9312 10548 9364 10600
rect 9680 10548 9732 10600
rect 6736 10480 6788 10532
rect 12256 10548 12308 10600
rect 12440 10591 12492 10600
rect 12440 10557 12449 10591
rect 12449 10557 12483 10591
rect 12483 10557 12492 10591
rect 12440 10548 12492 10557
rect 12992 10548 13044 10600
rect 13176 10548 13228 10600
rect 15016 10548 15068 10600
rect 15292 10548 15344 10600
rect 15936 10548 15988 10600
rect 16580 10548 16632 10600
rect 16856 10548 16908 10600
rect 18328 10548 18380 10600
rect 18696 10548 18748 10600
rect 18880 10548 18932 10600
rect 10968 10480 11020 10532
rect 11796 10480 11848 10532
rect 12164 10480 12216 10532
rect 13360 10480 13412 10532
rect 13728 10480 13780 10532
rect 1768 10412 1820 10464
rect 2136 10455 2188 10464
rect 2136 10421 2145 10455
rect 2145 10421 2179 10455
rect 2179 10421 2188 10455
rect 3608 10455 3660 10464
rect 2136 10412 2188 10421
rect 3608 10421 3617 10455
rect 3617 10421 3651 10455
rect 3651 10421 3660 10455
rect 3608 10412 3660 10421
rect 3976 10455 4028 10464
rect 3976 10421 3985 10455
rect 3985 10421 4019 10455
rect 4019 10421 4028 10455
rect 3976 10412 4028 10421
rect 5172 10455 5224 10464
rect 5172 10421 5181 10455
rect 5181 10421 5215 10455
rect 5215 10421 5224 10455
rect 5172 10412 5224 10421
rect 6184 10412 6236 10464
rect 7380 10412 7432 10464
rect 8668 10412 8720 10464
rect 8852 10455 8904 10464
rect 8852 10421 8861 10455
rect 8861 10421 8895 10455
rect 8895 10421 8904 10455
rect 8852 10412 8904 10421
rect 9220 10412 9272 10464
rect 9588 10412 9640 10464
rect 12716 10412 12768 10464
rect 12992 10412 13044 10464
rect 17868 10480 17920 10532
rect 20444 10480 20496 10532
rect 14188 10412 14240 10464
rect 15200 10412 15252 10464
rect 16488 10412 16540 10464
rect 16856 10412 16908 10464
rect 17224 10455 17276 10464
rect 17224 10421 17233 10455
rect 17233 10421 17267 10455
rect 17267 10421 17276 10455
rect 17224 10412 17276 10421
rect 17684 10412 17736 10464
rect 18972 10412 19024 10464
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 1768 10251 1820 10260
rect 1768 10217 1777 10251
rect 1777 10217 1811 10251
rect 1811 10217 1820 10251
rect 1768 10208 1820 10217
rect 1860 10208 1912 10260
rect 3056 10208 3108 10260
rect 3608 10208 3660 10260
rect 5172 10208 5224 10260
rect 3516 10140 3568 10192
rect 6000 10208 6052 10260
rect 6184 10251 6236 10260
rect 6184 10217 6193 10251
rect 6193 10217 6227 10251
rect 6227 10217 6236 10251
rect 6184 10208 6236 10217
rect 6092 10183 6144 10192
rect 2872 10072 2924 10124
rect 3884 10072 3936 10124
rect 6092 10149 6101 10183
rect 6101 10149 6135 10183
rect 6135 10149 6144 10183
rect 6092 10140 6144 10149
rect 5080 10072 5132 10124
rect 6644 10140 6696 10192
rect 7104 10140 7156 10192
rect 7656 10183 7708 10192
rect 7656 10149 7690 10183
rect 7690 10149 7708 10183
rect 7656 10140 7708 10149
rect 8208 10208 8260 10260
rect 10968 10208 11020 10260
rect 11152 10208 11204 10260
rect 12808 10208 12860 10260
rect 17684 10251 17736 10260
rect 17684 10217 17693 10251
rect 17693 10217 17727 10251
rect 17727 10217 17736 10251
rect 17684 10208 17736 10217
rect 7288 10115 7340 10124
rect 7288 10081 7297 10115
rect 7297 10081 7331 10115
rect 7331 10081 7340 10115
rect 7288 10072 7340 10081
rect 8208 10072 8260 10124
rect 9680 10115 9732 10124
rect 9680 10081 9689 10115
rect 9689 10081 9723 10115
rect 9723 10081 9732 10115
rect 9680 10072 9732 10081
rect 10508 10072 10560 10124
rect 10784 10072 10836 10124
rect 11980 10140 12032 10192
rect 13636 10140 13688 10192
rect 15200 10140 15252 10192
rect 19800 10208 19852 10260
rect 20076 10208 20128 10260
rect 20444 10208 20496 10260
rect 3608 10047 3660 10056
rect 3608 10013 3617 10047
rect 3617 10013 3651 10047
rect 3651 10013 3660 10047
rect 3608 10004 3660 10013
rect 4068 10047 4120 10056
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 6184 10004 6236 10056
rect 11060 10004 11112 10056
rect 11980 10047 12032 10056
rect 11980 10013 11989 10047
rect 11989 10013 12023 10047
rect 12023 10013 12032 10047
rect 11980 10004 12032 10013
rect 12808 10047 12860 10056
rect 12808 10013 12817 10047
rect 12817 10013 12851 10047
rect 12851 10013 12860 10047
rect 12808 10004 12860 10013
rect 14556 10115 14608 10124
rect 2780 9868 2832 9920
rect 5356 9936 5408 9988
rect 3976 9868 4028 9920
rect 7288 9936 7340 9988
rect 8668 9936 8720 9988
rect 9680 9936 9732 9988
rect 11704 9936 11756 9988
rect 12164 9936 12216 9988
rect 6920 9868 6972 9920
rect 7196 9868 7248 9920
rect 10876 9868 10928 9920
rect 11060 9868 11112 9920
rect 13360 9911 13412 9920
rect 13360 9877 13369 9911
rect 13369 9877 13403 9911
rect 13403 9877 13412 9911
rect 13360 9868 13412 9877
rect 14556 10081 14565 10115
rect 14565 10081 14599 10115
rect 14599 10081 14608 10115
rect 14556 10072 14608 10081
rect 14464 10004 14516 10056
rect 15292 10072 15344 10124
rect 15568 10004 15620 10056
rect 17684 10072 17736 10124
rect 17960 10072 18012 10124
rect 18420 10115 18472 10124
rect 18420 10081 18429 10115
rect 18429 10081 18463 10115
rect 18463 10081 18472 10115
rect 18420 10072 18472 10081
rect 22468 10140 22520 10192
rect 18880 10072 18932 10124
rect 19524 10072 19576 10124
rect 15844 10004 15896 10056
rect 16028 10004 16080 10056
rect 16764 10047 16816 10056
rect 16764 10013 16773 10047
rect 16773 10013 16807 10047
rect 16807 10013 16816 10047
rect 16764 10004 16816 10013
rect 16856 10047 16908 10056
rect 16856 10013 16865 10047
rect 16865 10013 16899 10047
rect 16899 10013 16908 10047
rect 17868 10047 17920 10056
rect 16856 10004 16908 10013
rect 17868 10013 17877 10047
rect 17877 10013 17911 10047
rect 17911 10013 17920 10047
rect 17868 10004 17920 10013
rect 18328 10004 18380 10056
rect 18696 10004 18748 10056
rect 14556 9868 14608 9920
rect 16120 9936 16172 9988
rect 16764 9868 16816 9920
rect 17040 9868 17092 9920
rect 19340 9868 19392 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 2136 9664 2188 9716
rect 2872 9707 2924 9716
rect 2872 9673 2881 9707
rect 2881 9673 2915 9707
rect 2915 9673 2924 9707
rect 2872 9664 2924 9673
rect 7196 9664 7248 9716
rect 8300 9664 8352 9716
rect 5356 9596 5408 9648
rect 2044 9528 2096 9580
rect 2780 9528 2832 9580
rect 3792 9528 3844 9580
rect 5816 9528 5868 9580
rect 10508 9639 10560 9648
rect 10508 9605 10517 9639
rect 10517 9605 10551 9639
rect 10551 9605 10560 9639
rect 10508 9596 10560 9605
rect 13176 9664 13228 9716
rect 14188 9664 14240 9716
rect 15292 9664 15344 9716
rect 15568 9664 15620 9716
rect 15844 9664 15896 9716
rect 16212 9596 16264 9648
rect 19248 9596 19300 9648
rect 2228 9503 2280 9512
rect 2228 9469 2237 9503
rect 2237 9469 2271 9503
rect 2271 9469 2280 9503
rect 2228 9460 2280 9469
rect 3700 9460 3752 9512
rect 4068 9460 4120 9512
rect 6184 9460 6236 9512
rect 6828 9503 6880 9512
rect 6828 9469 6837 9503
rect 6837 9469 6871 9503
rect 6871 9469 6880 9503
rect 6828 9460 6880 9469
rect 11060 9528 11112 9580
rect 7472 9460 7524 9512
rect 8208 9460 8260 9512
rect 10508 9460 10560 9512
rect 10876 9460 10928 9512
rect 12440 9503 12492 9512
rect 12440 9469 12449 9503
rect 12449 9469 12483 9503
rect 12483 9469 12492 9503
rect 12440 9460 12492 9469
rect 12992 9460 13044 9512
rect 3332 9367 3384 9376
rect 3332 9333 3341 9367
rect 3341 9333 3375 9367
rect 3375 9333 3384 9367
rect 3332 9324 3384 9333
rect 4068 9324 4120 9376
rect 5356 9324 5408 9376
rect 5448 9324 5500 9376
rect 6184 9324 6236 9376
rect 9588 9392 9640 9444
rect 10232 9392 10284 9444
rect 10508 9324 10560 9376
rect 11704 9392 11756 9444
rect 13176 9392 13228 9444
rect 16764 9571 16816 9580
rect 16764 9537 16773 9571
rect 16773 9537 16807 9571
rect 16807 9537 16816 9571
rect 16764 9528 16816 9537
rect 20352 9571 20404 9580
rect 15200 9460 15252 9512
rect 20352 9537 20361 9571
rect 20361 9537 20395 9571
rect 20395 9537 20404 9571
rect 20352 9528 20404 9537
rect 17408 9503 17460 9512
rect 17408 9469 17417 9503
rect 17417 9469 17451 9503
rect 17451 9469 17460 9503
rect 17408 9460 17460 9469
rect 17684 9460 17736 9512
rect 18144 9460 18196 9512
rect 19432 9460 19484 9512
rect 20720 9503 20772 9512
rect 20720 9469 20729 9503
rect 20729 9469 20763 9503
rect 20763 9469 20772 9503
rect 20720 9460 20772 9469
rect 15568 9392 15620 9444
rect 11152 9367 11204 9376
rect 11152 9333 11161 9367
rect 11161 9333 11195 9367
rect 11195 9333 11204 9367
rect 11152 9324 11204 9333
rect 13820 9367 13872 9376
rect 13820 9333 13829 9367
rect 13829 9333 13863 9367
rect 13863 9333 13872 9367
rect 13820 9324 13872 9333
rect 14188 9367 14240 9376
rect 14188 9333 14197 9367
rect 14197 9333 14231 9367
rect 14231 9333 14240 9367
rect 14188 9324 14240 9333
rect 14464 9324 14516 9376
rect 17224 9392 17276 9444
rect 18512 9392 18564 9444
rect 16028 9367 16080 9376
rect 16028 9333 16037 9367
rect 16037 9333 16071 9367
rect 16071 9333 16080 9367
rect 16028 9324 16080 9333
rect 16672 9367 16724 9376
rect 16672 9333 16681 9367
rect 16681 9333 16715 9367
rect 16715 9333 16724 9367
rect 16672 9324 16724 9333
rect 17868 9324 17920 9376
rect 19524 9324 19576 9376
rect 19708 9367 19760 9376
rect 19708 9333 19717 9367
rect 19717 9333 19751 9367
rect 19751 9333 19760 9367
rect 19708 9324 19760 9333
rect 20076 9367 20128 9376
rect 20076 9333 20085 9367
rect 20085 9333 20119 9367
rect 20119 9333 20128 9367
rect 20076 9324 20128 9333
rect 20168 9367 20220 9376
rect 20168 9333 20177 9367
rect 20177 9333 20211 9367
rect 20211 9333 20220 9367
rect 20168 9324 20220 9333
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 5080 9120 5132 9172
rect 5724 9120 5776 9172
rect 6368 9163 6420 9172
rect 4896 9052 4948 9104
rect 2596 9027 2648 9036
rect 2596 8993 2630 9027
rect 2630 8993 2648 9027
rect 2596 8984 2648 8993
rect 5172 8984 5224 9036
rect 1584 8916 1636 8968
rect 4344 8916 4396 8968
rect 5080 8916 5132 8968
rect 5816 9052 5868 9104
rect 6368 9129 6377 9163
rect 6377 9129 6411 9163
rect 6411 9129 6420 9163
rect 6368 9120 6420 9129
rect 6736 9120 6788 9172
rect 7380 9120 7432 9172
rect 8944 9120 8996 9172
rect 10232 9120 10284 9172
rect 11152 9120 11204 9172
rect 11704 9120 11756 9172
rect 13360 9120 13412 9172
rect 14556 9120 14608 9172
rect 6184 9052 6236 9104
rect 5632 8984 5684 9036
rect 6368 8984 6420 9036
rect 6552 8959 6604 8968
rect 6552 8925 6561 8959
rect 6561 8925 6595 8959
rect 6595 8925 6604 8959
rect 6552 8916 6604 8925
rect 8852 9052 8904 9104
rect 9588 9052 9640 9104
rect 11428 9052 11480 9104
rect 16028 9052 16080 9104
rect 16672 9120 16724 9172
rect 17960 9163 18012 9172
rect 17960 9129 17969 9163
rect 17969 9129 18003 9163
rect 18003 9129 18012 9163
rect 17960 9120 18012 9129
rect 19708 9120 19760 9172
rect 17868 9052 17920 9104
rect 18880 9052 18932 9104
rect 21180 9120 21232 9172
rect 20720 9052 20772 9104
rect 6736 8848 6788 8900
rect 9128 8984 9180 9036
rect 10784 8984 10836 9036
rect 11704 8984 11756 9036
rect 8852 8916 8904 8968
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 10232 8916 10284 8925
rect 10968 8916 11020 8968
rect 11244 8959 11296 8968
rect 11244 8925 11253 8959
rect 11253 8925 11287 8959
rect 11287 8925 11296 8959
rect 11244 8916 11296 8925
rect 11428 8959 11480 8968
rect 11428 8925 11437 8959
rect 11437 8925 11471 8959
rect 11471 8925 11480 8959
rect 11428 8916 11480 8925
rect 11980 8916 12032 8968
rect 12348 8959 12400 8968
rect 12348 8925 12357 8959
rect 12357 8925 12391 8959
rect 12391 8925 12400 8959
rect 12348 8916 12400 8925
rect 12256 8848 12308 8900
rect 12440 8848 12492 8900
rect 13268 8984 13320 9036
rect 15384 8984 15436 9036
rect 16672 8984 16724 9036
rect 19708 8984 19760 9036
rect 19984 9027 20036 9036
rect 19984 8993 19993 9027
rect 19993 8993 20027 9027
rect 20027 8993 20036 9027
rect 19984 8984 20036 8993
rect 15200 8916 15252 8968
rect 16856 8916 16908 8968
rect 18604 8959 18656 8968
rect 18604 8925 18613 8959
rect 18613 8925 18647 8959
rect 18647 8925 18656 8959
rect 18604 8916 18656 8925
rect 19248 8916 19300 8968
rect 19616 8959 19668 8968
rect 19616 8925 19625 8959
rect 19625 8925 19659 8959
rect 19659 8925 19668 8959
rect 19616 8916 19668 8925
rect 20352 8916 20404 8968
rect 13268 8848 13320 8900
rect 18788 8848 18840 8900
rect 18972 8891 19024 8900
rect 18972 8857 18981 8891
rect 18981 8857 19015 8891
rect 19015 8857 19024 8891
rect 18972 8848 19024 8857
rect 7380 8780 7432 8832
rect 8024 8780 8076 8832
rect 8392 8780 8444 8832
rect 8668 8780 8720 8832
rect 11152 8780 11204 8832
rect 13360 8780 13412 8832
rect 14280 8780 14332 8832
rect 14648 8780 14700 8832
rect 15200 8780 15252 8832
rect 15476 8780 15528 8832
rect 15568 8780 15620 8832
rect 16764 8780 16816 8832
rect 19984 8780 20036 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 3700 8576 3752 8628
rect 2596 8508 2648 8560
rect 1492 8372 1544 8424
rect 3700 8415 3752 8424
rect 3700 8381 3709 8415
rect 3709 8381 3743 8415
rect 3743 8381 3752 8415
rect 3700 8372 3752 8381
rect 9588 8576 9640 8628
rect 10232 8576 10284 8628
rect 13176 8576 13228 8628
rect 13820 8576 13872 8628
rect 15660 8576 15712 8628
rect 16488 8576 16540 8628
rect 17960 8576 18012 8628
rect 18604 8576 18656 8628
rect 18880 8576 18932 8628
rect 19432 8576 19484 8628
rect 6828 8508 6880 8560
rect 7012 8508 7064 8560
rect 9864 8508 9916 8560
rect 7288 8483 7340 8492
rect 2136 8304 2188 8356
rect 5172 8372 5224 8424
rect 6920 8372 6972 8424
rect 3976 8347 4028 8356
rect 3976 8313 4010 8347
rect 4010 8313 4028 8347
rect 3976 8304 4028 8313
rect 3884 8236 3936 8288
rect 7012 8304 7064 8356
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 7472 8483 7524 8492
rect 7472 8449 7481 8483
rect 7481 8449 7515 8483
rect 7515 8449 7524 8483
rect 7472 8440 7524 8449
rect 8024 8372 8076 8424
rect 8208 8372 8260 8424
rect 9864 8372 9916 8424
rect 8760 8304 8812 8356
rect 9128 8304 9180 8356
rect 11060 8508 11112 8560
rect 11612 8508 11664 8560
rect 12348 8508 12400 8560
rect 10324 8372 10376 8424
rect 10876 8440 10928 8492
rect 14004 8440 14056 8492
rect 14280 8440 14332 8492
rect 14648 8440 14700 8492
rect 15384 8440 15436 8492
rect 15568 8440 15620 8492
rect 15752 8440 15804 8492
rect 16764 8483 16816 8492
rect 16764 8449 16773 8483
rect 16773 8449 16807 8483
rect 16807 8449 16816 8483
rect 16764 8440 16816 8449
rect 17132 8508 17184 8560
rect 17684 8551 17736 8560
rect 17684 8517 17693 8551
rect 17693 8517 17727 8551
rect 17727 8517 17736 8551
rect 17684 8508 17736 8517
rect 18236 8440 18288 8492
rect 19340 8440 19392 8492
rect 20260 8508 20312 8560
rect 19616 8483 19668 8492
rect 19616 8449 19625 8483
rect 19625 8449 19659 8483
rect 19659 8449 19668 8483
rect 19616 8440 19668 8449
rect 10784 8372 10836 8424
rect 12072 8372 12124 8424
rect 13268 8372 13320 8424
rect 14188 8372 14240 8424
rect 17868 8415 17920 8424
rect 5724 8279 5776 8288
rect 5724 8245 5733 8279
rect 5733 8245 5767 8279
rect 5767 8245 5776 8279
rect 5724 8236 5776 8245
rect 6828 8279 6880 8288
rect 6828 8245 6837 8279
rect 6837 8245 6871 8279
rect 6871 8245 6880 8279
rect 6828 8236 6880 8245
rect 9312 8236 9364 8288
rect 9496 8236 9548 8288
rect 9864 8236 9916 8288
rect 15200 8304 15252 8356
rect 12440 8236 12492 8288
rect 12992 8236 13044 8288
rect 13912 8236 13964 8288
rect 15016 8236 15068 8288
rect 15568 8279 15620 8288
rect 15568 8245 15577 8279
rect 15577 8245 15611 8279
rect 15611 8245 15620 8279
rect 15568 8236 15620 8245
rect 16304 8304 16356 8356
rect 17868 8381 17877 8415
rect 17877 8381 17911 8415
rect 17911 8381 17920 8415
rect 17868 8372 17920 8381
rect 19432 8415 19484 8424
rect 19432 8381 19441 8415
rect 19441 8381 19475 8415
rect 19475 8381 19484 8415
rect 19432 8372 19484 8381
rect 19800 8372 19852 8424
rect 20536 8372 20588 8424
rect 17776 8304 17828 8356
rect 19708 8304 19760 8356
rect 20444 8347 20496 8356
rect 20444 8313 20453 8347
rect 20453 8313 20487 8347
rect 20487 8313 20496 8347
rect 20444 8304 20496 8313
rect 17592 8236 17644 8288
rect 18236 8236 18288 8288
rect 18420 8279 18472 8288
rect 18420 8245 18429 8279
rect 18429 8245 18463 8279
rect 18463 8245 18472 8279
rect 18420 8236 18472 8245
rect 19984 8236 20036 8288
rect 21364 8236 21416 8288
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 3056 8032 3108 8084
rect 3332 8032 3384 8084
rect 5724 8032 5776 8084
rect 6828 8032 6880 8084
rect 7012 8075 7064 8084
rect 7012 8041 7021 8075
rect 7021 8041 7055 8075
rect 7055 8041 7064 8075
rect 7012 8032 7064 8041
rect 7380 8075 7432 8084
rect 7380 8041 7389 8075
rect 7389 8041 7423 8075
rect 7423 8041 7432 8075
rect 7380 8032 7432 8041
rect 8668 8032 8720 8084
rect 10416 8032 10468 8084
rect 10784 8032 10836 8084
rect 11060 8032 11112 8084
rect 11704 8075 11756 8084
rect 11704 8041 11713 8075
rect 11713 8041 11747 8075
rect 11747 8041 11756 8075
rect 11704 8032 11756 8041
rect 13544 8032 13596 8084
rect 1676 7896 1728 7948
rect 2412 7896 2464 7948
rect 3976 7964 4028 8016
rect 3700 7896 3752 7948
rect 4896 7896 4948 7948
rect 5908 7964 5960 8016
rect 6736 7964 6788 8016
rect 8760 7964 8812 8016
rect 6920 7896 6972 7948
rect 9496 7896 9548 7948
rect 4160 7760 4212 7812
rect 7656 7828 7708 7880
rect 8116 7828 8168 7880
rect 9588 7828 9640 7880
rect 12532 7964 12584 8016
rect 10968 7896 11020 7948
rect 11612 7896 11664 7948
rect 13912 7964 13964 8016
rect 14464 7964 14516 8016
rect 15568 8032 15620 8084
rect 17776 8032 17828 8084
rect 17868 8032 17920 8084
rect 18972 8032 19024 8084
rect 20168 8032 20220 8084
rect 20996 8032 21048 8084
rect 10324 7871 10376 7880
rect 10324 7837 10333 7871
rect 10333 7837 10367 7871
rect 10367 7837 10376 7871
rect 10324 7828 10376 7837
rect 11980 7828 12032 7880
rect 1952 7692 2004 7744
rect 2412 7692 2464 7744
rect 4068 7692 4120 7744
rect 5908 7692 5960 7744
rect 6368 7692 6420 7744
rect 7380 7692 7432 7744
rect 8208 7735 8260 7744
rect 8208 7701 8217 7735
rect 8217 7701 8251 7735
rect 8251 7701 8260 7735
rect 8208 7692 8260 7701
rect 10416 7760 10468 7812
rect 11060 7760 11112 7812
rect 9864 7692 9916 7744
rect 10968 7692 11020 7744
rect 14004 7896 14056 7948
rect 12164 7828 12216 7880
rect 12440 7828 12492 7880
rect 13728 7828 13780 7880
rect 12716 7760 12768 7812
rect 15200 7896 15252 7948
rect 16396 7896 16448 7948
rect 16672 7896 16724 7948
rect 17684 7896 17736 7948
rect 17776 7896 17828 7948
rect 19064 7939 19116 7948
rect 15568 7828 15620 7880
rect 16764 7828 16816 7880
rect 19064 7905 19073 7939
rect 19073 7905 19107 7939
rect 19107 7905 19116 7939
rect 19064 7896 19116 7905
rect 19708 7896 19760 7948
rect 19340 7828 19392 7880
rect 19800 7828 19852 7880
rect 19892 7828 19944 7880
rect 15660 7760 15712 7812
rect 12992 7692 13044 7744
rect 13544 7692 13596 7744
rect 13728 7735 13780 7744
rect 13728 7701 13737 7735
rect 13737 7701 13771 7735
rect 13771 7701 13780 7735
rect 13728 7692 13780 7701
rect 14004 7692 14056 7744
rect 16948 7760 17000 7812
rect 18236 7760 18288 7812
rect 18512 7760 18564 7812
rect 18788 7760 18840 7812
rect 16304 7692 16356 7744
rect 16580 7692 16632 7744
rect 17684 7692 17736 7744
rect 19432 7692 19484 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 4160 7531 4212 7540
rect 4160 7497 4169 7531
rect 4169 7497 4203 7531
rect 4203 7497 4212 7531
rect 4160 7488 4212 7497
rect 4252 7488 4304 7540
rect 1952 7395 2004 7404
rect 1952 7361 1961 7395
rect 1961 7361 1995 7395
rect 1995 7361 2004 7395
rect 1952 7352 2004 7361
rect 2136 7395 2188 7404
rect 2136 7361 2145 7395
rect 2145 7361 2179 7395
rect 2179 7361 2188 7395
rect 2136 7352 2188 7361
rect 4896 7352 4948 7404
rect 5264 7352 5316 7404
rect 10048 7488 10100 7540
rect 10968 7488 11020 7540
rect 12440 7531 12492 7540
rect 12440 7497 12449 7531
rect 12449 7497 12483 7531
rect 12483 7497 12492 7531
rect 12440 7488 12492 7497
rect 13360 7488 13412 7540
rect 8760 7463 8812 7472
rect 8760 7429 8769 7463
rect 8769 7429 8803 7463
rect 8803 7429 8812 7463
rect 8760 7420 8812 7429
rect 9496 7463 9548 7472
rect 9496 7429 9505 7463
rect 9505 7429 9539 7463
rect 9539 7429 9548 7463
rect 9496 7420 9548 7429
rect 7288 7352 7340 7404
rect 9404 7395 9456 7404
rect 2412 7284 2464 7336
rect 1584 7216 1636 7268
rect 3700 7284 3752 7336
rect 7380 7327 7432 7336
rect 7380 7293 7389 7327
rect 7389 7293 7423 7327
rect 7423 7293 7432 7327
rect 7380 7284 7432 7293
rect 9404 7361 9413 7395
rect 9413 7361 9447 7395
rect 9447 7361 9456 7395
rect 11244 7420 11296 7472
rect 9404 7352 9456 7361
rect 10324 7352 10376 7404
rect 2872 7216 2924 7268
rect 4712 7216 4764 7268
rect 6276 7216 6328 7268
rect 7472 7216 7524 7268
rect 1492 7191 1544 7200
rect 1492 7157 1501 7191
rect 1501 7157 1535 7191
rect 1535 7157 1544 7191
rect 1492 7148 1544 7157
rect 4252 7148 4304 7200
rect 5356 7148 5408 7200
rect 5724 7191 5776 7200
rect 5724 7157 5733 7191
rect 5733 7157 5767 7191
rect 5767 7157 5776 7191
rect 5724 7148 5776 7157
rect 10692 7352 10744 7404
rect 10784 7352 10836 7404
rect 13176 7420 13228 7472
rect 12348 7352 12400 7404
rect 13268 7352 13320 7404
rect 13544 7488 13596 7540
rect 14372 7531 14424 7540
rect 14372 7497 14381 7531
rect 14381 7497 14415 7531
rect 14415 7497 14424 7531
rect 14372 7488 14424 7497
rect 14464 7488 14516 7540
rect 17408 7488 17460 7540
rect 20536 7488 20588 7540
rect 13636 7420 13688 7472
rect 15752 7420 15804 7472
rect 10508 7284 10560 7336
rect 11980 7284 12032 7336
rect 13176 7284 13228 7336
rect 14556 7352 14608 7404
rect 15936 7352 15988 7404
rect 16304 7352 16356 7404
rect 11244 7216 11296 7268
rect 9956 7148 10008 7200
rect 10508 7191 10560 7200
rect 10508 7157 10517 7191
rect 10517 7157 10551 7191
rect 10551 7157 10560 7191
rect 10508 7148 10560 7157
rect 10968 7148 11020 7200
rect 11796 7148 11848 7200
rect 12532 7148 12584 7200
rect 14096 7284 14148 7336
rect 15292 7284 15344 7336
rect 13912 7216 13964 7268
rect 14096 7148 14148 7200
rect 14556 7148 14608 7200
rect 15476 7216 15528 7268
rect 18972 7420 19024 7472
rect 17592 7395 17644 7404
rect 17592 7361 17601 7395
rect 17601 7361 17635 7395
rect 17635 7361 17644 7395
rect 17592 7352 17644 7361
rect 18696 7352 18748 7404
rect 16856 7284 16908 7336
rect 17776 7284 17828 7336
rect 18512 7284 18564 7336
rect 19248 7284 19300 7336
rect 19432 7284 19484 7336
rect 15016 7148 15068 7200
rect 15384 7191 15436 7200
rect 15384 7157 15393 7191
rect 15393 7157 15427 7191
rect 15427 7157 15436 7191
rect 15384 7148 15436 7157
rect 19064 7216 19116 7268
rect 16304 7148 16356 7200
rect 16764 7191 16816 7200
rect 16764 7157 16773 7191
rect 16773 7157 16807 7191
rect 16807 7157 16816 7191
rect 16764 7148 16816 7157
rect 16948 7191 17000 7200
rect 16948 7157 16957 7191
rect 16957 7157 16991 7191
rect 16991 7157 17000 7191
rect 16948 7148 17000 7157
rect 17960 7148 18012 7200
rect 18328 7148 18380 7200
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 4896 6987 4948 6996
rect 4896 6953 4905 6987
rect 4905 6953 4939 6987
rect 4939 6953 4948 6987
rect 4896 6944 4948 6953
rect 5908 6987 5960 6996
rect 5908 6953 5917 6987
rect 5917 6953 5951 6987
rect 5951 6953 5960 6987
rect 5908 6944 5960 6953
rect 6092 6944 6144 6996
rect 9404 6944 9456 6996
rect 2412 6919 2464 6928
rect 2412 6885 2421 6919
rect 2421 6885 2455 6919
rect 2455 6885 2464 6919
rect 2412 6876 2464 6885
rect 3976 6876 4028 6928
rect 11704 6944 11756 6996
rect 12348 6944 12400 6996
rect 12532 6944 12584 6996
rect 10876 6876 10928 6928
rect 7288 6851 7340 6860
rect 7288 6817 7297 6851
rect 7297 6817 7331 6851
rect 7331 6817 7340 6851
rect 7288 6808 7340 6817
rect 8300 6851 8352 6860
rect 8300 6817 8309 6851
rect 8309 6817 8343 6851
rect 8343 6817 8352 6851
rect 8300 6808 8352 6817
rect 8392 6851 8444 6860
rect 8392 6817 8401 6851
rect 8401 6817 8435 6851
rect 8435 6817 8444 6851
rect 8392 6808 8444 6817
rect 8668 6808 8720 6860
rect 10048 6851 10100 6860
rect 2872 6740 2924 6792
rect 3148 6740 3200 6792
rect 4620 6740 4672 6792
rect 3516 6672 3568 6724
rect 4896 6672 4948 6724
rect 5264 6740 5316 6792
rect 6092 6740 6144 6792
rect 6552 6740 6604 6792
rect 7656 6740 7708 6792
rect 8760 6740 8812 6792
rect 9772 6740 9824 6792
rect 10048 6817 10057 6851
rect 10057 6817 10091 6851
rect 10091 6817 10100 6851
rect 10048 6808 10100 6817
rect 10324 6808 10376 6860
rect 12440 6876 12492 6928
rect 13360 6919 13412 6928
rect 13360 6885 13369 6919
rect 13369 6885 13403 6919
rect 13403 6885 13412 6919
rect 13360 6876 13412 6885
rect 13728 6876 13780 6928
rect 13268 6808 13320 6860
rect 14372 6944 14424 6996
rect 17592 6944 17644 6996
rect 19432 6944 19484 6996
rect 15384 6876 15436 6928
rect 15844 6876 15896 6928
rect 19984 6876 20036 6928
rect 14372 6808 14424 6860
rect 15200 6808 15252 6860
rect 9864 6672 9916 6724
rect 5080 6604 5132 6656
rect 6092 6604 6144 6656
rect 6184 6604 6236 6656
rect 6736 6604 6788 6656
rect 8300 6604 8352 6656
rect 8760 6604 8812 6656
rect 9312 6604 9364 6656
rect 13084 6740 13136 6792
rect 13820 6740 13872 6792
rect 14832 6783 14884 6792
rect 14832 6749 14841 6783
rect 14841 6749 14875 6783
rect 14875 6749 14884 6783
rect 14832 6740 14884 6749
rect 16488 6808 16540 6860
rect 18512 6851 18564 6860
rect 18512 6817 18521 6851
rect 18521 6817 18555 6851
rect 18555 6817 18564 6851
rect 18512 6808 18564 6817
rect 16580 6783 16632 6792
rect 12716 6715 12768 6724
rect 12716 6681 12725 6715
rect 12725 6681 12759 6715
rect 12759 6681 12768 6715
rect 12716 6672 12768 6681
rect 12256 6604 12308 6656
rect 13268 6604 13320 6656
rect 14924 6604 14976 6656
rect 15384 6647 15436 6656
rect 15384 6613 15393 6647
rect 15393 6613 15427 6647
rect 15427 6613 15436 6647
rect 15384 6604 15436 6613
rect 16580 6749 16589 6783
rect 16589 6749 16623 6783
rect 16623 6749 16632 6783
rect 16580 6740 16632 6749
rect 18972 6740 19024 6792
rect 19248 6808 19300 6860
rect 20352 6808 20404 6860
rect 17592 6672 17644 6724
rect 18880 6672 18932 6724
rect 20444 6672 20496 6724
rect 21272 6672 21324 6724
rect 16856 6604 16908 6656
rect 19156 6604 19208 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 2872 6443 2924 6452
rect 2872 6409 2881 6443
rect 2881 6409 2915 6443
rect 2915 6409 2924 6443
rect 2872 6400 2924 6409
rect 3516 6443 3568 6452
rect 3516 6409 3525 6443
rect 3525 6409 3559 6443
rect 3559 6409 3568 6443
rect 3516 6400 3568 6409
rect 6184 6400 6236 6452
rect 4620 6332 4672 6384
rect 3148 6264 3200 6316
rect 5080 6307 5132 6316
rect 5080 6273 5089 6307
rect 5089 6273 5123 6307
rect 5123 6273 5132 6307
rect 5080 6264 5132 6273
rect 6092 6307 6144 6316
rect 6092 6273 6101 6307
rect 6101 6273 6135 6307
rect 6135 6273 6144 6307
rect 6092 6264 6144 6273
rect 6184 6307 6236 6316
rect 6184 6273 6193 6307
rect 6193 6273 6227 6307
rect 6227 6273 6236 6307
rect 6184 6264 6236 6273
rect 7104 6264 7156 6316
rect 7656 6264 7708 6316
rect 9404 6400 9456 6452
rect 12624 6400 12676 6452
rect 13084 6400 13136 6452
rect 13452 6400 13504 6452
rect 15200 6400 15252 6452
rect 15384 6400 15436 6452
rect 11796 6332 11848 6384
rect 14004 6332 14056 6384
rect 14648 6332 14700 6384
rect 16488 6400 16540 6452
rect 16856 6443 16908 6452
rect 16856 6409 16865 6443
rect 16865 6409 16899 6443
rect 16899 6409 16908 6443
rect 16856 6400 16908 6409
rect 17224 6400 17276 6452
rect 19156 6400 19208 6452
rect 20352 6443 20404 6452
rect 20352 6409 20361 6443
rect 20361 6409 20395 6443
rect 20395 6409 20404 6443
rect 20352 6400 20404 6409
rect 10140 6264 10192 6316
rect 11704 6264 11756 6316
rect 1584 6196 1636 6248
rect 5724 6196 5776 6248
rect 6644 6196 6696 6248
rect 8668 6196 8720 6248
rect 9128 6196 9180 6248
rect 11980 6264 12032 6316
rect 2320 6128 2372 6180
rect 6644 6060 6696 6112
rect 7288 6103 7340 6112
rect 7288 6069 7297 6103
rect 7297 6069 7331 6103
rect 7331 6069 7340 6103
rect 7288 6060 7340 6069
rect 10876 6128 10928 6180
rect 12440 6239 12492 6248
rect 12440 6205 12449 6239
rect 12449 6205 12483 6239
rect 12483 6205 12492 6239
rect 12440 6196 12492 6205
rect 12348 6128 12400 6180
rect 14280 6264 14332 6316
rect 15200 6307 15252 6316
rect 12716 6239 12768 6248
rect 12716 6205 12750 6239
rect 12750 6205 12768 6239
rect 12716 6196 12768 6205
rect 12992 6196 13044 6248
rect 13636 6128 13688 6180
rect 14280 6128 14332 6180
rect 14832 6128 14884 6180
rect 15200 6273 15209 6307
rect 15209 6273 15243 6307
rect 15243 6273 15252 6307
rect 15200 6264 15252 6273
rect 16488 6264 16540 6316
rect 16580 6196 16632 6248
rect 16672 6196 16724 6248
rect 17592 6196 17644 6248
rect 18972 6239 19024 6248
rect 18972 6205 18981 6239
rect 18981 6205 19015 6239
rect 19015 6205 19024 6239
rect 18972 6196 19024 6205
rect 21088 6264 21140 6316
rect 9404 6060 9456 6112
rect 9772 6060 9824 6112
rect 10968 6060 11020 6112
rect 13084 6060 13136 6112
rect 13820 6103 13872 6112
rect 13820 6069 13829 6103
rect 13829 6069 13863 6103
rect 13863 6069 13872 6103
rect 13820 6060 13872 6069
rect 14556 6103 14608 6112
rect 14556 6069 14565 6103
rect 14565 6069 14599 6103
rect 14599 6069 14608 6103
rect 14556 6060 14608 6069
rect 15200 6060 15252 6112
rect 16488 6128 16540 6180
rect 19340 6128 19392 6180
rect 16672 6060 16724 6112
rect 20996 6060 21048 6112
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 2320 5856 2372 5908
rect 3148 5899 3200 5908
rect 3148 5865 3157 5899
rect 3157 5865 3191 5899
rect 3191 5865 3200 5899
rect 3148 5856 3200 5865
rect 3700 5856 3752 5908
rect 4620 5856 4672 5908
rect 6184 5856 6236 5908
rect 6644 5899 6696 5908
rect 6644 5865 6653 5899
rect 6653 5865 6687 5899
rect 6687 5865 6696 5899
rect 6644 5856 6696 5865
rect 6736 5899 6788 5908
rect 6736 5865 6745 5899
rect 6745 5865 6779 5899
rect 6779 5865 6788 5899
rect 6736 5856 6788 5865
rect 7288 5856 7340 5908
rect 9312 5856 9364 5908
rect 11520 5856 11572 5908
rect 14464 5856 14516 5908
rect 16488 5856 16540 5908
rect 20720 5856 20772 5908
rect 2688 5788 2740 5840
rect 4068 5788 4120 5840
rect 7196 5788 7248 5840
rect 1584 5720 1636 5772
rect 4896 5720 4948 5772
rect 5816 5720 5868 5772
rect 7012 5720 7064 5772
rect 7380 5788 7432 5840
rect 8484 5788 8536 5840
rect 10692 5788 10744 5840
rect 13820 5788 13872 5840
rect 9772 5720 9824 5772
rect 12440 5720 12492 5772
rect 15200 5788 15252 5840
rect 17960 5788 18012 5840
rect 14464 5720 14516 5772
rect 15016 5720 15068 5772
rect 15384 5720 15436 5772
rect 16948 5720 17000 5772
rect 18052 5720 18104 5772
rect 18880 5720 18932 5772
rect 19892 5763 19944 5772
rect 19892 5729 19901 5763
rect 19901 5729 19935 5763
rect 19935 5729 19944 5763
rect 19892 5720 19944 5729
rect 2780 5652 2832 5704
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 6828 5695 6880 5704
rect 6828 5661 6837 5695
rect 6837 5661 6871 5695
rect 6871 5661 6880 5695
rect 6828 5652 6880 5661
rect 8484 5652 8536 5704
rect 9128 5652 9180 5704
rect 10784 5652 10836 5704
rect 11796 5652 11848 5704
rect 3424 5516 3476 5568
rect 6092 5516 6144 5568
rect 9404 5584 9456 5636
rect 10968 5584 11020 5636
rect 17316 5652 17368 5704
rect 19340 5652 19392 5704
rect 13820 5584 13872 5636
rect 20352 5652 20404 5704
rect 8208 5516 8260 5568
rect 8944 5516 8996 5568
rect 10784 5516 10836 5568
rect 10876 5516 10928 5568
rect 11980 5516 12032 5568
rect 13544 5516 13596 5568
rect 13728 5559 13780 5568
rect 13728 5525 13737 5559
rect 13737 5525 13771 5559
rect 13771 5525 13780 5559
rect 13728 5516 13780 5525
rect 14096 5516 14148 5568
rect 18788 5516 18840 5568
rect 19156 5516 19208 5568
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 2412 5312 2464 5364
rect 4068 5312 4120 5364
rect 12348 5312 12400 5364
rect 13360 5312 13412 5364
rect 14280 5355 14332 5364
rect 14280 5321 14289 5355
rect 14289 5321 14323 5355
rect 14323 5321 14332 5355
rect 14280 5312 14332 5321
rect 14556 5312 14608 5364
rect 17960 5312 18012 5364
rect 19340 5312 19392 5364
rect 20260 5312 20312 5364
rect 2320 5176 2372 5228
rect 3700 5219 3752 5228
rect 2688 5108 2740 5160
rect 3700 5185 3709 5219
rect 3709 5185 3743 5219
rect 3743 5185 3752 5219
rect 3700 5176 3752 5185
rect 7472 5219 7524 5228
rect 7472 5185 7481 5219
rect 7481 5185 7515 5219
rect 7515 5185 7524 5219
rect 7472 5176 7524 5185
rect 7656 5176 7708 5228
rect 8944 5176 8996 5228
rect 11796 5244 11848 5296
rect 14096 5244 14148 5296
rect 14188 5244 14240 5296
rect 18880 5244 18932 5296
rect 9680 5176 9732 5228
rect 9772 5176 9824 5228
rect 10876 5176 10928 5228
rect 11060 5176 11112 5228
rect 11980 5176 12032 5228
rect 12716 5176 12768 5228
rect 13636 5219 13688 5228
rect 13636 5185 13645 5219
rect 13645 5185 13679 5219
rect 13679 5185 13688 5219
rect 13636 5176 13688 5185
rect 15200 5176 15252 5228
rect 15844 5219 15896 5228
rect 15844 5185 15853 5219
rect 15853 5185 15887 5219
rect 15887 5185 15896 5219
rect 15844 5176 15896 5185
rect 17316 5176 17368 5228
rect 4160 5108 4212 5160
rect 5448 5108 5500 5160
rect 8208 5108 8260 5160
rect 9312 5108 9364 5160
rect 9404 5108 9456 5160
rect 10968 5151 11020 5160
rect 5816 5040 5868 5092
rect 7012 5040 7064 5092
rect 2412 5015 2464 5024
rect 2412 4981 2421 5015
rect 2421 4981 2455 5015
rect 2455 4981 2464 5015
rect 2412 4972 2464 4981
rect 3240 4972 3292 5024
rect 3516 5015 3568 5024
rect 3516 4981 3525 5015
rect 3525 4981 3559 5015
rect 3559 4981 3568 5015
rect 5724 5015 5776 5024
rect 3516 4972 3568 4981
rect 5724 4981 5733 5015
rect 5733 4981 5767 5015
rect 5767 4981 5776 5015
rect 5724 4972 5776 4981
rect 7196 5015 7248 5024
rect 7196 4981 7205 5015
rect 7205 4981 7239 5015
rect 7239 4981 7248 5015
rect 7196 4972 7248 4981
rect 7288 5015 7340 5024
rect 7288 4981 7297 5015
rect 7297 4981 7331 5015
rect 7331 4981 7340 5015
rect 7288 4972 7340 4981
rect 8392 4972 8444 5024
rect 10140 5040 10192 5092
rect 9128 4972 9180 5024
rect 9680 4972 9732 5024
rect 10968 5117 10977 5151
rect 10977 5117 11011 5151
rect 11011 5117 11020 5151
rect 10968 5108 11020 5117
rect 12440 5108 12492 5160
rect 14004 5108 14056 5160
rect 13636 5040 13688 5092
rect 12808 5015 12860 5024
rect 12808 4981 12817 5015
rect 12817 4981 12851 5015
rect 12851 4981 12860 5015
rect 12808 4972 12860 4981
rect 15476 5108 15528 5160
rect 15568 5108 15620 5160
rect 16120 5108 16172 5160
rect 16580 5108 16632 5160
rect 14188 5040 14240 5092
rect 15292 5040 15344 5092
rect 17960 5040 18012 5092
rect 18696 5108 18748 5160
rect 14280 4972 14332 5024
rect 15200 4972 15252 5024
rect 16856 4972 16908 5024
rect 17408 5015 17460 5024
rect 17408 4981 17417 5015
rect 17417 4981 17451 5015
rect 17451 4981 17460 5015
rect 17408 4972 17460 4981
rect 17592 4972 17644 5024
rect 18972 5040 19024 5092
rect 19432 5108 19484 5160
rect 19800 4972 19852 5024
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 2412 4768 2464 4820
rect 5448 4768 5500 4820
rect 7472 4768 7524 4820
rect 8392 4811 8444 4820
rect 8392 4777 8401 4811
rect 8401 4777 8435 4811
rect 8435 4777 8444 4811
rect 8392 4768 8444 4777
rect 9404 4768 9456 4820
rect 9680 4811 9732 4820
rect 9680 4777 9689 4811
rect 9689 4777 9723 4811
rect 9723 4777 9732 4811
rect 9680 4768 9732 4777
rect 10508 4768 10560 4820
rect 13820 4768 13872 4820
rect 14188 4811 14240 4820
rect 14188 4777 14197 4811
rect 14197 4777 14231 4811
rect 14231 4777 14240 4811
rect 14188 4768 14240 4777
rect 15844 4768 15896 4820
rect 17316 4768 17368 4820
rect 19432 4768 19484 4820
rect 19892 4768 19944 4820
rect 5816 4700 5868 4752
rect 2780 4632 2832 4684
rect 2964 4632 3016 4684
rect 6828 4700 6880 4752
rect 8300 4743 8352 4752
rect 2320 4564 2372 4616
rect 2688 4607 2740 4616
rect 2688 4573 2697 4607
rect 2697 4573 2731 4607
rect 2731 4573 2740 4607
rect 2688 4564 2740 4573
rect 2872 4607 2924 4616
rect 2872 4573 2881 4607
rect 2881 4573 2915 4607
rect 2915 4573 2924 4607
rect 2872 4564 2924 4573
rect 3608 4607 3660 4616
rect 3608 4573 3617 4607
rect 3617 4573 3651 4607
rect 3651 4573 3660 4607
rect 3608 4564 3660 4573
rect 4252 4564 4304 4616
rect 5724 4607 5776 4616
rect 5724 4573 5733 4607
rect 5733 4573 5767 4607
rect 5767 4573 5776 4607
rect 5724 4564 5776 4573
rect 2412 4496 2464 4548
rect 5080 4471 5132 4480
rect 5080 4437 5089 4471
rect 5089 4437 5123 4471
rect 5123 4437 5132 4471
rect 5080 4428 5132 4437
rect 6920 4632 6972 4684
rect 8300 4709 8309 4743
rect 8309 4709 8343 4743
rect 8343 4709 8352 4743
rect 8300 4700 8352 4709
rect 10324 4700 10376 4752
rect 11060 4700 11112 4752
rect 11704 4700 11756 4752
rect 11152 4632 11204 4684
rect 12440 4632 12492 4684
rect 13912 4700 13964 4752
rect 11704 4607 11756 4616
rect 9588 4496 9640 4548
rect 11704 4573 11713 4607
rect 11713 4573 11747 4607
rect 11747 4573 11756 4607
rect 11704 4564 11756 4573
rect 11980 4564 12032 4616
rect 12348 4564 12400 4616
rect 13268 4675 13320 4684
rect 13268 4641 13277 4675
rect 13277 4641 13311 4675
rect 13311 4641 13320 4675
rect 13268 4632 13320 4641
rect 14280 4632 14332 4684
rect 15936 4700 15988 4752
rect 16488 4700 16540 4752
rect 16948 4700 17000 4752
rect 15384 4632 15436 4684
rect 18696 4700 18748 4752
rect 10968 4496 11020 4548
rect 12992 4496 13044 4548
rect 13820 4496 13872 4548
rect 14556 4496 14608 4548
rect 19064 4496 19116 4548
rect 19340 4496 19392 4548
rect 20076 4607 20128 4616
rect 20076 4573 20085 4607
rect 20085 4573 20119 4607
rect 20119 4573 20128 4607
rect 20076 4564 20128 4573
rect 20260 4700 20312 4752
rect 20260 4564 20312 4616
rect 19984 4496 20036 4548
rect 7932 4471 7984 4480
rect 7932 4437 7941 4471
rect 7941 4437 7975 4471
rect 7975 4437 7984 4471
rect 7932 4428 7984 4437
rect 8300 4428 8352 4480
rect 8852 4428 8904 4480
rect 9128 4428 9180 4480
rect 11980 4428 12032 4480
rect 12900 4428 12952 4480
rect 15108 4428 15160 4480
rect 20444 4428 20496 4480
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 3516 4224 3568 4276
rect 4160 4156 4212 4208
rect 4344 4156 4396 4208
rect 3424 4088 3476 4140
rect 7288 4224 7340 4276
rect 10140 4267 10192 4276
rect 10140 4233 10149 4267
rect 10149 4233 10183 4267
rect 10183 4233 10192 4267
rect 10140 4224 10192 4233
rect 10968 4224 11020 4276
rect 13912 4224 13964 4276
rect 14004 4224 14056 4276
rect 16212 4224 16264 4276
rect 17960 4224 18012 4276
rect 19432 4224 19484 4276
rect 19616 4224 19668 4276
rect 19984 4224 20036 4276
rect 4896 4088 4948 4140
rect 5724 4156 5776 4208
rect 6920 4156 6972 4208
rect 11888 4156 11940 4208
rect 13820 4199 13872 4208
rect 13820 4165 13829 4199
rect 13829 4165 13863 4199
rect 13863 4165 13872 4199
rect 13820 4156 13872 4165
rect 2688 4020 2740 4072
rect 4712 4020 4764 4072
rect 2504 3952 2556 4004
rect 3148 3952 3200 4004
rect 3884 3952 3936 4004
rect 4160 3952 4212 4004
rect 4988 3952 5040 4004
rect 6092 4063 6144 4072
rect 6092 4029 6101 4063
rect 6101 4029 6135 4063
rect 6135 4029 6144 4063
rect 6092 4020 6144 4029
rect 10508 4088 10560 4140
rect 11704 4131 11756 4140
rect 6644 4020 6696 4072
rect 7932 4020 7984 4072
rect 8484 4063 8536 4072
rect 8484 4029 8493 4063
rect 8493 4029 8527 4063
rect 8527 4029 8536 4063
rect 8484 4020 8536 4029
rect 10140 4020 10192 4072
rect 11704 4097 11713 4131
rect 11713 4097 11747 4131
rect 11747 4097 11756 4131
rect 11704 4088 11756 4097
rect 11796 4088 11848 4140
rect 14464 4088 14516 4140
rect 5264 3995 5316 4004
rect 5264 3961 5273 3995
rect 5273 3961 5307 3995
rect 5307 3961 5316 3995
rect 5264 3952 5316 3961
rect 2412 3884 2464 3936
rect 2872 3884 2924 3936
rect 3516 3884 3568 3936
rect 3976 3884 4028 3936
rect 7196 3952 7248 4004
rect 7656 3952 7708 4004
rect 10048 3952 10100 4004
rect 10232 3952 10284 4004
rect 13820 4020 13872 4072
rect 14280 4020 14332 4072
rect 16488 4156 16540 4208
rect 15844 4131 15896 4140
rect 15844 4097 15853 4131
rect 15853 4097 15887 4131
rect 15887 4097 15896 4131
rect 15844 4088 15896 4097
rect 17776 4088 17828 4140
rect 17960 4088 18012 4140
rect 18696 4156 18748 4208
rect 16580 4020 16632 4072
rect 16672 4020 16724 4072
rect 20536 4088 20588 4140
rect 20260 4063 20312 4072
rect 20260 4029 20269 4063
rect 20269 4029 20303 4063
rect 20303 4029 20312 4063
rect 20260 4020 20312 4029
rect 6920 3884 6972 3936
rect 7380 3927 7432 3936
rect 7380 3893 7389 3927
rect 7389 3893 7423 3927
rect 7423 3893 7432 3927
rect 7380 3884 7432 3893
rect 8944 3884 8996 3936
rect 9312 3884 9364 3936
rect 10600 3884 10652 3936
rect 11244 3884 11296 3936
rect 12440 3884 12492 3936
rect 12624 3884 12676 3936
rect 19616 3952 19668 4004
rect 13728 3884 13780 3936
rect 14096 3927 14148 3936
rect 14096 3893 14105 3927
rect 14105 3893 14139 3927
rect 14139 3893 14148 3927
rect 14096 3884 14148 3893
rect 14280 3884 14332 3936
rect 15384 3884 15436 3936
rect 16580 3884 16632 3936
rect 17592 3927 17644 3936
rect 17592 3893 17601 3927
rect 17601 3893 17635 3927
rect 17635 3893 17644 3927
rect 17592 3884 17644 3893
rect 17776 3884 17828 3936
rect 18788 3884 18840 3936
rect 19892 3884 19944 3936
rect 20260 3884 20312 3936
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 2412 3680 2464 3732
rect 2964 3723 3016 3732
rect 2964 3689 2973 3723
rect 2973 3689 3007 3723
rect 3007 3689 3016 3723
rect 2964 3680 3016 3689
rect 3424 3723 3476 3732
rect 3424 3689 3433 3723
rect 3433 3689 3467 3723
rect 3467 3689 3476 3723
rect 3424 3680 3476 3689
rect 3608 3680 3660 3732
rect 5080 3680 5132 3732
rect 7012 3680 7064 3732
rect 7380 3723 7432 3732
rect 7380 3689 7389 3723
rect 7389 3689 7423 3723
rect 7423 3689 7432 3723
rect 7380 3680 7432 3689
rect 11520 3723 11572 3732
rect 4344 3612 4396 3664
rect 4896 3612 4948 3664
rect 9772 3612 9824 3664
rect 3056 3544 3108 3596
rect 2504 3476 2556 3528
rect 4712 3544 4764 3596
rect 5080 3544 5132 3596
rect 5540 3544 5592 3596
rect 5816 3544 5868 3596
rect 6828 3544 6880 3596
rect 3516 3519 3568 3528
rect 3516 3485 3525 3519
rect 3525 3485 3559 3519
rect 3559 3485 3568 3519
rect 8760 3544 8812 3596
rect 3516 3476 3568 3485
rect 8208 3476 8260 3528
rect 8392 3476 8444 3528
rect 9404 3544 9456 3596
rect 10232 3544 10284 3596
rect 11520 3689 11529 3723
rect 11529 3689 11563 3723
rect 11563 3689 11572 3723
rect 11520 3680 11572 3689
rect 11888 3723 11940 3732
rect 11888 3689 11897 3723
rect 11897 3689 11931 3723
rect 11931 3689 11940 3723
rect 11888 3680 11940 3689
rect 14004 3723 14056 3732
rect 11060 3655 11112 3664
rect 11060 3621 11069 3655
rect 11069 3621 11103 3655
rect 11103 3621 11112 3655
rect 11060 3612 11112 3621
rect 12900 3655 12952 3664
rect 12900 3621 12909 3655
rect 12909 3621 12943 3655
rect 12943 3621 12952 3655
rect 12900 3612 12952 3621
rect 14004 3689 14013 3723
rect 14013 3689 14047 3723
rect 14047 3689 14056 3723
rect 14004 3680 14056 3689
rect 15200 3680 15252 3732
rect 15384 3723 15436 3732
rect 15384 3689 15393 3723
rect 15393 3689 15427 3723
rect 15427 3689 15436 3723
rect 15384 3680 15436 3689
rect 15752 3680 15804 3732
rect 16120 3680 16172 3732
rect 17316 3723 17368 3732
rect 17316 3689 17325 3723
rect 17325 3689 17359 3723
rect 17359 3689 17368 3723
rect 17316 3680 17368 3689
rect 17408 3680 17460 3732
rect 19064 3680 19116 3732
rect 20076 3680 20128 3732
rect 14096 3612 14148 3664
rect 15108 3612 15160 3664
rect 17500 3612 17552 3664
rect 17960 3612 18012 3664
rect 11888 3544 11940 3596
rect 12992 3587 13044 3596
rect 12992 3553 13001 3587
rect 13001 3553 13035 3587
rect 13035 3553 13044 3587
rect 12992 3544 13044 3553
rect 13544 3544 13596 3596
rect 14556 3587 14608 3596
rect 14556 3553 14565 3587
rect 14565 3553 14599 3587
rect 14599 3553 14608 3587
rect 14556 3544 14608 3553
rect 15384 3544 15436 3596
rect 9312 3476 9364 3528
rect 5724 3340 5776 3392
rect 6644 3340 6696 3392
rect 10324 3519 10376 3528
rect 10324 3485 10333 3519
rect 10333 3485 10367 3519
rect 10367 3485 10376 3519
rect 10508 3519 10560 3528
rect 10324 3476 10376 3485
rect 10508 3485 10517 3519
rect 10517 3485 10551 3519
rect 10551 3485 10560 3519
rect 10508 3476 10560 3485
rect 11796 3476 11848 3528
rect 13728 3476 13780 3528
rect 14096 3519 14148 3528
rect 14096 3485 14105 3519
rect 14105 3485 14139 3519
rect 14139 3485 14148 3519
rect 14096 3476 14148 3485
rect 16488 3476 16540 3528
rect 17040 3544 17092 3596
rect 18512 3612 18564 3664
rect 19340 3612 19392 3664
rect 20812 3612 20864 3664
rect 19616 3544 19668 3596
rect 17316 3476 17368 3528
rect 17500 3519 17552 3528
rect 17500 3485 17509 3519
rect 17509 3485 17543 3519
rect 17543 3485 17552 3519
rect 17500 3476 17552 3485
rect 17960 3476 18012 3528
rect 18696 3476 18748 3528
rect 19340 3476 19392 3528
rect 19708 3476 19760 3528
rect 19800 3476 19852 3528
rect 20536 3476 20588 3528
rect 10600 3408 10652 3460
rect 11612 3408 11664 3460
rect 12532 3451 12584 3460
rect 12532 3417 12541 3451
rect 12541 3417 12575 3451
rect 12575 3417 12584 3451
rect 12532 3408 12584 3417
rect 14280 3408 14332 3460
rect 14832 3408 14884 3460
rect 10324 3340 10376 3392
rect 14004 3340 14056 3392
rect 17408 3340 17460 3392
rect 17592 3408 17644 3460
rect 19340 3340 19392 3392
rect 19432 3340 19484 3392
rect 19708 3340 19760 3392
rect 20444 3408 20496 3460
rect 21640 3408 21692 3460
rect 21180 3340 21232 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 2044 3136 2096 3188
rect 2688 3136 2740 3188
rect 2596 3000 2648 3052
rect 1492 2932 1544 2984
rect 3332 3136 3384 3188
rect 4252 3136 4304 3188
rect 4620 3068 4672 3120
rect 6092 3136 6144 3188
rect 7472 3136 7524 3188
rect 7564 3136 7616 3188
rect 8208 3179 8260 3188
rect 8208 3145 8217 3179
rect 8217 3145 8251 3179
rect 8251 3145 8260 3179
rect 8208 3136 8260 3145
rect 8760 3136 8812 3188
rect 10140 3179 10192 3188
rect 10140 3145 10149 3179
rect 10149 3145 10183 3179
rect 10183 3145 10192 3179
rect 10140 3136 10192 3145
rect 10692 3136 10744 3188
rect 11796 3179 11848 3188
rect 11796 3145 11805 3179
rect 11805 3145 11839 3179
rect 11839 3145 11848 3179
rect 11796 3136 11848 3145
rect 12440 3179 12492 3188
rect 12440 3145 12449 3179
rect 12449 3145 12483 3179
rect 12483 3145 12492 3179
rect 12440 3136 12492 3145
rect 13176 3136 13228 3188
rect 11888 3068 11940 3120
rect 13820 3068 13872 3120
rect 14648 3136 14700 3188
rect 15476 3179 15528 3188
rect 15476 3145 15485 3179
rect 15485 3145 15519 3179
rect 15519 3145 15528 3179
rect 15476 3136 15528 3145
rect 20628 3136 20680 3188
rect 5816 3000 5868 3052
rect 11612 3000 11664 3052
rect 12164 3000 12216 3052
rect 12992 3043 13044 3052
rect 12992 3009 13001 3043
rect 13001 3009 13035 3043
rect 13035 3009 13044 3043
rect 12992 3000 13044 3009
rect 14096 3000 14148 3052
rect 1032 2864 1084 2916
rect 2228 2864 2280 2916
rect 3148 2796 3200 2848
rect 3516 2864 3568 2916
rect 4160 2864 4212 2916
rect 5540 2864 5592 2916
rect 6000 2864 6052 2916
rect 8392 2932 8444 2984
rect 8484 2932 8536 2984
rect 11704 2932 11756 2984
rect 12900 2975 12952 2984
rect 12900 2941 12909 2975
rect 12909 2941 12943 2975
rect 12943 2941 12952 2975
rect 12900 2932 12952 2941
rect 7104 2907 7156 2916
rect 7104 2873 7138 2907
rect 7138 2873 7156 2907
rect 7104 2864 7156 2873
rect 7472 2864 7524 2916
rect 8668 2864 8720 2916
rect 9036 2907 9088 2916
rect 9036 2873 9070 2907
rect 9070 2873 9088 2907
rect 9036 2864 9088 2873
rect 10232 2864 10284 2916
rect 6276 2796 6328 2848
rect 8484 2796 8536 2848
rect 9404 2796 9456 2848
rect 14740 2932 14792 2984
rect 19524 3068 19576 3120
rect 15108 3043 15160 3052
rect 15108 3009 15117 3043
rect 15117 3009 15151 3043
rect 15151 3009 15160 3043
rect 15108 3000 15160 3009
rect 15292 3000 15344 3052
rect 16120 3043 16172 3052
rect 16120 3009 16129 3043
rect 16129 3009 16163 3043
rect 16163 3009 16172 3043
rect 16120 3000 16172 3009
rect 17500 3043 17552 3052
rect 17500 3009 17509 3043
rect 17509 3009 17543 3043
rect 17543 3009 17552 3043
rect 17500 3000 17552 3009
rect 17592 3000 17644 3052
rect 19340 3000 19392 3052
rect 19892 3043 19944 3052
rect 18328 2932 18380 2984
rect 19248 2932 19300 2984
rect 19892 3009 19901 3043
rect 19901 3009 19935 3043
rect 19935 3009 19944 3043
rect 19892 3000 19944 3009
rect 20536 3068 20588 3120
rect 19800 2975 19852 2984
rect 19800 2941 19809 2975
rect 19809 2941 19843 2975
rect 19843 2941 19852 2975
rect 19800 2932 19852 2941
rect 20260 2932 20312 2984
rect 14372 2864 14424 2916
rect 15016 2864 15068 2916
rect 15292 2864 15344 2916
rect 13544 2796 13596 2848
rect 13820 2839 13872 2848
rect 13820 2805 13829 2839
rect 13829 2805 13863 2839
rect 13863 2805 13872 2839
rect 13820 2796 13872 2805
rect 13912 2839 13964 2848
rect 13912 2805 13921 2839
rect 13921 2805 13955 2839
rect 13955 2805 13964 2839
rect 16764 2864 16816 2916
rect 17868 2864 17920 2916
rect 13912 2796 13964 2805
rect 16304 2796 16356 2848
rect 18512 2864 18564 2916
rect 22100 2796 22152 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 2228 2635 2280 2644
rect 2228 2601 2237 2635
rect 2237 2601 2271 2635
rect 2271 2601 2280 2635
rect 2228 2592 2280 2601
rect 2780 2635 2832 2644
rect 2780 2601 2789 2635
rect 2789 2601 2823 2635
rect 2823 2601 2832 2635
rect 2780 2592 2832 2601
rect 4712 2592 4764 2644
rect 1952 2524 2004 2576
rect 3148 2524 3200 2576
rect 3424 2567 3476 2576
rect 3424 2533 3433 2567
rect 3433 2533 3467 2567
rect 3467 2533 3476 2567
rect 3424 2524 3476 2533
rect 5172 2592 5224 2644
rect 6092 2592 6144 2644
rect 6920 2635 6972 2644
rect 6920 2601 6929 2635
rect 6929 2601 6963 2635
rect 6963 2601 6972 2635
rect 6920 2592 6972 2601
rect 10232 2635 10284 2644
rect 8300 2567 8352 2576
rect 8300 2533 8309 2567
rect 8309 2533 8343 2567
rect 8343 2533 8352 2567
rect 10232 2601 10241 2635
rect 10241 2601 10275 2635
rect 10275 2601 10284 2635
rect 10232 2592 10284 2601
rect 10692 2592 10744 2644
rect 10968 2592 11020 2644
rect 12348 2592 12400 2644
rect 12808 2592 12860 2644
rect 13452 2592 13504 2644
rect 13636 2592 13688 2644
rect 13912 2592 13964 2644
rect 8300 2524 8352 2533
rect 8760 2456 8812 2508
rect 10508 2524 10560 2576
rect 11796 2524 11848 2576
rect 3516 2431 3568 2440
rect 3516 2397 3525 2431
rect 3525 2397 3559 2431
rect 3559 2397 3568 2431
rect 3516 2388 3568 2397
rect 5724 2388 5776 2440
rect 6276 2431 6328 2440
rect 6276 2397 6285 2431
rect 6285 2397 6319 2431
rect 6319 2397 6328 2431
rect 6276 2388 6328 2397
rect 7104 2388 7156 2440
rect 7564 2431 7616 2440
rect 7564 2397 7573 2431
rect 7573 2397 7607 2431
rect 7607 2397 7616 2431
rect 7564 2388 7616 2397
rect 8392 2431 8444 2440
rect 8392 2397 8401 2431
rect 8401 2397 8435 2431
rect 8435 2397 8444 2431
rect 8392 2388 8444 2397
rect 10232 2456 10284 2508
rect 12992 2524 13044 2576
rect 15200 2592 15252 2644
rect 15660 2592 15712 2644
rect 15936 2635 15988 2644
rect 15936 2601 15945 2635
rect 15945 2601 15979 2635
rect 15979 2601 15988 2635
rect 15936 2592 15988 2601
rect 16028 2592 16080 2644
rect 16948 2635 17000 2644
rect 16948 2601 16957 2635
rect 16957 2601 16991 2635
rect 16991 2601 17000 2635
rect 16948 2592 17000 2601
rect 19064 2635 19116 2644
rect 19064 2601 19073 2635
rect 19073 2601 19107 2635
rect 19107 2601 19116 2635
rect 19064 2592 19116 2601
rect 19524 2635 19576 2644
rect 19524 2601 19533 2635
rect 19533 2601 19567 2635
rect 19567 2601 19576 2635
rect 19524 2592 19576 2601
rect 20444 2635 20496 2644
rect 15752 2524 15804 2576
rect 20444 2601 20453 2635
rect 20453 2601 20487 2635
rect 20487 2601 20496 2635
rect 20444 2592 20496 2601
rect 20536 2524 20588 2576
rect 3056 2320 3108 2372
rect 3148 2320 3200 2372
rect 10140 2388 10192 2440
rect 12256 2456 12308 2508
rect 13820 2456 13872 2508
rect 15108 2456 15160 2508
rect 17224 2456 17276 2508
rect 17316 2456 17368 2508
rect 17776 2456 17828 2508
rect 13360 2431 13412 2440
rect 1768 2295 1820 2304
rect 1768 2261 1777 2295
rect 1777 2261 1811 2295
rect 1811 2261 1820 2295
rect 1768 2252 1820 2261
rect 2964 2295 3016 2304
rect 2964 2261 2973 2295
rect 2973 2261 3007 2295
rect 3007 2261 3016 2295
rect 2964 2252 3016 2261
rect 9312 2320 9364 2372
rect 13360 2397 13369 2431
rect 13369 2397 13403 2431
rect 13403 2397 13412 2431
rect 13360 2388 13412 2397
rect 13912 2388 13964 2440
rect 15016 2388 15068 2440
rect 16120 2388 16172 2440
rect 16396 2320 16448 2372
rect 19340 2388 19392 2440
rect 20352 2388 20404 2440
rect 12624 2252 12676 2304
rect 14188 2252 14240 2304
rect 14924 2252 14976 2304
rect 20260 2320 20312 2372
rect 22560 2252 22612 2304
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 2872 2048 2924 2100
rect 3424 2048 3476 2100
rect 6276 2048 6328 2100
rect 20168 2048 20220 2100
rect 1768 1980 1820 2032
rect 15108 1980 15160 2032
rect 16856 1980 16908 2032
rect 18972 1980 19024 2032
rect 2964 1912 3016 1964
rect 15292 1912 15344 1964
rect 8760 1844 8812 1896
rect 15200 1844 15252 1896
rect 3056 1776 3108 1828
rect 3516 1776 3568 1828
rect 8392 1776 8444 1828
rect 10600 1776 10652 1828
rect 12072 1708 12124 1760
rect 1492 1640 1544 1692
rect 8852 1640 8904 1692
rect 10508 1640 10560 1692
rect 16672 1640 16724 1692
rect 2412 1572 2464 1624
rect 8300 1572 8352 1624
rect 3240 1300 3292 1352
rect 4988 1300 5040 1352
rect 16764 1300 16816 1352
rect 17960 1300 18012 1352
rect 572 1232 624 1284
rect 7656 1232 7708 1284
rect 13084 1096 13136 1148
rect 15384 1096 15436 1148
rect 19800 552 19852 604
rect 20996 552 21048 604
<< metal2 >>
rect 202 22320 258 22800
rect 662 22320 718 22800
rect 1122 22320 1178 22800
rect 1582 22320 1638 22800
rect 2042 22320 2098 22800
rect 2502 22320 2558 22800
rect 3054 22320 3110 22800
rect 3238 22536 3294 22545
rect 3238 22471 3294 22480
rect 216 16726 244 22320
rect 676 18766 704 22320
rect 1136 19242 1164 22320
rect 1124 19236 1176 19242
rect 1124 19178 1176 19184
rect 1596 19122 1624 22320
rect 1860 19916 1912 19922
rect 1860 19858 1912 19864
rect 1766 19680 1822 19689
rect 1766 19615 1822 19624
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 1504 19094 1624 19122
rect 664 18760 716 18766
rect 664 18702 716 18708
rect 1504 18154 1532 19094
rect 1582 19000 1638 19009
rect 1582 18935 1638 18944
rect 1596 18834 1624 18935
rect 1584 18828 1636 18834
rect 1584 18770 1636 18776
rect 1688 18465 1716 19246
rect 1780 18970 1808 19615
rect 1768 18964 1820 18970
rect 1768 18906 1820 18912
rect 1872 18902 1900 19858
rect 1860 18896 1912 18902
rect 1860 18838 1912 18844
rect 2056 18698 2084 22320
rect 2136 19916 2188 19922
rect 2136 19858 2188 19864
rect 2044 18692 2096 18698
rect 2044 18634 2096 18640
rect 1674 18456 1730 18465
rect 1674 18391 1730 18400
rect 1674 18320 1730 18329
rect 1674 18255 1730 18264
rect 1492 18148 1544 18154
rect 1492 18090 1544 18096
rect 1688 17882 1716 18255
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1582 17776 1638 17785
rect 1582 17711 1638 17720
rect 1400 17128 1452 17134
rect 1400 17070 1452 17076
rect 204 16720 256 16726
rect 204 16662 256 16668
rect 1412 16658 1440 17070
rect 1490 16824 1546 16833
rect 1596 16794 1624 17711
rect 1674 17368 1730 17377
rect 1674 17303 1730 17312
rect 1490 16759 1546 16768
rect 1584 16788 1636 16794
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1504 15706 1532 16759
rect 1584 16730 1636 16736
rect 1688 16250 1716 17303
rect 1676 16244 1728 16250
rect 1676 16186 1728 16192
rect 1676 16040 1728 16046
rect 1676 15982 1728 15988
rect 1492 15700 1544 15706
rect 1492 15642 1544 15648
rect 1584 15564 1636 15570
rect 1584 15506 1636 15512
rect 1492 14952 1544 14958
rect 1492 14894 1544 14900
rect 1504 14618 1532 14894
rect 1492 14612 1544 14618
rect 1492 14554 1544 14560
rect 1492 14476 1544 14482
rect 1492 14418 1544 14424
rect 1504 12986 1532 14418
rect 1492 12980 1544 12986
rect 1492 12922 1544 12928
rect 1596 12424 1624 15506
rect 1688 15026 1716 15982
rect 1780 15609 1808 18158
rect 2148 18034 2176 19858
rect 2516 18970 2544 22320
rect 3068 22234 3096 22320
rect 3056 22228 3108 22234
rect 3056 22170 3108 22176
rect 3054 22128 3110 22137
rect 3054 22063 3110 22072
rect 2962 21584 3018 21593
rect 2962 21519 3018 21528
rect 2870 21176 2926 21185
rect 2870 21111 2926 21120
rect 2778 20632 2834 20641
rect 2778 20567 2834 20576
rect 2792 19786 2820 20567
rect 2884 20058 2912 21111
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 2780 19780 2832 19786
rect 2780 19722 2832 19728
rect 2688 19304 2740 19310
rect 2872 19304 2924 19310
rect 2688 19246 2740 19252
rect 2778 19272 2834 19281
rect 2504 18964 2556 18970
rect 2504 18906 2556 18912
rect 2228 18828 2280 18834
rect 2228 18770 2280 18776
rect 2056 18006 2176 18034
rect 1952 17876 2004 17882
rect 1952 17818 2004 17824
rect 1964 17202 1992 17818
rect 1952 17196 2004 17202
rect 1952 17138 2004 17144
rect 1766 15600 1822 15609
rect 2056 15570 2084 18006
rect 2134 17368 2190 17377
rect 2134 17303 2190 17312
rect 2148 17202 2176 17303
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 2240 15586 2268 18770
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 2332 17814 2360 18158
rect 2320 17808 2372 17814
rect 2320 17750 2372 17756
rect 2318 17640 2374 17649
rect 2318 17575 2374 17584
rect 2332 16794 2360 17575
rect 2504 17128 2556 17134
rect 2504 17070 2556 17076
rect 2320 16788 2372 16794
rect 2320 16730 2372 16736
rect 2412 16788 2464 16794
rect 2412 16730 2464 16736
rect 2424 16590 2452 16730
rect 2412 16584 2464 16590
rect 2412 16526 2464 16532
rect 2516 16250 2544 17070
rect 2504 16244 2556 16250
rect 2504 16186 2556 16192
rect 2502 16008 2558 16017
rect 2502 15943 2504 15952
rect 2556 15943 2558 15952
rect 2504 15914 2556 15920
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 2596 15904 2648 15910
rect 2596 15846 2648 15852
rect 1766 15535 1822 15544
rect 2044 15564 2096 15570
rect 2240 15558 2360 15586
rect 2044 15506 2096 15512
rect 1676 15020 1728 15026
rect 1676 14962 1728 14968
rect 2044 14816 2096 14822
rect 2044 14758 2096 14764
rect 1768 14408 1820 14414
rect 1768 14350 1820 14356
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1504 12396 1624 12424
rect 1504 10606 1532 12396
rect 1688 10810 1716 12582
rect 1780 11218 1808 14350
rect 1860 13728 1912 13734
rect 1860 13670 1912 13676
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 1492 10600 1544 10606
rect 1492 10542 1544 10548
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1780 10266 1808 10406
rect 1872 10266 1900 13670
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1492 8424 1544 8430
rect 1596 8412 1624 8910
rect 1544 8384 1624 8412
rect 1492 8366 1544 8372
rect 1596 7274 1624 8384
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1584 7268 1636 7274
rect 1584 7210 1636 7216
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 570 3360 626 3369
rect 216 3318 570 3346
rect 216 480 244 3318
rect 570 3295 626 3304
rect 1504 2990 1532 7142
rect 1596 6254 1624 7210
rect 1584 6248 1636 6254
rect 1584 6190 1636 6196
rect 1596 5778 1624 6190
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 1688 5658 1716 7890
rect 1964 7834 1992 13330
rect 2056 9586 2084 14758
rect 2228 14272 2280 14278
rect 2228 14214 2280 14220
rect 2136 13796 2188 13802
rect 2136 13738 2188 13744
rect 2148 13394 2176 13738
rect 2136 13388 2188 13394
rect 2136 13330 2188 13336
rect 2148 12374 2176 13330
rect 2136 12368 2188 12374
rect 2136 12310 2188 12316
rect 2148 11626 2176 12310
rect 2136 11620 2188 11626
rect 2136 11562 2188 11568
rect 2148 11218 2176 11562
rect 2136 11212 2188 11218
rect 2136 11154 2188 11160
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 2148 9722 2176 10406
rect 2136 9716 2188 9722
rect 2136 9658 2188 9664
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 2240 9518 2268 14214
rect 2332 12442 2360 15558
rect 2424 15337 2452 15846
rect 2608 15706 2636 15846
rect 2596 15700 2648 15706
rect 2596 15642 2648 15648
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 2410 15328 2466 15337
rect 2410 15263 2466 15272
rect 2412 13864 2464 13870
rect 2412 13806 2464 13812
rect 2516 13818 2544 15438
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2608 14278 2636 14758
rect 2700 14657 2728 19246
rect 2872 19246 2924 19252
rect 2778 19207 2834 19216
rect 2792 18426 2820 19207
rect 2884 18873 2912 19246
rect 2976 19174 3004 21519
rect 3068 19310 3096 22063
rect 3146 20224 3202 20233
rect 3146 20159 3202 20168
rect 3160 19514 3188 20159
rect 3148 19508 3200 19514
rect 3148 19450 3200 19456
rect 3056 19304 3108 19310
rect 3056 19246 3108 19252
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 2870 18864 2926 18873
rect 2870 18799 2926 18808
rect 3056 18692 3108 18698
rect 3056 18634 3108 18640
rect 3068 18426 3096 18634
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 3056 18216 3108 18222
rect 3054 18184 3056 18193
rect 3108 18184 3110 18193
rect 3054 18119 3110 18128
rect 3252 18086 3280 22471
rect 3514 22320 3570 22800
rect 3974 22320 4030 22800
rect 4434 22320 4490 22800
rect 4894 22320 4950 22800
rect 5354 22320 5410 22800
rect 5906 22320 5962 22800
rect 6366 22320 6422 22800
rect 6826 22320 6882 22800
rect 7286 22320 7342 22800
rect 7746 22320 7802 22800
rect 8206 22320 8262 22800
rect 8758 22320 8814 22800
rect 9218 22320 9274 22800
rect 9678 22320 9734 22800
rect 10138 22320 10194 22800
rect 10598 22320 10654 22800
rect 11058 22320 11114 22800
rect 11610 22320 11666 22800
rect 12070 22320 12126 22800
rect 12530 22320 12586 22800
rect 12990 22320 13046 22800
rect 13450 22320 13506 22800
rect 13910 22320 13966 22800
rect 14462 22320 14518 22800
rect 14922 22320 14978 22800
rect 15382 22320 15438 22800
rect 15842 22320 15898 22800
rect 16302 22320 16358 22800
rect 16762 22320 16818 22800
rect 17314 22320 17370 22800
rect 17774 22320 17830 22800
rect 18234 22320 18290 22800
rect 18694 22320 18750 22800
rect 19062 22536 19118 22545
rect 19062 22471 19118 22480
rect 3332 20256 3384 20262
rect 3332 20198 3384 20204
rect 3344 20058 3372 20198
rect 3332 20052 3384 20058
rect 3332 19994 3384 20000
rect 3332 19916 3384 19922
rect 3332 19858 3384 19864
rect 3344 19514 3372 19858
rect 3332 19508 3384 19514
rect 3332 19450 3384 19456
rect 3528 19394 3556 22320
rect 3700 22228 3752 22234
rect 3700 22170 3752 22176
rect 3608 20324 3660 20330
rect 3608 20266 3660 20272
rect 3620 20058 3648 20266
rect 3608 20052 3660 20058
rect 3608 19994 3660 20000
rect 3344 19366 3556 19394
rect 3344 18816 3372 19366
rect 3516 19304 3568 19310
rect 3516 19246 3568 19252
rect 3424 18828 3476 18834
rect 3344 18788 3424 18816
rect 3240 18080 3292 18086
rect 3240 18022 3292 18028
rect 3344 17898 3372 18788
rect 3424 18770 3476 18776
rect 3528 18766 3556 19246
rect 3516 18760 3568 18766
rect 3516 18702 3568 18708
rect 3606 18728 3662 18737
rect 3424 18692 3476 18698
rect 3424 18634 3476 18640
rect 3436 18426 3464 18634
rect 3424 18420 3476 18426
rect 3424 18362 3476 18368
rect 3528 18272 3556 18702
rect 3606 18663 3608 18672
rect 3660 18663 3662 18672
rect 3608 18634 3660 18640
rect 3712 18426 3740 22170
rect 3988 19281 4016 22320
rect 4448 19802 4476 22320
rect 4264 19774 4476 19802
rect 3974 19272 4030 19281
rect 3974 19207 4030 19216
rect 3884 19168 3936 19174
rect 3790 19136 3846 19145
rect 3884 19110 3936 19116
rect 3976 19168 4028 19174
rect 3976 19110 4028 19116
rect 3790 19071 3846 19080
rect 3700 18420 3752 18426
rect 3700 18362 3752 18368
rect 3608 18284 3660 18290
rect 3252 17882 3372 17898
rect 3240 17876 3372 17882
rect 3292 17870 3372 17876
rect 3436 18244 3608 18272
rect 3240 17818 3292 17824
rect 3056 17740 3108 17746
rect 3056 17682 3108 17688
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 2792 17241 2820 17614
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 2778 17232 2834 17241
rect 2778 17167 2834 17176
rect 2884 17082 2912 17478
rect 2792 17054 2912 17082
rect 2962 17096 3018 17105
rect 2792 16794 2820 17054
rect 2962 17031 2964 17040
rect 3016 17031 3018 17040
rect 2964 17002 3016 17008
rect 2872 16992 2924 16998
rect 2872 16934 2924 16940
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 2792 15502 2820 16050
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 2884 14958 2912 16934
rect 2964 15020 3016 15026
rect 2964 14962 3016 14968
rect 2872 14952 2924 14958
rect 2872 14894 2924 14900
rect 2686 14648 2742 14657
rect 2686 14583 2742 14592
rect 2778 14512 2834 14521
rect 2778 14447 2834 14456
rect 2596 14272 2648 14278
rect 2596 14214 2648 14220
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2320 12300 2372 12306
rect 2320 12242 2372 12248
rect 2332 11558 2360 12242
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2332 10674 2360 11494
rect 2424 11286 2452 13806
rect 2516 13790 2728 13818
rect 2504 13728 2556 13734
rect 2504 13670 2556 13676
rect 2516 12442 2544 13670
rect 2504 12436 2556 12442
rect 2504 12378 2556 12384
rect 2596 12368 2648 12374
rect 2596 12310 2648 12316
rect 2504 12300 2556 12306
rect 2504 12242 2556 12248
rect 2412 11280 2464 11286
rect 2412 11222 2464 11228
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2320 10532 2372 10538
rect 2320 10474 2372 10480
rect 2228 9512 2280 9518
rect 2228 9454 2280 9460
rect 2136 8356 2188 8362
rect 2136 8298 2188 8304
rect 1964 7806 2084 7834
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 1964 7410 1992 7686
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1688 5630 1900 5658
rect 1492 2984 1544 2990
rect 1492 2926 1544 2932
rect 1032 2916 1084 2922
rect 1032 2858 1084 2864
rect 572 1284 624 1290
rect 572 1226 624 1232
rect 584 480 612 1226
rect 1044 480 1072 2858
rect 1872 2553 1900 5630
rect 2056 3194 2084 7806
rect 2148 7410 2176 8298
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 2332 7154 2360 10474
rect 2424 7954 2452 11222
rect 2412 7948 2464 7954
rect 2412 7890 2464 7896
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2424 7342 2452 7686
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2240 7126 2360 7154
rect 2240 4604 2268 7126
rect 2412 6928 2464 6934
rect 2412 6870 2464 6876
rect 2320 6180 2372 6186
rect 2320 6122 2372 6128
rect 2332 5914 2360 6122
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2332 5234 2360 5850
rect 2424 5370 2452 6870
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2412 5024 2464 5030
rect 2412 4966 2464 4972
rect 2424 4826 2452 4966
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2516 4706 2544 12242
rect 2608 11014 2636 12310
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 2608 10538 2636 10950
rect 2596 10532 2648 10538
rect 2596 10474 2648 10480
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2608 8566 2636 8978
rect 2596 8560 2648 8566
rect 2596 8502 2648 8508
rect 2424 4678 2544 4706
rect 2320 4616 2372 4622
rect 2240 4576 2320 4604
rect 2320 4558 2372 4564
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 2332 3097 2360 4558
rect 2424 4554 2452 4678
rect 2412 4548 2464 4554
rect 2412 4490 2464 4496
rect 2504 4004 2556 4010
rect 2504 3946 2556 3952
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 2424 3738 2452 3878
rect 2412 3732 2464 3738
rect 2412 3674 2464 3680
rect 2516 3534 2544 3946
rect 2504 3528 2556 3534
rect 2504 3470 2556 3476
rect 2318 3088 2374 3097
rect 2608 3058 2636 8502
rect 2700 7449 2728 13790
rect 2792 11354 2820 14447
rect 2976 14414 3004 14962
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 2976 14090 3004 14350
rect 2884 14074 3004 14090
rect 2872 14068 3004 14074
rect 2924 14062 3004 14068
rect 2872 14010 2924 14016
rect 2872 13388 2924 13394
rect 2872 13330 2924 13336
rect 2884 12850 2912 13330
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 2884 12442 2912 12786
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 2976 11898 3004 12582
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 3068 11642 3096 17682
rect 3436 17377 3464 18244
rect 3608 18226 3660 18232
rect 3804 18154 3832 19071
rect 3896 18290 3924 19110
rect 3884 18284 3936 18290
rect 3884 18226 3936 18232
rect 3792 18148 3844 18154
rect 3792 18090 3844 18096
rect 3516 17740 3568 17746
rect 3516 17682 3568 17688
rect 3422 17368 3478 17377
rect 3528 17338 3556 17682
rect 3608 17672 3660 17678
rect 3988 17649 4016 19110
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 4080 18222 4108 18906
rect 4264 18737 4292 19774
rect 4712 19712 4764 19718
rect 4712 19654 4764 19660
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 4724 19310 4752 19654
rect 4712 19304 4764 19310
rect 4764 19264 4844 19292
rect 4712 19246 4764 19252
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 4724 18970 4752 19110
rect 4712 18964 4764 18970
rect 4712 18906 4764 18912
rect 4344 18828 4396 18834
rect 4344 18770 4396 18776
rect 4250 18728 4306 18737
rect 4356 18698 4384 18770
rect 4250 18663 4306 18672
rect 4344 18692 4396 18698
rect 4344 18634 4396 18640
rect 4160 18624 4212 18630
rect 4212 18584 4292 18612
rect 4160 18566 4212 18572
rect 4068 18216 4120 18222
rect 4068 18158 4120 18164
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 4172 17814 4200 18022
rect 4264 17882 4292 18584
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4712 18284 4764 18290
rect 4632 18244 4712 18272
rect 4526 18184 4582 18193
rect 4526 18119 4528 18128
rect 4580 18119 4582 18128
rect 4528 18090 4580 18096
rect 4252 17876 4304 17882
rect 4252 17818 4304 17824
rect 4160 17808 4212 17814
rect 4160 17750 4212 17756
rect 4632 17678 4660 18244
rect 4712 18226 4764 18232
rect 4712 18148 4764 18154
rect 4712 18090 4764 18096
rect 4160 17672 4212 17678
rect 3608 17614 3660 17620
rect 3974 17640 4030 17649
rect 3620 17338 3648 17614
rect 4160 17614 4212 17620
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 3974 17575 4030 17584
rect 3422 17303 3478 17312
rect 3516 17332 3568 17338
rect 3148 17060 3200 17066
rect 3148 17002 3200 17008
rect 3160 16046 3188 17002
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 3344 16522 3372 16934
rect 3332 16516 3384 16522
rect 3436 16504 3464 17303
rect 3516 17274 3568 17280
rect 3608 17332 3660 17338
rect 3608 17274 3660 17280
rect 3620 16590 3648 17274
rect 4172 17270 4200 17614
rect 4724 17610 4752 18090
rect 4816 17746 4844 19264
rect 4908 19258 4936 22320
rect 5172 19916 5224 19922
rect 5172 19858 5224 19864
rect 4986 19272 5042 19281
rect 4908 19230 4986 19258
rect 4986 19207 5042 19216
rect 5184 18426 5212 19858
rect 5368 19802 5396 22320
rect 5724 20052 5776 20058
rect 5724 19994 5776 20000
rect 5368 19774 5488 19802
rect 5356 19712 5408 19718
rect 5356 19654 5408 19660
rect 5368 19310 5396 19654
rect 5356 19304 5408 19310
rect 5356 19246 5408 19252
rect 5264 18828 5316 18834
rect 5264 18770 5316 18776
rect 4988 18420 5040 18426
rect 4988 18362 5040 18368
rect 5172 18420 5224 18426
rect 5172 18362 5224 18368
rect 4896 18080 4948 18086
rect 4896 18022 4948 18028
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 4712 17604 4764 17610
rect 4712 17546 4764 17552
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 4160 17264 4212 17270
rect 4212 17224 4384 17252
rect 4160 17206 4212 17212
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 3608 16584 3660 16590
rect 3608 16526 3660 16532
rect 3436 16476 3556 16504
rect 3332 16458 3384 16464
rect 3422 16416 3478 16425
rect 3422 16351 3478 16360
rect 3330 16144 3386 16153
rect 3330 16079 3386 16088
rect 3148 16040 3200 16046
rect 3148 15982 3200 15988
rect 3160 15094 3188 15982
rect 3344 15706 3372 16079
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 3436 15162 3464 16351
rect 3528 15978 3556 16476
rect 3516 15972 3568 15978
rect 3516 15914 3568 15920
rect 3528 15502 3556 15914
rect 3700 15904 3752 15910
rect 3700 15846 3752 15852
rect 3974 15872 4030 15881
rect 3712 15638 3740 15846
rect 3974 15807 4030 15816
rect 3700 15632 3752 15638
rect 3700 15574 3752 15580
rect 3516 15496 3568 15502
rect 3516 15438 3568 15444
rect 3988 15434 4016 15807
rect 4172 15706 4200 16594
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4264 15638 4292 16730
rect 4356 16590 4384 17224
rect 4908 16998 4936 18022
rect 5000 17882 5028 18362
rect 4988 17876 5040 17882
rect 4988 17818 5040 17824
rect 5080 17672 5132 17678
rect 5080 17614 5132 17620
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4712 16720 4764 16726
rect 4712 16662 4764 16668
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4724 16250 4752 16662
rect 4712 16244 4764 16250
rect 4712 16186 4764 16192
rect 5092 15706 5120 17614
rect 5184 17066 5212 17614
rect 5276 17542 5304 18770
rect 5368 18766 5396 19246
rect 5356 18760 5408 18766
rect 5356 18702 5408 18708
rect 5356 18624 5408 18630
rect 5356 18566 5408 18572
rect 5264 17536 5316 17542
rect 5264 17478 5316 17484
rect 5276 17270 5304 17478
rect 5264 17264 5316 17270
rect 5264 17206 5316 17212
rect 5172 17060 5224 17066
rect 5172 17002 5224 17008
rect 5264 16584 5316 16590
rect 5264 16526 5316 16532
rect 5276 16114 5304 16526
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5368 15994 5396 18566
rect 5460 18442 5488 19774
rect 5630 19000 5686 19009
rect 5630 18935 5686 18944
rect 5644 18601 5672 18935
rect 5630 18592 5686 18601
rect 5630 18527 5686 18536
rect 5460 18414 5672 18442
rect 5540 18284 5592 18290
rect 5540 18226 5592 18232
rect 5552 17746 5580 18226
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 5460 16794 5488 17478
rect 5552 17338 5580 17682
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 5644 16561 5672 18414
rect 5736 16810 5764 19994
rect 5736 16782 5856 16810
rect 5630 16552 5686 16561
rect 5540 16516 5592 16522
rect 5630 16487 5686 16496
rect 5540 16458 5592 16464
rect 5276 15966 5396 15994
rect 5552 15978 5580 16458
rect 5540 15972 5592 15978
rect 5080 15700 5132 15706
rect 5080 15642 5132 15648
rect 4252 15632 4304 15638
rect 4252 15574 4304 15580
rect 4896 15564 4948 15570
rect 4948 15524 5028 15552
rect 4896 15506 4948 15512
rect 4066 15464 4122 15473
rect 3976 15428 4028 15434
rect 4066 15399 4122 15408
rect 3976 15370 4028 15376
rect 4080 15366 4108 15399
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 4250 15328 4306 15337
rect 4250 15263 4306 15272
rect 3424 15156 3476 15162
rect 3424 15098 3476 15104
rect 3976 15156 4028 15162
rect 4264 15144 4292 15263
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4264 15116 4660 15144
rect 3976 15098 4028 15104
rect 3148 15088 3200 15094
rect 3148 15030 3200 15036
rect 3424 14952 3476 14958
rect 3424 14894 3476 14900
rect 3516 14952 3568 14958
rect 3516 14894 3568 14900
rect 3148 14544 3200 14550
rect 3148 14486 3200 14492
rect 3160 12628 3188 14486
rect 3240 14476 3292 14482
rect 3240 14418 3292 14424
rect 3252 13530 3280 14418
rect 3330 13560 3386 13569
rect 3240 13524 3292 13530
rect 3330 13495 3386 13504
rect 3240 13466 3292 13472
rect 3240 12640 3292 12646
rect 3160 12600 3240 12628
rect 3240 12582 3292 12588
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 2976 11614 3096 11642
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2976 10810 3004 11614
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 3068 10266 3096 11494
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 2872 10124 2924 10130
rect 2872 10066 2924 10072
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2792 9586 2820 9862
rect 2884 9722 2912 10066
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 2686 7440 2742 7449
rect 2686 7375 2742 7384
rect 2872 7268 2924 7274
rect 2872 7210 2924 7216
rect 2884 6798 2912 7210
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 2884 6458 2912 6734
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 2688 5840 2740 5846
rect 2688 5782 2740 5788
rect 2700 5166 2728 5782
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2688 5160 2740 5166
rect 2688 5102 2740 5108
rect 2700 4622 2728 5102
rect 2792 4690 2820 5646
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 2688 4616 2740 4622
rect 2688 4558 2740 4564
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2778 4448 2834 4457
rect 2778 4383 2834 4392
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2700 3194 2728 4014
rect 2688 3188 2740 3194
rect 2688 3130 2740 3136
rect 2318 3023 2374 3032
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 2228 2916 2280 2922
rect 2228 2858 2280 2864
rect 2240 2650 2268 2858
rect 2792 2650 2820 4383
rect 2884 3942 2912 4558
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2976 3738 3004 4626
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 3068 3602 3096 8026
rect 3160 6798 3188 12242
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 3160 5914 3188 6258
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3252 5030 3280 12582
rect 3344 12442 3372 13495
rect 3332 12436 3384 12442
rect 3332 12378 3384 12384
rect 3436 10674 3464 14894
rect 3528 14550 3556 14894
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 3516 14544 3568 14550
rect 3516 14486 3568 14492
rect 3516 14340 3568 14346
rect 3516 14282 3568 14288
rect 3528 11898 3556 14282
rect 3792 14068 3844 14074
rect 3792 14010 3844 14016
rect 3606 13832 3662 13841
rect 3606 13767 3608 13776
rect 3660 13767 3662 13776
rect 3608 13738 3660 13744
rect 3620 13258 3648 13738
rect 3700 13728 3752 13734
rect 3700 13670 3752 13676
rect 3608 13252 3660 13258
rect 3608 13194 3660 13200
rect 3712 12850 3740 13670
rect 3700 12844 3752 12850
rect 3700 12786 3752 12792
rect 3700 12232 3752 12238
rect 3700 12174 3752 12180
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3514 11792 3570 11801
rect 3514 11727 3570 11736
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3344 8090 3372 9318
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 3436 5574 3464 10610
rect 3528 10198 3556 11727
rect 3620 11694 3648 12038
rect 3712 11830 3740 12174
rect 3700 11824 3752 11830
rect 3700 11766 3752 11772
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3712 11354 3740 11766
rect 3700 11348 3752 11354
rect 3700 11290 3752 11296
rect 3608 10464 3660 10470
rect 3608 10406 3660 10412
rect 3620 10266 3648 10406
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 3516 10192 3568 10198
rect 3516 10134 3568 10140
rect 3608 10056 3660 10062
rect 3712 10044 3740 11290
rect 3804 11218 3832 14010
rect 3896 11393 3924 14758
rect 3988 14414 4016 15098
rect 4066 14920 4122 14929
rect 4066 14855 4122 14864
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 3988 13870 4016 14350
rect 4080 14074 4108 14855
rect 4632 14822 4660 15116
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 4066 13968 4122 13977
rect 4066 13903 4068 13912
rect 4120 13903 4122 13912
rect 4068 13874 4120 13880
rect 3976 13864 4028 13870
rect 3976 13806 4028 13812
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 4080 12986 4108 13330
rect 4068 12980 4120 12986
rect 4068 12922 4120 12928
rect 3976 12912 4028 12918
rect 3976 12854 4028 12860
rect 3988 12617 4016 12854
rect 3974 12608 4030 12617
rect 3974 12543 4030 12552
rect 4172 12442 4200 14758
rect 4252 14544 4304 14550
rect 4632 14521 4660 14758
rect 4252 14486 4304 14492
rect 4618 14512 4674 14521
rect 4264 13734 4292 14486
rect 4618 14447 4674 14456
rect 4896 14476 4948 14482
rect 4896 14418 4948 14424
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4816 13870 4844 14214
rect 4528 13864 4580 13870
rect 4528 13806 4580 13812
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 4252 13728 4304 13734
rect 4252 13670 4304 13676
rect 4540 13258 4568 13806
rect 4816 13326 4844 13806
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4528 13252 4580 13258
rect 4528 13194 4580 13200
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4250 13016 4306 13025
rect 4388 13008 4684 13028
rect 4250 12951 4252 12960
rect 4304 12951 4306 12960
rect 4252 12922 4304 12928
rect 4816 12850 4844 13262
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 4252 12776 4304 12782
rect 4908 12730 4936 14418
rect 4252 12718 4304 12724
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4264 11762 4292 12718
rect 4540 12702 4936 12730
rect 4540 12170 4568 12702
rect 4710 12608 4766 12617
rect 4710 12543 4766 12552
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 4250 11520 4306 11529
rect 4250 11455 4306 11464
rect 3882 11384 3938 11393
rect 3882 11319 3938 11328
rect 3792 11212 3844 11218
rect 3792 11154 3844 11160
rect 3804 10742 3832 11154
rect 3792 10736 3844 10742
rect 3792 10678 3844 10684
rect 3660 10016 3740 10044
rect 3608 9998 3660 10004
rect 3804 9586 3832 10678
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3896 9761 3924 10066
rect 3988 9926 4016 10406
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 3976 9920 4028 9926
rect 3976 9862 4028 9868
rect 3882 9752 3938 9761
rect 3882 9687 3938 9696
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 4080 9518 4108 9998
rect 4264 9602 4292 11455
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4264 9574 4384 9602
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 3712 8634 3740 9454
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 4080 8809 4108 9318
rect 4356 8974 4384 9574
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 4066 8800 4122 8809
rect 4066 8735 4122 8744
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 3712 8430 3740 8570
rect 3700 8424 3752 8430
rect 3700 8366 3752 8372
rect 3712 7954 3740 8366
rect 3976 8356 4028 8362
rect 3976 8298 4028 8304
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3700 7948 3752 7954
rect 3700 7890 3752 7896
rect 3712 7342 3740 7890
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3516 6724 3568 6730
rect 3516 6666 3568 6672
rect 3528 6458 3556 6666
rect 3516 6452 3568 6458
rect 3516 6394 3568 6400
rect 3700 5908 3752 5914
rect 3700 5850 3752 5856
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3712 5234 3740 5850
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 3056 3596 3108 3602
rect 3056 3538 3108 3544
rect 3068 3505 3096 3538
rect 3054 3496 3110 3505
rect 3054 3431 3110 3440
rect 3160 2854 3188 3946
rect 3148 2848 3200 2854
rect 3148 2790 3200 2796
rect 2228 2644 2280 2650
rect 2228 2586 2280 2592
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 1952 2576 2004 2582
rect 1858 2544 1914 2553
rect 1952 2518 2004 2524
rect 3148 2576 3200 2582
rect 3148 2518 3200 2524
rect 1858 2479 1914 2488
rect 1768 2304 1820 2310
rect 1768 2246 1820 2252
rect 1780 2038 1808 2246
rect 1768 2032 1820 2038
rect 1768 1974 1820 1980
rect 1492 1692 1544 1698
rect 1492 1634 1544 1640
rect 1504 480 1532 1634
rect 1964 480 1992 2518
rect 3160 2378 3188 2518
rect 3056 2372 3108 2378
rect 3056 2314 3108 2320
rect 3148 2372 3200 2378
rect 3148 2314 3200 2320
rect 2964 2304 3016 2310
rect 2964 2246 3016 2252
rect 2872 2100 2924 2106
rect 2872 2042 2924 2048
rect 2412 1624 2464 1630
rect 2412 1566 2464 1572
rect 2424 480 2452 1566
rect 2884 480 2912 2042
rect 2976 1970 3004 2246
rect 2964 1964 3016 1970
rect 2964 1906 3016 1912
rect 3068 1834 3096 2314
rect 3252 2145 3280 4966
rect 3528 4282 3556 4966
rect 3608 4616 3660 4622
rect 3608 4558 3660 4564
rect 3516 4276 3568 4282
rect 3516 4218 3568 4224
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3436 3738 3464 4082
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3528 3534 3556 3878
rect 3620 3738 3648 4558
rect 3896 4010 3924 8230
rect 3988 8022 4016 8298
rect 4066 8256 4122 8265
rect 4066 8191 4122 8200
rect 3976 8016 4028 8022
rect 3976 7958 4028 7964
rect 3974 7848 4030 7857
rect 3974 7783 4030 7792
rect 3988 6934 4016 7783
rect 4080 7750 4108 8191
rect 4160 7812 4212 7818
rect 4160 7754 4212 7760
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 4172 7546 4200 7754
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4264 7426 4292 7482
rect 4724 7460 4752 12543
rect 5000 12322 5028 15524
rect 5172 15088 5224 15094
rect 5092 15048 5172 15076
rect 5092 12442 5120 15048
rect 5172 15030 5224 15036
rect 5172 13456 5224 13462
rect 5172 13398 5224 13404
rect 5184 12714 5212 13398
rect 5276 12889 5304 15966
rect 5540 15914 5592 15920
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5460 15162 5488 15506
rect 5540 15496 5592 15502
rect 5540 15438 5592 15444
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 5448 14884 5500 14890
rect 5448 14826 5500 14832
rect 5356 14612 5408 14618
rect 5356 14554 5408 14560
rect 5262 12880 5318 12889
rect 5262 12815 5318 12824
rect 5172 12708 5224 12714
rect 5172 12650 5224 12656
rect 5262 12608 5318 12617
rect 5262 12543 5318 12552
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 5000 12294 5212 12322
rect 4896 12164 4948 12170
rect 4896 12106 4948 12112
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4080 7398 4292 7426
rect 4448 7432 4752 7460
rect 4080 7313 4108 7398
rect 4448 7324 4476 7432
rect 4066 7304 4122 7313
rect 4066 7239 4122 7248
rect 4172 7296 4476 7324
rect 4618 7304 4674 7313
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 4172 6780 4200 7296
rect 4618 7239 4674 7248
rect 4712 7268 4764 7274
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 3988 6752 4200 6780
rect 3884 4004 3936 4010
rect 3884 3946 3936 3952
rect 3988 3942 4016 6752
rect 4066 5944 4122 5953
rect 4066 5879 4122 5888
rect 4080 5846 4108 5879
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 4068 5704 4120 5710
rect 4120 5664 4200 5692
rect 4068 5646 4120 5652
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4080 5001 4108 5306
rect 4172 5166 4200 5664
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 4264 5012 4292 7142
rect 4632 6798 4660 7239
rect 4816 7256 4844 11834
rect 4908 10606 4936 12106
rect 4988 11824 5040 11830
rect 4988 11766 5040 11772
rect 5000 11150 5028 11766
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5092 11354 5120 11494
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 5184 11257 5212 12294
rect 5170 11248 5226 11257
rect 5170 11183 5226 11192
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 4896 10600 4948 10606
rect 4948 10560 5028 10588
rect 4896 10542 4948 10548
rect 4896 9104 4948 9110
rect 4896 9046 4948 9052
rect 4908 7954 4936 9046
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 4908 7410 4936 7890
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 4764 7228 4844 7256
rect 4712 7210 4764 7216
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4620 6384 4672 6390
rect 4620 6326 4672 6332
rect 4632 5914 4660 6326
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4066 4992 4122 5001
rect 4066 4927 4122 4936
rect 4172 4984 4292 5012
rect 4172 4214 4200 4984
rect 4252 4616 4304 4622
rect 4252 4558 4304 4564
rect 4160 4208 4212 4214
rect 4160 4150 4212 4156
rect 4066 4040 4122 4049
rect 4066 3975 4122 3984
rect 4160 4004 4212 4010
rect 3976 3936 4028 3942
rect 3698 3904 3754 3913
rect 3976 3878 4028 3884
rect 3698 3839 3754 3848
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 3238 2136 3294 2145
rect 3238 2071 3294 2080
rect 3056 1828 3108 1834
rect 3056 1770 3108 1776
rect 3240 1352 3292 1358
rect 3240 1294 3292 1300
rect 3252 649 3280 1294
rect 3238 640 3294 649
rect 3238 575 3294 584
rect 3344 480 3372 3130
rect 3528 2922 3556 3470
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 3424 2576 3476 2582
rect 3424 2518 3476 2524
rect 3436 2106 3464 2518
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 3424 2100 3476 2106
rect 3424 2042 3476 2048
rect 3528 1834 3556 2382
rect 3516 1828 3568 1834
rect 3516 1770 3568 1776
rect 3712 480 3740 3839
rect 202 0 258 480
rect 570 0 626 480
rect 1030 0 1086 480
rect 1490 0 1546 480
rect 1950 0 2006 480
rect 2410 0 2466 480
rect 2870 0 2926 480
rect 3330 0 3386 480
rect 3698 0 3754 480
rect 3988 241 4016 3878
rect 4080 3097 4108 3975
rect 4160 3946 4212 3952
rect 4066 3088 4122 3097
rect 4172 3074 4200 3946
rect 4264 3194 4292 4558
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4344 4208 4396 4214
rect 4344 4150 4396 4156
rect 4356 3670 4384 4150
rect 4724 4078 4752 7210
rect 4894 7032 4950 7041
rect 4894 6967 4896 6976
rect 4948 6967 4950 6976
rect 4896 6938 4948 6944
rect 4896 6724 4948 6730
rect 4896 6666 4948 6672
rect 4908 5778 4936 6666
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 4908 4146 4936 5714
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 5000 4010 5028 10560
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5184 10266 5212 10406
rect 5172 10260 5224 10266
rect 5172 10202 5224 10208
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 5092 9178 5120 10066
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5172 9036 5224 9042
rect 5172 8978 5224 8984
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 5092 7313 5120 8910
rect 5184 8430 5212 8978
rect 5172 8424 5224 8430
rect 5172 8366 5224 8372
rect 5276 7868 5304 12543
rect 5368 11898 5396 14554
rect 5460 12782 5488 14826
rect 5552 14600 5580 15438
rect 5644 15144 5672 16487
rect 5828 16017 5856 16782
rect 5814 16008 5870 16017
rect 5814 15943 5870 15952
rect 5644 15116 5856 15144
rect 5552 14572 5764 14600
rect 5538 14512 5594 14521
rect 5538 14447 5540 14456
rect 5592 14447 5594 14456
rect 5632 14476 5684 14482
rect 5540 14418 5592 14424
rect 5632 14418 5684 14424
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5552 13530 5580 14214
rect 5644 13734 5672 14418
rect 5632 13728 5684 13734
rect 5632 13670 5684 13676
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5644 13274 5672 13670
rect 5736 13433 5764 14572
rect 5828 14521 5856 15116
rect 5814 14512 5870 14521
rect 5814 14447 5870 14456
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5722 13424 5778 13433
rect 5828 13394 5856 13670
rect 5722 13359 5778 13368
rect 5816 13388 5868 13394
rect 5816 13330 5868 13336
rect 5724 13320 5776 13326
rect 5644 13268 5724 13274
rect 5644 13262 5776 13268
rect 5644 13246 5764 13262
rect 5644 12850 5672 13246
rect 5920 13138 5948 22320
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 6196 18426 6224 18702
rect 6380 18442 6408 22320
rect 6460 19304 6512 19310
rect 6460 19246 6512 19252
rect 6472 18766 6500 19246
rect 6736 19236 6788 19242
rect 6736 19178 6788 19184
rect 6748 18834 6776 19178
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 6736 18692 6788 18698
rect 6736 18634 6788 18640
rect 6184 18420 6236 18426
rect 6380 18414 6592 18442
rect 6184 18362 6236 18368
rect 6276 18216 6328 18222
rect 5828 13110 5948 13138
rect 6012 18176 6276 18204
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5448 12776 5500 12782
rect 5446 12744 5448 12753
rect 5500 12744 5502 12753
rect 5446 12679 5502 12688
rect 5448 12300 5500 12306
rect 5448 12242 5500 12248
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5460 11762 5488 12242
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5828 11336 5856 13110
rect 5906 13016 5962 13025
rect 5906 12951 5962 12960
rect 5736 11308 5856 11336
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5356 10736 5408 10742
rect 5356 10678 5408 10684
rect 5368 9994 5396 10678
rect 5644 10674 5672 11154
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5356 9988 5408 9994
rect 5356 9930 5408 9936
rect 5356 9648 5408 9654
rect 5356 9590 5408 9596
rect 5368 9382 5396 9590
rect 5460 9382 5488 10610
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5354 8528 5410 8537
rect 5354 8463 5410 8472
rect 5184 7840 5304 7868
rect 5078 7304 5134 7313
rect 5078 7239 5134 7248
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 5092 6322 5120 6598
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 4988 4004 5040 4010
rect 4988 3946 5040 3952
rect 5092 3738 5120 4422
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 4344 3664 4396 3670
rect 4344 3606 4396 3612
rect 4896 3664 4948 3670
rect 4948 3624 5028 3652
rect 4896 3606 4948 3612
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 4620 3120 4672 3126
rect 4172 3046 4384 3074
rect 4620 3062 4672 3068
rect 4066 3023 4122 3032
rect 4160 2916 4212 2922
rect 4160 2858 4212 2864
rect 4172 480 4200 2858
rect 4356 2292 4384 3046
rect 4264 2264 4384 2292
rect 4632 2292 4660 3062
rect 4724 2650 4752 3538
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4632 2264 4752 2292
rect 4264 1193 4292 2264
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4724 1442 4752 2264
rect 4632 1414 4752 1442
rect 4250 1184 4306 1193
rect 4250 1119 4306 1128
rect 4632 480 4660 1414
rect 5000 1358 5028 3624
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 4988 1352 5040 1358
rect 4988 1294 5040 1300
rect 5092 480 5120 3538
rect 5184 2650 5212 7840
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5276 6798 5304 7346
rect 5368 7206 5396 8463
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5460 5166 5488 9318
rect 5736 9178 5764 11308
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5828 9586 5856 11154
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 5632 9036 5684 9042
rect 5552 8996 5632 9024
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5460 4729 5488 4762
rect 5446 4720 5502 4729
rect 5446 4655 5502 4664
rect 5264 4004 5316 4010
rect 5264 3946 5316 3952
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5276 1601 5304 3946
rect 5552 3602 5580 8996
rect 5632 8978 5684 8984
rect 5736 8786 5764 9114
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 5828 8888 5856 9046
rect 5920 8956 5948 12951
rect 6012 10810 6040 18176
rect 6276 18158 6328 18164
rect 6460 18080 6512 18086
rect 6460 18022 6512 18028
rect 6472 16590 6500 18022
rect 6564 17785 6592 18414
rect 6748 18193 6776 18634
rect 6840 18329 6868 22320
rect 7300 20346 7328 22320
rect 7116 20318 7328 20346
rect 7380 20392 7432 20398
rect 7380 20334 7432 20340
rect 6920 19916 6972 19922
rect 6920 19858 6972 19864
rect 6826 18320 6882 18329
rect 6826 18255 6882 18264
rect 6734 18184 6790 18193
rect 6734 18119 6790 18128
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6550 17776 6606 17785
rect 6550 17711 6606 17720
rect 6644 17536 6696 17542
rect 6644 17478 6696 17484
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 6460 16584 6512 16590
rect 6460 16526 6512 16532
rect 6184 16448 6236 16454
rect 6184 16390 6236 16396
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 6196 16182 6224 16390
rect 6184 16176 6236 16182
rect 6184 16118 6236 16124
rect 6090 16008 6146 16017
rect 6090 15943 6146 15952
rect 6104 15337 6132 15943
rect 6196 15570 6224 16118
rect 6472 16046 6500 16390
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 6368 15360 6420 15366
rect 6090 15328 6146 15337
rect 6368 15302 6420 15308
rect 6090 15263 6146 15272
rect 6104 14890 6132 15263
rect 6380 15162 6408 15302
rect 6368 15156 6420 15162
rect 6368 15098 6420 15104
rect 6564 15094 6592 17138
rect 6184 15088 6236 15094
rect 6184 15030 6236 15036
rect 6552 15088 6604 15094
rect 6552 15030 6604 15036
rect 6092 14884 6144 14890
rect 6092 14826 6144 14832
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 6104 12986 6132 13806
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6196 12646 6224 15030
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6276 13864 6328 13870
rect 6276 13806 6328 13812
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 6092 11076 6144 11082
rect 6092 11018 6144 11024
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 6012 10266 6040 10610
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 6104 10198 6132 11018
rect 6184 10464 6236 10470
rect 6184 10406 6236 10412
rect 6196 10266 6224 10406
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 6092 10192 6144 10198
rect 6092 10134 6144 10140
rect 6184 10056 6236 10062
rect 6090 10024 6146 10033
rect 6184 9998 6236 10004
rect 6090 9959 6146 9968
rect 5920 8928 6040 8956
rect 5828 8860 5948 8888
rect 5736 8758 5856 8786
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5736 8090 5764 8230
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5736 6254 5764 7142
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 5828 5778 5856 8758
rect 5920 8022 5948 8860
rect 6012 8537 6040 8928
rect 5998 8528 6054 8537
rect 5998 8463 6054 8472
rect 6104 8378 6132 9959
rect 6196 9518 6224 9998
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 6196 9382 6224 9454
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6196 9110 6224 9318
rect 6184 9104 6236 9110
rect 6184 9046 6236 9052
rect 6012 8350 6132 8378
rect 5908 8016 5960 8022
rect 5908 7958 5960 7964
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5920 7002 5948 7686
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5816 5092 5868 5098
rect 5816 5034 5868 5040
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5736 4622 5764 4966
rect 5828 4758 5856 5034
rect 5816 4752 5868 4758
rect 5816 4694 5868 4700
rect 5724 4616 5776 4622
rect 5724 4558 5776 4564
rect 5736 4214 5764 4558
rect 5724 4208 5776 4214
rect 5724 4150 5776 4156
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5736 3398 5764 4150
rect 5828 3602 5856 4694
rect 5920 3641 5948 6938
rect 5906 3632 5962 3641
rect 5816 3596 5868 3602
rect 5906 3567 5962 3576
rect 5816 3538 5868 3544
rect 5724 3392 5776 3398
rect 5724 3334 5776 3340
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 5262 1592 5318 1601
rect 5262 1527 5318 1536
rect 5552 480 5580 2858
rect 5736 2446 5764 3334
rect 5828 3058 5856 3538
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 5920 2802 5948 3567
rect 6012 2922 6040 8350
rect 6288 7274 6316 13806
rect 6366 12744 6422 12753
rect 6366 12679 6422 12688
rect 6380 9178 6408 12679
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 6366 9072 6422 9081
rect 6366 9007 6368 9016
rect 6420 9007 6422 9016
rect 6368 8978 6420 8984
rect 6366 8664 6422 8673
rect 6366 8599 6422 8608
rect 6380 7750 6408 8599
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6276 7268 6328 7274
rect 6276 7210 6328 7216
rect 6090 7032 6146 7041
rect 6090 6967 6092 6976
rect 6144 6967 6146 6976
rect 6092 6938 6144 6944
rect 6092 6792 6144 6798
rect 6090 6760 6092 6769
rect 6144 6760 6146 6769
rect 6090 6695 6146 6704
rect 6092 6656 6144 6662
rect 6092 6598 6144 6604
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 6104 6322 6132 6598
rect 6196 6458 6224 6598
rect 6184 6452 6236 6458
rect 6184 6394 6236 6400
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6196 5914 6224 6258
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 6104 4078 6132 5510
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 6000 2916 6052 2922
rect 6000 2858 6052 2864
rect 6104 2802 6132 3130
rect 6276 2848 6328 2854
rect 5920 2774 6040 2802
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 6012 480 6040 2774
rect 6104 2796 6276 2802
rect 6104 2790 6328 2796
rect 6104 2774 6316 2790
rect 6104 2650 6132 2774
rect 6092 2644 6144 2650
rect 6092 2586 6144 2592
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 6288 2106 6316 2382
rect 6276 2100 6328 2106
rect 6276 2042 6328 2048
rect 6472 480 6500 14418
rect 6564 11937 6592 14758
rect 6656 14385 6684 17478
rect 6734 16688 6790 16697
rect 6840 16674 6868 17818
rect 6932 17202 6960 19858
rect 7116 17649 7144 20318
rect 7392 20210 7420 20334
rect 7208 20182 7420 20210
rect 7102 17640 7158 17649
rect 7102 17575 7158 17584
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 6920 17060 6972 17066
rect 6920 17002 6972 17008
rect 6790 16646 6868 16674
rect 6734 16623 6736 16632
rect 6788 16623 6790 16632
rect 6736 16594 6788 16600
rect 6734 16280 6790 16289
rect 6932 16250 6960 17002
rect 7024 16250 7052 17070
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 7116 16794 7144 16934
rect 7104 16788 7156 16794
rect 7104 16730 7156 16736
rect 7104 16584 7156 16590
rect 7104 16526 7156 16532
rect 6734 16215 6790 16224
rect 6920 16244 6972 16250
rect 6642 14376 6698 14385
rect 6642 14311 6698 14320
rect 6656 12918 6684 14311
rect 6644 12912 6696 12918
rect 6644 12854 6696 12860
rect 6748 12186 6776 16215
rect 6920 16186 6972 16192
rect 7012 16244 7064 16250
rect 7012 16186 7064 16192
rect 7116 16182 7144 16526
rect 7104 16176 7156 16182
rect 7104 16118 7156 16124
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 7012 16108 7064 16114
rect 7012 16050 7064 16056
rect 6840 15706 6868 16050
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 6932 14890 6960 15846
rect 7024 15502 7052 16050
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 7116 15638 7144 15846
rect 7104 15632 7156 15638
rect 7104 15574 7156 15580
rect 7012 15496 7064 15502
rect 7012 15438 7064 15444
rect 6920 14884 6972 14890
rect 6920 14826 6972 14832
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6840 14618 6868 14758
rect 6918 14648 6974 14657
rect 6828 14612 6880 14618
rect 6918 14583 6920 14592
rect 6828 14554 6880 14560
rect 6972 14583 6974 14592
rect 6920 14554 6972 14560
rect 7024 14498 7052 15438
rect 7208 15314 7236 20182
rect 7760 20074 7788 22320
rect 8220 20398 8248 22320
rect 8208 20392 8260 20398
rect 8208 20334 8260 20340
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 7392 20046 7788 20074
rect 7288 19168 7340 19174
rect 7286 19136 7288 19145
rect 7340 19136 7342 19145
rect 7286 19071 7342 19080
rect 7288 18964 7340 18970
rect 7288 18906 7340 18912
rect 7300 17882 7328 18906
rect 7288 17876 7340 17882
rect 7288 17818 7340 17824
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 6840 14470 7052 14498
rect 7116 15286 7236 15314
rect 6840 13870 6868 14470
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6840 12714 6868 13806
rect 6932 13530 6960 14214
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6828 12708 6880 12714
rect 6828 12650 6880 12656
rect 6932 12594 6960 13126
rect 6656 12158 6776 12186
rect 6840 12566 6960 12594
rect 6550 11928 6606 11937
rect 6550 11863 6606 11872
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6564 9058 6592 10746
rect 6656 10713 6684 12158
rect 6736 12096 6788 12102
rect 6840 12084 6868 12566
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 6788 12056 6868 12084
rect 6920 12096 6972 12102
rect 6736 12038 6788 12044
rect 6920 12038 6972 12044
rect 6748 11150 6776 12038
rect 6932 11762 6960 12038
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6828 11552 6880 11558
rect 6828 11494 6880 11500
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6840 10810 6868 11494
rect 6932 11286 6960 11698
rect 6920 11280 6972 11286
rect 6920 11222 6972 11228
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6642 10704 6698 10713
rect 6642 10639 6698 10648
rect 6656 10198 6684 10639
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6644 10192 6696 10198
rect 6644 10134 6696 10140
rect 6748 9178 6776 10474
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 6564 9030 6684 9058
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6564 8809 6592 8910
rect 6550 8800 6606 8809
rect 6550 8735 6606 8744
rect 6550 8528 6606 8537
rect 6550 8463 6606 8472
rect 6564 6798 6592 8463
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6564 6361 6592 6734
rect 6550 6352 6606 6361
rect 6550 6287 6606 6296
rect 6656 6254 6684 9030
rect 6736 8900 6788 8906
rect 6736 8842 6788 8848
rect 6748 8022 6776 8842
rect 6840 8566 6868 9454
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6932 8430 6960 9862
rect 7024 8566 7052 12378
rect 7116 11558 7144 15286
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 7208 13530 7236 15098
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 7208 12986 7236 13330
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7196 12708 7248 12714
rect 7196 12650 7248 12656
rect 7208 12306 7236 12650
rect 7300 12442 7328 15982
rect 7392 13802 7420 20046
rect 8024 19984 8076 19990
rect 8024 19926 8076 19932
rect 7748 19916 7800 19922
rect 7748 19858 7800 19864
rect 7470 19544 7526 19553
rect 7470 19479 7526 19488
rect 7484 18737 7512 19479
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 7564 19236 7616 19242
rect 7564 19178 7616 19184
rect 7470 18728 7526 18737
rect 7470 18663 7526 18672
rect 7472 18080 7524 18086
rect 7470 18048 7472 18057
rect 7524 18048 7526 18057
rect 7470 17983 7526 17992
rect 7472 17740 7524 17746
rect 7472 17682 7524 17688
rect 7484 16794 7512 17682
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 7576 16454 7604 19178
rect 7668 18970 7696 19246
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 7654 18728 7710 18737
rect 7654 18663 7710 18672
rect 7668 18086 7696 18663
rect 7656 18080 7708 18086
rect 7656 18022 7708 18028
rect 7760 17882 7788 19858
rect 8036 19514 8064 19926
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 8116 19712 8168 19718
rect 8116 19654 8168 19660
rect 8024 19508 8076 19514
rect 8024 19450 8076 19456
rect 8128 19242 8156 19654
rect 8116 19236 8168 19242
rect 8116 19178 8168 19184
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 8220 18970 8248 19790
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8312 19514 8340 19654
rect 8300 19508 8352 19514
rect 8300 19450 8352 19456
rect 8668 19168 8720 19174
rect 8390 19136 8446 19145
rect 8668 19110 8720 19116
rect 8390 19071 8446 19080
rect 8208 18964 8260 18970
rect 8208 18906 8260 18912
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 8116 18420 8168 18426
rect 8116 18362 8168 18368
rect 8128 18290 8156 18362
rect 8312 18290 8340 18770
rect 8404 18601 8432 19071
rect 8680 18834 8708 19110
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 8390 18592 8446 18601
rect 8390 18527 8446 18536
rect 8668 18420 8720 18426
rect 8668 18362 8720 18368
rect 8390 18320 8446 18329
rect 8116 18284 8168 18290
rect 8116 18226 8168 18232
rect 8300 18284 8352 18290
rect 8390 18255 8446 18264
rect 8300 18226 8352 18232
rect 8208 18080 8260 18086
rect 8208 18022 8260 18028
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 7840 17808 7892 17814
rect 7840 17750 7892 17756
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 7760 17542 7788 17614
rect 7748 17536 7800 17542
rect 7748 17478 7800 17484
rect 7852 17338 7880 17750
rect 8220 17338 8248 18022
rect 8298 17640 8354 17649
rect 8298 17575 8354 17584
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 7748 17060 7800 17066
rect 7748 17002 7800 17008
rect 7656 16720 7708 16726
rect 7656 16662 7708 16668
rect 7564 16448 7616 16454
rect 7564 16390 7616 16396
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 7484 15162 7512 16186
rect 7576 16046 7604 16390
rect 7564 16040 7616 16046
rect 7564 15982 7616 15988
rect 7668 15162 7696 16662
rect 7760 16046 7788 17002
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8220 16250 8248 16594
rect 8116 16244 8168 16250
rect 8116 16186 8168 16192
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8128 16153 8156 16186
rect 8114 16144 8170 16153
rect 8114 16079 8170 16088
rect 7748 16040 7800 16046
rect 7748 15982 7800 15988
rect 7760 15706 7788 15982
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 7930 15192 7986 15201
rect 7472 15156 7524 15162
rect 7472 15098 7524 15104
rect 7656 15156 7708 15162
rect 7930 15127 7986 15136
rect 7656 15098 7708 15104
rect 7564 15088 7616 15094
rect 7564 15030 7616 15036
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7484 14414 7512 14962
rect 7576 14618 7604 15030
rect 7656 14952 7708 14958
rect 7654 14920 7656 14929
rect 7708 14920 7710 14929
rect 7944 14890 7972 15127
rect 8220 15026 8248 15642
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 7654 14855 7710 14864
rect 7932 14884 7984 14890
rect 7932 14826 7984 14832
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7562 14512 7618 14521
rect 7562 14447 7618 14456
rect 7838 14512 7894 14521
rect 7838 14447 7840 14456
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 7484 13841 7512 14350
rect 7470 13832 7526 13841
rect 7380 13796 7432 13802
rect 7470 13767 7526 13776
rect 7380 13738 7432 13744
rect 7576 13138 7604 14447
rect 7892 14447 7894 14456
rect 7840 14418 7892 14424
rect 8312 13954 8340 17575
rect 8404 15473 8432 18255
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8496 16658 8524 16934
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8390 15464 8446 15473
rect 8390 15399 8446 15408
rect 8404 14414 8432 15399
rect 8588 15162 8616 16730
rect 8576 15156 8628 15162
rect 8576 15098 8628 15104
rect 8576 14816 8628 14822
rect 8576 14758 8628 14764
rect 8588 14550 8616 14758
rect 8576 14544 8628 14550
rect 8576 14486 8628 14492
rect 8680 14482 8708 18362
rect 8668 14476 8720 14482
rect 8668 14418 8720 14424
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8208 13932 8260 13938
rect 8312 13926 8616 13954
rect 8208 13874 8260 13880
rect 8220 13734 8248 13874
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 8300 13728 8352 13734
rect 8300 13670 8352 13676
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7576 13110 7696 13138
rect 7562 13016 7618 13025
rect 7562 12951 7618 12960
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 7196 12164 7248 12170
rect 7196 12106 7248 12112
rect 7208 11830 7236 12106
rect 7196 11824 7248 11830
rect 7196 11766 7248 11772
rect 7104 11552 7156 11558
rect 7156 11512 7236 11540
rect 7104 11494 7156 11500
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 7012 8560 7064 8566
rect 7012 8502 7064 8508
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6840 8090 6868 8230
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6736 8016 6788 8022
rect 6736 7958 6788 7964
rect 6932 7954 6960 8366
rect 7012 8356 7064 8362
rect 7012 8298 7064 8304
rect 7024 8090 7052 8298
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6644 6248 6696 6254
rect 6644 6190 6696 6196
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6656 5914 6684 6054
rect 6748 5914 6776 6598
rect 7116 6322 7144 10134
rect 7208 9926 7236 11512
rect 7392 11354 7420 12718
rect 7380 11348 7432 11354
rect 7300 11308 7380 11336
rect 7300 10130 7328 11308
rect 7380 11290 7432 11296
rect 7380 11008 7432 11014
rect 7380 10950 7432 10956
rect 7392 10656 7420 10950
rect 7472 10668 7524 10674
rect 7392 10628 7472 10656
rect 7472 10610 7524 10616
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7300 9738 7328 9930
rect 7208 9722 7328 9738
rect 7196 9716 7328 9722
rect 7248 9710 7328 9716
rect 7196 9658 7248 9664
rect 7392 9178 7420 10406
rect 7484 9518 7512 10610
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7380 9172 7432 9178
rect 7380 9114 7432 9120
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7470 8800 7526 8809
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7300 8378 7328 8434
rect 7208 8350 7328 8378
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7208 6202 7236 8350
rect 7392 8090 7420 8774
rect 7470 8735 7526 8744
rect 7484 8498 7512 8735
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7300 6866 7328 7346
rect 7392 7342 7420 7686
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7288 6860 7340 6866
rect 7288 6802 7340 6808
rect 7116 6174 7236 6202
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 7012 5772 7064 5778
rect 7012 5714 7064 5720
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6840 4758 6868 5646
rect 7024 5098 7052 5714
rect 7012 5092 7064 5098
rect 7012 5034 7064 5040
rect 6828 4752 6880 4758
rect 6828 4694 6880 4700
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6656 3398 6684 4014
rect 6840 3602 6868 4694
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6932 4214 6960 4626
rect 6920 4208 6972 4214
rect 6920 4150 6972 4156
rect 6932 4026 6960 4150
rect 6932 3998 7052 4026
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 6734 3360 6790 3369
rect 6734 3295 6790 3304
rect 6748 1034 6776 3295
rect 6932 2650 6960 3878
rect 7024 3738 7052 3998
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 7116 3369 7144 6174
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7300 5914 7328 6054
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7392 5846 7420 7278
rect 7472 7268 7524 7274
rect 7472 7210 7524 7216
rect 7196 5840 7248 5846
rect 7194 5808 7196 5817
rect 7380 5840 7432 5846
rect 7248 5808 7250 5817
rect 7380 5782 7432 5788
rect 7194 5743 7250 5752
rect 7484 5234 7512 7210
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7288 5024 7340 5030
rect 7288 4966 7340 4972
rect 7208 4010 7236 4966
rect 7300 4282 7328 4966
rect 7484 4826 7512 5170
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7196 4004 7248 4010
rect 7196 3946 7248 3952
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7392 3738 7420 3878
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7576 3516 7604 12951
rect 7668 11898 7696 13110
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7668 11354 7696 11698
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7668 10198 7696 11290
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 7654 10024 7710 10033
rect 7654 9959 7710 9968
rect 7668 7886 7696 9959
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7668 6322 7696 6734
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7668 5234 7696 6258
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7656 4004 7708 4010
rect 7656 3946 7708 3952
rect 7300 3488 7604 3516
rect 7102 3360 7158 3369
rect 7102 3295 7158 3304
rect 7104 2916 7156 2922
rect 7104 2858 7156 2864
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 7116 2446 7144 2858
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 6748 1006 6868 1034
rect 6840 480 6868 1006
rect 7300 480 7328 3488
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 7484 2922 7512 3130
rect 7472 2916 7524 2922
rect 7472 2858 7524 2864
rect 7576 2446 7604 3130
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7668 1290 7696 3946
rect 7656 1284 7708 1290
rect 7656 1226 7708 1232
rect 7760 480 7788 13466
rect 8220 12714 8248 13670
rect 8312 13530 8340 13670
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8404 13462 8432 13806
rect 8588 13734 8616 13926
rect 8576 13728 8628 13734
rect 8576 13670 8628 13676
rect 8392 13456 8444 13462
rect 8392 13398 8444 13404
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8496 12986 8524 13262
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8588 12918 8616 13670
rect 8576 12912 8628 12918
rect 8576 12854 8628 12860
rect 8772 12764 8800 22320
rect 9232 19938 9260 22320
rect 9692 20466 9720 22320
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9772 20052 9824 20058
rect 9772 19994 9824 20000
rect 8852 19916 8904 19922
rect 9232 19910 9352 19938
rect 8852 19858 8904 19864
rect 8864 18426 8892 19858
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 9220 19848 9272 19854
rect 9220 19790 9272 19796
rect 8956 18970 8984 19790
rect 9128 19236 9180 19242
rect 9128 19178 9180 19184
rect 8944 18964 8996 18970
rect 8944 18906 8996 18912
rect 9034 18864 9090 18873
rect 9034 18799 9090 18808
rect 9048 18426 9076 18799
rect 9140 18766 9168 19178
rect 9232 19174 9260 19790
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 8852 18420 8904 18426
rect 8852 18362 8904 18368
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 9140 18290 9168 18702
rect 9036 18284 9088 18290
rect 9036 18226 9088 18232
rect 9128 18284 9180 18290
rect 9128 18226 9180 18232
rect 9048 17678 9076 18226
rect 8944 17672 8996 17678
rect 8944 17614 8996 17620
rect 9036 17672 9088 17678
rect 9036 17614 9088 17620
rect 8956 17338 8984 17614
rect 9140 17610 9168 18226
rect 9232 17678 9260 19110
rect 9220 17672 9272 17678
rect 9220 17614 9272 17620
rect 9128 17604 9180 17610
rect 9128 17546 9180 17552
rect 8944 17332 8996 17338
rect 8944 17274 8996 17280
rect 9140 17202 9168 17546
rect 9218 17504 9274 17513
rect 9218 17439 9274 17448
rect 9232 17338 9260 17439
rect 9220 17332 9272 17338
rect 9220 17274 9272 17280
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 8852 17060 8904 17066
rect 8852 17002 8904 17008
rect 8588 12736 8800 12764
rect 8864 16232 8892 17002
rect 9140 16794 9168 17138
rect 9128 16788 9180 16794
rect 9128 16730 9180 16736
rect 9128 16652 9180 16658
rect 9128 16594 9180 16600
rect 8944 16244 8996 16250
rect 8864 16204 8944 16232
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 7932 12368 7984 12374
rect 7932 12310 7984 12316
rect 7840 12300 7892 12306
rect 7840 12242 7892 12248
rect 7852 11762 7880 12242
rect 7944 12209 7972 12310
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 7930 12200 7986 12209
rect 7930 12135 7986 12144
rect 8036 11898 8064 12242
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 8220 11150 8248 12650
rect 8300 12640 8352 12646
rect 8298 12608 8300 12617
rect 8352 12608 8354 12617
rect 8298 12543 8354 12552
rect 8390 12336 8446 12345
rect 8390 12271 8446 12280
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 8312 11014 8340 11834
rect 8404 11558 8432 12271
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 8116 10600 8168 10606
rect 8114 10568 8116 10577
rect 8168 10568 8170 10577
rect 8114 10503 8170 10512
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 8220 10266 8248 10610
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8220 9518 8248 10066
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8036 8430 8064 8774
rect 8220 8430 8248 9454
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8128 7188 8156 7822
rect 8220 7750 8248 8366
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8128 7160 8248 7188
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 8220 5658 8248 7160
rect 8312 6866 8340 9658
rect 8404 9058 8432 11494
rect 8496 11354 8524 11494
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8496 9194 8524 10950
rect 8588 10033 8616 12736
rect 8760 12164 8812 12170
rect 8760 12106 8812 12112
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8680 11694 8708 12038
rect 8772 11801 8800 12106
rect 8758 11792 8814 11801
rect 8758 11727 8814 11736
rect 8668 11688 8720 11694
rect 8668 11630 8720 11636
rect 8758 11520 8814 11529
rect 8758 11455 8814 11464
rect 8772 11286 8800 11455
rect 8760 11280 8812 11286
rect 8760 11222 8812 11228
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8574 10024 8630 10033
rect 8680 9994 8708 10406
rect 8574 9959 8630 9968
rect 8668 9988 8720 9994
rect 8668 9930 8720 9936
rect 8496 9166 8708 9194
rect 8404 9030 8616 9058
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8404 7528 8432 8774
rect 8404 7500 8524 7528
rect 8390 7440 8446 7449
rect 8390 7375 8446 7384
rect 8404 6866 8432 7375
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8128 5630 8248 5658
rect 8128 5012 8156 5630
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8220 5166 8248 5510
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8128 4984 8248 5012
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 8220 4865 8248 4984
rect 8206 4856 8262 4865
rect 8206 4791 8262 4800
rect 8312 4758 8340 6598
rect 8496 5930 8524 7500
rect 8404 5902 8524 5930
rect 8404 5137 8432 5902
rect 8484 5840 8536 5846
rect 8484 5782 8536 5788
rect 8496 5710 8524 5782
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8390 5128 8446 5137
rect 8390 5063 8446 5072
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 8404 4826 8432 4966
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 7944 4078 7972 4422
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8220 3194 8248 3470
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8312 3074 8340 4422
rect 8496 4078 8524 5646
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 8220 3046 8340 3074
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 8220 480 8248 3046
rect 8404 2990 8432 3470
rect 8496 2990 8524 4014
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8588 2802 8616 9030
rect 8680 8838 8708 9166
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8772 8480 8800 11222
rect 8864 10713 8892 16204
rect 8944 16186 8996 16192
rect 9034 16008 9090 16017
rect 9034 15943 9090 15952
rect 9048 15570 9076 15943
rect 9036 15564 9088 15570
rect 9036 15506 9088 15512
rect 9140 15450 9168 16594
rect 9048 15422 9168 15450
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 8944 15156 8996 15162
rect 8944 15098 8996 15104
rect 8956 13161 8984 15098
rect 8942 13152 8998 13161
rect 8942 13087 8998 13096
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 8956 11762 8984 12922
rect 9048 11898 9076 15422
rect 9232 15337 9260 15438
rect 9218 15328 9274 15337
rect 9218 15263 9274 15272
rect 9324 15144 9352 19910
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 9496 18692 9548 18698
rect 9496 18634 9548 18640
rect 9588 18692 9640 18698
rect 9588 18634 9640 18640
rect 9508 18426 9536 18634
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 9496 18420 9548 18426
rect 9496 18362 9548 18368
rect 9416 17678 9444 18362
rect 9496 18080 9548 18086
rect 9494 18048 9496 18057
rect 9548 18048 9550 18057
rect 9494 17983 9550 17992
rect 9404 17672 9456 17678
rect 9404 17614 9456 17620
rect 9416 17377 9444 17614
rect 9402 17368 9458 17377
rect 9402 17303 9458 17312
rect 9404 17060 9456 17066
rect 9404 17002 9456 17008
rect 9140 15116 9352 15144
rect 9140 14618 9168 15116
rect 9218 15056 9274 15065
rect 9218 14991 9274 15000
rect 9312 15020 9364 15026
rect 9232 14822 9260 14991
rect 9312 14962 9364 14968
rect 9324 14822 9352 14962
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 9140 14113 9168 14554
rect 9126 14104 9182 14113
rect 9232 14074 9260 14758
rect 9126 14039 9182 14048
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9128 13728 9180 13734
rect 9128 13670 9180 13676
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 9140 11642 9168 13670
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9232 12986 9260 13262
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9218 12472 9274 12481
rect 9218 12407 9274 12416
rect 9232 11762 9260 12407
rect 9324 12209 9352 14758
rect 9310 12200 9366 12209
rect 9310 12135 9366 12144
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 8956 11614 9168 11642
rect 9220 11620 9272 11626
rect 8850 10704 8906 10713
rect 8850 10639 8906 10648
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8864 9110 8892 10406
rect 8956 9178 8984 11614
rect 9220 11562 9272 11568
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9036 11280 9088 11286
rect 9036 11222 9088 11228
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 8852 9104 8904 9110
rect 8852 9046 8904 9052
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8864 8809 8892 8910
rect 8850 8800 8906 8809
rect 8850 8735 8906 8744
rect 8772 8452 8892 8480
rect 8760 8356 8812 8362
rect 8760 8298 8812 8304
rect 8666 8120 8722 8129
rect 8666 8055 8668 8064
rect 8720 8055 8722 8064
rect 8668 8026 8720 8032
rect 8772 8022 8800 8298
rect 8760 8016 8812 8022
rect 8760 7958 8812 7964
rect 8772 7478 8800 7958
rect 8760 7472 8812 7478
rect 8760 7414 8812 7420
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8680 6254 8708 6802
rect 8760 6792 8812 6798
rect 8758 6760 8760 6769
rect 8812 6760 8814 6769
rect 8758 6695 8814 6704
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8772 3754 8800 6598
rect 8864 4486 8892 8452
rect 8956 5574 8984 9114
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 8956 3942 8984 5170
rect 9048 4298 9076 11222
rect 9140 10606 9168 11494
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 9232 10470 9260 11562
rect 9324 10606 9352 11834
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9310 10432 9366 10441
rect 9310 10367 9366 10376
rect 9324 10010 9352 10367
rect 9232 9982 9352 10010
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 9140 8945 9168 8978
rect 9126 8936 9182 8945
rect 9126 8871 9182 8880
rect 9128 8356 9180 8362
rect 9128 8298 9180 8304
rect 9140 6338 9168 8298
rect 9232 6905 9260 9982
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 9218 6896 9274 6905
rect 9218 6831 9274 6840
rect 9324 6662 9352 8230
rect 9416 7410 9444 17002
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9508 15434 9536 16934
rect 9600 16436 9628 18634
rect 9692 18630 9720 19858
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9692 18290 9720 18362
rect 9784 18358 9812 19994
rect 9864 19984 9916 19990
rect 9864 19926 9916 19932
rect 9956 19984 10008 19990
rect 9956 19926 10008 19932
rect 9772 18352 9824 18358
rect 9772 18294 9824 18300
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9876 17218 9904 19926
rect 9968 18426 9996 19926
rect 10046 19136 10102 19145
rect 10046 19071 10102 19080
rect 9956 18420 10008 18426
rect 9956 18362 10008 18368
rect 10060 18068 10088 19071
rect 10152 18193 10180 22320
rect 10232 20392 10284 20398
rect 10232 20334 10284 20340
rect 10244 19446 10272 20334
rect 10508 19916 10560 19922
rect 10508 19858 10560 19864
rect 10416 19848 10468 19854
rect 10416 19790 10468 19796
rect 10428 19718 10456 19790
rect 10416 19712 10468 19718
rect 10416 19654 10468 19660
rect 10322 19544 10378 19553
rect 10322 19479 10378 19488
rect 10232 19440 10284 19446
rect 10232 19382 10284 19388
rect 10232 19168 10284 19174
rect 10230 19136 10232 19145
rect 10284 19136 10286 19145
rect 10230 19071 10286 19080
rect 10336 18873 10364 19479
rect 10416 19304 10468 19310
rect 10416 19246 10468 19252
rect 10322 18864 10378 18873
rect 10322 18799 10378 18808
rect 10230 18456 10286 18465
rect 10428 18426 10456 19246
rect 10230 18391 10286 18400
rect 10416 18420 10468 18426
rect 10138 18184 10194 18193
rect 10138 18119 10194 18128
rect 10244 18068 10272 18391
rect 10416 18362 10468 18368
rect 10416 18080 10468 18086
rect 10060 18040 10180 18068
rect 10244 18040 10416 18068
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 9784 17190 9904 17218
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9692 16726 9720 16934
rect 9680 16720 9732 16726
rect 9680 16662 9732 16668
rect 9680 16448 9732 16454
rect 9600 16408 9680 16436
rect 9680 16390 9732 16396
rect 9692 16046 9720 16390
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9600 15745 9628 15982
rect 9586 15736 9642 15745
rect 9692 15706 9720 15982
rect 9586 15671 9642 15680
rect 9680 15700 9732 15706
rect 9496 15428 9548 15434
rect 9496 15370 9548 15376
rect 9508 13734 9536 15370
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 9600 13274 9628 15671
rect 9680 15642 9732 15648
rect 9692 15570 9720 15642
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9784 15450 9812 17190
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9956 17128 10008 17134
rect 9956 17070 10008 17076
rect 9692 15422 9812 15450
rect 9692 13852 9720 15422
rect 9770 15328 9826 15337
rect 9770 15263 9826 15272
rect 9784 15026 9812 15263
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 9876 14906 9904 17070
rect 9784 14878 9904 14906
rect 9784 14822 9812 14878
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 9772 13864 9824 13870
rect 9692 13824 9772 13852
rect 9772 13806 9824 13812
rect 9876 13394 9904 13942
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 9600 13246 9812 13274
rect 9680 13184 9732 13190
rect 9586 13152 9642 13161
rect 9680 13126 9732 13132
rect 9586 13087 9642 13096
rect 9600 12356 9628 13087
rect 9692 12442 9720 13126
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9508 12328 9628 12356
rect 9508 8294 9536 12328
rect 9784 12288 9812 13246
rect 9600 12260 9812 12288
rect 9600 11558 9628 12260
rect 9772 12096 9824 12102
rect 9678 12064 9734 12073
rect 9772 12038 9824 12044
rect 9678 11999 9734 12008
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9600 11286 9628 11494
rect 9588 11280 9640 11286
rect 9588 11222 9640 11228
rect 9692 11218 9720 11999
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9586 10840 9642 10849
rect 9586 10775 9642 10784
rect 9600 10470 9628 10775
rect 9784 10742 9812 12038
rect 9876 11762 9904 13330
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9772 10736 9824 10742
rect 9772 10678 9824 10684
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9692 10130 9720 10542
rect 9770 10160 9826 10169
rect 9680 10124 9732 10130
rect 9770 10095 9826 10104
rect 9680 10066 9732 10072
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 9588 9444 9640 9450
rect 9588 9386 9640 9392
rect 9600 9110 9628 9386
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 9600 8634 9628 9046
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9508 7478 9536 7890
rect 9600 7886 9628 8570
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9404 6996 9456 7002
rect 9404 6938 9456 6944
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9416 6458 9444 6938
rect 9586 6896 9642 6905
rect 9586 6831 9642 6840
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9140 6310 9260 6338
rect 9128 6248 9180 6254
rect 9128 6190 9180 6196
rect 9140 5710 9168 6190
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9140 4486 9168 4966
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 9048 4270 9168 4298
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8680 3726 8800 3754
rect 8680 2922 8708 3726
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8772 3194 8800 3538
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8668 2916 8720 2922
rect 8668 2858 8720 2864
rect 8772 2802 8800 3130
rect 9034 2952 9090 2961
rect 9034 2887 9036 2896
rect 9088 2887 9090 2896
rect 9036 2858 9088 2864
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 8312 1630 8340 2518
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8404 1834 8432 2382
rect 8496 2009 8524 2790
rect 8588 2774 8708 2802
rect 8772 2774 8892 2802
rect 8482 2000 8538 2009
rect 8482 1935 8538 1944
rect 8392 1828 8444 1834
rect 8392 1770 8444 1776
rect 8300 1624 8352 1630
rect 8300 1566 8352 1572
rect 8680 480 8708 2774
rect 8760 2508 8812 2514
rect 8760 2450 8812 2456
rect 8772 1902 8800 2450
rect 8760 1896 8812 1902
rect 8760 1838 8812 1844
rect 8864 1698 8892 2774
rect 8852 1692 8904 1698
rect 8852 1634 8904 1640
rect 9140 480 9168 4270
rect 9232 3505 9260 6310
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9324 5166 9352 5850
rect 9416 5642 9444 6054
rect 9404 5636 9456 5642
rect 9404 5578 9456 5584
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9416 4826 9444 5102
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9600 4554 9628 6831
rect 9692 6202 9720 9930
rect 9784 6798 9812 10095
rect 9876 8673 9904 11290
rect 9862 8664 9918 8673
rect 9862 8599 9918 8608
rect 9864 8560 9916 8566
rect 9862 8528 9864 8537
rect 9916 8528 9918 8537
rect 9862 8463 9918 8472
rect 9864 8424 9916 8430
rect 9862 8392 9864 8401
rect 9916 8392 9918 8401
rect 9862 8327 9918 8336
rect 9864 8288 9916 8294
rect 9862 8256 9864 8265
rect 9916 8256 9918 8265
rect 9862 8191 9918 8200
rect 9862 8120 9918 8129
rect 9862 8055 9918 8064
rect 9876 7750 9904 8055
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9968 7206 9996 17070
rect 10060 15978 10088 17682
rect 10048 15972 10100 15978
rect 10048 15914 10100 15920
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 10060 13274 10088 14418
rect 10152 14396 10180 18040
rect 10416 18022 10468 18028
rect 10520 17814 10548 19858
rect 10508 17808 10560 17814
rect 10508 17750 10560 17756
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10520 17202 10548 17478
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 10416 16652 10468 16658
rect 10416 16594 10468 16600
rect 10428 15706 10456 16594
rect 10520 15881 10548 17138
rect 10506 15872 10562 15881
rect 10506 15807 10562 15816
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 10244 14618 10272 14758
rect 10336 14618 10364 15098
rect 10232 14612 10284 14618
rect 10232 14554 10284 14560
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 10232 14408 10284 14414
rect 10152 14368 10232 14396
rect 10232 14350 10284 14356
rect 10060 13246 10180 13274
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 10060 12714 10088 13126
rect 10152 12714 10180 13246
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 10140 12708 10192 12714
rect 10140 12650 10192 12656
rect 10152 11354 10180 12650
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10140 11212 10192 11218
rect 10140 11154 10192 11160
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 10060 7546 10088 11086
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 10048 6860 10100 6866
rect 9968 6820 10048 6848
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9864 6724 9916 6730
rect 9864 6666 9916 6672
rect 9876 6633 9904 6666
rect 9862 6624 9918 6633
rect 9862 6559 9918 6568
rect 9692 6174 9904 6202
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9784 5778 9812 6054
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9784 5234 9812 5714
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9692 5114 9720 5170
rect 9692 5086 9812 5114
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9692 4826 9720 4966
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9324 3534 9352 3878
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9312 3528 9364 3534
rect 9218 3496 9274 3505
rect 9312 3470 9364 3476
rect 9218 3431 9274 3440
rect 9324 2378 9352 3470
rect 9416 2854 9444 3538
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 9312 2372 9364 2378
rect 9312 2314 9364 2320
rect 9600 480 9628 4490
rect 9784 3670 9812 5086
rect 9876 5001 9904 6174
rect 9862 4992 9918 5001
rect 9862 4927 9918 4936
rect 9772 3664 9824 3670
rect 9678 3632 9734 3641
rect 9772 3606 9824 3612
rect 9678 3567 9734 3576
rect 9692 2417 9720 3567
rect 9876 2904 9904 4927
rect 9968 3097 9996 6820
rect 10048 6802 10100 6808
rect 10152 6322 10180 11154
rect 10244 10169 10272 14350
rect 10428 13870 10456 15642
rect 10520 15570 10548 15807
rect 10508 15564 10560 15570
rect 10508 15506 10560 15512
rect 10506 15192 10562 15201
rect 10506 15127 10562 15136
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 10322 13016 10378 13025
rect 10322 12951 10378 12960
rect 10520 12968 10548 15127
rect 10612 13138 10640 22320
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 10692 19848 10744 19854
rect 10692 19790 10744 19796
rect 10704 13462 10732 19790
rect 10782 19408 10838 19417
rect 10782 19343 10838 19352
rect 10796 19310 10824 19343
rect 10784 19304 10836 19310
rect 10784 19246 10836 19252
rect 10796 17746 10824 19246
rect 10784 17740 10836 17746
rect 10784 17682 10836 17688
rect 10888 17626 10916 20402
rect 10968 18964 11020 18970
rect 10968 18906 11020 18912
rect 10980 18290 11008 18906
rect 10968 18284 11020 18290
rect 10968 18226 11020 18232
rect 10796 17598 10916 17626
rect 10692 13456 10744 13462
rect 10692 13398 10744 13404
rect 10612 13110 10732 13138
rect 10336 12850 10364 12951
rect 10520 12940 10640 12968
rect 10414 12880 10470 12889
rect 10324 12844 10376 12850
rect 10414 12815 10470 12824
rect 10508 12844 10560 12850
rect 10324 12786 10376 12792
rect 10322 12744 10378 12753
rect 10322 12679 10378 12688
rect 10336 12458 10364 12679
rect 10428 12646 10456 12815
rect 10508 12786 10560 12792
rect 10416 12640 10468 12646
rect 10416 12582 10468 12588
rect 10336 12430 10456 12458
rect 10324 11212 10376 11218
rect 10324 11154 10376 11160
rect 10230 10160 10286 10169
rect 10230 10095 10286 10104
rect 10232 9444 10284 9450
rect 10232 9386 10284 9392
rect 10244 9178 10272 9386
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10244 8634 10272 8910
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10336 8514 10364 11154
rect 10428 10713 10456 12430
rect 10520 11014 10548 12786
rect 10508 11008 10560 11014
rect 10508 10950 10560 10956
rect 10414 10704 10470 10713
rect 10414 10639 10470 10648
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10414 9752 10470 9761
rect 10414 9687 10470 9696
rect 10244 8486 10364 8514
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10046 6080 10102 6089
rect 10046 6015 10102 6024
rect 10060 4010 10088 6015
rect 10140 5092 10192 5098
rect 10140 5034 10192 5040
rect 10152 4282 10180 5034
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 10244 4162 10272 8486
rect 10324 8424 10376 8430
rect 10324 8366 10376 8372
rect 10336 7886 10364 8366
rect 10428 8090 10456 9687
rect 10520 9654 10548 10066
rect 10508 9648 10560 9654
rect 10508 9590 10560 9596
rect 10520 9518 10548 9590
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10520 8945 10548 9318
rect 10506 8936 10562 8945
rect 10506 8871 10562 8880
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10336 7410 10364 7822
rect 10428 7818 10456 8026
rect 10416 7812 10468 7818
rect 10416 7754 10468 7760
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10520 7342 10548 8871
rect 10612 8072 10640 12940
rect 10704 12850 10732 13110
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10704 10588 10732 12582
rect 10796 11150 10824 17598
rect 10966 16688 11022 16697
rect 10966 16623 11022 16632
rect 10980 16153 11008 16623
rect 10966 16144 11022 16153
rect 10966 16079 11022 16088
rect 10876 15972 10928 15978
rect 10876 15914 10928 15920
rect 10888 15434 10916 15914
rect 10968 15564 11020 15570
rect 10968 15506 11020 15512
rect 10876 15428 10928 15434
rect 10876 15370 10928 15376
rect 10888 12850 10916 15370
rect 10980 15201 11008 15506
rect 10966 15192 11022 15201
rect 10966 15127 11022 15136
rect 10968 15020 11020 15026
rect 10968 14962 11020 14968
rect 10980 14414 11008 14962
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 10968 13388 11020 13394
rect 10968 13330 11020 13336
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10980 11830 11008 13330
rect 11072 12306 11100 22320
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 11256 19145 11284 19246
rect 11428 19236 11480 19242
rect 11428 19178 11480 19184
rect 11242 19136 11298 19145
rect 11242 19071 11298 19080
rect 11440 18970 11468 19178
rect 11428 18964 11480 18970
rect 11428 18906 11480 18912
rect 11152 18896 11204 18902
rect 11152 18838 11204 18844
rect 11164 17338 11192 18838
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 11624 17270 11652 22320
rect 12084 19938 12112 22320
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 11992 19910 12112 19938
rect 11704 19848 11756 19854
rect 11704 19790 11756 19796
rect 11716 19242 11744 19790
rect 11704 19236 11756 19242
rect 11704 19178 11756 19184
rect 11702 19136 11758 19145
rect 11702 19071 11758 19080
rect 11716 18834 11744 19071
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11428 17264 11480 17270
rect 11428 17206 11480 17212
rect 11612 17264 11664 17270
rect 11612 17206 11664 17212
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11164 16250 11192 16594
rect 11440 16522 11468 17206
rect 11518 17096 11574 17105
rect 11518 17031 11574 17040
rect 11532 16726 11560 17031
rect 11520 16720 11572 16726
rect 11520 16662 11572 16668
rect 11428 16516 11480 16522
rect 11428 16458 11480 16464
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11164 14958 11192 15438
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11152 14952 11204 14958
rect 11624 14929 11652 17206
rect 11716 16794 11744 17682
rect 11704 16788 11756 16794
rect 11704 16730 11756 16736
rect 11702 16416 11758 16425
rect 11702 16351 11758 16360
rect 11152 14894 11204 14900
rect 11610 14920 11666 14929
rect 11610 14855 11666 14864
rect 11152 14816 11204 14822
rect 11150 14784 11152 14793
rect 11204 14784 11206 14793
rect 11150 14719 11206 14728
rect 11334 14784 11390 14793
rect 11334 14719 11390 14728
rect 11348 14550 11376 14719
rect 11336 14544 11388 14550
rect 11336 14486 11388 14492
rect 11716 14346 11744 16351
rect 11704 14340 11756 14346
rect 11704 14282 11756 14288
rect 11612 14272 11664 14278
rect 11808 14249 11836 18158
rect 11900 16794 11928 19858
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11886 16552 11942 16561
rect 11886 16487 11942 16496
rect 11900 16454 11928 16487
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 11886 16280 11942 16289
rect 11886 16215 11942 16224
rect 11900 15706 11928 16215
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11612 14214 11664 14220
rect 11794 14240 11850 14249
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 11164 13190 11192 13806
rect 11624 13569 11652 14214
rect 11794 14175 11850 14184
rect 11702 14104 11758 14113
rect 11702 14039 11758 14048
rect 11610 13560 11666 13569
rect 11610 13495 11666 13504
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11164 12424 11192 13126
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11520 12912 11572 12918
rect 11520 12854 11572 12860
rect 11164 12396 11284 12424
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 10968 11824 11020 11830
rect 10968 11766 11020 11772
rect 11072 11354 11100 12242
rect 11152 12164 11204 12170
rect 11256 12152 11284 12396
rect 11532 12345 11560 12854
rect 11716 12832 11744 14039
rect 11808 12918 11836 14175
rect 11796 12912 11848 12918
rect 11796 12854 11848 12860
rect 11624 12804 11744 12832
rect 11624 12646 11652 12804
rect 11702 12744 11758 12753
rect 11702 12679 11758 12688
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11518 12336 11574 12345
rect 11518 12271 11574 12280
rect 11336 12164 11388 12170
rect 11256 12124 11336 12152
rect 11152 12106 11204 12112
rect 11336 12106 11388 12112
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 10704 10560 10824 10588
rect 10690 10296 10746 10305
rect 10690 10231 10746 10240
rect 10704 8401 10732 10231
rect 10796 10130 10824 10560
rect 10968 10532 11020 10538
rect 10968 10474 11020 10480
rect 10874 10296 10930 10305
rect 10980 10266 11008 10474
rect 11072 10441 11100 11086
rect 11058 10432 11114 10441
rect 11058 10367 11114 10376
rect 10874 10231 10930 10240
rect 10968 10260 11020 10266
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 10796 9042 10824 10066
rect 10888 9926 10916 10231
rect 10968 10202 11020 10208
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10888 8498 10916 9454
rect 10980 8974 11008 10202
rect 11072 10062 11100 10367
rect 11164 10266 11192 12106
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11624 11812 11652 12582
rect 11716 12322 11744 12679
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11808 12442 11836 12582
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 11716 12294 11836 12322
rect 11704 12164 11756 12170
rect 11704 12106 11756 12112
rect 11334 11792 11390 11801
rect 11334 11727 11390 11736
rect 11532 11784 11652 11812
rect 11348 11286 11376 11727
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 11532 11150 11560 11784
rect 11612 11620 11664 11626
rect 11612 11562 11664 11568
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11624 10742 11652 11562
rect 11612 10736 11664 10742
rect 11612 10678 11664 10684
rect 11152 10260 11204 10266
rect 11152 10202 11204 10208
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11072 9586 11100 9862
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11058 9480 11114 9489
rect 11058 9415 11114 9424
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 11072 8650 11100 9415
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 11242 9344 11298 9353
rect 11164 9178 11192 9318
rect 11242 9279 11298 9288
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 11256 8974 11284 9279
rect 11428 9104 11480 9110
rect 11428 9046 11480 9052
rect 11440 8974 11468 9046
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 10980 8622 11100 8650
rect 10876 8492 10928 8498
rect 10876 8434 10928 8440
rect 10784 8424 10836 8430
rect 10690 8392 10746 8401
rect 10784 8366 10836 8372
rect 10690 8327 10746 8336
rect 10796 8090 10824 8366
rect 10784 8084 10836 8090
rect 10612 8044 10732 8072
rect 10598 7984 10654 7993
rect 10598 7919 10654 7928
rect 10508 7336 10560 7342
rect 10508 7278 10560 7284
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10324 6860 10376 6866
rect 10324 6802 10376 6808
rect 10336 6769 10364 6802
rect 10322 6760 10378 6769
rect 10322 6695 10378 6704
rect 10520 4826 10548 7142
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 10324 4752 10376 4758
rect 10324 4694 10376 4700
rect 10336 4457 10364 4694
rect 10322 4448 10378 4457
rect 10322 4383 10378 4392
rect 10506 4176 10562 4185
rect 10244 4134 10364 4162
rect 10140 4072 10192 4078
rect 10336 4049 10364 4134
rect 10506 4111 10508 4120
rect 10560 4111 10562 4120
rect 10508 4082 10560 4088
rect 10140 4014 10192 4020
rect 10322 4040 10378 4049
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 10152 3194 10180 4014
rect 10232 4004 10284 4010
rect 10322 3975 10378 3984
rect 10232 3946 10284 3952
rect 10244 3602 10272 3946
rect 10612 3942 10640 7919
rect 10704 7410 10732 8044
rect 10980 8072 11008 8622
rect 11060 8560 11112 8566
rect 11060 8502 11112 8508
rect 11072 8090 11100 8502
rect 10784 8026 10836 8032
rect 10888 8044 11008 8072
rect 11060 8084 11112 8090
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10704 6769 10732 7346
rect 10690 6760 10746 6769
rect 10690 6695 10746 6704
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 9954 3088 10010 3097
rect 9954 3023 10010 3032
rect 10244 2922 10272 3538
rect 10324 3528 10376 3534
rect 10508 3528 10560 3534
rect 10324 3470 10376 3476
rect 10506 3496 10508 3505
rect 10560 3496 10562 3505
rect 10336 3398 10364 3470
rect 10506 3431 10562 3440
rect 10600 3460 10652 3466
rect 10600 3402 10652 3408
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 10232 2916 10284 2922
rect 9876 2876 9996 2904
rect 9678 2408 9734 2417
rect 9678 2343 9734 2352
rect 9968 480 9996 2876
rect 10232 2858 10284 2864
rect 10230 2816 10286 2825
rect 10230 2751 10286 2760
rect 10244 2650 10272 2751
rect 10414 2680 10470 2689
rect 10232 2644 10284 2650
rect 10414 2615 10470 2624
rect 10232 2586 10284 2592
rect 10138 2544 10194 2553
rect 10244 2514 10272 2586
rect 10138 2479 10194 2488
rect 10232 2508 10284 2514
rect 10152 2446 10180 2479
rect 10232 2450 10284 2456
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 10428 480 10456 2615
rect 10508 2576 10560 2582
rect 10508 2518 10560 2524
rect 10520 1698 10548 2518
rect 10612 1834 10640 3402
rect 10704 3194 10732 5782
rect 10796 5710 10824 7346
rect 10888 6934 10916 8044
rect 11060 8026 11112 8032
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 10980 7857 11008 7890
rect 10966 7848 11022 7857
rect 10966 7783 11022 7792
rect 11060 7812 11112 7818
rect 11060 7754 11112 7760
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10980 7546 11008 7686
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10876 6928 10928 6934
rect 10876 6870 10928 6876
rect 10980 6633 11008 7142
rect 10966 6624 11022 6633
rect 10966 6559 11022 6568
rect 10876 6180 10928 6186
rect 10876 6122 10928 6128
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10888 5574 10916 6122
rect 10968 6112 11020 6118
rect 10966 6080 10968 6089
rect 11020 6080 11022 6089
rect 10966 6015 11022 6024
rect 11072 5681 11100 7754
rect 11164 6089 11192 8774
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11624 8566 11652 10678
rect 11716 9994 11744 12106
rect 11808 11694 11836 12294
rect 11900 12288 11928 15438
rect 11992 14822 12020 19910
rect 12440 19848 12492 19854
rect 12440 19790 12492 19796
rect 12452 19514 12480 19790
rect 12348 19508 12400 19514
rect 12348 19450 12400 19456
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12254 19408 12310 19417
rect 12360 19394 12388 19450
rect 12360 19366 12480 19394
rect 12254 19343 12310 19352
rect 12268 19292 12296 19343
rect 12348 19304 12400 19310
rect 12268 19264 12348 19292
rect 12348 19246 12400 19252
rect 12256 19168 12308 19174
rect 12256 19110 12308 19116
rect 12162 19000 12218 19009
rect 12072 18964 12124 18970
rect 12162 18935 12218 18944
rect 12072 18906 12124 18912
rect 12084 17660 12112 18906
rect 12176 17882 12204 18935
rect 12268 18766 12296 19110
rect 12452 18970 12480 19366
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 12268 18290 12296 18702
rect 12438 18320 12494 18329
rect 12256 18284 12308 18290
rect 12544 18306 12572 22320
rect 12900 19712 12952 19718
rect 12900 19654 12952 19660
rect 12714 19272 12770 19281
rect 12714 19207 12770 19216
rect 12728 18578 12756 19207
rect 12806 18592 12862 18601
rect 12728 18550 12806 18578
rect 12806 18527 12862 18536
rect 12544 18278 12756 18306
rect 12438 18255 12494 18264
rect 12256 18226 12308 18232
rect 12164 17876 12216 17882
rect 12164 17818 12216 17824
rect 12256 17672 12308 17678
rect 12084 17632 12256 17660
rect 12256 17614 12308 17620
rect 12346 17640 12402 17649
rect 12162 17232 12218 17241
rect 12268 17202 12296 17614
rect 12346 17575 12402 17584
rect 12162 17167 12218 17176
rect 12256 17196 12308 17202
rect 12072 16652 12124 16658
rect 12072 16594 12124 16600
rect 11980 14816 12032 14822
rect 11980 14758 12032 14764
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 11992 12356 12020 14554
rect 12084 12714 12112 16594
rect 12176 14618 12204 17167
rect 12256 17138 12308 17144
rect 12256 16108 12308 16114
rect 12256 16050 12308 16056
rect 12268 15881 12296 16050
rect 12360 15910 12388 17575
rect 12452 16998 12480 18255
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12532 18148 12584 18154
rect 12532 18090 12584 18096
rect 12544 17921 12572 18090
rect 12530 17912 12586 17921
rect 12530 17847 12586 17856
rect 12636 17542 12664 18158
rect 12624 17536 12676 17542
rect 12530 17504 12586 17513
rect 12624 17478 12676 17484
rect 12530 17439 12586 17448
rect 12544 17134 12572 17439
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12636 16590 12664 17478
rect 12728 16640 12756 18278
rect 12820 18193 12848 18527
rect 12806 18184 12862 18193
rect 12806 18119 12862 18128
rect 12799 18080 12851 18086
rect 12912 18068 12940 19654
rect 13004 19281 13032 22320
rect 13464 20210 13492 22320
rect 13464 20182 13676 20210
rect 13268 20052 13320 20058
rect 13268 19994 13320 20000
rect 13084 19304 13136 19310
rect 12990 19272 13046 19281
rect 13084 19246 13136 19252
rect 12990 19207 13046 19216
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 13004 18766 13032 19110
rect 12992 18760 13044 18766
rect 13096 18737 13124 19246
rect 13176 19236 13228 19242
rect 13176 19178 13228 19184
rect 12992 18702 13044 18708
rect 13082 18728 13138 18737
rect 13082 18663 13138 18672
rect 13188 18630 13216 19178
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 13280 18442 13308 19994
rect 13452 19916 13504 19922
rect 13452 19858 13504 19864
rect 13358 19272 13414 19281
rect 13358 19207 13414 19216
rect 13372 18766 13400 19207
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13188 18414 13308 18442
rect 13084 18080 13136 18086
rect 12912 18040 13084 18068
rect 12799 18022 12851 18028
rect 13084 18022 13136 18028
rect 12820 17882 12848 18022
rect 12808 17876 12860 17882
rect 12808 17818 12860 17824
rect 13084 17808 13136 17814
rect 13084 17750 13136 17756
rect 12728 16612 12940 16640
rect 12532 16584 12584 16590
rect 12530 16552 12532 16561
rect 12624 16584 12676 16590
rect 12584 16552 12586 16561
rect 12440 16516 12492 16522
rect 12624 16526 12676 16532
rect 12714 16552 12770 16561
rect 12530 16487 12586 16496
rect 12714 16487 12770 16496
rect 12440 16458 12492 16464
rect 12452 16046 12480 16458
rect 12624 16244 12676 16250
rect 12624 16186 12676 16192
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 12348 15904 12400 15910
rect 12254 15872 12310 15881
rect 12348 15846 12400 15852
rect 12532 15904 12584 15910
rect 12532 15846 12584 15852
rect 12254 15807 12310 15816
rect 12268 15502 12296 15807
rect 12544 15706 12572 15846
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12440 15564 12492 15570
rect 12360 15524 12440 15552
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 12360 14929 12388 15524
rect 12440 15506 12492 15512
rect 12530 15464 12586 15473
rect 12530 15399 12586 15408
rect 12440 15360 12492 15366
rect 12438 15328 12440 15337
rect 12492 15328 12494 15337
rect 12438 15263 12494 15272
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12346 14920 12402 14929
rect 12346 14855 12402 14864
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 12164 14612 12216 14618
rect 12164 14554 12216 14560
rect 12268 13705 12296 14758
rect 12452 13938 12480 14962
rect 12544 14958 12572 15399
rect 12532 14952 12584 14958
rect 12532 14894 12584 14900
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12544 14482 12572 14758
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12348 13728 12400 13734
rect 12254 13696 12310 13705
rect 12348 13670 12400 13676
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12544 13682 12572 14418
rect 12636 14260 12664 16186
rect 12728 15910 12756 16487
rect 12808 16244 12860 16250
rect 12808 16186 12860 16192
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12820 15638 12848 16186
rect 12808 15632 12860 15638
rect 12808 15574 12860 15580
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12714 15192 12770 15201
rect 12714 15127 12716 15136
rect 12768 15127 12770 15136
rect 12716 15098 12768 15104
rect 12714 14920 12770 14929
rect 12714 14855 12770 14864
rect 12728 14618 12756 14855
rect 12716 14612 12768 14618
rect 12716 14554 12768 14560
rect 12716 14272 12768 14278
rect 12636 14232 12716 14260
rect 12636 13938 12664 14232
rect 12716 14214 12768 14220
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12820 13870 12848 15302
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12254 13631 12310 13640
rect 12268 13190 12296 13631
rect 12360 13394 12388 13670
rect 12452 13530 12480 13670
rect 12544 13654 12664 13682
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12636 13462 12664 13654
rect 12624 13456 12676 13462
rect 12624 13398 12676 13404
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 12254 12880 12310 12889
rect 12254 12815 12310 12824
rect 12072 12708 12124 12714
rect 12072 12650 12124 12656
rect 11992 12328 12204 12356
rect 11900 12260 12020 12288
rect 11886 12200 11942 12209
rect 11886 12135 11942 12144
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11796 11552 11848 11558
rect 11796 11494 11848 11500
rect 11808 10674 11836 11494
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11796 10532 11848 10538
rect 11796 10474 11848 10480
rect 11704 9988 11756 9994
rect 11704 9930 11756 9936
rect 11704 9444 11756 9450
rect 11704 9386 11756 9392
rect 11716 9178 11744 9386
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11612 8560 11664 8566
rect 11612 8502 11664 8508
rect 11716 8090 11744 8978
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11244 7472 11296 7478
rect 11244 7414 11296 7420
rect 11256 7274 11284 7414
rect 11244 7268 11296 7274
rect 11244 7210 11296 7216
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11518 6352 11574 6361
rect 11518 6287 11574 6296
rect 11150 6080 11206 6089
rect 11150 6015 11206 6024
rect 11532 5914 11560 6287
rect 11520 5908 11572 5914
rect 11520 5850 11572 5856
rect 11150 5808 11206 5817
rect 11150 5743 11206 5752
rect 11058 5672 11114 5681
rect 10968 5636 11020 5642
rect 11058 5607 11114 5616
rect 10968 5578 11020 5584
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10876 5568 10928 5574
rect 10876 5510 10928 5516
rect 10796 3913 10824 5510
rect 10888 5234 10916 5510
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 10980 5166 11008 5578
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 10968 5160 11020 5166
rect 10874 5128 10930 5137
rect 10968 5102 11020 5108
rect 10874 5063 10930 5072
rect 10782 3904 10838 3913
rect 10782 3839 10838 3848
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10704 2650 10732 3130
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 10600 1828 10652 1834
rect 10600 1770 10652 1776
rect 10508 1692 10560 1698
rect 10508 1634 10560 1640
rect 10888 480 10916 5063
rect 11072 4758 11100 5170
rect 11060 4752 11112 4758
rect 11060 4694 11112 4700
rect 11164 4690 11192 5743
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 10968 4548 11020 4554
rect 10968 4490 11020 4496
rect 10980 4282 11008 4490
rect 11058 4448 11114 4457
rect 11058 4383 11114 4392
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 11072 3670 11100 4383
rect 11164 4049 11192 4626
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11150 4040 11206 4049
rect 11150 3975 11206 3984
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11060 3664 11112 3670
rect 11060 3606 11112 3612
rect 11256 3448 11284 3878
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11532 3641 11560 3674
rect 11518 3632 11574 3641
rect 11518 3567 11574 3576
rect 11624 3466 11652 7890
rect 11808 7206 11836 10474
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11716 6322 11744 6938
rect 11794 6488 11850 6497
rect 11794 6423 11850 6432
rect 11808 6390 11836 6423
rect 11796 6384 11848 6390
rect 11796 6326 11848 6332
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11796 5704 11848 5710
rect 11794 5672 11796 5681
rect 11848 5672 11850 5681
rect 11794 5607 11850 5616
rect 11702 5400 11758 5409
rect 11702 5335 11758 5344
rect 11716 5137 11744 5335
rect 11796 5296 11848 5302
rect 11796 5238 11848 5244
rect 11702 5128 11758 5137
rect 11702 5063 11758 5072
rect 11704 4752 11756 4758
rect 11704 4694 11756 4700
rect 11716 4622 11744 4694
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11716 4146 11744 4558
rect 11808 4146 11836 5238
rect 11900 4298 11928 12135
rect 11992 11098 12020 12260
rect 12070 12200 12126 12209
rect 12070 12135 12126 12144
rect 12084 11801 12112 12135
rect 12070 11792 12126 11801
rect 12070 11727 12126 11736
rect 11992 11070 12112 11098
rect 11980 11008 12032 11014
rect 11980 10950 12032 10956
rect 11992 10198 12020 10950
rect 11980 10192 12032 10198
rect 11980 10134 12032 10140
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 11992 8974 12020 9998
rect 12084 9081 12112 11070
rect 12176 10538 12204 12328
rect 12268 11801 12296 12815
rect 12254 11792 12310 11801
rect 12254 11727 12310 11736
rect 12256 11688 12308 11694
rect 12256 11630 12308 11636
rect 12268 11150 12296 11630
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12256 10600 12308 10606
rect 12256 10542 12308 10548
rect 12164 10532 12216 10538
rect 12164 10474 12216 10480
rect 12268 10441 12296 10542
rect 12254 10432 12310 10441
rect 12254 10367 12310 10376
rect 12164 9988 12216 9994
rect 12164 9930 12216 9936
rect 12070 9072 12126 9081
rect 12070 9007 12126 9016
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 11992 7886 12020 8910
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 11992 6322 12020 7278
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 11992 5234 12020 5510
rect 11980 5228 12032 5234
rect 11980 5170 12032 5176
rect 11978 4856 12034 4865
rect 11978 4791 12034 4800
rect 11992 4622 12020 4791
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11980 4480 12032 4486
rect 11978 4448 11980 4457
rect 12032 4448 12034 4457
rect 11978 4383 12034 4392
rect 11900 4270 12020 4298
rect 11888 4208 11940 4214
rect 11888 4150 11940 4156
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 11164 3420 11284 3448
rect 11612 3460 11664 3466
rect 11164 2666 11192 3420
rect 11612 3402 11664 3408
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11612 3052 11664 3058
rect 11612 2994 11664 3000
rect 10968 2644 11020 2650
rect 11072 2638 11192 2666
rect 11072 2632 11100 2638
rect 11020 2604 11100 2632
rect 10968 2586 11020 2592
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11624 1306 11652 2994
rect 11716 2990 11744 4082
rect 11900 3738 11928 4150
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11808 3194 11836 3470
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 11808 2582 11836 3130
rect 11900 3126 11928 3538
rect 11888 3120 11940 3126
rect 11888 3062 11940 3068
rect 11796 2576 11848 2582
rect 11796 2518 11848 2524
rect 11900 2428 11928 3062
rect 11348 1278 11652 1306
rect 11808 2400 11928 2428
rect 11348 480 11376 1278
rect 11808 480 11836 2400
rect 11992 1442 12020 4270
rect 12084 1766 12112 8366
rect 12176 7886 12204 9930
rect 12360 8974 12388 13330
rect 12452 12646 12480 13330
rect 12532 12844 12584 12850
rect 12636 12832 12664 13398
rect 12716 13252 12768 13258
rect 12716 13194 12768 13200
rect 12584 12804 12664 12832
rect 12532 12786 12584 12792
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12544 11694 12572 12786
rect 12728 12730 12756 13194
rect 12806 13016 12862 13025
rect 12806 12951 12862 12960
rect 12636 12702 12756 12730
rect 12636 12306 12664 12702
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12624 12300 12676 12306
rect 12624 12242 12676 12248
rect 12728 12152 12756 12582
rect 12820 12374 12848 12951
rect 12808 12368 12860 12374
rect 12808 12310 12860 12316
rect 12912 12186 12940 16612
rect 13096 15638 13124 17750
rect 13188 15994 13216 18414
rect 13268 18352 13320 18358
rect 13268 18294 13320 18300
rect 13280 17814 13308 18294
rect 13268 17808 13320 17814
rect 13268 17750 13320 17756
rect 13372 17134 13400 18702
rect 13464 18698 13492 19858
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 13452 18692 13504 18698
rect 13452 18634 13504 18640
rect 13556 18426 13584 19790
rect 13544 18420 13596 18426
rect 13544 18362 13596 18368
rect 13452 18352 13504 18358
rect 13452 18294 13504 18300
rect 13464 18057 13492 18294
rect 13450 18048 13506 18057
rect 13450 17983 13506 17992
rect 13452 17876 13504 17882
rect 13452 17818 13504 17824
rect 13464 17513 13492 17818
rect 13544 17808 13596 17814
rect 13544 17750 13596 17756
rect 13450 17504 13506 17513
rect 13450 17439 13506 17448
rect 13556 17377 13584 17750
rect 13542 17368 13598 17377
rect 13542 17303 13598 17312
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13266 16688 13322 16697
rect 13372 16658 13400 17070
rect 13452 17060 13504 17066
rect 13452 17002 13504 17008
rect 13464 16833 13492 17002
rect 13450 16824 13506 16833
rect 13450 16759 13506 16768
rect 13266 16623 13268 16632
rect 13320 16623 13322 16632
rect 13360 16652 13412 16658
rect 13268 16594 13320 16600
rect 13360 16594 13412 16600
rect 13648 16114 13676 20182
rect 13924 20040 13952 22320
rect 14476 20058 14504 22320
rect 14936 20369 14964 22320
rect 14922 20360 14978 20369
rect 14922 20295 14978 20304
rect 15396 20262 15424 22320
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 14464 20052 14516 20058
rect 13924 20012 14044 20040
rect 13728 19848 13780 19854
rect 13728 19790 13780 19796
rect 13740 19514 13768 19790
rect 13728 19508 13780 19514
rect 13780 19468 13860 19496
rect 13728 19450 13780 19456
rect 13726 19136 13782 19145
rect 13726 19071 13782 19080
rect 13740 18426 13768 19071
rect 13832 18902 13860 19468
rect 13820 18896 13872 18902
rect 13820 18838 13872 18844
rect 13728 18420 13780 18426
rect 13728 18362 13780 18368
rect 13912 18284 13964 18290
rect 13912 18226 13964 18232
rect 13726 18048 13782 18057
rect 13726 17983 13782 17992
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13188 15966 13308 15994
rect 13176 15904 13228 15910
rect 13176 15846 13228 15852
rect 13084 15632 13136 15638
rect 13084 15574 13136 15580
rect 13188 15094 13216 15846
rect 13176 15088 13228 15094
rect 13176 15030 13228 15036
rect 12992 14544 13044 14550
rect 12992 14486 13044 14492
rect 13004 14249 13032 14486
rect 12990 14240 13046 14249
rect 12990 14175 13046 14184
rect 13084 13796 13136 13802
rect 13084 13738 13136 13744
rect 13096 13530 13124 13738
rect 13084 13524 13136 13530
rect 13084 13466 13136 13472
rect 13082 13288 13138 13297
rect 13082 13223 13138 13232
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 13004 12714 13032 13126
rect 12992 12708 13044 12714
rect 12992 12650 13044 12656
rect 12912 12158 13032 12186
rect 12728 12124 12848 12152
rect 12714 12064 12770 12073
rect 12714 11999 12770 12008
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12532 11076 12584 11082
rect 12532 11018 12584 11024
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12452 9518 12480 10542
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12348 8968 12400 8974
rect 12254 8936 12310 8945
rect 12348 8910 12400 8916
rect 12438 8936 12494 8945
rect 12254 8871 12256 8880
rect 12308 8871 12310 8880
rect 12438 8871 12440 8880
rect 12256 8842 12308 8848
rect 12492 8871 12494 8880
rect 12440 8842 12492 8848
rect 12438 8800 12494 8809
rect 12438 8735 12494 8744
rect 12348 8560 12400 8566
rect 12348 8502 12400 8508
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12360 7410 12388 8502
rect 12452 8294 12480 8735
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12544 8022 12572 11018
rect 12622 10840 12678 10849
rect 12622 10775 12678 10784
rect 12532 8016 12584 8022
rect 12532 7958 12584 7964
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12452 7546 12480 7822
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12162 7168 12218 7177
rect 12162 7103 12218 7112
rect 12176 3058 12204 7103
rect 12360 7002 12388 7346
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12544 7002 12572 7142
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12440 6928 12492 6934
rect 12440 6870 12492 6876
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12164 3052 12216 3058
rect 12164 2994 12216 3000
rect 12268 2514 12296 6598
rect 12452 6254 12480 6870
rect 12636 6458 12664 10775
rect 12728 10470 12756 11999
rect 12820 11626 12848 12124
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12808 11620 12860 11626
rect 12808 11562 12860 11568
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12728 9602 12756 10406
rect 12820 10266 12848 11290
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12820 9897 12848 9998
rect 12806 9888 12862 9897
rect 12806 9823 12862 9832
rect 12728 9574 12848 9602
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 12728 6730 12756 7754
rect 12716 6724 12768 6730
rect 12716 6666 12768 6672
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12728 6254 12756 6666
rect 12440 6248 12492 6254
rect 12346 6216 12402 6225
rect 12440 6190 12492 6196
rect 12716 6248 12768 6254
rect 12716 6190 12768 6196
rect 12346 6151 12348 6160
rect 12400 6151 12402 6160
rect 12348 6122 12400 6128
rect 12346 6080 12402 6089
rect 12346 6015 12402 6024
rect 12360 5658 12388 6015
rect 12452 5778 12480 6190
rect 12440 5772 12492 5778
rect 12492 5732 12664 5760
rect 12440 5714 12492 5720
rect 12530 5672 12586 5681
rect 12360 5630 12480 5658
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12360 4865 12388 5306
rect 12452 5166 12480 5630
rect 12530 5607 12586 5616
rect 12544 5273 12572 5607
rect 12530 5264 12586 5273
rect 12530 5199 12586 5208
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12530 5128 12586 5137
rect 12530 5063 12586 5072
rect 12346 4856 12402 4865
rect 12346 4791 12402 4800
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 12360 4321 12388 4558
rect 12346 4312 12402 4321
rect 12346 4247 12402 4256
rect 12452 4185 12480 4626
rect 12438 4176 12494 4185
rect 12438 4111 12494 4120
rect 12544 4026 12572 5063
rect 12360 3998 12572 4026
rect 12360 2961 12388 3998
rect 12636 3942 12664 5732
rect 12728 5234 12756 6190
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12820 5114 12848 9574
rect 12728 5086 12848 5114
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12452 3194 12480 3878
rect 12530 3768 12586 3777
rect 12530 3703 12586 3712
rect 12544 3466 12572 3703
rect 12532 3460 12584 3466
rect 12532 3402 12584 3408
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12346 2952 12402 2961
rect 12346 2887 12402 2896
rect 12360 2650 12388 2887
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 12256 2508 12308 2514
rect 12256 2450 12308 2456
rect 12636 2310 12664 3878
rect 12624 2304 12676 2310
rect 12624 2246 12676 2252
rect 12072 1760 12124 1766
rect 12072 1702 12124 1708
rect 11992 1414 12296 1442
rect 12268 480 12296 1414
rect 12728 480 12756 5086
rect 12808 5024 12860 5030
rect 12808 4966 12860 4972
rect 12820 2650 12848 4966
rect 12912 4593 12940 12038
rect 13004 11558 13032 12158
rect 13096 12073 13124 13223
rect 13188 12889 13216 15030
rect 13280 15026 13308 15966
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 13266 14240 13322 14249
rect 13266 14175 13322 14184
rect 13280 13938 13308 14175
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 13174 12880 13230 12889
rect 13174 12815 13230 12824
rect 13280 12238 13308 13874
rect 13372 13734 13400 16050
rect 13452 15904 13504 15910
rect 13452 15846 13504 15852
rect 13544 15904 13596 15910
rect 13544 15846 13596 15852
rect 13464 13870 13492 15846
rect 13556 15502 13584 15846
rect 13634 15736 13690 15745
rect 13634 15671 13636 15680
rect 13688 15671 13690 15680
rect 13636 15642 13688 15648
rect 13544 15496 13596 15502
rect 13740 15450 13768 17983
rect 13924 17921 13952 18226
rect 13910 17912 13966 17921
rect 13910 17847 13966 17856
rect 13912 17740 13964 17746
rect 13912 17682 13964 17688
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13832 17202 13860 17614
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 13818 16280 13874 16289
rect 13818 16215 13874 16224
rect 13832 15978 13860 16215
rect 13820 15972 13872 15978
rect 13820 15914 13872 15920
rect 13924 15609 13952 17682
rect 14016 16425 14044 20012
rect 14464 19994 14516 20000
rect 14280 19916 14332 19922
rect 14280 19858 14332 19864
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 14188 19712 14240 19718
rect 14188 19654 14240 19660
rect 14096 18896 14148 18902
rect 14096 18838 14148 18844
rect 14108 18290 14136 18838
rect 14096 18284 14148 18290
rect 14096 18226 14148 18232
rect 14200 18170 14228 19654
rect 14292 19553 14320 19858
rect 14372 19848 14424 19854
rect 14648 19848 14700 19854
rect 14372 19790 14424 19796
rect 14568 19808 14648 19836
rect 14278 19544 14334 19553
rect 14278 19479 14334 19488
rect 14384 19417 14412 19790
rect 14464 19780 14516 19786
rect 14464 19722 14516 19728
rect 14370 19408 14426 19417
rect 14370 19343 14426 19352
rect 14476 19310 14504 19722
rect 14464 19304 14516 19310
rect 14464 19246 14516 19252
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14108 18142 14228 18170
rect 14002 16416 14058 16425
rect 14002 16351 14058 16360
rect 14004 15972 14056 15978
rect 14004 15914 14056 15920
rect 13910 15600 13966 15609
rect 13910 15535 13966 15544
rect 13544 15438 13596 15444
rect 13648 15422 13768 15450
rect 14016 15434 14044 15914
rect 14004 15428 14056 15434
rect 13542 14784 13598 14793
rect 13542 14719 13598 14728
rect 13556 14006 13584 14719
rect 13544 14000 13596 14006
rect 13544 13942 13596 13948
rect 13648 13954 13676 15422
rect 14004 15370 14056 15376
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13728 14884 13780 14890
rect 13728 14826 13780 14832
rect 13740 14278 13768 14826
rect 13832 14618 13860 15302
rect 13912 14952 13964 14958
rect 13912 14894 13964 14900
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13728 14272 13780 14278
rect 13726 14240 13728 14249
rect 13780 14240 13782 14249
rect 13726 14175 13782 14184
rect 13924 14113 13952 14894
rect 14004 14408 14056 14414
rect 14004 14350 14056 14356
rect 13910 14104 13966 14113
rect 13910 14039 13966 14048
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 13452 13388 13504 13394
rect 13452 13330 13504 13336
rect 13360 13320 13412 13326
rect 13358 13288 13360 13297
rect 13412 13288 13414 13297
rect 13358 13223 13414 13232
rect 13360 12300 13412 12306
rect 13360 12242 13412 12248
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13372 12102 13400 12242
rect 13464 12220 13492 13330
rect 13556 12753 13584 13942
rect 13648 13926 13768 13954
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 13542 12744 13598 12753
rect 13542 12679 13598 12688
rect 13648 12442 13676 13806
rect 13740 13462 13768 13926
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 13726 13288 13782 13297
rect 13726 13223 13782 13232
rect 13740 13190 13768 13223
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13544 12232 13596 12238
rect 13464 12192 13544 12220
rect 13544 12174 13596 12180
rect 13360 12096 13412 12102
rect 13082 12064 13138 12073
rect 13360 12038 13412 12044
rect 13450 12064 13506 12073
rect 13082 11999 13138 12008
rect 13450 11999 13506 12008
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 12992 11552 13044 11558
rect 13044 11512 13216 11540
rect 12992 11494 13044 11500
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 13004 10849 13032 11086
rect 12990 10840 13046 10849
rect 12990 10775 13046 10784
rect 12990 10704 13046 10713
rect 12990 10639 13046 10648
rect 13004 10606 13032 10639
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 13004 9518 13032 10406
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 12992 8288 13044 8294
rect 13096 8265 13124 11154
rect 13188 10810 13216 11512
rect 13266 11520 13322 11529
rect 13266 11455 13322 11464
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 13176 10600 13228 10606
rect 13176 10542 13228 10548
rect 13188 9722 13216 10542
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 13176 9444 13228 9450
rect 13176 9386 13228 9392
rect 13188 8922 13216 9386
rect 13280 9042 13308 11455
rect 13372 11150 13400 11834
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13372 10538 13400 11086
rect 13360 10532 13412 10538
rect 13360 10474 13412 10480
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 13372 9178 13400 9862
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13188 8906 13308 8922
rect 13188 8900 13320 8906
rect 13188 8894 13268 8900
rect 13268 8842 13320 8848
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 12992 8230 13044 8236
rect 13082 8256 13138 8265
rect 13004 8106 13032 8230
rect 13082 8191 13138 8200
rect 13004 8078 13124 8106
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 13004 6905 13032 7686
rect 12990 6896 13046 6905
rect 12990 6831 13046 6840
rect 13096 6798 13124 8078
rect 13188 7478 13216 8570
rect 13280 8430 13308 8842
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13176 7472 13228 7478
rect 13176 7414 13228 7420
rect 13280 7410 13308 8366
rect 13372 7721 13400 8774
rect 13358 7712 13414 7721
rect 13358 7647 13414 7656
rect 13358 7576 13414 7585
rect 13358 7511 13360 7520
rect 13412 7511 13414 7520
rect 13464 7528 13492 11999
rect 13556 8090 13584 12174
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13648 11218 13676 12038
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13740 10674 13768 12650
rect 13832 11354 13860 13670
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 13924 13297 13952 13330
rect 13910 13288 13966 13297
rect 13910 13223 13966 13232
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 13924 12374 13952 13126
rect 14016 12986 14044 14350
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 13912 12368 13964 12374
rect 13912 12310 13964 12316
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13728 10532 13780 10538
rect 13728 10474 13780 10480
rect 13636 10192 13688 10198
rect 13636 10134 13688 10140
rect 13544 8084 13596 8090
rect 13544 8026 13596 8032
rect 13556 7750 13584 8026
rect 13648 7993 13676 10134
rect 13634 7984 13690 7993
rect 13634 7919 13690 7928
rect 13740 7886 13768 10474
rect 13832 9738 13860 11018
rect 13924 11014 13952 11494
rect 14016 11354 14044 12718
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 14002 10976 14058 10985
rect 13924 10713 13952 10950
rect 14002 10911 14058 10920
rect 13910 10704 13966 10713
rect 13910 10639 13966 10648
rect 13823 9710 13860 9738
rect 13823 9636 13851 9710
rect 13823 9608 13860 9636
rect 13832 9602 13860 9608
rect 13832 9574 13952 9602
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13832 8634 13860 9318
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13924 8294 13952 9574
rect 14016 8498 14044 10911
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13912 8016 13964 8022
rect 13912 7958 13964 7964
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13544 7540 13596 7546
rect 13360 7482 13412 7488
rect 13464 7500 13544 7528
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 13188 6905 13216 7278
rect 13174 6896 13230 6905
rect 13280 6866 13308 7346
rect 13464 7188 13492 7500
rect 13544 7482 13596 7488
rect 13636 7472 13688 7478
rect 13636 7414 13688 7420
rect 13464 7160 13584 7188
rect 13360 6928 13412 6934
rect 13360 6870 13412 6876
rect 13174 6831 13230 6840
rect 13268 6860 13320 6866
rect 13268 6802 13320 6808
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 13096 6458 13124 6734
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 13174 6216 13230 6225
rect 13004 5137 13032 6190
rect 13174 6151 13230 6160
rect 13084 6112 13136 6118
rect 13084 6054 13136 6060
rect 12990 5128 13046 5137
rect 12990 5063 13046 5072
rect 12898 4584 12954 4593
rect 12898 4519 12954 4528
rect 12992 4548 13044 4554
rect 12992 4490 13044 4496
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 12912 3670 12940 4422
rect 12900 3664 12952 3670
rect 12900 3606 12952 3612
rect 13004 3602 13032 4490
rect 12992 3596 13044 3602
rect 12992 3538 13044 3544
rect 12898 3496 12954 3505
rect 12898 3431 12954 3440
rect 12912 2990 12940 3431
rect 12992 3052 13044 3058
rect 12992 2994 13044 3000
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 13004 2582 13032 2994
rect 12992 2576 13044 2582
rect 12992 2518 13044 2524
rect 13096 1154 13124 6054
rect 13188 4570 13216 6151
rect 13280 4690 13308 6598
rect 13372 5370 13400 6870
rect 13556 6497 13584 7160
rect 13542 6488 13598 6497
rect 13452 6452 13504 6458
rect 13542 6423 13598 6432
rect 13452 6394 13504 6400
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13464 5216 13492 6394
rect 13648 6304 13676 7414
rect 13740 6934 13768 7686
rect 13924 7274 13952 7958
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 14016 7750 14044 7890
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 14108 7342 14136 18142
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 14200 17882 14228 18022
rect 14188 17876 14240 17882
rect 14188 17818 14240 17824
rect 14188 17332 14240 17338
rect 14292 17320 14320 18022
rect 14240 17292 14320 17320
rect 14188 17274 14240 17280
rect 14188 17196 14240 17202
rect 14188 17138 14240 17144
rect 14200 16658 14228 17138
rect 14384 17134 14412 18226
rect 14462 17504 14518 17513
rect 14462 17439 14518 17448
rect 14280 17128 14332 17134
rect 14280 17070 14332 17076
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 14188 16652 14240 16658
rect 14188 16594 14240 16600
rect 14200 16289 14228 16594
rect 14186 16280 14242 16289
rect 14186 16215 14242 16224
rect 14292 15366 14320 17070
rect 14384 16726 14412 17070
rect 14372 16720 14424 16726
rect 14372 16662 14424 16668
rect 14370 16416 14426 16425
rect 14370 16351 14426 16360
rect 14384 15638 14412 16351
rect 14476 16250 14504 17439
rect 14464 16244 14516 16250
rect 14464 16186 14516 16192
rect 14464 16040 14516 16046
rect 14464 15982 14516 15988
rect 14372 15632 14424 15638
rect 14372 15574 14424 15580
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14292 15162 14320 15302
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 14186 14104 14242 14113
rect 14186 14039 14188 14048
rect 14240 14039 14242 14048
rect 14188 14010 14240 14016
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 14200 13841 14228 13874
rect 14186 13832 14242 13841
rect 14186 13767 14242 13776
rect 14188 13456 14240 13462
rect 14188 13398 14240 13404
rect 14200 12986 14228 13398
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 14292 12782 14320 14758
rect 14384 14657 14412 15574
rect 14370 14648 14426 14657
rect 14370 14583 14426 14592
rect 14476 13190 14504 15982
rect 14464 13184 14516 13190
rect 14464 13126 14516 13132
rect 14568 13002 14596 19808
rect 14648 19790 14700 19796
rect 15016 19304 15068 19310
rect 15016 19246 15068 19252
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 15028 18737 15056 19246
rect 15108 19168 15160 19174
rect 15108 19110 15160 19116
rect 15014 18728 15070 18737
rect 15014 18663 15070 18672
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 15028 17678 15056 18566
rect 15120 18193 15148 19110
rect 15212 18329 15240 19858
rect 15384 19848 15436 19854
rect 15384 19790 15436 19796
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 15198 18320 15254 18329
rect 15198 18255 15254 18264
rect 15106 18184 15162 18193
rect 15106 18119 15162 18128
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 15108 17808 15160 17814
rect 15108 17750 15160 17756
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 15016 17128 15068 17134
rect 15016 17070 15068 17076
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 15028 16794 15056 17070
rect 15016 16788 15068 16794
rect 15016 16730 15068 16736
rect 14924 16448 14976 16454
rect 14924 16390 14976 16396
rect 14936 16289 14964 16390
rect 14646 16280 14702 16289
rect 14646 16215 14648 16224
rect 14700 16215 14702 16224
rect 14922 16280 14978 16289
rect 14922 16215 14978 16224
rect 14648 16186 14700 16192
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 15016 15564 15068 15570
rect 15016 15506 15068 15512
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 14924 14476 14976 14482
rect 14924 14418 14976 14424
rect 14936 13977 14964 14418
rect 14922 13968 14978 13977
rect 14922 13903 14978 13912
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 15028 13462 15056 15506
rect 15120 14890 15148 17750
rect 15212 16250 15240 18022
rect 15304 17882 15332 18770
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15200 16244 15252 16250
rect 15200 16186 15252 16192
rect 15396 16130 15424 19790
rect 15476 19168 15528 19174
rect 15476 19110 15528 19116
rect 15488 18193 15516 19110
rect 15660 18828 15712 18834
rect 15660 18770 15712 18776
rect 15568 18284 15620 18290
rect 15568 18226 15620 18232
rect 15474 18184 15530 18193
rect 15474 18119 15530 18128
rect 15476 18080 15528 18086
rect 15476 18022 15528 18028
rect 15212 16102 15424 16130
rect 15108 14884 15160 14890
rect 15108 14826 15160 14832
rect 15016 13456 15068 13462
rect 15016 13398 15068 13404
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14384 12974 14596 13002
rect 14280 12776 14332 12782
rect 14186 12744 14242 12753
rect 14280 12718 14332 12724
rect 14186 12679 14242 12688
rect 14200 12238 14228 12679
rect 14188 12232 14240 12238
rect 14240 12192 14320 12220
rect 14188 12174 14240 12180
rect 14186 12064 14242 12073
rect 14186 11999 14242 12008
rect 14200 11393 14228 11999
rect 14186 11384 14242 11393
rect 14186 11319 14242 11328
rect 14292 11150 14320 12192
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14186 10704 14242 10713
rect 14186 10639 14242 10648
rect 14280 10668 14332 10674
rect 14200 10470 14228 10639
rect 14280 10610 14332 10616
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14200 10305 14228 10406
rect 14186 10296 14242 10305
rect 14186 10231 14242 10240
rect 14200 9722 14228 10231
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14200 8430 14228 9318
rect 14292 8838 14320 10610
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 14188 8424 14240 8430
rect 14188 8366 14240 8372
rect 14292 8242 14320 8434
rect 14200 8214 14320 8242
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 13912 7268 13964 7274
rect 13912 7210 13964 7216
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 13728 6928 13780 6934
rect 13728 6870 13780 6876
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 13556 6276 13676 6304
rect 13556 5574 13584 6276
rect 13636 6180 13688 6186
rect 13636 6122 13688 6128
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13648 5234 13676 6122
rect 13832 6118 13860 6734
rect 14004 6384 14056 6390
rect 14004 6326 14056 6332
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13832 5846 13860 6054
rect 13910 5944 13966 5953
rect 13910 5879 13966 5888
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13372 5188 13492 5216
rect 13636 5228 13688 5234
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13188 4542 13308 4570
rect 13174 4176 13230 4185
rect 13174 4111 13230 4120
rect 13188 3369 13216 4111
rect 13174 3360 13230 3369
rect 13174 3295 13230 3304
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 13188 3097 13216 3130
rect 13174 3088 13230 3097
rect 13174 3023 13230 3032
rect 13174 2952 13230 2961
rect 13174 2887 13230 2896
rect 13084 1148 13136 1154
rect 13084 1090 13136 1096
rect 13188 480 13216 2887
rect 13280 1442 13308 4542
rect 13372 2446 13400 5188
rect 13636 5170 13688 5176
rect 13450 5128 13506 5137
rect 13450 5063 13506 5072
rect 13636 5092 13688 5098
rect 13464 2650 13492 5063
rect 13636 5034 13688 5040
rect 13542 4720 13598 4729
rect 13542 4655 13598 4664
rect 13556 3602 13584 4655
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 13542 2952 13598 2961
rect 13542 2887 13598 2896
rect 13556 2854 13584 2887
rect 13544 2848 13596 2854
rect 13544 2790 13596 2796
rect 13648 2650 13676 5034
rect 13740 3942 13768 5510
rect 13832 4826 13860 5578
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13924 4758 13952 5879
rect 14016 5166 14044 6326
rect 14108 5574 14136 7142
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 14200 5302 14228 8214
rect 14384 7698 14412 12974
rect 14464 12776 14516 12782
rect 14660 12753 14688 13262
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 14936 12753 14964 13126
rect 14464 12718 14516 12724
rect 14646 12744 14702 12753
rect 14476 10062 14504 12718
rect 14646 12679 14702 12688
rect 14922 12744 14978 12753
rect 14922 12679 14978 12688
rect 15016 12708 15068 12714
rect 15016 12650 15068 12656
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 15028 12238 15056 12650
rect 15120 12617 15148 13330
rect 15106 12608 15162 12617
rect 15106 12543 15162 12552
rect 15106 12472 15162 12481
rect 15106 12407 15162 12416
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 15016 12232 15068 12238
rect 15016 12174 15068 12180
rect 14660 12073 14688 12174
rect 14740 12164 14792 12170
rect 14740 12106 14792 12112
rect 14646 12064 14702 12073
rect 14646 11999 14702 12008
rect 14752 11762 14780 12106
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 14556 11280 14608 11286
rect 14556 11222 14608 11228
rect 14568 10130 14596 11222
rect 15028 11150 15056 12174
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 14660 10985 14688 11086
rect 14646 10976 14702 10985
rect 14646 10911 14702 10920
rect 15016 10600 15068 10606
rect 15014 10568 15016 10577
rect 15068 10568 15070 10577
rect 15014 10503 15070 10512
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14476 9217 14504 9318
rect 14462 9208 14518 9217
rect 14568 9178 14596 9862
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 14462 9143 14518 9152
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14462 8936 14518 8945
rect 14462 8871 14518 8880
rect 14476 8129 14504 8871
rect 14462 8120 14518 8129
rect 14462 8055 14518 8064
rect 14464 8016 14516 8022
rect 14464 7958 14516 7964
rect 14476 7721 14504 7958
rect 14292 7670 14412 7698
rect 14462 7712 14518 7721
rect 14292 6322 14320 7670
rect 14462 7647 14518 7656
rect 14462 7576 14518 7585
rect 14372 7540 14424 7546
rect 14462 7511 14464 7520
rect 14372 7482 14424 7488
rect 14516 7511 14518 7520
rect 14464 7482 14516 7488
rect 14384 7002 14412 7482
rect 14568 7410 14596 9114
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14660 8498 14688 8774
rect 15028 8673 15056 10503
rect 15014 8664 15070 8673
rect 15014 8599 15070 8608
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 15014 8392 15070 8401
rect 15014 8327 15070 8336
rect 15028 8294 15056 8327
rect 15016 8288 15068 8294
rect 15016 8230 15068 8236
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 14556 7404 14608 7410
rect 15120 7392 15148 12407
rect 15212 11898 15240 16102
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 15396 15881 15424 15982
rect 15382 15872 15438 15881
rect 15382 15807 15438 15816
rect 15384 15088 15436 15094
rect 15384 15030 15436 15036
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15304 14618 15332 14758
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15396 14482 15424 15030
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 15304 13870 15332 14350
rect 15488 14056 15516 18022
rect 15580 16998 15608 18226
rect 15672 18057 15700 18770
rect 15752 18760 15804 18766
rect 15750 18728 15752 18737
rect 15804 18728 15806 18737
rect 15750 18663 15806 18672
rect 15752 18420 15804 18426
rect 15752 18362 15804 18368
rect 15658 18048 15714 18057
rect 15658 17983 15714 17992
rect 15660 17740 15712 17746
rect 15660 17682 15712 17688
rect 15568 16992 15620 16998
rect 15568 16934 15620 16940
rect 15580 16658 15608 16934
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15580 15502 15608 16594
rect 15568 15496 15620 15502
rect 15568 15438 15620 15444
rect 15672 14278 15700 17682
rect 15764 15337 15792 18362
rect 15856 17513 15884 22320
rect 16316 20330 16344 22320
rect 16672 20460 16724 20466
rect 16672 20402 16724 20408
rect 16304 20324 16356 20330
rect 16304 20266 16356 20272
rect 16212 19372 16264 19378
rect 16212 19314 16264 19320
rect 15936 19304 15988 19310
rect 15936 19246 15988 19252
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 15948 17898 15976 19246
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 16040 18057 16068 18566
rect 16026 18048 16082 18057
rect 16026 17983 16082 17992
rect 15948 17870 16068 17898
rect 15936 17740 15988 17746
rect 15936 17682 15988 17688
rect 15842 17504 15898 17513
rect 15842 17439 15898 17448
rect 15844 16720 15896 16726
rect 15844 16662 15896 16668
rect 15856 16114 15884 16662
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 15844 15904 15896 15910
rect 15844 15846 15896 15852
rect 15856 15706 15884 15846
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 15750 15328 15806 15337
rect 15750 15263 15806 15272
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15396 14028 15516 14056
rect 15292 13864 15344 13870
rect 15292 13806 15344 13812
rect 15304 12986 15332 13806
rect 15396 13394 15424 14028
rect 15474 13968 15530 13977
rect 15474 13903 15530 13912
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15488 13326 15516 13903
rect 15764 13802 15792 14758
rect 15752 13796 15804 13802
rect 15752 13738 15804 13744
rect 15856 13682 15884 15642
rect 15948 14113 15976 17682
rect 15934 14104 15990 14113
rect 15934 14039 15990 14048
rect 15672 13654 15884 13682
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15384 13252 15436 13258
rect 15384 13194 15436 13200
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15304 12442 15332 12922
rect 15396 12782 15424 13194
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 15304 12306 15332 12378
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15488 11914 15516 13126
rect 15580 12102 15608 13330
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15200 11892 15252 11898
rect 15488 11886 15608 11914
rect 15200 11834 15252 11840
rect 15474 11792 15530 11801
rect 15474 11727 15530 11736
rect 15488 11558 15516 11727
rect 15580 11694 15608 11886
rect 15559 11688 15611 11694
rect 15559 11630 15611 11636
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15304 11354 15332 11494
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15580 11150 15608 11494
rect 15672 11354 15700 13654
rect 16040 13546 16068 17870
rect 15764 13518 16068 13546
rect 15764 11778 15792 13518
rect 15936 13388 15988 13394
rect 15936 13330 15988 13336
rect 15948 12986 15976 13330
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 15936 12640 15988 12646
rect 16040 12628 16068 13262
rect 15988 12600 16068 12628
rect 15936 12582 15988 12588
rect 15948 12306 15976 12582
rect 15936 12300 15988 12306
rect 15936 12242 15988 12248
rect 16028 12300 16080 12306
rect 16028 12242 16080 12248
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 15764 11750 15884 11778
rect 15948 11762 15976 12038
rect 15752 11688 15804 11694
rect 15752 11630 15804 11636
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 15660 11212 15712 11218
rect 15764 11200 15792 11630
rect 15712 11172 15792 11200
rect 15660 11154 15712 11160
rect 15568 11144 15620 11150
rect 15382 11112 15438 11121
rect 15568 11086 15620 11092
rect 15382 11047 15438 11056
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 15212 10470 15240 10678
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15198 10296 15254 10305
rect 15198 10231 15254 10240
rect 15212 10198 15240 10231
rect 15200 10192 15252 10198
rect 15200 10134 15252 10140
rect 15304 10130 15332 10542
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 15212 8974 15240 9454
rect 15200 8968 15252 8974
rect 15200 8910 15252 8916
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 15212 8362 15240 8774
rect 15200 8356 15252 8362
rect 15200 8298 15252 8304
rect 15200 7948 15252 7954
rect 15200 7890 15252 7896
rect 14556 7346 14608 7352
rect 14660 7364 15148 7392
rect 14660 7290 14688 7364
rect 14476 7262 14688 7290
rect 14372 6996 14424 7002
rect 14372 6938 14424 6944
rect 14372 6860 14424 6866
rect 14372 6802 14424 6808
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 14280 6180 14332 6186
rect 14280 6122 14332 6128
rect 14292 5370 14320 6122
rect 14280 5364 14332 5370
rect 14280 5306 14332 5312
rect 14096 5296 14148 5302
rect 14096 5238 14148 5244
rect 14188 5296 14240 5302
rect 14188 5238 14240 5244
rect 14004 5160 14056 5166
rect 14004 5102 14056 5108
rect 13912 4752 13964 4758
rect 13912 4694 13964 4700
rect 14108 4706 14136 5238
rect 14188 5092 14240 5098
rect 14188 5034 14240 5040
rect 14200 4826 14228 5034
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 14292 4865 14320 4966
rect 14278 4856 14334 4865
rect 14188 4820 14240 4826
rect 14278 4791 14334 4800
rect 14188 4762 14240 4768
rect 14108 4678 14228 4706
rect 13820 4548 13872 4554
rect 13820 4490 13872 4496
rect 13832 4214 13860 4490
rect 14002 4448 14058 4457
rect 14002 4383 14058 4392
rect 14016 4282 14044 4383
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 13820 4208 13872 4214
rect 13820 4150 13872 4156
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 13740 3534 13768 3878
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13726 3224 13782 3233
rect 13726 3159 13782 3168
rect 13740 2972 13768 3159
rect 13832 3126 13860 4014
rect 13924 3233 13952 4218
rect 14096 3936 14148 3942
rect 14002 3904 14058 3913
rect 14096 3878 14148 3884
rect 14002 3839 14058 3848
rect 14016 3738 14044 3839
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 14108 3670 14136 3878
rect 14096 3664 14148 3670
rect 14096 3606 14148 3612
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 13910 3224 13966 3233
rect 13910 3159 13966 3168
rect 13820 3120 13872 3126
rect 13820 3062 13872 3068
rect 13740 2944 13952 2972
rect 13924 2854 13952 2944
rect 13820 2848 13872 2854
rect 13818 2816 13820 2825
rect 13912 2848 13964 2854
rect 13872 2816 13874 2825
rect 13912 2790 13964 2796
rect 13818 2751 13874 2760
rect 13452 2644 13504 2650
rect 13452 2586 13504 2592
rect 13636 2644 13688 2650
rect 13636 2586 13688 2592
rect 13832 2514 13860 2751
rect 13910 2680 13966 2689
rect 13910 2615 13912 2624
rect 13964 2615 13966 2624
rect 13912 2586 13964 2592
rect 13910 2544 13966 2553
rect 13820 2508 13872 2514
rect 13910 2479 13966 2488
rect 13820 2450 13872 2456
rect 13924 2446 13952 2479
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 13280 1414 13584 1442
rect 13556 480 13584 1414
rect 14016 480 14044 3334
rect 14108 3058 14136 3470
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 14200 2310 14228 4678
rect 14280 4684 14332 4690
rect 14280 4626 14332 4632
rect 14292 4078 14320 4626
rect 14280 4072 14332 4078
rect 14280 4014 14332 4020
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 14292 3466 14320 3878
rect 14280 3460 14332 3466
rect 14280 3402 14332 3408
rect 14384 3346 14412 6802
rect 14476 5914 14504 7262
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 14568 6984 14596 7142
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 14568 6956 14688 6984
rect 14660 6390 14688 6956
rect 14832 6792 14884 6798
rect 14832 6734 14884 6740
rect 14648 6384 14700 6390
rect 14648 6326 14700 6332
rect 14844 6186 14872 6734
rect 14924 6656 14976 6662
rect 14924 6598 14976 6604
rect 14936 6497 14964 6598
rect 14922 6488 14978 6497
rect 14922 6423 14978 6432
rect 14832 6180 14884 6186
rect 14832 6122 14884 6128
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 15028 6066 15056 7142
rect 15212 6984 15240 7890
rect 15304 7342 15332 9658
rect 15396 9489 15424 11047
rect 15750 10976 15806 10985
rect 15750 10911 15806 10920
rect 15764 10441 15792 10911
rect 15750 10432 15806 10441
rect 15750 10367 15806 10376
rect 15568 10056 15620 10062
rect 15620 10016 15700 10044
rect 15568 9998 15620 10004
rect 15568 9716 15620 9722
rect 15568 9658 15620 9664
rect 15580 9602 15608 9658
rect 15488 9574 15608 9602
rect 15382 9480 15438 9489
rect 15382 9415 15438 9424
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 15396 8650 15424 8978
rect 15488 8838 15516 9574
rect 15568 9444 15620 9450
rect 15568 9386 15620 9392
rect 15580 8838 15608 9386
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15396 8622 15516 8650
rect 15384 8492 15436 8498
rect 15384 8434 15436 8440
rect 15396 8265 15424 8434
rect 15382 8256 15438 8265
rect 15382 8191 15438 8200
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15488 7274 15516 8622
rect 15580 8498 15608 8774
rect 15672 8634 15700 10016
rect 15764 8809 15792 10367
rect 15856 10169 15884 11750
rect 15936 11756 15988 11762
rect 15936 11698 15988 11704
rect 15948 10606 15976 11698
rect 16040 10849 16068 12242
rect 16026 10840 16082 10849
rect 16026 10775 16082 10784
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 15842 10160 15898 10169
rect 15842 10095 15898 10104
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 15856 9722 15884 9998
rect 15934 9888 15990 9897
rect 15934 9823 15990 9832
rect 15844 9716 15896 9722
rect 15844 9658 15896 9664
rect 15750 8800 15806 8809
rect 15750 8735 15806 8744
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15764 8498 15792 8735
rect 15568 8492 15620 8498
rect 15568 8434 15620 8440
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 15568 8288 15620 8294
rect 15568 8230 15620 8236
rect 15580 8090 15608 8230
rect 15568 8084 15620 8090
rect 15568 8026 15620 8032
rect 15948 7936 15976 9823
rect 16040 9382 16068 9998
rect 16132 9994 16160 19246
rect 16224 18766 16252 19314
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 16224 17898 16252 18702
rect 16304 18624 16356 18630
rect 16304 18566 16356 18572
rect 16316 18057 16344 18566
rect 16488 18148 16540 18154
rect 16488 18090 16540 18096
rect 16302 18048 16358 18057
rect 16302 17983 16358 17992
rect 16224 17870 16344 17898
rect 16212 17128 16264 17134
rect 16212 17070 16264 17076
rect 16224 16454 16252 17070
rect 16212 16448 16264 16454
rect 16212 16390 16264 16396
rect 16224 15434 16252 16390
rect 16212 15428 16264 15434
rect 16212 15370 16264 15376
rect 16224 14890 16252 15370
rect 16212 14884 16264 14890
rect 16212 14826 16264 14832
rect 16210 13288 16266 13297
rect 16210 13223 16266 13232
rect 16224 12073 16252 13223
rect 16210 12064 16266 12073
rect 16210 11999 16266 12008
rect 16316 11642 16344 17870
rect 16500 16674 16528 18090
rect 16592 17882 16620 19246
rect 16684 18970 16712 20402
rect 16776 19281 16804 22320
rect 17328 19938 17356 22320
rect 17788 20398 17816 22320
rect 18248 20890 18276 22320
rect 18708 21706 18736 22320
rect 18970 22128 19026 22137
rect 18970 22063 19026 22072
rect 18616 21678 18736 21706
rect 18510 21176 18566 21185
rect 18510 21111 18566 21120
rect 17880 20862 18276 20890
rect 17776 20392 17828 20398
rect 17776 20334 17828 20340
rect 16960 19910 17356 19938
rect 17408 19916 17460 19922
rect 16762 19272 16818 19281
rect 16762 19207 16818 19216
rect 16672 18964 16724 18970
rect 16672 18906 16724 18912
rect 16672 18760 16724 18766
rect 16672 18702 16724 18708
rect 16684 18601 16712 18702
rect 16670 18592 16726 18601
rect 16670 18527 16726 18536
rect 16960 18426 16988 19910
rect 17408 19858 17460 19864
rect 17040 19848 17092 19854
rect 17040 19790 17092 19796
rect 16948 18420 17000 18426
rect 16948 18362 17000 18368
rect 16764 18352 16816 18358
rect 16764 18294 16816 18300
rect 16776 17882 16804 18294
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 16960 18193 16988 18226
rect 16946 18184 17002 18193
rect 16946 18119 17002 18128
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 16764 17876 16816 17882
rect 16764 17818 16816 17824
rect 16580 17740 16632 17746
rect 16580 17682 16632 17688
rect 16764 17740 16816 17746
rect 16764 17682 16816 17688
rect 16592 16697 16620 17682
rect 16408 16646 16528 16674
rect 16578 16688 16634 16697
rect 16408 15473 16436 16646
rect 16578 16623 16634 16632
rect 16580 16516 16632 16522
rect 16580 16458 16632 16464
rect 16488 15904 16540 15910
rect 16488 15846 16540 15852
rect 16394 15464 16450 15473
rect 16394 15399 16450 15408
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16408 12442 16436 13126
rect 16500 12714 16528 15846
rect 16592 15638 16620 16458
rect 16670 16280 16726 16289
rect 16670 16215 16726 16224
rect 16684 16046 16712 16215
rect 16672 16040 16724 16046
rect 16672 15982 16724 15988
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16684 15706 16712 15846
rect 16672 15700 16724 15706
rect 16672 15642 16724 15648
rect 16580 15632 16632 15638
rect 16580 15574 16632 15580
rect 16776 15366 16804 17682
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 16868 17134 16896 17614
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 16948 17128 17000 17134
rect 16948 17070 17000 17076
rect 16868 16794 16896 17070
rect 16856 16788 16908 16794
rect 16856 16730 16908 16736
rect 16856 16448 16908 16454
rect 16856 16390 16908 16396
rect 16764 15360 16816 15366
rect 16764 15302 16816 15308
rect 16868 15162 16896 16390
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 16672 15088 16724 15094
rect 16672 15030 16724 15036
rect 16684 14929 16712 15030
rect 16764 15020 16816 15026
rect 16764 14962 16816 14968
rect 16670 14920 16726 14929
rect 16670 14855 16726 14864
rect 16580 14000 16632 14006
rect 16580 13942 16632 13948
rect 16488 12708 16540 12714
rect 16488 12650 16540 12656
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16224 11614 16344 11642
rect 16120 9988 16172 9994
rect 16120 9930 16172 9936
rect 16118 9888 16174 9897
rect 16118 9823 16174 9832
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 16040 9110 16068 9318
rect 16028 9104 16080 9110
rect 16028 9046 16080 9052
rect 15856 7908 15976 7936
rect 15568 7880 15620 7886
rect 15568 7822 15620 7828
rect 15476 7268 15528 7274
rect 15476 7210 15528 7216
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15120 6956 15240 6984
rect 15120 6225 15148 6956
rect 15396 6934 15424 7142
rect 15384 6928 15436 6934
rect 15384 6870 15436 6876
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 15212 6458 15240 6802
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 15396 6458 15424 6598
rect 15200 6452 15252 6458
rect 15200 6394 15252 6400
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 15200 6316 15252 6322
rect 15252 6276 15424 6304
rect 15200 6258 15252 6264
rect 15106 6216 15162 6225
rect 15106 6151 15162 6160
rect 15200 6112 15252 6118
rect 15106 6080 15162 6089
rect 14464 5908 14516 5914
rect 14464 5850 14516 5856
rect 14462 5808 14518 5817
rect 14462 5743 14464 5752
rect 14516 5743 14518 5752
rect 14464 5714 14516 5720
rect 14568 5370 14596 6054
rect 15028 6038 15106 6066
rect 14684 6012 14980 6032
rect 15200 6054 15252 6060
rect 15106 6015 15162 6024
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 15106 5944 15162 5953
rect 15106 5879 15162 5888
rect 15016 5772 15068 5778
rect 15016 5714 15068 5720
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 14556 4548 14608 4554
rect 14556 4490 14608 4496
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14476 3448 14504 4082
rect 14568 3602 14596 4490
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 14556 3596 14608 3602
rect 14556 3538 14608 3544
rect 14832 3460 14884 3466
rect 14476 3420 14596 3448
rect 14384 3318 14504 3346
rect 14372 2916 14424 2922
rect 14372 2858 14424 2864
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 14384 2009 14412 2858
rect 14370 2000 14426 2009
rect 14370 1935 14426 1944
rect 14476 480 14504 3318
rect 14568 2961 14596 3420
rect 14832 3402 14884 3408
rect 14646 3224 14702 3233
rect 14646 3159 14648 3168
rect 14700 3159 14702 3168
rect 14648 3130 14700 3136
rect 14740 2984 14792 2990
rect 14554 2952 14610 2961
rect 14844 2972 14872 3402
rect 14792 2944 14872 2972
rect 14740 2926 14792 2932
rect 15028 2922 15056 5714
rect 15120 4570 15148 5879
rect 15212 5846 15240 6054
rect 15200 5840 15252 5846
rect 15200 5782 15252 5788
rect 15212 5234 15240 5782
rect 15396 5778 15424 6276
rect 15384 5772 15436 5778
rect 15384 5714 15436 5720
rect 15290 5264 15346 5273
rect 15200 5228 15252 5234
rect 15290 5199 15346 5208
rect 15200 5170 15252 5176
rect 15304 5098 15332 5199
rect 15292 5092 15344 5098
rect 15292 5034 15344 5040
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15212 4842 15240 4966
rect 15212 4814 15332 4842
rect 15120 4542 15240 4570
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 15120 3670 15148 4422
rect 15212 3738 15240 4542
rect 15200 3732 15252 3738
rect 15200 3674 15252 3680
rect 15108 3664 15160 3670
rect 15108 3606 15160 3612
rect 15304 3058 15332 4814
rect 15396 4690 15424 5714
rect 15580 5166 15608 7822
rect 15660 7812 15712 7818
rect 15660 7754 15712 7760
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15568 5160 15620 5166
rect 15568 5102 15620 5108
rect 15384 4684 15436 4690
rect 15384 4626 15436 4632
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 15396 3738 15424 3878
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15384 3596 15436 3602
rect 15384 3538 15436 3544
rect 15108 3052 15160 3058
rect 15108 2994 15160 3000
rect 15292 3052 15344 3058
rect 15292 2994 15344 3000
rect 14554 2887 14610 2896
rect 15016 2916 15068 2922
rect 15016 2858 15068 2864
rect 15120 2802 15148 2994
rect 15292 2916 15344 2922
rect 15292 2858 15344 2864
rect 15028 2774 15148 2802
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 15028 2446 15056 2774
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15108 2508 15160 2514
rect 15108 2450 15160 2456
rect 15016 2440 15068 2446
rect 15016 2382 15068 2388
rect 14924 2304 14976 2310
rect 14924 2246 14976 2252
rect 14936 480 14964 2246
rect 15120 2038 15148 2450
rect 15108 2032 15160 2038
rect 15108 1974 15160 1980
rect 15212 1902 15240 2586
rect 15304 1970 15332 2858
rect 15396 2417 15424 3538
rect 15488 3194 15516 5102
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 15672 2650 15700 7754
rect 15752 7472 15804 7478
rect 15752 7414 15804 7420
rect 15764 4026 15792 7414
rect 15856 6934 15884 7908
rect 16026 7712 16082 7721
rect 16026 7647 16082 7656
rect 15936 7404 15988 7410
rect 15936 7346 15988 7352
rect 15844 6928 15896 6934
rect 15842 6896 15844 6905
rect 15896 6896 15898 6905
rect 15842 6831 15898 6840
rect 15844 5228 15896 5234
rect 15844 5170 15896 5176
rect 15856 4826 15884 5170
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 15856 4146 15884 4762
rect 15948 4758 15976 7346
rect 15936 4752 15988 4758
rect 15936 4694 15988 4700
rect 15844 4140 15896 4146
rect 15844 4082 15896 4088
rect 15764 3998 15884 4026
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15660 2644 15712 2650
rect 15660 2586 15712 2592
rect 15764 2582 15792 3674
rect 15752 2576 15804 2582
rect 15752 2518 15804 2524
rect 15382 2408 15438 2417
rect 15382 2343 15438 2352
rect 15292 1964 15344 1970
rect 15292 1906 15344 1912
rect 15200 1896 15252 1902
rect 15200 1838 15252 1844
rect 15384 1148 15436 1154
rect 15384 1090 15436 1096
rect 15396 480 15424 1090
rect 15856 480 15884 3998
rect 15934 2680 15990 2689
rect 16040 2650 16068 7647
rect 16132 5166 16160 9823
rect 16224 9654 16252 11614
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16302 11384 16358 11393
rect 16408 11354 16436 11494
rect 16302 11319 16358 11328
rect 16396 11348 16448 11354
rect 16212 9648 16264 9654
rect 16212 9590 16264 9596
rect 16316 9466 16344 11319
rect 16396 11290 16448 11296
rect 16500 11234 16528 12650
rect 16592 12594 16620 13942
rect 16776 13802 16804 14962
rect 16856 14884 16908 14890
rect 16856 14826 16908 14832
rect 16764 13796 16816 13802
rect 16764 13738 16816 13744
rect 16672 13728 16724 13734
rect 16672 13670 16724 13676
rect 16762 13696 16818 13705
rect 16684 12850 16712 13670
rect 16762 13631 16818 13640
rect 16776 13433 16804 13631
rect 16762 13424 16818 13433
rect 16762 13359 16764 13368
rect 16816 13359 16818 13368
rect 16764 13330 16816 13336
rect 16672 12844 16724 12850
rect 16724 12804 16804 12832
rect 16672 12786 16724 12792
rect 16592 12566 16712 12594
rect 16684 11558 16712 12566
rect 16776 11762 16804 12804
rect 16868 12306 16896 14826
rect 16960 14482 16988 17070
rect 17052 16017 17080 19790
rect 17132 19372 17184 19378
rect 17132 19314 17184 19320
rect 17144 17864 17172 19314
rect 17314 18456 17370 18465
rect 17314 18391 17370 18400
rect 17328 18290 17356 18391
rect 17316 18284 17368 18290
rect 17316 18226 17368 18232
rect 17224 18080 17276 18086
rect 17222 18048 17224 18057
rect 17276 18048 17278 18057
rect 17222 17983 17278 17992
rect 17144 17836 17264 17864
rect 17132 17740 17184 17746
rect 17132 17682 17184 17688
rect 17144 16998 17172 17682
rect 17132 16992 17184 16998
rect 17132 16934 17184 16940
rect 17132 16720 17184 16726
rect 17130 16688 17132 16697
rect 17184 16688 17186 16697
rect 17130 16623 17186 16632
rect 17132 16244 17184 16250
rect 17132 16186 17184 16192
rect 17038 16008 17094 16017
rect 17038 15943 17094 15952
rect 17040 15360 17092 15366
rect 17040 15302 17092 15308
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 17052 14414 17080 15302
rect 17040 14408 17092 14414
rect 17040 14350 17092 14356
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 16946 13832 17002 13841
rect 16946 13767 16948 13776
rect 17000 13767 17002 13776
rect 16948 13738 17000 13744
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16960 13161 16988 13330
rect 16946 13152 17002 13161
rect 16946 13087 17002 13096
rect 16946 12472 17002 12481
rect 16946 12407 16948 12416
rect 17000 12407 17002 12416
rect 16948 12378 17000 12384
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16854 11792 16910 11801
rect 16764 11756 16816 11762
rect 16854 11727 16856 11736
rect 16764 11698 16816 11704
rect 16908 11727 16910 11736
rect 16856 11698 16908 11704
rect 17052 11642 17080 14214
rect 17144 13530 17172 16186
rect 17236 15094 17264 17836
rect 17316 17332 17368 17338
rect 17316 17274 17368 17280
rect 17328 16969 17356 17274
rect 17314 16960 17370 16969
rect 17314 16895 17370 16904
rect 17420 16794 17448 19858
rect 17880 19417 17908 20862
rect 17960 19984 18012 19990
rect 17960 19926 18012 19932
rect 17866 19408 17922 19417
rect 17866 19343 17922 19352
rect 17972 18902 18000 19926
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 18050 19408 18106 19417
rect 18050 19343 18106 19352
rect 17776 18896 17828 18902
rect 17960 18896 18012 18902
rect 17776 18838 17828 18844
rect 17866 18864 17922 18873
rect 17592 18760 17644 18766
rect 17592 18702 17644 18708
rect 17500 18352 17552 18358
rect 17500 18294 17552 18300
rect 17408 16788 17460 16794
rect 17408 16730 17460 16736
rect 17316 16584 17368 16590
rect 17316 16526 17368 16532
rect 17224 15088 17276 15094
rect 17224 15030 17276 15036
rect 17224 13728 17276 13734
rect 17224 13670 17276 13676
rect 17132 13524 17184 13530
rect 17132 13466 17184 13472
rect 17130 13424 17186 13433
rect 17130 13359 17186 13368
rect 17144 11694 17172 13359
rect 17236 13025 17264 13670
rect 17222 13016 17278 13025
rect 17222 12951 17278 12960
rect 17224 12776 17276 12782
rect 17224 12718 17276 12724
rect 16868 11614 17080 11642
rect 17132 11688 17184 11694
rect 17132 11630 17184 11636
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16580 11348 16632 11354
rect 16632 11308 16712 11336
rect 16580 11290 16632 11296
rect 16408 11206 16528 11234
rect 16580 11212 16632 11218
rect 16408 9761 16436 11206
rect 16580 11154 16632 11160
rect 16488 11076 16540 11082
rect 16488 11018 16540 11024
rect 16500 10985 16528 11018
rect 16486 10976 16542 10985
rect 16486 10911 16542 10920
rect 16592 10810 16620 11154
rect 16580 10804 16632 10810
rect 16580 10746 16632 10752
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16488 10464 16540 10470
rect 16488 10406 16540 10412
rect 16394 9752 16450 9761
rect 16394 9687 16450 9696
rect 16224 9438 16344 9466
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 16132 3738 16160 5102
rect 16224 5001 16252 9438
rect 16302 8800 16358 8809
rect 16302 8735 16358 8744
rect 16316 8362 16344 8735
rect 16500 8634 16528 10406
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16304 8356 16356 8362
rect 16304 8298 16356 8304
rect 16316 7857 16344 8298
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16302 7848 16358 7857
rect 16302 7783 16358 7792
rect 16304 7744 16356 7750
rect 16304 7686 16356 7692
rect 16316 7410 16344 7686
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16210 4992 16266 5001
rect 16210 4927 16266 4936
rect 16212 4276 16264 4282
rect 16212 4218 16264 4224
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 15934 2615 15936 2624
rect 15988 2615 15990 2624
rect 16028 2644 16080 2650
rect 15936 2586 15988 2592
rect 16028 2586 16080 2592
rect 16132 2446 16160 2994
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 16224 626 16252 4218
rect 16316 2854 16344 7142
rect 16304 2848 16356 2854
rect 16304 2790 16356 2796
rect 16408 2378 16436 7890
rect 16592 7750 16620 10542
rect 16684 9466 16712 11308
rect 16770 11144 16822 11150
rect 16770 11086 16822 11092
rect 16776 10577 16804 11086
rect 16868 10606 16896 11614
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16856 10600 16908 10606
rect 16762 10568 16818 10577
rect 16856 10542 16908 10548
rect 16762 10503 16818 10512
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 16868 10062 16896 10406
rect 16764 10056 16816 10062
rect 16762 10024 16764 10033
rect 16856 10056 16908 10062
rect 16816 10024 16818 10033
rect 16856 9998 16908 10004
rect 16762 9959 16818 9968
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 16776 9586 16804 9862
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16684 9438 16804 9466
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16684 9178 16712 9318
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 16684 8650 16712 8978
rect 16776 8838 16804 9438
rect 16868 8974 16896 9998
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 16684 8622 16804 8650
rect 16776 8498 16804 8622
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16672 7948 16724 7954
rect 16672 7890 16724 7896
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 16500 6458 16528 6802
rect 16580 6792 16632 6798
rect 16684 6780 16712 7890
rect 16776 7886 16804 8434
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 16960 7818 16988 11494
rect 17236 11234 17264 12718
rect 17328 12646 17356 16526
rect 17408 15632 17460 15638
rect 17408 15574 17460 15580
rect 17420 14958 17448 15574
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17420 13938 17448 14758
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17316 12640 17368 12646
rect 17314 12608 17316 12617
rect 17368 12608 17370 12617
rect 17314 12543 17370 12552
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17040 11212 17092 11218
rect 17040 11154 17092 11160
rect 17144 11206 17264 11234
rect 17052 10985 17080 11154
rect 17038 10976 17094 10985
rect 17038 10911 17094 10920
rect 17040 9920 17092 9926
rect 17040 9862 17092 9868
rect 16948 7812 17000 7818
rect 16948 7754 17000 7760
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16764 7200 16816 7206
rect 16762 7168 16764 7177
rect 16816 7168 16818 7177
rect 16762 7103 16818 7112
rect 16632 6752 16712 6780
rect 16868 6746 16896 7278
rect 16948 7200 17000 7206
rect 16948 7142 17000 7148
rect 16580 6734 16632 6740
rect 16488 6452 16540 6458
rect 16488 6394 16540 6400
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16500 6186 16528 6258
rect 16592 6254 16620 6734
rect 16776 6718 16896 6746
rect 16670 6488 16726 6497
rect 16670 6423 16726 6432
rect 16684 6254 16712 6423
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16672 6248 16724 6254
rect 16672 6190 16724 6196
rect 16488 6180 16540 6186
rect 16488 6122 16540 6128
rect 16500 5914 16528 6122
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16488 5908 16540 5914
rect 16488 5850 16540 5856
rect 16580 5160 16632 5166
rect 16578 5128 16580 5137
rect 16632 5128 16634 5137
rect 16578 5063 16634 5072
rect 16488 4752 16540 4758
rect 16488 4694 16540 4700
rect 16500 4214 16528 4694
rect 16488 4208 16540 4214
rect 16684 4196 16712 6054
rect 16488 4150 16540 4156
rect 16592 4168 16712 4196
rect 16500 3534 16528 4150
rect 16592 4078 16620 4168
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16672 4072 16724 4078
rect 16672 4014 16724 4020
rect 16580 3936 16632 3942
rect 16578 3904 16580 3913
rect 16632 3904 16634 3913
rect 16578 3839 16634 3848
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 16396 2372 16448 2378
rect 16396 2314 16448 2320
rect 16592 2009 16620 3839
rect 16578 2000 16634 2009
rect 16578 1935 16634 1944
rect 16684 1850 16712 4014
rect 16776 2922 16804 6718
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 16868 6458 16896 6598
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16960 5778 16988 7142
rect 16948 5772 17000 5778
rect 16948 5714 17000 5720
rect 16946 5536 17002 5545
rect 16946 5471 17002 5480
rect 16856 5024 16908 5030
rect 16856 4966 16908 4972
rect 16764 2916 16816 2922
rect 16764 2858 16816 2864
rect 16868 2038 16896 4966
rect 16960 4758 16988 5471
rect 16948 4752 17000 4758
rect 16948 4694 17000 4700
rect 17052 3602 17080 9862
rect 17144 8650 17172 11206
rect 17328 11121 17356 11290
rect 17420 11150 17448 13874
rect 17408 11144 17460 11150
rect 17314 11112 17370 11121
rect 17408 11086 17460 11092
rect 17314 11047 17370 11056
rect 17316 11008 17368 11014
rect 17316 10950 17368 10956
rect 17224 10736 17276 10742
rect 17222 10704 17224 10713
rect 17276 10704 17278 10713
rect 17222 10639 17278 10648
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17236 9450 17264 10406
rect 17328 10305 17356 10950
rect 17420 10674 17448 11086
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17314 10296 17370 10305
rect 17314 10231 17370 10240
rect 17314 10024 17370 10033
rect 17314 9959 17370 9968
rect 17224 9444 17276 9450
rect 17224 9386 17276 9392
rect 17328 8945 17356 9959
rect 17406 9888 17462 9897
rect 17406 9823 17462 9832
rect 17420 9518 17448 9823
rect 17408 9512 17460 9518
rect 17408 9454 17460 9460
rect 17314 8936 17370 8945
rect 17314 8871 17370 8880
rect 17144 8622 17264 8650
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 16946 2680 17002 2689
rect 16946 2615 16948 2624
rect 17000 2615 17002 2624
rect 16948 2586 17000 2592
rect 16856 2032 16908 2038
rect 16856 1974 16908 1980
rect 16684 1822 16804 1850
rect 16672 1692 16724 1698
rect 16672 1634 16724 1640
rect 16224 598 16344 626
rect 16316 480 16344 598
rect 16684 480 16712 1634
rect 16776 1358 16804 1822
rect 16764 1352 16816 1358
rect 16764 1294 16816 1300
rect 17144 480 17172 8502
rect 17236 6458 17264 8622
rect 17420 7546 17448 9454
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 17224 6452 17276 6458
rect 17224 6394 17276 6400
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 17328 5234 17356 5646
rect 17316 5228 17368 5234
rect 17316 5170 17368 5176
rect 17328 4826 17356 5170
rect 17408 5024 17460 5030
rect 17408 4966 17460 4972
rect 17316 4820 17368 4826
rect 17316 4762 17368 4768
rect 17222 4312 17278 4321
rect 17222 4247 17278 4256
rect 17236 2632 17264 4247
rect 17314 3768 17370 3777
rect 17420 3738 17448 4966
rect 17314 3703 17316 3712
rect 17368 3703 17370 3712
rect 17408 3732 17460 3738
rect 17316 3674 17368 3680
rect 17408 3674 17460 3680
rect 17512 3670 17540 18294
rect 17604 12617 17632 18702
rect 17684 18624 17736 18630
rect 17684 18566 17736 18572
rect 17590 12608 17646 12617
rect 17590 12543 17646 12552
rect 17590 12336 17646 12345
rect 17590 12271 17646 12280
rect 17604 11898 17632 12271
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17590 11792 17646 11801
rect 17696 11778 17724 18566
rect 17788 17785 17816 18838
rect 17960 18838 18012 18844
rect 17866 18799 17868 18808
rect 17920 18799 17922 18808
rect 17868 18770 17920 18776
rect 18064 18714 18092 19343
rect 18420 19304 18472 19310
rect 18420 19246 18472 19252
rect 18432 18873 18460 19246
rect 18524 19174 18552 21111
rect 18616 19825 18644 21678
rect 18694 21584 18750 21593
rect 18694 21519 18750 21528
rect 18602 19816 18658 19825
rect 18602 19751 18658 19760
rect 18602 19272 18658 19281
rect 18602 19207 18658 19216
rect 18512 19168 18564 19174
rect 18512 19110 18564 19116
rect 18616 18970 18644 19207
rect 18708 19174 18736 21519
rect 18984 20058 19012 22063
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 18880 19916 18932 19922
rect 18880 19858 18932 19864
rect 18788 19712 18840 19718
rect 18788 19654 18840 19660
rect 18696 19168 18748 19174
rect 18696 19110 18748 19116
rect 18604 18964 18656 18970
rect 18604 18906 18656 18912
rect 18418 18864 18474 18873
rect 18694 18864 18750 18873
rect 18418 18799 18474 18808
rect 18604 18828 18656 18834
rect 18694 18799 18750 18808
rect 18604 18770 18656 18776
rect 17972 18686 18092 18714
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 17866 18184 17922 18193
rect 17866 18119 17922 18128
rect 17774 17776 17830 17785
rect 17774 17711 17830 17720
rect 17776 17672 17828 17678
rect 17776 17614 17828 17620
rect 17788 16794 17816 17614
rect 17880 17338 17908 18119
rect 17972 17649 18000 18686
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 18236 18352 18288 18358
rect 18236 18294 18288 18300
rect 18052 18080 18104 18086
rect 18050 18048 18052 18057
rect 18104 18048 18106 18057
rect 18050 17983 18106 17992
rect 17958 17640 18014 17649
rect 17958 17575 18014 17584
rect 18248 17524 18276 18294
rect 17972 17496 18276 17524
rect 17972 17338 18000 17496
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 17868 17332 17920 17338
rect 17868 17274 17920 17280
rect 17960 17332 18012 17338
rect 17960 17274 18012 17280
rect 17866 16824 17922 16833
rect 17776 16788 17828 16794
rect 17866 16759 17922 16768
rect 17776 16730 17828 16736
rect 17774 16688 17830 16697
rect 17774 16623 17776 16632
rect 17828 16623 17830 16632
rect 17776 16594 17828 16600
rect 17776 16516 17828 16522
rect 17776 16458 17828 16464
rect 17788 16114 17816 16458
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17774 15464 17830 15473
rect 17774 15399 17830 15408
rect 17788 12617 17816 15399
rect 17880 14618 17908 16759
rect 17972 16425 18000 17274
rect 18420 17264 18472 17270
rect 18420 17206 18472 17212
rect 18328 17060 18380 17066
rect 18328 17002 18380 17008
rect 18052 16992 18104 16998
rect 18144 16992 18196 16998
rect 18052 16934 18104 16940
rect 18142 16960 18144 16969
rect 18340 16969 18368 17002
rect 18196 16960 18198 16969
rect 18064 16726 18092 16934
rect 18142 16895 18198 16904
rect 18326 16960 18382 16969
rect 18326 16895 18382 16904
rect 18236 16788 18288 16794
rect 18236 16730 18288 16736
rect 18052 16720 18104 16726
rect 18052 16662 18104 16668
rect 18248 16561 18276 16730
rect 18432 16590 18460 17206
rect 18524 16794 18552 18702
rect 18616 18222 18644 18770
rect 18708 18426 18736 18799
rect 18696 18420 18748 18426
rect 18696 18362 18748 18368
rect 18800 18329 18828 19654
rect 18892 19446 18920 19858
rect 18972 19780 19024 19786
rect 18972 19722 19024 19728
rect 18880 19440 18932 19446
rect 18880 19382 18932 19388
rect 18880 19168 18932 19174
rect 18880 19110 18932 19116
rect 18786 18320 18842 18329
rect 18786 18255 18842 18264
rect 18604 18216 18656 18222
rect 18604 18158 18656 18164
rect 18696 18148 18748 18154
rect 18696 18090 18748 18096
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 18510 16688 18566 16697
rect 18510 16623 18512 16632
rect 18564 16623 18566 16632
rect 18512 16594 18564 16600
rect 18420 16584 18472 16590
rect 18234 16552 18290 16561
rect 18420 16526 18472 16532
rect 18234 16487 18290 16496
rect 17958 16416 18014 16425
rect 18510 16416 18566 16425
rect 17958 16351 18014 16360
rect 18116 16348 18412 16368
rect 18510 16351 18566 16360
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 18524 16250 18552 16351
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 17960 15360 18012 15366
rect 17960 15302 18012 15308
rect 18512 15360 18564 15366
rect 18512 15302 18564 15308
rect 17972 15026 18000 15302
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 18052 15088 18104 15094
rect 18052 15030 18104 15036
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17958 14920 18014 14929
rect 17958 14855 18014 14864
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17880 13870 17908 14214
rect 17972 14074 18000 14855
rect 18064 14657 18092 15030
rect 18524 15026 18552 15302
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18050 14648 18106 14657
rect 18050 14583 18106 14592
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 18418 13968 18474 13977
rect 18418 13903 18474 13912
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17880 13190 17908 13806
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 18328 13796 18380 13802
rect 18328 13738 18380 13744
rect 17972 13530 18000 13738
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 18340 13326 18368 13738
rect 18432 13462 18460 13903
rect 18420 13456 18472 13462
rect 18420 13398 18472 13404
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 17868 13184 17920 13190
rect 17868 13126 17920 13132
rect 17880 12986 17908 13126
rect 17868 12980 17920 12986
rect 17868 12922 17920 12928
rect 17972 12900 18000 13262
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 18616 12900 18644 18022
rect 17972 12872 18184 12900
rect 17960 12708 18012 12714
rect 17960 12650 18012 12656
rect 18052 12708 18104 12714
rect 18052 12650 18104 12656
rect 17774 12608 17830 12617
rect 17774 12543 17830 12552
rect 17868 12436 17920 12442
rect 17868 12378 17920 12384
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17788 11898 17816 12174
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17696 11750 17816 11778
rect 17590 11727 17646 11736
rect 17604 8294 17632 11727
rect 17684 11688 17736 11694
rect 17682 11656 17684 11665
rect 17736 11656 17738 11665
rect 17682 11591 17738 11600
rect 17682 11248 17738 11257
rect 17682 11183 17684 11192
rect 17736 11183 17738 11192
rect 17684 11154 17736 11160
rect 17684 10464 17736 10470
rect 17684 10406 17736 10412
rect 17696 10266 17724 10406
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17684 10124 17736 10130
rect 17684 10066 17736 10072
rect 17696 9518 17724 10066
rect 17684 9512 17736 9518
rect 17684 9454 17736 9460
rect 17696 8566 17724 9454
rect 17684 8560 17736 8566
rect 17684 8502 17736 8508
rect 17592 8288 17644 8294
rect 17592 8230 17644 8236
rect 17696 7954 17724 8502
rect 17788 8362 17816 11750
rect 17880 10674 17908 12378
rect 17972 11218 18000 12650
rect 18064 12306 18092 12650
rect 18156 12306 18184 12872
rect 18432 12872 18644 12900
rect 18328 12708 18380 12714
rect 18328 12650 18380 12656
rect 18340 12481 18368 12650
rect 18326 12472 18382 12481
rect 18432 12442 18460 12872
rect 18708 12696 18736 18090
rect 18788 17672 18840 17678
rect 18788 17614 18840 17620
rect 18800 16794 18828 17614
rect 18892 17105 18920 19110
rect 18984 17785 19012 19722
rect 18970 17776 19026 17785
rect 18970 17711 19026 17720
rect 18972 17672 19024 17678
rect 18972 17614 19024 17620
rect 18878 17096 18934 17105
rect 18878 17031 18934 17040
rect 18880 16992 18932 16998
rect 18880 16934 18932 16940
rect 18788 16788 18840 16794
rect 18788 16730 18840 16736
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18800 16114 18828 16526
rect 18788 16108 18840 16114
rect 18788 16050 18840 16056
rect 18788 15496 18840 15502
rect 18788 15438 18840 15444
rect 18800 14346 18828 15438
rect 18788 14340 18840 14346
rect 18788 14282 18840 14288
rect 18786 13968 18842 13977
rect 18786 13903 18842 13912
rect 18800 13530 18828 13903
rect 18788 13524 18840 13530
rect 18788 13466 18840 13472
rect 18786 13152 18842 13161
rect 18786 13087 18842 13096
rect 18616 12668 18736 12696
rect 18326 12407 18382 12416
rect 18420 12436 18472 12442
rect 18420 12378 18472 12384
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 18144 12300 18196 12306
rect 18144 12242 18196 12248
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 18512 11008 18564 11014
rect 18512 10950 18564 10956
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 18524 10674 18552 10950
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 18512 10668 18564 10674
rect 18512 10610 18564 10616
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 17868 10532 17920 10538
rect 17868 10474 17920 10480
rect 17880 10062 17908 10474
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17880 9217 17908 9318
rect 17866 9208 17922 9217
rect 17972 9178 18000 10066
rect 18340 10062 18368 10542
rect 18524 10282 18552 10610
rect 18616 10452 18644 12668
rect 18694 12608 18750 12617
rect 18694 12543 18750 12552
rect 18708 10606 18736 12543
rect 18800 11506 18828 13087
rect 18892 13025 18920 16934
rect 18984 13734 19012 17614
rect 19076 16658 19104 22471
rect 19154 22320 19210 22800
rect 19614 22320 19670 22800
rect 20166 22320 20222 22800
rect 20626 22320 20682 22800
rect 21086 22320 21142 22800
rect 21546 22320 21602 22800
rect 22006 22320 22062 22800
rect 22466 22320 22522 22800
rect 19168 18306 19196 22320
rect 19246 20632 19302 20641
rect 19246 20567 19302 20576
rect 19260 20058 19288 20567
rect 19338 20224 19394 20233
rect 19338 20159 19394 20168
rect 19248 20052 19300 20058
rect 19248 19994 19300 20000
rect 19352 19514 19380 20159
rect 19430 19680 19486 19689
rect 19430 19615 19486 19624
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 19340 19236 19392 19242
rect 19340 19178 19392 19184
rect 19246 18456 19302 18465
rect 19352 18426 19380 19178
rect 19444 18970 19472 19615
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 19628 18902 19656 22320
rect 20076 19916 20128 19922
rect 20076 19858 20128 19864
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19904 19417 19932 19654
rect 19890 19408 19946 19417
rect 19890 19343 19946 19352
rect 19708 19168 19760 19174
rect 19708 19110 19760 19116
rect 19892 19168 19944 19174
rect 19892 19110 19944 19116
rect 19616 18896 19668 18902
rect 19616 18838 19668 18844
rect 19246 18391 19248 18400
rect 19300 18391 19302 18400
rect 19340 18420 19392 18426
rect 19248 18362 19300 18368
rect 19340 18362 19392 18368
rect 19616 18420 19668 18426
rect 19616 18362 19668 18368
rect 19168 18278 19288 18306
rect 19156 18216 19208 18222
rect 19156 18158 19208 18164
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 19168 15722 19196 18158
rect 19260 17241 19288 18278
rect 19524 18284 19576 18290
rect 19524 18226 19576 18232
rect 19340 18148 19392 18154
rect 19340 18090 19392 18096
rect 19352 17610 19380 18090
rect 19432 18080 19484 18086
rect 19432 18022 19484 18028
rect 19340 17604 19392 17610
rect 19340 17546 19392 17552
rect 19246 17232 19302 17241
rect 19246 17167 19302 17176
rect 19340 17196 19392 17202
rect 19340 17138 19392 17144
rect 19248 17128 19300 17134
rect 19352 17082 19380 17138
rect 19300 17076 19380 17082
rect 19248 17070 19380 17076
rect 19260 17054 19380 17070
rect 19248 16992 19300 16998
rect 19340 16992 19392 16998
rect 19248 16934 19300 16940
rect 19338 16960 19340 16969
rect 19392 16960 19394 16969
rect 19076 15694 19196 15722
rect 19076 14822 19104 15694
rect 19156 15564 19208 15570
rect 19156 15506 19208 15512
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 19168 14618 19196 15506
rect 19260 15094 19288 16934
rect 19338 16895 19394 16904
rect 19444 15722 19472 18022
rect 19352 15694 19472 15722
rect 19352 15366 19380 15694
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 19340 15360 19392 15366
rect 19340 15302 19392 15308
rect 19444 15162 19472 15506
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 19248 15088 19300 15094
rect 19248 15030 19300 15036
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19156 14612 19208 14618
rect 19156 14554 19208 14560
rect 19246 14512 19302 14521
rect 19352 14498 19380 14962
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19444 14618 19472 14758
rect 19432 14612 19484 14618
rect 19432 14554 19484 14560
rect 19352 14470 19472 14498
rect 19246 14447 19302 14456
rect 19064 14408 19116 14414
rect 19064 14350 19116 14356
rect 19260 14362 19288 14447
rect 19444 14414 19472 14470
rect 19432 14408 19484 14414
rect 18972 13728 19024 13734
rect 18972 13670 19024 13676
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 18878 13016 18934 13025
rect 18878 12951 18934 12960
rect 18984 11540 19012 13330
rect 19076 12102 19104 14350
rect 19260 14334 19380 14362
rect 19432 14350 19484 14356
rect 19248 14272 19300 14278
rect 19248 14214 19300 14220
rect 19260 12696 19288 14214
rect 19352 13274 19380 14334
rect 19444 14074 19472 14350
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19430 13832 19486 13841
rect 19430 13767 19432 13776
rect 19484 13767 19486 13776
rect 19432 13738 19484 13744
rect 19444 13394 19472 13738
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 19352 13246 19472 13274
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19352 13025 19380 13126
rect 19338 13016 19394 13025
rect 19338 12951 19394 12960
rect 19168 12668 19288 12696
rect 19168 12617 19196 12668
rect 19154 12608 19210 12617
rect 19444 12594 19472 13246
rect 19536 12986 19564 18226
rect 19628 17814 19656 18362
rect 19720 18057 19748 19110
rect 19800 18624 19852 18630
rect 19800 18566 19852 18572
rect 19812 18193 19840 18566
rect 19798 18184 19854 18193
rect 19798 18119 19854 18128
rect 19800 18080 19852 18086
rect 19706 18048 19762 18057
rect 19800 18022 19852 18028
rect 19706 17983 19762 17992
rect 19812 17882 19840 18022
rect 19904 17921 19932 19110
rect 19984 18828 20036 18834
rect 19984 18770 20036 18776
rect 19890 17912 19946 17921
rect 19800 17876 19852 17882
rect 19890 17847 19946 17856
rect 19800 17818 19852 17824
rect 19996 17814 20024 18770
rect 19616 17808 19668 17814
rect 19616 17750 19668 17756
rect 19984 17808 20036 17814
rect 19984 17750 20036 17756
rect 19708 17740 19760 17746
rect 19708 17682 19760 17688
rect 19800 17740 19852 17746
rect 19800 17682 19852 17688
rect 19720 16590 19748 17682
rect 19616 16584 19668 16590
rect 19616 16526 19668 16532
rect 19708 16584 19760 16590
rect 19708 16526 19760 16532
rect 19628 16250 19656 16526
rect 19616 16244 19668 16250
rect 19616 16186 19668 16192
rect 19616 15904 19668 15910
rect 19616 15846 19668 15852
rect 19628 15609 19656 15846
rect 19708 15632 19760 15638
rect 19614 15600 19670 15609
rect 19708 15574 19760 15580
rect 19614 15535 19670 15544
rect 19616 15360 19668 15366
rect 19616 15302 19668 15308
rect 19628 14890 19656 15302
rect 19616 14884 19668 14890
rect 19616 14826 19668 14832
rect 19614 14376 19670 14385
rect 19614 14311 19616 14320
rect 19668 14311 19670 14320
rect 19616 14282 19668 14288
rect 19720 14074 19748 15574
rect 19708 14068 19760 14074
rect 19708 14010 19760 14016
rect 19614 13968 19670 13977
rect 19614 13903 19670 13912
rect 19628 13802 19656 13903
rect 19616 13796 19668 13802
rect 19616 13738 19668 13744
rect 19812 13546 19840 17682
rect 19984 17672 20036 17678
rect 19984 17614 20036 17620
rect 19996 16794 20024 17614
rect 19984 16788 20036 16794
rect 19984 16730 20036 16736
rect 20088 16153 20116 19858
rect 20180 19310 20208 22320
rect 20444 19848 20496 19854
rect 20364 19808 20444 19836
rect 20364 19378 20392 19808
rect 20444 19790 20496 19796
rect 20352 19372 20404 19378
rect 20352 19314 20404 19320
rect 20168 19304 20220 19310
rect 20168 19246 20220 19252
rect 20168 19168 20220 19174
rect 20168 19110 20220 19116
rect 20180 18465 20208 19110
rect 20364 18766 20392 19314
rect 20640 19242 20668 22320
rect 20996 19916 21048 19922
rect 20996 19858 21048 19864
rect 20628 19236 20680 19242
rect 20628 19178 20680 19184
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 20352 18760 20404 18766
rect 20916 18737 20944 19110
rect 20352 18702 20404 18708
rect 20902 18728 20958 18737
rect 20166 18456 20222 18465
rect 20166 18391 20222 18400
rect 20364 18358 20392 18702
rect 20902 18663 20958 18672
rect 20352 18352 20404 18358
rect 20352 18294 20404 18300
rect 20168 17740 20220 17746
rect 20168 17682 20220 17688
rect 20180 17338 20208 17682
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20074 16144 20130 16153
rect 20074 16079 20130 16088
rect 20364 15994 20392 18294
rect 20720 18148 20772 18154
rect 20720 18090 20772 18096
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20548 16590 20576 17138
rect 20536 16584 20588 16590
rect 20536 16526 20588 16532
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20180 15966 20392 15994
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 19904 13841 19932 14758
rect 19890 13832 19946 13841
rect 19890 13767 19946 13776
rect 19892 13728 19944 13734
rect 19892 13670 19944 13676
rect 19628 13518 19840 13546
rect 19524 12980 19576 12986
rect 19524 12922 19576 12928
rect 19154 12543 19210 12552
rect 19260 12566 19472 12594
rect 19154 12472 19210 12481
rect 19154 12407 19156 12416
rect 19208 12407 19210 12416
rect 19156 12378 19208 12384
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 19156 11892 19208 11898
rect 19156 11834 19208 11840
rect 18984 11512 19104 11540
rect 18800 11478 18920 11506
rect 18786 11384 18842 11393
rect 18786 11319 18788 11328
rect 18840 11319 18842 11328
rect 18788 11290 18840 11296
rect 18892 11234 18920 11478
rect 18800 11206 18920 11234
rect 18800 11150 18828 11206
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18880 11144 18932 11150
rect 18880 11086 18932 11092
rect 18788 11008 18840 11014
rect 18788 10950 18840 10956
rect 18696 10600 18748 10606
rect 18800 10577 18828 10950
rect 18892 10606 18920 11086
rect 18880 10600 18932 10606
rect 18696 10542 18748 10548
rect 18786 10568 18842 10577
rect 18880 10542 18932 10548
rect 18786 10503 18842 10512
rect 18616 10424 18828 10452
rect 18524 10254 18644 10282
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 18328 10056 18380 10062
rect 18432 10033 18460 10066
rect 18328 9998 18380 10004
rect 18418 10024 18474 10033
rect 18418 9959 18474 9968
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 17866 9143 17922 9152
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 17868 9104 17920 9110
rect 17868 9046 17920 9052
rect 17880 8430 17908 9046
rect 18156 8820 18184 9454
rect 18512 9444 18564 9450
rect 18512 9386 18564 9392
rect 17972 8792 18184 8820
rect 17972 8634 18000 8792
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 18234 8528 18290 8537
rect 18234 8463 18236 8472
rect 18288 8463 18290 8472
rect 18236 8434 18288 8440
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 17776 8356 17828 8362
rect 17776 8298 17828 8304
rect 18236 8288 18288 8294
rect 18236 8230 18288 8236
rect 18420 8288 18472 8294
rect 18420 8230 18472 8236
rect 17776 8084 17828 8090
rect 17776 8026 17828 8032
rect 17868 8084 17920 8090
rect 17868 8026 17920 8032
rect 17788 7954 17816 8026
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 17684 7744 17736 7750
rect 17684 7686 17736 7692
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17604 7002 17632 7346
rect 17592 6996 17644 7002
rect 17592 6938 17644 6944
rect 17592 6724 17644 6730
rect 17592 6666 17644 6672
rect 17604 6633 17632 6666
rect 17590 6624 17646 6633
rect 17590 6559 17646 6568
rect 17592 6248 17644 6254
rect 17592 6190 17644 6196
rect 17604 6089 17632 6190
rect 17590 6080 17646 6089
rect 17590 6015 17646 6024
rect 17590 5400 17646 5409
rect 17590 5335 17646 5344
rect 17604 5030 17632 5335
rect 17592 5024 17644 5030
rect 17592 4966 17644 4972
rect 17592 3936 17644 3942
rect 17592 3878 17644 3884
rect 17500 3664 17552 3670
rect 17500 3606 17552 3612
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 17328 2961 17356 3470
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 17314 2952 17370 2961
rect 17420 2938 17448 3334
rect 17512 3058 17540 3470
rect 17604 3466 17632 3878
rect 17592 3460 17644 3466
rect 17592 3402 17644 3408
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17592 3052 17644 3058
rect 17592 2994 17644 3000
rect 17604 2938 17632 2994
rect 17420 2910 17632 2938
rect 17314 2887 17370 2896
rect 17696 2836 17724 7686
rect 17776 7336 17828 7342
rect 17776 7278 17828 7284
rect 17788 4146 17816 7278
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17788 3233 17816 3878
rect 17774 3224 17830 3233
rect 17774 3159 17830 3168
rect 17774 3088 17830 3097
rect 17774 3023 17830 3032
rect 17604 2808 17724 2836
rect 17236 2604 17356 2632
rect 17222 2544 17278 2553
rect 17328 2514 17356 2604
rect 17222 2479 17224 2488
rect 17276 2479 17278 2488
rect 17316 2508 17368 2514
rect 17224 2450 17276 2456
rect 17316 2450 17368 2456
rect 17604 480 17632 2808
rect 17788 2514 17816 3023
rect 17880 2922 17908 8026
rect 18248 7818 18276 8230
rect 18432 7993 18460 8230
rect 18418 7984 18474 7993
rect 18418 7919 18474 7928
rect 18524 7818 18552 9386
rect 18616 8974 18644 10254
rect 18696 10056 18748 10062
rect 18696 9998 18748 10004
rect 18604 8968 18656 8974
rect 18604 8910 18656 8916
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 18236 7812 18288 7818
rect 18236 7754 18288 7760
rect 18512 7812 18564 7818
rect 18512 7754 18564 7760
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 18524 7342 18552 7754
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 17960 7200 18012 7206
rect 17960 7142 18012 7148
rect 18328 7200 18380 7206
rect 18328 7142 18380 7148
rect 17972 5846 18000 7142
rect 18340 6769 18368 7142
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 18326 6760 18382 6769
rect 18326 6695 18382 6704
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 17960 5840 18012 5846
rect 17960 5782 18012 5788
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 18064 5658 18092 5714
rect 17972 5630 18092 5658
rect 17972 5370 18000 5630
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17960 5092 18012 5098
rect 17960 5034 18012 5040
rect 17972 4282 18000 5034
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 17960 4276 18012 4282
rect 17960 4218 18012 4224
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 17972 3670 18000 4082
rect 18524 3670 18552 6802
rect 17960 3664 18012 3670
rect 18512 3664 18564 3670
rect 18012 3624 18092 3652
rect 17960 3606 18012 3612
rect 17960 3528 18012 3534
rect 18064 3505 18092 3624
rect 18512 3606 18564 3612
rect 17960 3470 18012 3476
rect 18050 3496 18106 3505
rect 17868 2916 17920 2922
rect 17868 2858 17920 2864
rect 17776 2508 17828 2514
rect 17776 2450 17828 2456
rect 17972 1601 18000 3470
rect 18050 3431 18106 3440
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 18616 3097 18644 8570
rect 18708 7585 18736 9998
rect 18800 9489 18828 10424
rect 18892 10130 18920 10542
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 18880 10124 18932 10130
rect 18880 10066 18932 10072
rect 18878 10024 18934 10033
rect 18878 9959 18934 9968
rect 18892 9625 18920 9959
rect 18878 9616 18934 9625
rect 18878 9551 18934 9560
rect 18786 9480 18842 9489
rect 18786 9415 18842 9424
rect 18800 8906 18828 9415
rect 18880 9104 18932 9110
rect 18880 9046 18932 9052
rect 18788 8900 18840 8906
rect 18788 8842 18840 8848
rect 18892 8634 18920 9046
rect 18984 8906 19012 10406
rect 18972 8900 19024 8906
rect 18972 8842 19024 8848
rect 18970 8800 19026 8809
rect 18970 8735 19026 8744
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 18786 8256 18842 8265
rect 18786 8191 18842 8200
rect 18800 7818 18828 8191
rect 18984 8090 19012 8735
rect 18972 8084 19024 8090
rect 18972 8026 19024 8032
rect 18788 7812 18840 7818
rect 18788 7754 18840 7760
rect 18694 7576 18750 7585
rect 18694 7511 18750 7520
rect 18984 7478 19012 8026
rect 19076 7954 19104 11512
rect 19064 7948 19116 7954
rect 19064 7890 19116 7896
rect 18972 7472 19024 7478
rect 18972 7414 19024 7420
rect 18696 7404 18748 7410
rect 18696 7346 18748 7352
rect 18708 5166 18736 7346
rect 18984 7177 19012 7414
rect 19076 7274 19104 7890
rect 19064 7268 19116 7274
rect 19064 7210 19116 7216
rect 18970 7168 19026 7177
rect 18970 7103 19026 7112
rect 18878 6896 18934 6905
rect 18878 6831 18934 6840
rect 18892 6730 18920 6831
rect 18972 6792 19024 6798
rect 18972 6734 19024 6740
rect 18880 6724 18932 6730
rect 18880 6666 18932 6672
rect 18984 6254 19012 6734
rect 18972 6248 19024 6254
rect 18972 6190 19024 6196
rect 18878 5808 18934 5817
rect 18878 5743 18880 5752
rect 18932 5743 18934 5752
rect 18880 5714 18932 5720
rect 18788 5568 18840 5574
rect 18788 5510 18840 5516
rect 18800 5409 18828 5510
rect 18786 5400 18842 5409
rect 18786 5335 18842 5344
rect 18880 5296 18932 5302
rect 18880 5238 18932 5244
rect 18696 5160 18748 5166
rect 18696 5102 18748 5108
rect 18708 4758 18736 5102
rect 18696 4752 18748 4758
rect 18696 4694 18748 4700
rect 18708 4214 18736 4694
rect 18696 4208 18748 4214
rect 18696 4150 18748 4156
rect 18708 3534 18736 4150
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18800 3641 18828 3878
rect 18892 3777 18920 5238
rect 18984 5098 19012 6190
rect 19076 5386 19104 7210
rect 19168 6746 19196 11834
rect 19260 9654 19288 12566
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19352 11354 19380 12242
rect 19628 11898 19656 13518
rect 19708 13388 19760 13394
rect 19904 13376 19932 13670
rect 19708 13330 19760 13336
rect 19812 13348 19932 13376
rect 19616 11892 19668 11898
rect 19616 11834 19668 11840
rect 19616 11620 19668 11626
rect 19720 11608 19748 13330
rect 19812 12442 19840 13348
rect 19892 13184 19944 13190
rect 19890 13152 19892 13161
rect 19944 13152 19946 13161
rect 19890 13087 19946 13096
rect 19890 12880 19946 12889
rect 19890 12815 19946 12824
rect 19904 12617 19932 12815
rect 19890 12608 19946 12617
rect 19890 12543 19946 12552
rect 19800 12436 19852 12442
rect 19800 12378 19852 12384
rect 19800 11824 19852 11830
rect 19798 11792 19800 11801
rect 19852 11792 19854 11801
rect 19798 11727 19854 11736
rect 19668 11580 19748 11608
rect 19616 11562 19668 11568
rect 19812 11558 19840 11727
rect 19800 11552 19852 11558
rect 19800 11494 19852 11500
rect 19340 11348 19392 11354
rect 19340 11290 19392 11296
rect 19800 10260 19852 10266
rect 19800 10202 19852 10208
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 19338 10024 19394 10033
rect 19338 9959 19394 9968
rect 19352 9926 19380 9959
rect 19340 9920 19392 9926
rect 19340 9862 19392 9868
rect 19248 9648 19300 9654
rect 19248 9590 19300 9596
rect 19432 9512 19484 9518
rect 19432 9454 19484 9460
rect 19338 9344 19394 9353
rect 19338 9279 19394 9288
rect 19248 8968 19300 8974
rect 19246 8936 19248 8945
rect 19300 8936 19302 8945
rect 19246 8871 19302 8880
rect 19352 8809 19380 9279
rect 19338 8800 19394 8809
rect 19338 8735 19394 8744
rect 19444 8634 19472 9454
rect 19536 9382 19564 10066
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19708 9376 19760 9382
rect 19708 9318 19760 9324
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 19430 8528 19486 8537
rect 19340 8492 19392 8498
rect 19430 8463 19486 8472
rect 19340 8434 19392 8440
rect 19352 7886 19380 8434
rect 19444 8430 19472 8463
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19432 7744 19484 7750
rect 19432 7686 19484 7692
rect 19444 7342 19472 7686
rect 19248 7336 19300 7342
rect 19248 7278 19300 7284
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 19260 6866 19288 7278
rect 19444 7002 19472 7278
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19248 6860 19300 6866
rect 19248 6802 19300 6808
rect 19168 6718 19472 6746
rect 19156 6656 19208 6662
rect 19208 6616 19288 6644
rect 19156 6598 19208 6604
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 19168 5574 19196 6394
rect 19156 5568 19208 5574
rect 19156 5510 19208 5516
rect 19076 5358 19196 5386
rect 18972 5092 19024 5098
rect 18972 5034 19024 5040
rect 19064 4548 19116 4554
rect 19064 4490 19116 4496
rect 18970 4040 19026 4049
rect 18970 3975 19026 3984
rect 18878 3768 18934 3777
rect 18878 3703 18934 3712
rect 18786 3632 18842 3641
rect 18786 3567 18842 3576
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 18984 3233 19012 3975
rect 19076 3738 19104 4490
rect 19064 3732 19116 3738
rect 19064 3674 19116 3680
rect 18970 3224 19026 3233
rect 18970 3159 19026 3168
rect 18326 3088 18382 3097
rect 18326 3023 18382 3032
rect 18602 3088 18658 3097
rect 18602 3023 18658 3032
rect 18340 2990 18368 3023
rect 18328 2984 18380 2990
rect 19076 2972 19104 3674
rect 18328 2926 18380 2932
rect 18800 2944 19104 2972
rect 18512 2916 18564 2922
rect 18512 2858 18564 2864
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 18050 1864 18106 1873
rect 18050 1799 18106 1808
rect 17958 1592 18014 1601
rect 17958 1527 18014 1536
rect 17960 1352 18012 1358
rect 17960 1294 18012 1300
rect 17972 1193 18000 1294
rect 17958 1184 18014 1193
rect 17958 1119 18014 1128
rect 18064 480 18092 1799
rect 18524 480 18552 2858
rect 18800 2417 18828 2944
rect 18878 2816 18934 2825
rect 18878 2751 18934 2760
rect 18786 2408 18842 2417
rect 18786 2343 18842 2352
rect 3974 232 4030 241
rect 3974 167 4030 176
rect 4158 0 4214 480
rect 4618 0 4674 480
rect 5078 0 5134 480
rect 5538 0 5594 480
rect 5998 0 6054 480
rect 6458 0 6514 480
rect 6826 0 6882 480
rect 7286 0 7342 480
rect 7746 0 7802 480
rect 8206 0 8262 480
rect 8666 0 8722 480
rect 9126 0 9182 480
rect 9586 0 9642 480
rect 9954 0 10010 480
rect 10414 0 10470 480
rect 10874 0 10930 480
rect 11334 0 11390 480
rect 11794 0 11850 480
rect 12254 0 12310 480
rect 12714 0 12770 480
rect 13174 0 13230 480
rect 13542 0 13598 480
rect 14002 0 14058 480
rect 14462 0 14518 480
rect 14922 0 14978 480
rect 15382 0 15438 480
rect 15842 0 15898 480
rect 16302 0 16358 480
rect 16670 0 16726 480
rect 17130 0 17186 480
rect 17590 0 17646 480
rect 18050 0 18106 480
rect 18510 0 18566 480
rect 18892 241 18920 2751
rect 19064 2644 19116 2650
rect 19064 2586 19116 2592
rect 19076 2553 19104 2586
rect 19062 2544 19118 2553
rect 19062 2479 19118 2488
rect 18972 2032 19024 2038
rect 18972 1974 19024 1980
rect 18984 480 19012 1974
rect 19168 649 19196 5358
rect 19260 4128 19288 6616
rect 19340 6180 19392 6186
rect 19340 6122 19392 6128
rect 19352 5710 19380 6122
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19352 5370 19380 5646
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19444 5250 19472 6718
rect 19352 5222 19472 5250
rect 19352 4554 19380 5222
rect 19432 5160 19484 5166
rect 19432 5102 19484 5108
rect 19444 4826 19472 5102
rect 19432 4820 19484 4826
rect 19432 4762 19484 4768
rect 19340 4548 19392 4554
rect 19340 4490 19392 4496
rect 19444 4282 19472 4762
rect 19432 4276 19484 4282
rect 19432 4218 19484 4224
rect 19260 4100 19472 4128
rect 19340 3664 19392 3670
rect 19338 3632 19340 3641
rect 19392 3632 19394 3641
rect 19338 3567 19394 3576
rect 19340 3528 19392 3534
rect 19246 3496 19302 3505
rect 19340 3470 19392 3476
rect 19246 3431 19302 3440
rect 19260 2990 19288 3431
rect 19352 3398 19380 3470
rect 19444 3398 19472 4100
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19536 3210 19564 9318
rect 19720 9178 19748 9318
rect 19708 9172 19760 9178
rect 19708 9114 19760 9120
rect 19708 9036 19760 9042
rect 19708 8978 19760 8984
rect 19616 8968 19668 8974
rect 19616 8910 19668 8916
rect 19628 8498 19656 8910
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 19720 8362 19748 8978
rect 19812 8430 19840 10202
rect 19800 8424 19852 8430
rect 19800 8366 19852 8372
rect 19708 8356 19760 8362
rect 19708 8298 19760 8304
rect 19708 7948 19760 7954
rect 19708 7890 19760 7896
rect 19614 4312 19670 4321
rect 19614 4247 19616 4256
rect 19668 4247 19670 4256
rect 19616 4218 19668 4224
rect 19628 4010 19656 4218
rect 19616 4004 19668 4010
rect 19616 3946 19668 3952
rect 19616 3596 19668 3602
rect 19616 3538 19668 3544
rect 19628 3233 19656 3538
rect 19720 3534 19748 7890
rect 19812 7886 19840 8366
rect 19904 7886 19932 12543
rect 19996 9042 20024 15846
rect 20076 15496 20128 15502
rect 20076 15438 20128 15444
rect 20088 15162 20116 15438
rect 20076 15156 20128 15162
rect 20076 15098 20128 15104
rect 20180 14906 20208 15966
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 20352 15904 20404 15910
rect 20352 15846 20404 15852
rect 20088 14878 20208 14906
rect 20088 10266 20116 14878
rect 20168 14816 20220 14822
rect 20166 14784 20168 14793
rect 20220 14784 20222 14793
rect 20166 14719 20222 14728
rect 20168 14476 20220 14482
rect 20168 14418 20220 14424
rect 20180 11218 20208 14418
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 20076 9376 20128 9382
rect 20076 9318 20128 9324
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 19984 9036 20036 9042
rect 19984 8978 20036 8984
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 19996 8294 20024 8774
rect 19984 8288 20036 8294
rect 19984 8230 20036 8236
rect 19800 7880 19852 7886
rect 19800 7822 19852 7828
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 19984 6928 20036 6934
rect 19984 6870 20036 6876
rect 19892 5772 19944 5778
rect 19892 5714 19944 5720
rect 19800 5024 19852 5030
rect 19800 4966 19852 4972
rect 19812 3534 19840 4966
rect 19904 4826 19932 5714
rect 19892 4820 19944 4826
rect 19892 4762 19944 4768
rect 19996 4706 20024 6870
rect 20088 6066 20116 9318
rect 20180 8090 20208 9318
rect 20272 8650 20300 15846
rect 20364 15337 20392 15846
rect 20350 15328 20406 15337
rect 20350 15263 20406 15272
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 20364 12646 20392 14350
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 20364 9586 20392 12582
rect 20456 10538 20484 16050
rect 20548 12306 20576 16526
rect 20628 16040 20680 16046
rect 20628 15982 20680 15988
rect 20536 12300 20588 12306
rect 20536 12242 20588 12248
rect 20536 11620 20588 11626
rect 20536 11562 20588 11568
rect 20444 10532 20496 10538
rect 20444 10474 20496 10480
rect 20456 10266 20484 10474
rect 20444 10260 20496 10266
rect 20444 10202 20496 10208
rect 20352 9580 20404 9586
rect 20352 9522 20404 9528
rect 20364 8974 20392 9522
rect 20352 8968 20404 8974
rect 20548 8956 20576 11562
rect 20640 11286 20668 15982
rect 20732 11694 20760 18090
rect 20904 17536 20956 17542
rect 20904 17478 20956 17484
rect 20916 17202 20944 17478
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 20812 17060 20864 17066
rect 20812 17002 20864 17008
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20628 11280 20680 11286
rect 20628 11222 20680 11228
rect 20732 11234 20760 11494
rect 20824 11354 20852 17002
rect 20904 16652 20956 16658
rect 20904 16594 20956 16600
rect 20916 16182 20944 16594
rect 20904 16176 20956 16182
rect 20904 16118 20956 16124
rect 20904 13728 20956 13734
rect 20904 13670 20956 13676
rect 20916 13569 20944 13670
rect 20902 13560 20958 13569
rect 20902 13495 20958 13504
rect 20904 13456 20956 13462
rect 20904 13398 20956 13404
rect 20916 12986 20944 13398
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 20640 10810 20668 11222
rect 20732 11206 20852 11234
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 20720 9512 20772 9518
rect 20720 9454 20772 9460
rect 20732 9110 20760 9454
rect 20720 9104 20772 9110
rect 20720 9046 20772 9052
rect 20548 8928 20760 8956
rect 20352 8910 20404 8916
rect 20272 8622 20668 8650
rect 20260 8560 20312 8566
rect 20260 8502 20312 8508
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20088 6038 20208 6066
rect 19904 4678 20024 4706
rect 19904 3942 19932 4678
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 19984 4548 20036 4554
rect 19984 4490 20036 4496
rect 19996 4282 20024 4490
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 19892 3936 19944 3942
rect 19892 3878 19944 3884
rect 20088 3738 20116 4558
rect 20076 3732 20128 3738
rect 20076 3674 20128 3680
rect 19708 3528 19760 3534
rect 19708 3470 19760 3476
rect 19800 3528 19852 3534
rect 19800 3470 19852 3476
rect 19708 3392 19760 3398
rect 19708 3334 19760 3340
rect 19352 3182 19564 3210
rect 19614 3224 19670 3233
rect 19352 3058 19380 3182
rect 19614 3159 19670 3168
rect 19524 3120 19576 3126
rect 19524 3062 19576 3068
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19248 2984 19300 2990
rect 19248 2926 19300 2932
rect 19352 2446 19380 2994
rect 19536 2650 19564 3062
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 19720 2530 19748 3334
rect 19890 3224 19946 3233
rect 19890 3159 19946 3168
rect 19798 3088 19854 3097
rect 19904 3058 19932 3159
rect 19798 3023 19854 3032
rect 19892 3052 19944 3058
rect 19812 2990 19840 3023
rect 19892 2994 19944 3000
rect 19800 2984 19852 2990
rect 19800 2926 19852 2932
rect 19444 2502 19748 2530
rect 19340 2440 19392 2446
rect 19340 2382 19392 2388
rect 19154 640 19210 649
rect 19154 575 19210 584
rect 19444 480 19472 2502
rect 20180 2106 20208 6038
rect 20272 5522 20300 8502
rect 20536 8424 20588 8430
rect 20536 8366 20588 8372
rect 20444 8356 20496 8362
rect 20444 8298 20496 8304
rect 20352 6860 20404 6866
rect 20352 6802 20404 6808
rect 20364 6458 20392 6802
rect 20456 6730 20484 8298
rect 20548 7546 20576 8366
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20444 6724 20496 6730
rect 20444 6666 20496 6672
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 20364 5710 20392 6394
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 20272 5494 20392 5522
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 20272 4758 20300 5306
rect 20260 4752 20312 4758
rect 20260 4694 20312 4700
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 20272 4078 20300 4558
rect 20260 4072 20312 4078
rect 20260 4014 20312 4020
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 20272 2990 20300 3878
rect 20260 2984 20312 2990
rect 20260 2926 20312 2932
rect 20364 2446 20392 5494
rect 20444 4480 20496 4486
rect 20444 4422 20496 4428
rect 20456 3466 20484 4422
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 20548 3534 20576 4082
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20444 3460 20496 3466
rect 20444 3402 20496 3408
rect 20640 3194 20668 8622
rect 20732 7857 20760 8928
rect 20718 7848 20774 7857
rect 20718 7783 20774 7792
rect 20720 5908 20772 5914
rect 20720 5850 20772 5856
rect 20628 3188 20680 3194
rect 20628 3130 20680 3136
rect 20536 3120 20588 3126
rect 20536 3062 20588 3068
rect 20442 2680 20498 2689
rect 20442 2615 20444 2624
rect 20496 2615 20498 2624
rect 20444 2586 20496 2592
rect 20548 2582 20576 3062
rect 20536 2576 20588 2582
rect 20536 2518 20588 2524
rect 20352 2440 20404 2446
rect 20352 2382 20404 2388
rect 20260 2372 20312 2378
rect 20260 2314 20312 2320
rect 20168 2100 20220 2106
rect 20168 2042 20220 2048
rect 19800 604 19852 610
rect 19800 546 19852 552
rect 19812 480 19840 546
rect 20272 480 20300 2314
rect 20732 480 20760 5850
rect 20824 4457 20852 11206
rect 21008 8090 21036 19858
rect 21100 15065 21128 22320
rect 21272 19304 21324 19310
rect 21272 19246 21324 19252
rect 21180 16176 21232 16182
rect 21180 16118 21232 16124
rect 21086 15056 21142 15065
rect 21086 14991 21142 15000
rect 21088 13864 21140 13870
rect 21088 13806 21140 13812
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 21100 6322 21128 13806
rect 21192 13297 21220 16118
rect 21178 13288 21234 13297
rect 21178 13223 21234 13232
rect 21192 9178 21220 13223
rect 21284 11082 21312 19246
rect 21560 18698 21588 22320
rect 21548 18692 21600 18698
rect 21548 18634 21600 18640
rect 22020 18426 22048 22320
rect 22008 18420 22060 18426
rect 22008 18362 22060 18368
rect 21454 17368 21510 17377
rect 21454 17303 21510 17312
rect 21364 16720 21416 16726
rect 21364 16662 21416 16668
rect 21376 15706 21404 16662
rect 21364 15700 21416 15706
rect 21364 15642 21416 15648
rect 21362 13968 21418 13977
rect 21362 13903 21418 13912
rect 21376 11393 21404 13903
rect 21468 11898 21496 17303
rect 21456 11892 21508 11898
rect 21456 11834 21508 11840
rect 21362 11384 21418 11393
rect 21362 11319 21418 11328
rect 21272 11076 21324 11082
rect 21272 11018 21324 11024
rect 22480 10198 22508 22320
rect 22468 10192 22520 10198
rect 22468 10134 22520 10140
rect 21180 9172 21232 9178
rect 21180 9114 21232 9120
rect 21364 8288 21416 8294
rect 21364 8230 21416 8236
rect 21272 6724 21324 6730
rect 21272 6666 21324 6672
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 20996 6112 21048 6118
rect 20996 6054 21048 6060
rect 20810 4448 20866 4457
rect 20810 4383 20866 4392
rect 20812 3664 20864 3670
rect 20812 3606 20864 3612
rect 20824 3505 20852 3606
rect 20810 3496 20866 3505
rect 20810 3431 20866 3440
rect 21008 610 21036 6054
rect 21180 3392 21232 3398
rect 21180 3334 21232 3340
rect 20996 604 21048 610
rect 20996 546 21048 552
rect 21192 480 21220 3334
rect 21284 1601 21312 6666
rect 21270 1592 21326 1601
rect 21270 1527 21326 1536
rect 21376 1193 21404 8230
rect 21640 3460 21692 3466
rect 21640 3402 21692 3408
rect 21362 1184 21418 1193
rect 21362 1119 21418 1128
rect 21652 480 21680 3402
rect 22100 2848 22152 2854
rect 22100 2790 22152 2796
rect 22112 480 22140 2790
rect 22560 2304 22612 2310
rect 22560 2246 22612 2252
rect 22572 480 22600 2246
rect 18878 232 18934 241
rect 18878 167 18934 176
rect 18970 0 19026 480
rect 19430 0 19486 480
rect 19798 0 19854 480
rect 20258 0 20314 480
rect 20718 0 20774 480
rect 21178 0 21234 480
rect 21638 0 21694 480
rect 22098 0 22154 480
rect 22558 0 22614 480
<< via2 >>
rect 3238 22480 3294 22536
rect 1766 19624 1822 19680
rect 1582 18944 1638 19000
rect 1674 18400 1730 18456
rect 1674 18264 1730 18320
rect 1582 17720 1638 17776
rect 1490 16768 1546 16824
rect 1674 17312 1730 17368
rect 3054 22072 3110 22128
rect 2962 21528 3018 21584
rect 2870 21120 2926 21176
rect 2778 20576 2834 20632
rect 1766 15544 1822 15600
rect 2134 17312 2190 17368
rect 2318 17584 2374 17640
rect 2502 15972 2558 16008
rect 2502 15952 2504 15972
rect 2504 15952 2556 15972
rect 2556 15952 2558 15972
rect 570 3304 626 3360
rect 2410 15272 2466 15328
rect 2778 19216 2834 19272
rect 3146 20168 3202 20224
rect 2870 18808 2926 18864
rect 3054 18164 3056 18184
rect 3056 18164 3108 18184
rect 3108 18164 3110 18184
rect 3054 18128 3110 18164
rect 19062 22480 19118 22536
rect 3606 18692 3662 18728
rect 3606 18672 3608 18692
rect 3608 18672 3660 18692
rect 3660 18672 3662 18692
rect 3974 19216 4030 19272
rect 3790 19080 3846 19136
rect 2778 17176 2834 17232
rect 2962 17060 3018 17096
rect 2962 17040 2964 17060
rect 2964 17040 3016 17060
rect 3016 17040 3018 17060
rect 2686 14592 2742 14648
rect 2778 14456 2834 14512
rect 2318 3032 2374 3088
rect 3422 17312 3478 17368
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4250 18672 4306 18728
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4526 18148 4582 18184
rect 4526 18128 4528 18148
rect 4528 18128 4580 18148
rect 4580 18128 4582 18148
rect 3974 17584 4030 17640
rect 4986 19216 5042 19272
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 3422 16360 3478 16416
rect 3330 16088 3386 16144
rect 3974 15816 4030 15872
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 5630 18944 5686 19000
rect 5630 18536 5686 18592
rect 5630 16496 5686 16552
rect 4066 15408 4122 15464
rect 4250 15272 4306 15328
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 3330 13504 3386 13560
rect 2686 7384 2742 7440
rect 2778 4392 2834 4448
rect 3606 13796 3662 13832
rect 3606 13776 3608 13796
rect 3608 13776 3660 13796
rect 3660 13776 3662 13796
rect 3514 11736 3570 11792
rect 4066 14864 4122 14920
rect 4066 13932 4122 13968
rect 4066 13912 4068 13932
rect 4068 13912 4120 13932
rect 4120 13912 4122 13932
rect 3974 12552 4030 12608
rect 4618 14456 4674 14512
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4250 12980 4306 13016
rect 4250 12960 4252 12980
rect 4252 12960 4304 12980
rect 4304 12960 4306 12980
rect 4710 12552 4766 12608
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4250 11464 4306 11520
rect 3882 11328 3938 11384
rect 3882 9696 3938 9752
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4066 8744 4122 8800
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 3054 3440 3110 3496
rect 1858 2488 1914 2544
rect 4066 8200 4122 8256
rect 3974 7792 4030 7848
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 5262 12824 5318 12880
rect 5262 12552 5318 12608
rect 4066 7248 4122 7304
rect 4618 7248 4674 7304
rect 4066 5888 4122 5944
rect 5170 11192 5226 11248
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4066 4936 4122 4992
rect 4066 3984 4122 4040
rect 3698 3848 3754 3904
rect 3238 2080 3294 2136
rect 3238 584 3294 640
rect 4066 3032 4122 3088
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4894 6996 4950 7032
rect 4894 6976 4896 6996
rect 4896 6976 4948 6996
rect 4948 6976 4950 6996
rect 5814 15952 5870 16008
rect 5538 14476 5594 14512
rect 5538 14456 5540 14476
rect 5540 14456 5592 14476
rect 5592 14456 5594 14476
rect 5814 14456 5870 14512
rect 5722 13368 5778 13424
rect 5446 12724 5448 12744
rect 5448 12724 5500 12744
rect 5500 12724 5502 12744
rect 5446 12688 5502 12724
rect 5906 12960 5962 13016
rect 5354 8472 5410 8528
rect 5078 7248 5134 7304
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 4250 1128 4306 1184
rect 5446 4664 5502 4720
rect 6826 18264 6882 18320
rect 6734 18128 6790 18184
rect 6550 17720 6606 17776
rect 6090 15952 6146 16008
rect 6090 15272 6146 15328
rect 6090 9968 6146 10024
rect 5998 8472 6054 8528
rect 5906 3576 5962 3632
rect 5262 1536 5318 1592
rect 6366 12688 6422 12744
rect 6366 9036 6422 9072
rect 6366 9016 6368 9036
rect 6368 9016 6420 9036
rect 6420 9016 6422 9036
rect 6366 8608 6422 8664
rect 6090 6996 6146 7032
rect 6090 6976 6092 6996
rect 6092 6976 6144 6996
rect 6144 6976 6146 6996
rect 6090 6740 6092 6760
rect 6092 6740 6144 6760
rect 6144 6740 6146 6760
rect 6090 6704 6146 6740
rect 6734 16652 6790 16688
rect 7102 17584 7158 17640
rect 6734 16632 6736 16652
rect 6736 16632 6788 16652
rect 6788 16632 6790 16652
rect 6734 16224 6790 16280
rect 6642 14320 6698 14376
rect 6918 14612 6974 14648
rect 6918 14592 6920 14612
rect 6920 14592 6972 14612
rect 6972 14592 6974 14612
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 7286 19116 7288 19136
rect 7288 19116 7340 19136
rect 7340 19116 7342 19136
rect 7286 19080 7342 19116
rect 6550 11872 6606 11928
rect 6642 10648 6698 10704
rect 6550 8744 6606 8800
rect 6550 8472 6606 8528
rect 6550 6296 6606 6352
rect 7470 19488 7526 19544
rect 7470 18672 7526 18728
rect 7470 18028 7472 18048
rect 7472 18028 7524 18048
rect 7524 18028 7526 18048
rect 7470 17992 7526 18028
rect 7654 18672 7710 18728
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 8390 19080 8446 19136
rect 8390 18536 8446 18592
rect 8390 18264 8446 18320
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 8298 17584 8354 17640
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 8114 16088 8170 16144
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7930 15136 7986 15192
rect 7654 14900 7656 14920
rect 7656 14900 7708 14920
rect 7708 14900 7710 14920
rect 7654 14864 7710 14900
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 7562 14456 7618 14512
rect 7838 14476 7894 14512
rect 7838 14456 7840 14476
rect 7840 14456 7892 14476
rect 7892 14456 7894 14476
rect 7470 13776 7526 13832
rect 8390 15408 8446 15464
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7562 12960 7618 13016
rect 7470 8744 7526 8800
rect 6734 3304 6790 3360
rect 7194 5788 7196 5808
rect 7196 5788 7248 5808
rect 7248 5788 7250 5808
rect 7194 5752 7250 5788
rect 7654 9968 7710 10024
rect 7102 3304 7158 3360
rect 9034 18808 9090 18864
rect 9218 17448 9274 17504
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7930 12144 7986 12200
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 8298 12588 8300 12608
rect 8300 12588 8352 12608
rect 8352 12588 8354 12608
rect 8298 12552 8354 12588
rect 8390 12280 8446 12336
rect 8114 10548 8116 10568
rect 8116 10548 8168 10568
rect 8168 10548 8170 10568
rect 8114 10512 8170 10548
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 8758 11736 8814 11792
rect 8758 11464 8814 11520
rect 8574 9968 8630 10024
rect 8390 7384 8446 7440
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 8206 4800 8262 4856
rect 8390 5072 8446 5128
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 9034 15952 9090 16008
rect 8942 13096 8998 13152
rect 9218 15272 9274 15328
rect 9494 18028 9496 18048
rect 9496 18028 9548 18048
rect 9548 18028 9550 18048
rect 9494 17992 9550 18028
rect 9402 17312 9458 17368
rect 9218 15000 9274 15056
rect 9126 14048 9182 14104
rect 9218 12416 9274 12472
rect 9310 12144 9366 12200
rect 8850 10648 8906 10704
rect 8850 8744 8906 8800
rect 8666 8084 8722 8120
rect 8666 8064 8668 8084
rect 8668 8064 8720 8084
rect 8720 8064 8722 8084
rect 8758 6740 8760 6760
rect 8760 6740 8812 6760
rect 8812 6740 8814 6760
rect 8758 6704 8814 6740
rect 9310 10376 9366 10432
rect 9126 8880 9182 8936
rect 9218 6840 9274 6896
rect 10046 19080 10102 19136
rect 10322 19488 10378 19544
rect 10230 19116 10232 19136
rect 10232 19116 10284 19136
rect 10284 19116 10286 19136
rect 10230 19080 10286 19116
rect 10322 18808 10378 18864
rect 10230 18400 10286 18456
rect 10138 18128 10194 18184
rect 9586 15680 9642 15736
rect 9770 15272 9826 15328
rect 9586 13096 9642 13152
rect 9678 12008 9734 12064
rect 9586 10784 9642 10840
rect 9770 10104 9826 10160
rect 9586 6840 9642 6896
rect 9034 2916 9090 2952
rect 9034 2896 9036 2916
rect 9036 2896 9088 2916
rect 9088 2896 9090 2916
rect 8482 1944 8538 2000
rect 9862 8608 9918 8664
rect 9862 8508 9864 8528
rect 9864 8508 9916 8528
rect 9916 8508 9918 8528
rect 9862 8472 9918 8508
rect 9862 8372 9864 8392
rect 9864 8372 9916 8392
rect 9916 8372 9918 8392
rect 9862 8336 9918 8372
rect 9862 8236 9864 8256
rect 9864 8236 9916 8256
rect 9916 8236 9918 8256
rect 9862 8200 9918 8236
rect 9862 8064 9918 8120
rect 10506 15816 10562 15872
rect 9862 6568 9918 6624
rect 9218 3440 9274 3496
rect 9862 4936 9918 4992
rect 9678 3576 9734 3632
rect 10506 15136 10562 15192
rect 10322 12960 10378 13016
rect 10782 19352 10838 19408
rect 10414 12824 10470 12880
rect 10322 12688 10378 12744
rect 10230 10104 10286 10160
rect 10414 10648 10470 10704
rect 10414 9696 10470 9752
rect 10046 6024 10102 6080
rect 10506 8880 10562 8936
rect 10966 16632 11022 16688
rect 10966 16088 11022 16144
rect 10966 15136 11022 15192
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 11242 19080 11298 19136
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 11702 19080 11758 19136
rect 11518 17040 11574 17096
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11702 16360 11758 16416
rect 11610 14864 11666 14920
rect 11150 14764 11152 14784
rect 11152 14764 11204 14784
rect 11204 14764 11206 14784
rect 11150 14728 11206 14764
rect 11334 14728 11390 14784
rect 11886 16496 11942 16552
rect 11886 16224 11942 16280
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11794 14184 11850 14240
rect 11702 14048 11758 14104
rect 11610 13504 11666 13560
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11702 12688 11758 12744
rect 11518 12280 11574 12336
rect 10690 10240 10746 10296
rect 10874 10240 10930 10296
rect 11058 10376 11114 10432
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11334 11736 11390 11792
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11058 9424 11114 9480
rect 11242 9288 11298 9344
rect 10690 8336 10746 8392
rect 10598 7928 10654 7984
rect 10322 6704 10378 6760
rect 10322 4392 10378 4448
rect 10506 4140 10562 4176
rect 10506 4120 10508 4140
rect 10508 4120 10560 4140
rect 10560 4120 10562 4140
rect 10322 3984 10378 4040
rect 10690 6704 10746 6760
rect 9954 3032 10010 3088
rect 10506 3476 10508 3496
rect 10508 3476 10560 3496
rect 10560 3476 10562 3496
rect 10506 3440 10562 3476
rect 9678 2352 9734 2408
rect 10230 2760 10286 2816
rect 10414 2624 10470 2680
rect 10138 2488 10194 2544
rect 10966 7792 11022 7848
rect 10966 6568 11022 6624
rect 10966 6060 10968 6080
rect 10968 6060 11020 6080
rect 11020 6060 11022 6080
rect 10966 6024 11022 6060
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 12254 19352 12310 19408
rect 12162 18944 12218 19000
rect 12438 18264 12494 18320
rect 12714 19216 12770 19272
rect 12806 18536 12862 18592
rect 12162 17176 12218 17232
rect 12346 17584 12402 17640
rect 12530 17856 12586 17912
rect 12530 17448 12586 17504
rect 12806 18128 12862 18184
rect 12990 19216 13046 19272
rect 13082 18672 13138 18728
rect 13358 19216 13414 19272
rect 12530 16532 12532 16552
rect 12532 16532 12584 16552
rect 12584 16532 12586 16552
rect 12530 16496 12586 16532
rect 12714 16496 12770 16552
rect 12254 15816 12310 15872
rect 12530 15408 12586 15464
rect 12438 15308 12440 15328
rect 12440 15308 12492 15328
rect 12492 15308 12494 15328
rect 12438 15272 12494 15308
rect 12346 14864 12402 14920
rect 12254 13640 12310 13696
rect 12714 15156 12770 15192
rect 12714 15136 12716 15156
rect 12716 15136 12768 15156
rect 12768 15136 12770 15156
rect 12714 14864 12770 14920
rect 12254 12824 12310 12880
rect 11886 12144 11942 12200
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 11518 6296 11574 6352
rect 11150 6024 11206 6080
rect 11150 5752 11206 5808
rect 11058 5616 11114 5672
rect 10874 5072 10930 5128
rect 10782 3848 10838 3904
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 11058 4392 11114 4448
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 11150 3984 11206 4040
rect 11518 3576 11574 3632
rect 11794 6432 11850 6488
rect 11794 5652 11796 5672
rect 11796 5652 11848 5672
rect 11848 5652 11850 5672
rect 11794 5616 11850 5652
rect 11702 5344 11758 5400
rect 11702 5072 11758 5128
rect 12070 12144 12126 12200
rect 12070 11736 12126 11792
rect 12254 11736 12310 11792
rect 12254 10376 12310 10432
rect 12070 9016 12126 9072
rect 11978 4800 12034 4856
rect 11978 4428 11980 4448
rect 11980 4428 12032 4448
rect 12032 4428 12034 4448
rect 11978 4392 12034 4428
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 12806 12960 12862 13016
rect 13450 17992 13506 18048
rect 13450 17448 13506 17504
rect 13542 17312 13598 17368
rect 13266 16652 13322 16688
rect 13450 16768 13506 16824
rect 13266 16632 13268 16652
rect 13268 16632 13320 16652
rect 13320 16632 13322 16652
rect 14922 20304 14978 20360
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 13726 19080 13782 19136
rect 13726 17992 13782 18048
rect 12990 14184 13046 14240
rect 13082 13232 13138 13288
rect 12714 12008 12770 12064
rect 12254 8900 12310 8936
rect 12254 8880 12256 8900
rect 12256 8880 12308 8900
rect 12308 8880 12310 8900
rect 12438 8900 12494 8936
rect 12438 8880 12440 8900
rect 12440 8880 12492 8900
rect 12492 8880 12494 8900
rect 12438 8744 12494 8800
rect 12622 10784 12678 10840
rect 12162 7112 12218 7168
rect 12806 9832 12862 9888
rect 12346 6180 12402 6216
rect 12346 6160 12348 6180
rect 12348 6160 12400 6180
rect 12400 6160 12402 6180
rect 12346 6024 12402 6080
rect 12530 5616 12586 5672
rect 12530 5208 12586 5264
rect 12530 5072 12586 5128
rect 12346 4800 12402 4856
rect 12346 4256 12402 4312
rect 12438 4120 12494 4176
rect 12530 3712 12586 3768
rect 12346 2896 12402 2952
rect 13266 14184 13322 14240
rect 13174 12824 13230 12880
rect 13634 15700 13690 15736
rect 13634 15680 13636 15700
rect 13636 15680 13688 15700
rect 13688 15680 13690 15700
rect 13910 17856 13966 17912
rect 13818 16224 13874 16280
rect 14278 19488 14334 19544
rect 14370 19352 14426 19408
rect 14002 16360 14058 16416
rect 13910 15544 13966 15600
rect 13542 14728 13598 14784
rect 13726 14220 13728 14240
rect 13728 14220 13780 14240
rect 13780 14220 13782 14240
rect 13726 14184 13782 14220
rect 13910 14048 13966 14104
rect 13358 13268 13360 13288
rect 13360 13268 13412 13288
rect 13412 13268 13414 13288
rect 13358 13232 13414 13268
rect 13542 12688 13598 12744
rect 13726 13232 13782 13288
rect 13082 12008 13138 12064
rect 13450 12008 13506 12064
rect 12990 10784 13046 10840
rect 12990 10648 13046 10704
rect 13266 11464 13322 11520
rect 13082 8200 13138 8256
rect 12990 6840 13046 6896
rect 13358 7656 13414 7712
rect 13358 7540 13414 7576
rect 13358 7520 13360 7540
rect 13360 7520 13412 7540
rect 13412 7520 13414 7540
rect 13910 13232 13966 13288
rect 13634 7928 13690 7984
rect 14002 10920 14058 10976
rect 13910 10648 13966 10704
rect 13174 6840 13230 6896
rect 13174 6160 13230 6216
rect 12990 5072 13046 5128
rect 12898 4528 12954 4584
rect 12898 3440 12954 3496
rect 13542 6432 13598 6488
rect 14462 17448 14518 17504
rect 14186 16224 14242 16280
rect 14370 16360 14426 16416
rect 14186 14068 14242 14104
rect 14186 14048 14188 14068
rect 14188 14048 14240 14068
rect 14240 14048 14242 14068
rect 14186 13776 14242 13832
rect 14370 14592 14426 14648
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 15014 18672 15070 18728
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 15198 18264 15254 18320
rect 15106 18128 15162 18184
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14646 16244 14702 16280
rect 14646 16224 14648 16244
rect 14648 16224 14700 16244
rect 14700 16224 14702 16244
rect 14922 16224 14978 16280
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 14922 13912 14978 13968
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 15474 18128 15530 18184
rect 14186 12688 14242 12744
rect 14186 12008 14242 12064
rect 14186 11328 14242 11384
rect 14186 10648 14242 10704
rect 14186 10240 14242 10296
rect 13910 5888 13966 5944
rect 13174 4120 13230 4176
rect 13174 3304 13230 3360
rect 13174 3032 13230 3088
rect 13174 2896 13230 2952
rect 13450 5072 13506 5128
rect 13542 4664 13598 4720
rect 13542 2896 13598 2952
rect 14646 12688 14702 12744
rect 14922 12688 14978 12744
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 15106 12552 15162 12608
rect 15106 12416 15162 12472
rect 14646 12008 14702 12064
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 14646 10920 14702 10976
rect 15014 10548 15016 10568
rect 15016 10548 15068 10568
rect 15068 10548 15070 10568
rect 15014 10512 15070 10548
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14462 9152 14518 9208
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 14462 8880 14518 8936
rect 14462 8064 14518 8120
rect 14462 7656 14518 7712
rect 14462 7540 14518 7576
rect 14462 7520 14464 7540
rect 14464 7520 14516 7540
rect 14516 7520 14518 7540
rect 15014 8608 15070 8664
rect 15014 8336 15070 8392
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 15382 15816 15438 15872
rect 15750 18708 15752 18728
rect 15752 18708 15804 18728
rect 15804 18708 15806 18728
rect 15750 18672 15806 18708
rect 15658 17992 15714 18048
rect 16026 17992 16082 18048
rect 15842 17448 15898 17504
rect 15750 15272 15806 15328
rect 15474 13912 15530 13968
rect 15934 14048 15990 14104
rect 15474 11736 15530 11792
rect 15382 11056 15438 11112
rect 15198 10240 15254 10296
rect 14278 4800 14334 4856
rect 14002 4392 14058 4448
rect 13726 3168 13782 3224
rect 14002 3848 14058 3904
rect 13910 3168 13966 3224
rect 13818 2796 13820 2816
rect 13820 2796 13872 2816
rect 13872 2796 13874 2816
rect 13818 2760 13874 2796
rect 13910 2644 13966 2680
rect 13910 2624 13912 2644
rect 13912 2624 13964 2644
rect 13964 2624 13966 2644
rect 13910 2488 13966 2544
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14922 6432 14978 6488
rect 15750 10920 15806 10976
rect 15750 10376 15806 10432
rect 15382 9424 15438 9480
rect 15382 8200 15438 8256
rect 16026 10784 16082 10840
rect 15842 10104 15898 10160
rect 15934 9832 15990 9888
rect 15750 8744 15806 8800
rect 16302 17992 16358 18048
rect 16210 13232 16266 13288
rect 16210 12008 16266 12064
rect 18970 22072 19026 22128
rect 18510 21120 18566 21176
rect 16762 19216 16818 19272
rect 16670 18536 16726 18592
rect 16946 18128 17002 18184
rect 16578 16632 16634 16688
rect 16394 15408 16450 15464
rect 16670 16224 16726 16280
rect 16670 14864 16726 14920
rect 16118 9832 16174 9888
rect 15106 6160 15162 6216
rect 14462 5772 14518 5808
rect 14462 5752 14464 5772
rect 14464 5752 14516 5772
rect 14516 5752 14518 5772
rect 15106 6024 15162 6080
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 15106 5888 15162 5944
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 14370 1944 14426 2000
rect 14646 3188 14702 3224
rect 14646 3168 14648 3188
rect 14648 3168 14700 3188
rect 14700 3168 14702 3188
rect 14554 2896 14610 2952
rect 15290 5208 15346 5264
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 16026 7656 16082 7712
rect 15842 6876 15844 6896
rect 15844 6876 15896 6896
rect 15896 6876 15898 6896
rect 15842 6840 15898 6876
rect 15382 2352 15438 2408
rect 15934 2644 15990 2680
rect 16302 11328 16358 11384
rect 16762 13640 16818 13696
rect 16762 13388 16818 13424
rect 16762 13368 16764 13388
rect 16764 13368 16816 13388
rect 16816 13368 16818 13388
rect 17314 18400 17370 18456
rect 17222 18028 17224 18048
rect 17224 18028 17276 18048
rect 17276 18028 17278 18048
rect 17222 17992 17278 18028
rect 17130 16668 17132 16688
rect 17132 16668 17184 16688
rect 17184 16668 17186 16688
rect 17130 16632 17186 16668
rect 17038 15952 17094 16008
rect 16946 13796 17002 13832
rect 16946 13776 16948 13796
rect 16948 13776 17000 13796
rect 17000 13776 17002 13796
rect 16946 13096 17002 13152
rect 16946 12436 17002 12472
rect 16946 12416 16948 12436
rect 16948 12416 17000 12436
rect 17000 12416 17002 12436
rect 16854 11756 16910 11792
rect 16854 11736 16856 11756
rect 16856 11736 16908 11756
rect 16908 11736 16910 11756
rect 17314 16904 17370 16960
rect 17866 19352 17922 19408
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 18050 19352 18106 19408
rect 17130 13368 17186 13424
rect 17222 12960 17278 13016
rect 16486 10920 16542 10976
rect 16394 9696 16450 9752
rect 16302 8744 16358 8800
rect 16302 7792 16358 7848
rect 16210 4936 16266 4992
rect 15934 2624 15936 2644
rect 15936 2624 15988 2644
rect 15988 2624 15990 2644
rect 16762 10512 16818 10568
rect 16762 10004 16764 10024
rect 16764 10004 16816 10024
rect 16816 10004 16818 10024
rect 16762 9968 16818 10004
rect 17314 12588 17316 12608
rect 17316 12588 17368 12608
rect 17368 12588 17370 12608
rect 17314 12552 17370 12588
rect 17038 10920 17094 10976
rect 16762 7148 16764 7168
rect 16764 7148 16816 7168
rect 16816 7148 16818 7168
rect 16762 7112 16818 7148
rect 16670 6432 16726 6488
rect 16578 5108 16580 5128
rect 16580 5108 16632 5128
rect 16632 5108 16634 5128
rect 16578 5072 16634 5108
rect 16578 3884 16580 3904
rect 16580 3884 16632 3904
rect 16632 3884 16634 3904
rect 16578 3848 16634 3884
rect 16578 1944 16634 2000
rect 16946 5480 17002 5536
rect 17314 11056 17370 11112
rect 17222 10684 17224 10704
rect 17224 10684 17276 10704
rect 17276 10684 17278 10704
rect 17222 10648 17278 10684
rect 17314 10240 17370 10296
rect 17314 9968 17370 10024
rect 17406 9832 17462 9888
rect 17314 8880 17370 8936
rect 16946 2644 17002 2680
rect 16946 2624 16948 2644
rect 16948 2624 17000 2644
rect 17000 2624 17002 2644
rect 17222 4256 17278 4312
rect 17314 3732 17370 3768
rect 17314 3712 17316 3732
rect 17316 3712 17368 3732
rect 17368 3712 17370 3732
rect 17590 12552 17646 12608
rect 17590 12280 17646 12336
rect 17590 11736 17646 11792
rect 17866 18828 17922 18864
rect 17866 18808 17868 18828
rect 17868 18808 17920 18828
rect 17920 18808 17922 18828
rect 18694 21528 18750 21584
rect 18602 19760 18658 19816
rect 18602 19216 18658 19272
rect 18418 18808 18474 18864
rect 18694 18808 18750 18864
rect 17866 18128 17922 18184
rect 17774 17720 17830 17776
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 18050 18028 18052 18048
rect 18052 18028 18104 18048
rect 18104 18028 18106 18048
rect 18050 17992 18106 18028
rect 17958 17584 18014 17640
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 17866 16768 17922 16824
rect 17774 16652 17830 16688
rect 17774 16632 17776 16652
rect 17776 16632 17828 16652
rect 17828 16632 17830 16652
rect 17774 15408 17830 15464
rect 18142 16940 18144 16960
rect 18144 16940 18196 16960
rect 18196 16940 18198 16960
rect 18142 16904 18198 16940
rect 18326 16904 18382 16960
rect 18786 18264 18842 18320
rect 18510 16652 18566 16688
rect 18510 16632 18512 16652
rect 18512 16632 18564 16652
rect 18564 16632 18566 16652
rect 18234 16496 18290 16552
rect 17958 16360 18014 16416
rect 18510 16360 18566 16416
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 17958 14864 18014 14920
rect 18050 14592 18106 14648
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18418 13912 18474 13968
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 17774 12552 17830 12608
rect 17682 11636 17684 11656
rect 17684 11636 17736 11656
rect 17736 11636 17738 11656
rect 17682 11600 17738 11636
rect 17682 11212 17738 11248
rect 17682 11192 17684 11212
rect 17684 11192 17736 11212
rect 17736 11192 17738 11212
rect 18326 12416 18382 12472
rect 18970 17720 19026 17776
rect 18878 17040 18934 17096
rect 18786 13912 18842 13968
rect 18786 13096 18842 13152
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 17866 9152 17922 9208
rect 18694 12552 18750 12608
rect 19246 20576 19302 20632
rect 19338 20168 19394 20224
rect 19430 19624 19486 19680
rect 19246 18420 19302 18456
rect 19890 19352 19946 19408
rect 19246 18400 19248 18420
rect 19248 18400 19300 18420
rect 19300 18400 19302 18420
rect 19246 17176 19302 17232
rect 19338 16940 19340 16960
rect 19340 16940 19392 16960
rect 19392 16940 19394 16960
rect 19338 16904 19394 16940
rect 19246 14456 19302 14512
rect 18878 12960 18934 13016
rect 19430 13796 19486 13832
rect 19430 13776 19432 13796
rect 19432 13776 19484 13796
rect 19484 13776 19486 13796
rect 19338 12960 19394 13016
rect 19154 12552 19210 12608
rect 19798 18128 19854 18184
rect 19706 17992 19762 18048
rect 19890 17856 19946 17912
rect 19614 15544 19670 15600
rect 19614 14340 19670 14376
rect 19614 14320 19616 14340
rect 19616 14320 19668 14340
rect 19668 14320 19670 14340
rect 19614 13912 19670 13968
rect 20166 18400 20222 18456
rect 20902 18672 20958 18728
rect 20074 16088 20130 16144
rect 19890 13776 19946 13832
rect 19154 12436 19210 12472
rect 19154 12416 19156 12436
rect 19156 12416 19208 12436
rect 19208 12416 19210 12436
rect 18786 11348 18842 11384
rect 18786 11328 18788 11348
rect 18788 11328 18840 11348
rect 18840 11328 18842 11348
rect 18786 10512 18842 10568
rect 18418 9968 18474 10024
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 18234 8492 18290 8528
rect 18234 8472 18236 8492
rect 18236 8472 18288 8492
rect 18288 8472 18290 8492
rect 17590 6568 17646 6624
rect 17590 6024 17646 6080
rect 17590 5344 17646 5400
rect 17314 2896 17370 2952
rect 17774 3168 17830 3224
rect 17774 3032 17830 3088
rect 17222 2508 17278 2544
rect 17222 2488 17224 2508
rect 17224 2488 17276 2508
rect 17276 2488 17278 2508
rect 18418 7928 18474 7984
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 18326 6704 18382 6760
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 18050 3440 18106 3496
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 18878 9968 18934 10024
rect 18878 9560 18934 9616
rect 18786 9424 18842 9480
rect 18970 8744 19026 8800
rect 18786 8200 18842 8256
rect 18694 7520 18750 7576
rect 18970 7112 19026 7168
rect 18878 6840 18934 6896
rect 18878 5772 18934 5808
rect 18878 5752 18880 5772
rect 18880 5752 18932 5772
rect 18932 5752 18934 5772
rect 18786 5344 18842 5400
rect 19890 13132 19892 13152
rect 19892 13132 19944 13152
rect 19944 13132 19946 13152
rect 19890 13096 19946 13132
rect 19890 12824 19946 12880
rect 19890 12552 19946 12608
rect 19798 11772 19800 11792
rect 19800 11772 19852 11792
rect 19852 11772 19854 11792
rect 19798 11736 19854 11772
rect 19338 9968 19394 10024
rect 19338 9288 19394 9344
rect 19246 8916 19248 8936
rect 19248 8916 19300 8936
rect 19300 8916 19302 8936
rect 19246 8880 19302 8916
rect 19338 8744 19394 8800
rect 19430 8472 19486 8528
rect 18970 3984 19026 4040
rect 18878 3712 18934 3768
rect 18786 3576 18842 3632
rect 18970 3168 19026 3224
rect 18326 3032 18382 3088
rect 18602 3032 18658 3088
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 18050 1808 18106 1864
rect 17958 1536 18014 1592
rect 17958 1128 18014 1184
rect 18878 2760 18934 2816
rect 18786 2352 18842 2408
rect 3974 176 4030 232
rect 19062 2488 19118 2544
rect 19338 3612 19340 3632
rect 19340 3612 19392 3632
rect 19392 3612 19394 3632
rect 19338 3576 19394 3612
rect 19246 3440 19302 3496
rect 19614 4276 19670 4312
rect 19614 4256 19616 4276
rect 19616 4256 19668 4276
rect 19668 4256 19670 4276
rect 20166 14764 20168 14784
rect 20168 14764 20220 14784
rect 20220 14764 20222 14784
rect 20166 14728 20222 14764
rect 20350 15272 20406 15328
rect 20902 13504 20958 13560
rect 19614 3168 19670 3224
rect 19890 3168 19946 3224
rect 19798 3032 19854 3088
rect 19154 584 19210 640
rect 20718 7792 20774 7848
rect 20442 2644 20498 2680
rect 20442 2624 20444 2644
rect 20444 2624 20496 2644
rect 20496 2624 20498 2644
rect 21086 15000 21142 15056
rect 21178 13232 21234 13288
rect 21454 17312 21510 17368
rect 21362 13912 21418 13968
rect 21362 11328 21418 11384
rect 20810 4392 20866 4448
rect 20810 3440 20866 3496
rect 21270 1536 21326 1592
rect 21362 1128 21418 1184
rect 18878 176 18934 232
<< metal3 >>
rect 0 22538 480 22568
rect 3233 22538 3299 22541
rect 0 22536 3299 22538
rect 0 22480 3238 22536
rect 3294 22480 3299 22536
rect 0 22478 3299 22480
rect 0 22448 480 22478
rect 3233 22475 3299 22478
rect 19057 22538 19123 22541
rect 22320 22538 22800 22568
rect 19057 22536 22800 22538
rect 19057 22480 19062 22536
rect 19118 22480 22800 22536
rect 19057 22478 22800 22480
rect 19057 22475 19123 22478
rect 22320 22448 22800 22478
rect 0 22130 480 22160
rect 3049 22130 3115 22133
rect 0 22128 3115 22130
rect 0 22072 3054 22128
rect 3110 22072 3115 22128
rect 0 22070 3115 22072
rect 0 22040 480 22070
rect 3049 22067 3115 22070
rect 18965 22130 19031 22133
rect 22320 22130 22800 22160
rect 18965 22128 22800 22130
rect 18965 22072 18970 22128
rect 19026 22072 22800 22128
rect 18965 22070 22800 22072
rect 18965 22067 19031 22070
rect 22320 22040 22800 22070
rect 0 21586 480 21616
rect 2957 21586 3023 21589
rect 0 21584 3023 21586
rect 0 21528 2962 21584
rect 3018 21528 3023 21584
rect 0 21526 3023 21528
rect 0 21496 480 21526
rect 2957 21523 3023 21526
rect 18689 21586 18755 21589
rect 22320 21586 22800 21616
rect 18689 21584 22800 21586
rect 18689 21528 18694 21584
rect 18750 21528 22800 21584
rect 18689 21526 22800 21528
rect 18689 21523 18755 21526
rect 22320 21496 22800 21526
rect 0 21178 480 21208
rect 2865 21178 2931 21181
rect 0 21176 2931 21178
rect 0 21120 2870 21176
rect 2926 21120 2931 21176
rect 0 21118 2931 21120
rect 0 21088 480 21118
rect 2865 21115 2931 21118
rect 18505 21178 18571 21181
rect 22320 21178 22800 21208
rect 18505 21176 22800 21178
rect 18505 21120 18510 21176
rect 18566 21120 22800 21176
rect 18505 21118 22800 21120
rect 18505 21115 18571 21118
rect 22320 21088 22800 21118
rect 0 20634 480 20664
rect 2773 20634 2839 20637
rect 0 20632 2839 20634
rect 0 20576 2778 20632
rect 2834 20576 2839 20632
rect 0 20574 2839 20576
rect 0 20544 480 20574
rect 2773 20571 2839 20574
rect 19241 20634 19307 20637
rect 22320 20634 22800 20664
rect 19241 20632 22800 20634
rect 19241 20576 19246 20632
rect 19302 20576 22800 20632
rect 19241 20574 22800 20576
rect 19241 20571 19307 20574
rect 22320 20544 22800 20574
rect 13854 20300 13860 20364
rect 13924 20362 13930 20364
rect 14917 20362 14983 20365
rect 13924 20360 14983 20362
rect 13924 20304 14922 20360
rect 14978 20304 14983 20360
rect 13924 20302 14983 20304
rect 13924 20300 13930 20302
rect 14917 20299 14983 20302
rect 0 20226 480 20256
rect 3141 20226 3207 20229
rect 0 20224 3207 20226
rect 0 20168 3146 20224
rect 3202 20168 3207 20224
rect 0 20166 3207 20168
rect 0 20136 480 20166
rect 3141 20163 3207 20166
rect 19333 20226 19399 20229
rect 22320 20226 22800 20256
rect 19333 20224 22800 20226
rect 19333 20168 19338 20224
rect 19394 20168 22800 20224
rect 19333 20166 22800 20168
rect 19333 20163 19399 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 22320 20136 22800 20166
rect 14672 20095 14992 20096
rect 13670 19756 13676 19820
rect 13740 19818 13746 19820
rect 18597 19818 18663 19821
rect 13740 19816 18663 19818
rect 13740 19760 18602 19816
rect 18658 19760 18663 19816
rect 13740 19758 18663 19760
rect 13740 19756 13746 19758
rect 18597 19755 18663 19758
rect 0 19682 480 19712
rect 1761 19682 1827 19685
rect 0 19680 1827 19682
rect 0 19624 1766 19680
rect 1822 19624 1827 19680
rect 0 19622 1827 19624
rect 0 19592 480 19622
rect 1761 19619 1827 19622
rect 19425 19682 19491 19685
rect 22320 19682 22800 19712
rect 19425 19680 22800 19682
rect 19425 19624 19430 19680
rect 19486 19624 22800 19680
rect 19425 19622 22800 19624
rect 19425 19619 19491 19622
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 22320 19592 22800 19622
rect 18104 19551 18424 19552
rect 7465 19546 7531 19549
rect 10317 19546 10383 19549
rect 14273 19548 14339 19549
rect 14222 19546 14228 19548
rect 7465 19544 10383 19546
rect 7465 19488 7470 19544
rect 7526 19488 10322 19544
rect 10378 19488 10383 19544
rect 7465 19486 10383 19488
rect 14182 19486 14228 19546
rect 14292 19544 14339 19548
rect 14334 19488 14339 19544
rect 7465 19483 7531 19486
rect 10317 19483 10383 19486
rect 14222 19484 14228 19486
rect 14292 19484 14339 19488
rect 14273 19483 14339 19484
rect 10777 19410 10843 19413
rect 12249 19410 12315 19413
rect 14365 19412 14431 19413
rect 10777 19408 13370 19410
rect 10777 19352 10782 19408
rect 10838 19352 12254 19408
rect 12310 19352 13370 19408
rect 10777 19350 13370 19352
rect 10777 19347 10843 19350
rect 12249 19347 12315 19350
rect 0 19274 480 19304
rect 13310 19277 13370 19350
rect 14365 19408 14412 19412
rect 14476 19410 14482 19412
rect 17861 19410 17927 19413
rect 18045 19410 18111 19413
rect 14365 19352 14370 19408
rect 14365 19348 14412 19352
rect 14476 19350 14522 19410
rect 17861 19408 18111 19410
rect 17861 19352 17866 19408
rect 17922 19352 18050 19408
rect 18106 19352 18111 19408
rect 17861 19350 18111 19352
rect 14476 19348 14482 19350
rect 14365 19347 14431 19348
rect 17861 19347 17927 19350
rect 18045 19347 18111 19350
rect 19885 19412 19951 19413
rect 19885 19408 19932 19412
rect 19996 19410 20002 19412
rect 19885 19352 19890 19408
rect 19885 19348 19932 19352
rect 19996 19350 20042 19410
rect 19996 19348 20002 19350
rect 19885 19347 19951 19348
rect 2773 19274 2839 19277
rect 0 19272 2839 19274
rect 0 19216 2778 19272
rect 2834 19216 2839 19272
rect 0 19214 2839 19216
rect 0 19184 480 19214
rect 2773 19211 2839 19214
rect 3969 19274 4035 19277
rect 4102 19274 4108 19276
rect 3969 19272 4108 19274
rect 3969 19216 3974 19272
rect 4030 19216 4108 19272
rect 3969 19214 4108 19216
rect 3969 19211 4035 19214
rect 4102 19212 4108 19214
rect 4172 19212 4178 19276
rect 4981 19274 5047 19277
rect 12709 19274 12775 19277
rect 12985 19276 13051 19277
rect 4981 19272 12775 19274
rect 4981 19216 4986 19272
rect 5042 19216 12714 19272
rect 12770 19216 12775 19272
rect 4981 19214 12775 19216
rect 4981 19211 5047 19214
rect 12709 19211 12775 19214
rect 12934 19212 12940 19276
rect 13004 19274 13051 19276
rect 13004 19272 13096 19274
rect 13046 19216 13096 19272
rect 13004 19214 13096 19216
rect 13310 19272 13419 19277
rect 16757 19274 16823 19277
rect 13310 19216 13358 19272
rect 13414 19216 13419 19272
rect 13310 19214 13419 19216
rect 13004 19212 13051 19214
rect 12985 19211 13051 19212
rect 13353 19211 13419 19214
rect 13862 19272 16823 19274
rect 13862 19216 16762 19272
rect 16818 19216 16823 19272
rect 13862 19214 16823 19216
rect 3785 19138 3851 19141
rect 7281 19138 7347 19141
rect 3785 19136 7347 19138
rect 3785 19080 3790 19136
rect 3846 19080 7286 19136
rect 7342 19080 7347 19136
rect 3785 19078 7347 19080
rect 3785 19075 3851 19078
rect 7281 19075 7347 19078
rect 8385 19138 8451 19141
rect 10041 19138 10107 19141
rect 8385 19136 10107 19138
rect 8385 19080 8390 19136
rect 8446 19080 10046 19136
rect 10102 19080 10107 19136
rect 8385 19078 10107 19080
rect 8385 19075 8451 19078
rect 10041 19075 10107 19078
rect 10225 19138 10291 19141
rect 11237 19138 11303 19141
rect 10225 19136 11303 19138
rect 10225 19080 10230 19136
rect 10286 19080 11242 19136
rect 11298 19080 11303 19136
rect 10225 19078 11303 19080
rect 10225 19075 10291 19078
rect 11237 19075 11303 19078
rect 11697 19138 11763 19141
rect 13721 19138 13787 19141
rect 11697 19136 13787 19138
rect 11697 19080 11702 19136
rect 11758 19080 13726 19136
rect 13782 19080 13787 19136
rect 11697 19078 13787 19080
rect 11697 19075 11763 19078
rect 13721 19075 13787 19078
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 1577 19002 1643 19005
rect 5625 19002 5691 19005
rect 1577 19000 5691 19002
rect 1577 18944 1582 19000
rect 1638 18944 5630 19000
rect 5686 18944 5691 19000
rect 1577 18942 5691 18944
rect 1577 18939 1643 18942
rect 5625 18939 5691 18942
rect 12157 19002 12223 19005
rect 13862 19002 13922 19214
rect 16757 19211 16823 19214
rect 18597 19274 18663 19277
rect 22320 19274 22800 19304
rect 18597 19272 22800 19274
rect 18597 19216 18602 19272
rect 18658 19216 22800 19272
rect 18597 19214 22800 19216
rect 18597 19211 18663 19214
rect 22320 19184 22800 19214
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 12157 19000 13922 19002
rect 12157 18944 12162 19000
rect 12218 18944 13922 19000
rect 12157 18942 13922 18944
rect 12157 18939 12223 18942
rect 2865 18866 2931 18869
rect 9029 18866 9095 18869
rect 2865 18864 9095 18866
rect 2865 18808 2870 18864
rect 2926 18808 9034 18864
rect 9090 18808 9095 18864
rect 2865 18806 9095 18808
rect 2865 18803 2931 18806
rect 9029 18803 9095 18806
rect 10317 18866 10383 18869
rect 17861 18866 17927 18869
rect 10317 18864 17927 18866
rect 10317 18808 10322 18864
rect 10378 18808 17866 18864
rect 17922 18808 17927 18864
rect 10317 18806 17927 18808
rect 10317 18803 10383 18806
rect 17861 18803 17927 18806
rect 18413 18866 18479 18869
rect 18689 18866 18755 18869
rect 18413 18864 18755 18866
rect 18413 18808 18418 18864
rect 18474 18808 18694 18864
rect 18750 18808 18755 18864
rect 18413 18806 18755 18808
rect 18413 18803 18479 18806
rect 18689 18803 18755 18806
rect 0 18730 480 18760
rect 3601 18730 3667 18733
rect 0 18728 3667 18730
rect 0 18672 3606 18728
rect 3662 18672 3667 18728
rect 0 18670 3667 18672
rect 0 18640 480 18670
rect 3601 18667 3667 18670
rect 4245 18730 4311 18733
rect 4838 18730 4844 18732
rect 4245 18728 4844 18730
rect 4245 18672 4250 18728
rect 4306 18672 4844 18728
rect 4245 18670 4844 18672
rect 4245 18667 4311 18670
rect 4838 18668 4844 18670
rect 4908 18730 4914 18732
rect 7465 18730 7531 18733
rect 4908 18728 7531 18730
rect 4908 18672 7470 18728
rect 7526 18672 7531 18728
rect 4908 18670 7531 18672
rect 4908 18668 4914 18670
rect 7465 18667 7531 18670
rect 7649 18730 7715 18733
rect 13077 18730 13143 18733
rect 7649 18728 13143 18730
rect 7649 18672 7654 18728
rect 7710 18672 13082 18728
rect 13138 18672 13143 18728
rect 7649 18670 13143 18672
rect 7649 18667 7715 18670
rect 13077 18667 13143 18670
rect 15009 18730 15075 18733
rect 15142 18730 15148 18732
rect 15009 18728 15148 18730
rect 15009 18672 15014 18728
rect 15070 18672 15148 18728
rect 15009 18670 15148 18672
rect 15009 18667 15075 18670
rect 15142 18668 15148 18670
rect 15212 18668 15218 18732
rect 15745 18730 15811 18733
rect 15878 18730 15884 18732
rect 15745 18728 15884 18730
rect 15745 18672 15750 18728
rect 15806 18672 15884 18728
rect 15745 18670 15884 18672
rect 15745 18667 15811 18670
rect 15878 18668 15884 18670
rect 15948 18730 15954 18732
rect 18822 18730 18828 18732
rect 15948 18670 18828 18730
rect 15948 18668 15954 18670
rect 18822 18668 18828 18670
rect 18892 18668 18898 18732
rect 20897 18730 20963 18733
rect 22320 18730 22800 18760
rect 20897 18728 22800 18730
rect 20897 18672 20902 18728
rect 20958 18672 22800 18728
rect 20897 18670 22800 18672
rect 20897 18667 20963 18670
rect 22320 18640 22800 18670
rect 5625 18594 5691 18597
rect 8385 18594 8451 18597
rect 5625 18592 8451 18594
rect 5625 18536 5630 18592
rect 5686 18536 8390 18592
rect 8446 18536 8451 18592
rect 5625 18534 8451 18536
rect 5625 18531 5691 18534
rect 8385 18531 8451 18534
rect 12801 18594 12867 18597
rect 16665 18594 16731 18597
rect 12801 18592 16731 18594
rect 12801 18536 12806 18592
rect 12862 18536 16670 18592
rect 16726 18536 16731 18592
rect 12801 18534 16731 18536
rect 12801 18531 12867 18534
rect 16665 18531 16731 18534
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 1669 18458 1735 18461
rect 9254 18458 9260 18460
rect 1669 18456 4308 18458
rect 1669 18400 1674 18456
rect 1730 18400 4308 18456
rect 1669 18398 4308 18400
rect 1669 18395 1735 18398
rect 0 18322 480 18352
rect 1669 18322 1735 18325
rect 0 18320 1735 18322
rect 0 18264 1674 18320
rect 1730 18264 1735 18320
rect 0 18262 1735 18264
rect 4248 18322 4308 18398
rect 6686 18398 9260 18458
rect 6686 18322 6746 18398
rect 9254 18396 9260 18398
rect 9324 18458 9330 18460
rect 10225 18458 10291 18461
rect 17309 18458 17375 18461
rect 19241 18460 19307 18461
rect 19190 18458 19196 18460
rect 9324 18456 10291 18458
rect 9324 18400 10230 18456
rect 10286 18400 10291 18456
rect 9324 18398 10291 18400
rect 9324 18396 9330 18398
rect 10225 18395 10291 18398
rect 11654 18456 17375 18458
rect 11654 18400 17314 18456
rect 17370 18400 17375 18456
rect 11654 18398 17375 18400
rect 19150 18398 19196 18458
rect 19260 18456 19307 18460
rect 19302 18400 19307 18456
rect 4248 18262 6746 18322
rect 6821 18322 6887 18325
rect 8385 18322 8451 18325
rect 6821 18320 8451 18322
rect 6821 18264 6826 18320
rect 6882 18264 8390 18320
rect 8446 18264 8451 18320
rect 6821 18262 8451 18264
rect 0 18232 480 18262
rect 1669 18259 1735 18262
rect 6821 18259 6887 18262
rect 8385 18259 8451 18262
rect 8518 18260 8524 18324
rect 8588 18322 8594 18324
rect 11654 18322 11714 18398
rect 17309 18395 17375 18398
rect 19190 18396 19196 18398
rect 19260 18396 19307 18400
rect 19374 18396 19380 18460
rect 19444 18458 19450 18460
rect 20161 18458 20227 18461
rect 19444 18456 20227 18458
rect 19444 18400 20166 18456
rect 20222 18400 20227 18456
rect 19444 18398 20227 18400
rect 19444 18396 19450 18398
rect 19241 18395 19307 18396
rect 20161 18395 20227 18398
rect 8588 18262 11714 18322
rect 12433 18322 12499 18325
rect 15193 18322 15259 18325
rect 15510 18322 15516 18324
rect 12433 18320 15516 18322
rect 12433 18264 12438 18320
rect 12494 18264 15198 18320
rect 15254 18264 15516 18320
rect 12433 18262 15516 18264
rect 8588 18260 8594 18262
rect 12433 18259 12499 18262
rect 15193 18259 15259 18262
rect 15510 18260 15516 18262
rect 15580 18260 15586 18324
rect 18781 18322 18847 18325
rect 22320 18322 22800 18352
rect 18781 18320 22800 18322
rect 18781 18264 18786 18320
rect 18842 18264 22800 18320
rect 18781 18262 22800 18264
rect 18781 18259 18847 18262
rect 22320 18232 22800 18262
rect 3049 18186 3115 18189
rect 4521 18186 4587 18189
rect 3049 18184 4587 18186
rect 3049 18128 3054 18184
rect 3110 18128 4526 18184
rect 4582 18128 4587 18184
rect 3049 18126 4587 18128
rect 3049 18123 3115 18126
rect 4521 18123 4587 18126
rect 6729 18186 6795 18189
rect 10133 18188 10199 18189
rect 10133 18186 10180 18188
rect 6729 18184 9506 18186
rect 6729 18128 6734 18184
rect 6790 18128 9506 18184
rect 6729 18126 9506 18128
rect 10088 18184 10180 18186
rect 10088 18128 10138 18184
rect 10088 18126 10180 18128
rect 6729 18123 6795 18126
rect 9446 18053 9506 18126
rect 10133 18124 10180 18126
rect 10244 18124 10250 18188
rect 12801 18186 12867 18189
rect 13486 18186 13492 18188
rect 12801 18184 13492 18186
rect 12801 18128 12806 18184
rect 12862 18128 13492 18184
rect 12801 18126 13492 18128
rect 10133 18123 10199 18124
rect 12801 18123 12867 18126
rect 13486 18124 13492 18126
rect 13556 18124 13562 18188
rect 14038 18124 14044 18188
rect 14108 18186 14114 18188
rect 15101 18186 15167 18189
rect 14108 18184 15167 18186
rect 14108 18128 15106 18184
rect 15162 18128 15167 18184
rect 14108 18126 15167 18128
rect 14108 18124 14114 18126
rect 15101 18123 15167 18126
rect 15326 18124 15332 18188
rect 15396 18186 15402 18188
rect 15469 18186 15535 18189
rect 15396 18184 15535 18186
rect 15396 18128 15474 18184
rect 15530 18128 15535 18184
rect 15396 18126 15535 18128
rect 15396 18124 15402 18126
rect 15469 18123 15535 18126
rect 16941 18186 17007 18189
rect 17166 18186 17172 18188
rect 16941 18184 17172 18186
rect 16941 18128 16946 18184
rect 17002 18128 17172 18184
rect 16941 18126 17172 18128
rect 16941 18123 17007 18126
rect 17166 18124 17172 18126
rect 17236 18186 17242 18188
rect 17861 18186 17927 18189
rect 17236 18184 17927 18186
rect 17236 18128 17866 18184
rect 17922 18128 17927 18184
rect 17236 18126 17927 18128
rect 17236 18124 17242 18126
rect 17861 18123 17927 18126
rect 19793 18186 19859 18189
rect 20478 18186 20484 18188
rect 19793 18184 20484 18186
rect 19793 18128 19798 18184
rect 19854 18128 20484 18184
rect 19793 18126 20484 18128
rect 19793 18123 19859 18126
rect 20478 18124 20484 18126
rect 20548 18124 20554 18188
rect 7465 18052 7531 18053
rect 7414 17988 7420 18052
rect 7484 18050 7531 18052
rect 9446 18050 9555 18053
rect 13445 18050 13511 18053
rect 7484 18048 7576 18050
rect 7526 17992 7576 18048
rect 7484 17990 7576 17992
rect 9446 18048 13511 18050
rect 9446 17992 9494 18048
rect 9550 17992 13450 18048
rect 13506 17992 13511 18048
rect 9446 17990 13511 17992
rect 7484 17988 7531 17990
rect 7465 17987 7531 17988
rect 9489 17987 9555 17990
rect 13445 17987 13511 17990
rect 13721 18050 13787 18053
rect 15653 18052 15719 18053
rect 16021 18052 16087 18053
rect 13854 18050 13860 18052
rect 13721 18048 13860 18050
rect 13721 17992 13726 18048
rect 13782 17992 13860 18048
rect 13721 17990 13860 17992
rect 13721 17987 13787 17990
rect 13854 17988 13860 17990
rect 13924 17988 13930 18052
rect 15653 18048 15700 18052
rect 15764 18050 15770 18052
rect 15653 17992 15658 18048
rect 15653 17988 15700 17992
rect 15764 17990 15810 18050
rect 16021 18048 16068 18052
rect 16132 18050 16138 18052
rect 16297 18050 16363 18053
rect 16430 18050 16436 18052
rect 16021 17992 16026 18048
rect 15764 17988 15770 17990
rect 16021 17988 16068 17992
rect 16132 17990 16178 18050
rect 16297 18048 16436 18050
rect 16297 17992 16302 18048
rect 16358 17992 16436 18048
rect 16297 17990 16436 17992
rect 16132 17988 16138 17990
rect 15653 17987 15719 17988
rect 16021 17987 16087 17988
rect 16297 17987 16363 17990
rect 16430 17988 16436 17990
rect 16500 17988 16506 18052
rect 16614 17988 16620 18052
rect 16684 18050 16690 18052
rect 17217 18050 17283 18053
rect 16684 18048 17283 18050
rect 16684 17992 17222 18048
rect 17278 17992 17283 18048
rect 16684 17990 17283 17992
rect 16684 17988 16690 17990
rect 17217 17987 17283 17990
rect 17902 17988 17908 18052
rect 17972 18050 17978 18052
rect 18045 18050 18111 18053
rect 17972 18048 18111 18050
rect 17972 17992 18050 18048
rect 18106 17992 18111 18048
rect 17972 17990 18111 17992
rect 17972 17988 17978 17990
rect 18045 17987 18111 17990
rect 19701 18052 19767 18053
rect 19701 18048 19748 18052
rect 19812 18050 19818 18052
rect 19701 17992 19706 18048
rect 19701 17988 19748 17992
rect 19812 17990 19858 18050
rect 19812 17988 19818 17990
rect 19701 17987 19767 17988
rect 7808 17984 8128 17985
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 12525 17914 12591 17917
rect 13905 17914 13971 17917
rect 12525 17912 13971 17914
rect 12525 17856 12530 17912
rect 12586 17856 13910 17912
rect 13966 17856 13971 17912
rect 12525 17854 13971 17856
rect 12525 17851 12591 17854
rect 13905 17851 13971 17854
rect 19558 17852 19564 17916
rect 19628 17914 19634 17916
rect 19885 17914 19951 17917
rect 19628 17912 19951 17914
rect 19628 17856 19890 17912
rect 19946 17856 19951 17912
rect 19628 17854 19951 17856
rect 19628 17852 19634 17854
rect 19885 17851 19951 17854
rect 0 17778 480 17808
rect 1577 17778 1643 17781
rect 0 17776 1643 17778
rect 0 17720 1582 17776
rect 1638 17720 1643 17776
rect 0 17718 1643 17720
rect 0 17688 480 17718
rect 1577 17715 1643 17718
rect 6545 17778 6611 17781
rect 12750 17778 12756 17780
rect 6545 17776 12756 17778
rect 6545 17720 6550 17776
rect 6606 17720 12756 17776
rect 6545 17718 12756 17720
rect 6545 17715 6611 17718
rect 12750 17716 12756 17718
rect 12820 17778 12826 17780
rect 17769 17778 17835 17781
rect 12820 17776 17835 17778
rect 12820 17720 17774 17776
rect 17830 17720 17835 17776
rect 12820 17718 17835 17720
rect 12820 17716 12826 17718
rect 17769 17715 17835 17718
rect 18965 17778 19031 17781
rect 22320 17778 22800 17808
rect 18965 17776 22800 17778
rect 18965 17720 18970 17776
rect 19026 17720 22800 17776
rect 18965 17718 22800 17720
rect 18965 17715 19031 17718
rect 22320 17688 22800 17718
rect 2313 17642 2379 17645
rect 3969 17642 4035 17645
rect 7097 17642 7163 17645
rect 8293 17642 8359 17645
rect 2313 17640 4860 17642
rect 2313 17584 2318 17640
rect 2374 17584 3974 17640
rect 4030 17584 4860 17640
rect 2313 17582 4860 17584
rect 2313 17579 2379 17582
rect 3969 17579 4035 17582
rect 4800 17506 4860 17582
rect 7097 17640 8359 17642
rect 7097 17584 7102 17640
rect 7158 17584 8298 17640
rect 8354 17584 8359 17640
rect 7097 17582 8359 17584
rect 7097 17579 7163 17582
rect 8293 17579 8359 17582
rect 12341 17642 12407 17645
rect 17953 17642 18019 17645
rect 12341 17640 18019 17642
rect 12341 17584 12346 17640
rect 12402 17584 17958 17640
rect 18014 17584 18019 17640
rect 12341 17582 18019 17584
rect 12341 17579 12407 17582
rect 17953 17579 18019 17582
rect 9213 17506 9279 17509
rect 4800 17504 9279 17506
rect 4800 17448 9218 17504
rect 9274 17448 9279 17504
rect 4800 17446 9279 17448
rect 9213 17443 9279 17446
rect 12525 17506 12591 17509
rect 13118 17506 13124 17508
rect 12525 17504 13124 17506
rect 12525 17448 12530 17504
rect 12586 17448 13124 17504
rect 12525 17446 13124 17448
rect 12525 17443 12591 17446
rect 13118 17444 13124 17446
rect 13188 17506 13194 17508
rect 13445 17506 13511 17509
rect 14457 17506 14523 17509
rect 15837 17506 15903 17509
rect 13188 17504 13738 17506
rect 13188 17448 13450 17504
rect 13506 17448 13738 17504
rect 13188 17446 13738 17448
rect 13188 17444 13194 17446
rect 13445 17443 13511 17446
rect 4376 17440 4696 17441
rect 0 17370 480 17400
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 1669 17370 1735 17373
rect 0 17368 1735 17370
rect 0 17312 1674 17368
rect 1730 17312 1735 17368
rect 0 17310 1735 17312
rect 0 17280 480 17310
rect 1669 17307 1735 17310
rect 2129 17370 2195 17373
rect 3417 17370 3483 17373
rect 2129 17368 3483 17370
rect 2129 17312 2134 17368
rect 2190 17312 3422 17368
rect 3478 17312 3483 17368
rect 2129 17310 3483 17312
rect 2129 17307 2195 17310
rect 3417 17307 3483 17310
rect 9397 17372 9463 17373
rect 9397 17368 9444 17372
rect 9508 17370 9514 17372
rect 13537 17370 13603 17373
rect 9397 17312 9402 17368
rect 9397 17308 9444 17312
rect 9508 17310 9554 17370
rect 12022 17368 13603 17370
rect 12022 17312 13542 17368
rect 13598 17312 13603 17368
rect 12022 17310 13603 17312
rect 13678 17370 13738 17446
rect 14457 17504 15903 17506
rect 14457 17448 14462 17504
rect 14518 17448 15842 17504
rect 15898 17448 15903 17504
rect 14457 17446 15903 17448
rect 14457 17443 14523 17446
rect 15837 17443 15903 17446
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 16982 17370 16988 17372
rect 13678 17310 16988 17370
rect 9508 17308 9514 17310
rect 9397 17307 9463 17308
rect 2773 17234 2839 17237
rect 11646 17234 11652 17236
rect 2773 17232 11652 17234
rect 2773 17176 2778 17232
rect 2834 17176 11652 17232
rect 2773 17174 11652 17176
rect 2773 17171 2839 17174
rect 11646 17172 11652 17174
rect 11716 17234 11722 17236
rect 12022 17234 12082 17310
rect 13537 17307 13603 17310
rect 16982 17308 16988 17310
rect 17052 17308 17058 17372
rect 21449 17370 21515 17373
rect 22320 17370 22800 17400
rect 21449 17368 22800 17370
rect 21449 17312 21454 17368
rect 21510 17312 22800 17368
rect 21449 17310 22800 17312
rect 21449 17307 21515 17310
rect 22320 17280 22800 17310
rect 11716 17174 12082 17234
rect 12157 17234 12223 17237
rect 19241 17234 19307 17237
rect 12157 17232 19307 17234
rect 12157 17176 12162 17232
rect 12218 17176 19246 17232
rect 19302 17176 19307 17232
rect 12157 17174 19307 17176
rect 11716 17172 11722 17174
rect 12157 17171 12223 17174
rect 19241 17171 19307 17174
rect 2957 17098 3023 17101
rect 11513 17098 11579 17101
rect 18873 17098 18939 17101
rect 2957 17096 11392 17098
rect 2957 17040 2962 17096
rect 3018 17040 11392 17096
rect 2957 17038 11392 17040
rect 2957 17035 3023 17038
rect 11332 16962 11392 17038
rect 11513 17096 18939 17098
rect 11513 17040 11518 17096
rect 11574 17040 18878 17096
rect 18934 17040 18939 17096
rect 11513 17038 18939 17040
rect 11513 17035 11579 17038
rect 18873 17035 18939 17038
rect 12198 16962 12204 16964
rect 11332 16902 12204 16962
rect 12198 16900 12204 16902
rect 12268 16900 12274 16964
rect 17309 16962 17375 16965
rect 18137 16962 18203 16965
rect 17309 16960 18203 16962
rect 17309 16904 17314 16960
rect 17370 16904 18142 16960
rect 18198 16904 18203 16960
rect 17309 16902 18203 16904
rect 17309 16899 17375 16902
rect 18137 16899 18203 16902
rect 18321 16962 18387 16965
rect 19333 16962 19399 16965
rect 18321 16960 19399 16962
rect 18321 16904 18326 16960
rect 18382 16904 19338 16960
rect 19394 16904 19399 16960
rect 18321 16902 19399 16904
rect 18321 16899 18387 16902
rect 19333 16899 19399 16902
rect 7808 16896 8128 16897
rect 0 16826 480 16856
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 16831 14992 16832
rect 1485 16826 1551 16829
rect 13445 16826 13511 16829
rect 0 16824 1551 16826
rect 0 16768 1490 16824
rect 1546 16768 1551 16824
rect 0 16766 1551 16768
rect 0 16736 480 16766
rect 1485 16763 1551 16766
rect 10734 16824 13511 16826
rect 10734 16768 13450 16824
rect 13506 16768 13511 16824
rect 10734 16766 13511 16768
rect 6729 16690 6795 16693
rect 10734 16690 10794 16766
rect 13445 16763 13511 16766
rect 17861 16826 17927 16829
rect 22320 16826 22800 16856
rect 17861 16824 22800 16826
rect 17861 16768 17866 16824
rect 17922 16768 22800 16824
rect 17861 16766 22800 16768
rect 17861 16763 17927 16766
rect 22320 16736 22800 16766
rect 6729 16688 10794 16690
rect 6729 16632 6734 16688
rect 6790 16632 10794 16688
rect 6729 16630 10794 16632
rect 10961 16690 11027 16693
rect 13261 16690 13327 16693
rect 15878 16690 15884 16692
rect 10961 16688 12772 16690
rect 10961 16632 10966 16688
rect 11022 16632 12772 16688
rect 10961 16630 12772 16632
rect 6729 16627 6795 16630
rect 10961 16627 11027 16630
rect 12712 16557 12772 16630
rect 13261 16688 15884 16690
rect 13261 16632 13266 16688
rect 13322 16632 15884 16688
rect 13261 16630 15884 16632
rect 13261 16627 13327 16630
rect 15878 16628 15884 16630
rect 15948 16628 15954 16692
rect 16573 16688 16639 16693
rect 16573 16632 16578 16688
rect 16634 16632 16639 16688
rect 16573 16627 16639 16632
rect 17125 16690 17191 16693
rect 17769 16692 17835 16693
rect 17718 16690 17724 16692
rect 17125 16688 17724 16690
rect 17788 16690 17835 16692
rect 18505 16690 18571 16693
rect 18638 16690 18644 16692
rect 17788 16688 17880 16690
rect 17125 16632 17130 16688
rect 17186 16632 17724 16688
rect 17830 16632 17880 16688
rect 17125 16630 17724 16632
rect 17125 16627 17191 16630
rect 17718 16628 17724 16630
rect 17788 16630 17880 16632
rect 18505 16688 18644 16690
rect 18505 16632 18510 16688
rect 18566 16632 18644 16688
rect 18505 16630 18644 16632
rect 17788 16628 17835 16630
rect 17769 16627 17835 16628
rect 18505 16627 18571 16630
rect 18638 16628 18644 16630
rect 18708 16628 18714 16692
rect 5625 16554 5691 16557
rect 11881 16554 11947 16557
rect 5625 16552 11947 16554
rect 5625 16496 5630 16552
rect 5686 16496 11886 16552
rect 11942 16496 11947 16552
rect 5625 16494 11947 16496
rect 5625 16491 5691 16494
rect 11881 16491 11947 16494
rect 12198 16492 12204 16556
rect 12268 16554 12274 16556
rect 12525 16554 12591 16557
rect 12268 16552 12591 16554
rect 12268 16496 12530 16552
rect 12586 16496 12591 16552
rect 12268 16494 12591 16496
rect 12268 16492 12274 16494
rect 12525 16491 12591 16494
rect 12709 16554 12775 16557
rect 16576 16554 16636 16627
rect 12709 16552 16636 16554
rect 12709 16496 12714 16552
rect 12770 16496 16636 16552
rect 12709 16494 16636 16496
rect 12709 16491 12775 16494
rect 16798 16492 16804 16556
rect 16868 16554 16874 16556
rect 18229 16554 18295 16557
rect 16868 16552 18295 16554
rect 16868 16496 18234 16552
rect 18290 16496 18295 16552
rect 16868 16494 18295 16496
rect 16868 16492 16874 16494
rect 18229 16491 18295 16494
rect 0 16418 480 16448
rect 3417 16418 3483 16421
rect 0 16416 3483 16418
rect 0 16360 3422 16416
rect 3478 16360 3483 16416
rect 0 16358 3483 16360
rect 0 16328 480 16358
rect 3417 16355 3483 16358
rect 11697 16418 11763 16421
rect 13997 16418 14063 16421
rect 11697 16416 14063 16418
rect 11697 16360 11702 16416
rect 11758 16360 14002 16416
rect 14058 16360 14063 16416
rect 11697 16358 14063 16360
rect 11697 16355 11763 16358
rect 13997 16355 14063 16358
rect 14365 16418 14431 16421
rect 17953 16418 18019 16421
rect 14365 16416 18019 16418
rect 14365 16360 14370 16416
rect 14426 16360 17958 16416
rect 18014 16360 18019 16416
rect 14365 16358 18019 16360
rect 14365 16355 14431 16358
rect 17953 16355 18019 16358
rect 18505 16418 18571 16421
rect 22320 16418 22800 16448
rect 18505 16416 22800 16418
rect 18505 16360 18510 16416
rect 18566 16360 22800 16416
rect 18505 16358 22800 16360
rect 18505 16355 18571 16358
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 22320 16328 22800 16358
rect 18104 16287 18424 16288
rect 6729 16282 6795 16285
rect 11881 16282 11947 16285
rect 13813 16282 13879 16285
rect 4800 16280 11162 16282
rect 4800 16224 6734 16280
rect 6790 16224 11162 16280
rect 4800 16222 11162 16224
rect 3325 16146 3391 16149
rect 4800 16146 4860 16222
rect 6729 16219 6795 16222
rect 3325 16144 4860 16146
rect 3325 16088 3330 16144
rect 3386 16088 4860 16144
rect 3325 16086 4860 16088
rect 8109 16146 8175 16149
rect 10961 16146 11027 16149
rect 8109 16144 11027 16146
rect 8109 16088 8114 16144
rect 8170 16088 10966 16144
rect 11022 16088 11027 16144
rect 8109 16086 11027 16088
rect 11102 16146 11162 16222
rect 11881 16280 13879 16282
rect 11881 16224 11886 16280
rect 11942 16224 13818 16280
rect 13874 16224 13879 16280
rect 11881 16222 13879 16224
rect 11881 16219 11947 16222
rect 13813 16219 13879 16222
rect 14181 16282 14247 16285
rect 14641 16282 14707 16285
rect 14181 16280 14707 16282
rect 14181 16224 14186 16280
rect 14242 16224 14646 16280
rect 14702 16224 14707 16280
rect 14181 16222 14707 16224
rect 14181 16219 14247 16222
rect 14641 16219 14707 16222
rect 14917 16282 14983 16285
rect 16665 16282 16731 16285
rect 14917 16280 16731 16282
rect 14917 16224 14922 16280
rect 14978 16224 16670 16280
rect 16726 16224 16731 16280
rect 14917 16222 16731 16224
rect 14917 16219 14983 16222
rect 16665 16219 16731 16222
rect 20069 16146 20135 16149
rect 11102 16144 20135 16146
rect 11102 16088 20074 16144
rect 20130 16088 20135 16144
rect 11102 16086 20135 16088
rect 3325 16083 3391 16086
rect 8109 16083 8175 16086
rect 10961 16083 11027 16086
rect 20069 16083 20135 16086
rect 2497 16010 2563 16013
rect 5809 16010 5875 16013
rect 6085 16010 6151 16013
rect 2497 16008 6151 16010
rect 2497 15952 2502 16008
rect 2558 15952 5814 16008
rect 5870 15952 6090 16008
rect 6146 15952 6151 16008
rect 2497 15950 6151 15952
rect 2497 15947 2563 15950
rect 5809 15947 5875 15950
rect 6085 15947 6151 15950
rect 9029 16010 9095 16013
rect 17033 16010 17099 16013
rect 9029 16008 17099 16010
rect 9029 15952 9034 16008
rect 9090 15952 17038 16008
rect 17094 15952 17099 16008
rect 9029 15950 17099 15952
rect 9029 15947 9095 15950
rect 17033 15947 17099 15950
rect 0 15874 480 15904
rect 3969 15874 4035 15877
rect 0 15872 4035 15874
rect 0 15816 3974 15872
rect 4030 15816 4035 15872
rect 0 15814 4035 15816
rect 0 15784 480 15814
rect 3969 15811 4035 15814
rect 10501 15874 10567 15877
rect 12249 15874 12315 15877
rect 10501 15872 12315 15874
rect 10501 15816 10506 15872
rect 10562 15816 12254 15872
rect 12310 15816 12315 15872
rect 10501 15814 12315 15816
rect 10501 15811 10567 15814
rect 12249 15811 12315 15814
rect 12566 15812 12572 15876
rect 12636 15874 12642 15876
rect 15377 15874 15443 15877
rect 22320 15874 22800 15904
rect 12636 15814 14106 15874
rect 12636 15812 12642 15814
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 9581 15738 9647 15741
rect 13629 15738 13695 15741
rect 9581 15736 13695 15738
rect 9581 15680 9586 15736
rect 9642 15680 13634 15736
rect 13690 15680 13695 15736
rect 9581 15678 13695 15680
rect 9581 15675 9647 15678
rect 13629 15675 13695 15678
rect 1761 15602 1827 15605
rect 9622 15602 9628 15604
rect 1761 15600 9628 15602
rect 1761 15544 1766 15600
rect 1822 15544 9628 15600
rect 1761 15542 9628 15544
rect 1761 15539 1827 15542
rect 9622 15540 9628 15542
rect 9692 15602 9698 15604
rect 13905 15602 13971 15605
rect 9692 15600 13971 15602
rect 9692 15544 13910 15600
rect 13966 15544 13971 15600
rect 9692 15542 13971 15544
rect 14046 15602 14106 15814
rect 15377 15872 22800 15874
rect 15377 15816 15382 15872
rect 15438 15816 22800 15872
rect 15377 15814 22800 15816
rect 15377 15811 15443 15814
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 22320 15784 22800 15814
rect 14672 15743 14992 15744
rect 16246 15602 16252 15604
rect 14046 15542 16252 15602
rect 9692 15540 9698 15542
rect 13905 15539 13971 15542
rect 16246 15540 16252 15542
rect 16316 15602 16322 15604
rect 19609 15602 19675 15605
rect 16316 15600 19675 15602
rect 16316 15544 19614 15600
rect 19670 15544 19675 15600
rect 16316 15542 19675 15544
rect 16316 15540 16322 15542
rect 19609 15539 19675 15542
rect 0 15466 480 15496
rect 4061 15466 4127 15469
rect 0 15464 4127 15466
rect 0 15408 4066 15464
rect 4122 15408 4127 15464
rect 0 15406 4127 15408
rect 0 15376 480 15406
rect 4061 15403 4127 15406
rect 8385 15466 8451 15469
rect 12382 15466 12388 15468
rect 8385 15464 12388 15466
rect 8385 15408 8390 15464
rect 8446 15408 12388 15464
rect 8385 15406 12388 15408
rect 8385 15403 8451 15406
rect 12382 15404 12388 15406
rect 12452 15404 12458 15468
rect 12525 15466 12591 15469
rect 16389 15466 16455 15469
rect 12525 15464 16455 15466
rect 12525 15408 12530 15464
rect 12586 15408 16394 15464
rect 16450 15408 16455 15464
rect 12525 15406 16455 15408
rect 12525 15403 12591 15406
rect 16389 15403 16455 15406
rect 17769 15466 17835 15469
rect 22320 15466 22800 15496
rect 17769 15464 22800 15466
rect 17769 15408 17774 15464
rect 17830 15408 22800 15464
rect 17769 15406 22800 15408
rect 17769 15403 17835 15406
rect 22320 15376 22800 15406
rect 2405 15330 2471 15333
rect 4245 15330 4311 15333
rect 2405 15328 4311 15330
rect 2405 15272 2410 15328
rect 2466 15272 4250 15328
rect 4306 15272 4311 15328
rect 2405 15270 4311 15272
rect 2405 15267 2471 15270
rect 4245 15267 4311 15270
rect 6085 15330 6151 15333
rect 8518 15330 8524 15332
rect 6085 15328 8524 15330
rect 6085 15272 6090 15328
rect 6146 15272 8524 15328
rect 6085 15270 8524 15272
rect 6085 15267 6151 15270
rect 8518 15268 8524 15270
rect 8588 15268 8594 15332
rect 9213 15330 9279 15333
rect 9765 15330 9831 15333
rect 9213 15328 9831 15330
rect 9213 15272 9218 15328
rect 9274 15272 9770 15328
rect 9826 15272 9831 15328
rect 9213 15270 9831 15272
rect 9213 15267 9279 15270
rect 9765 15267 9831 15270
rect 12433 15330 12499 15333
rect 15745 15330 15811 15333
rect 20345 15332 20411 15333
rect 20294 15330 20300 15332
rect 12433 15328 15811 15330
rect 12433 15272 12438 15328
rect 12494 15272 15750 15328
rect 15806 15272 15811 15328
rect 12433 15270 15811 15272
rect 20254 15270 20300 15330
rect 20364 15328 20411 15332
rect 20406 15272 20411 15328
rect 12433 15267 12499 15270
rect 15745 15267 15811 15270
rect 20294 15268 20300 15270
rect 20364 15268 20411 15272
rect 20345 15267 20411 15268
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 7925 15194 7991 15197
rect 10501 15194 10567 15197
rect 10961 15194 11027 15197
rect 7925 15192 11027 15194
rect 7925 15136 7930 15192
rect 7986 15136 10506 15192
rect 10562 15136 10966 15192
rect 11022 15136 11027 15192
rect 7925 15134 11027 15136
rect 7925 15131 7991 15134
rect 10501 15131 10567 15134
rect 10961 15131 11027 15134
rect 12709 15194 12775 15197
rect 12709 15192 16130 15194
rect 12709 15136 12714 15192
rect 12770 15136 16130 15192
rect 12709 15134 16130 15136
rect 12709 15131 12775 15134
rect 9213 15058 9279 15061
rect 15326 15058 15332 15060
rect 9213 15056 15332 15058
rect 9213 15000 9218 15056
rect 9274 15000 15332 15056
rect 9213 14998 15332 15000
rect 9213 14995 9279 14998
rect 15326 14996 15332 14998
rect 15396 15058 15402 15060
rect 15878 15058 15884 15060
rect 15396 14998 15884 15058
rect 15396 14996 15402 14998
rect 15878 14996 15884 14998
rect 15948 14996 15954 15060
rect 16070 15058 16130 15134
rect 21081 15058 21147 15061
rect 16070 15056 21147 15058
rect 16070 15000 21086 15056
rect 21142 15000 21147 15056
rect 16070 14998 21147 15000
rect 21081 14995 21147 14998
rect 0 14922 480 14952
rect 4061 14922 4127 14925
rect 0 14920 4127 14922
rect 0 14864 4066 14920
rect 4122 14864 4127 14920
rect 0 14862 4127 14864
rect 0 14832 480 14862
rect 4061 14859 4127 14862
rect 7649 14922 7715 14925
rect 10542 14922 10548 14924
rect 7649 14920 10548 14922
rect 7649 14864 7654 14920
rect 7710 14864 10548 14920
rect 7649 14862 10548 14864
rect 7649 14859 7715 14862
rect 10542 14860 10548 14862
rect 10612 14922 10618 14924
rect 11605 14922 11671 14925
rect 10612 14920 11671 14922
rect 10612 14864 11610 14920
rect 11666 14864 11671 14920
rect 10612 14862 11671 14864
rect 10612 14860 10618 14862
rect 11605 14859 11671 14862
rect 11830 14860 11836 14924
rect 11900 14922 11906 14924
rect 12341 14922 12407 14925
rect 11900 14920 12407 14922
rect 11900 14864 12346 14920
rect 12402 14864 12407 14920
rect 11900 14862 12407 14864
rect 11900 14860 11906 14862
rect 12341 14859 12407 14862
rect 12709 14922 12775 14925
rect 16665 14922 16731 14925
rect 12709 14920 16731 14922
rect 12709 14864 12714 14920
rect 12770 14864 16670 14920
rect 16726 14864 16731 14920
rect 12709 14862 16731 14864
rect 12709 14859 12775 14862
rect 16665 14859 16731 14862
rect 17953 14922 18019 14925
rect 22320 14922 22800 14952
rect 17953 14920 22800 14922
rect 17953 14864 17958 14920
rect 18014 14864 22800 14920
rect 17953 14862 22800 14864
rect 17953 14859 18019 14862
rect 22320 14832 22800 14862
rect 9990 14724 9996 14788
rect 10060 14786 10066 14788
rect 11145 14786 11211 14789
rect 10060 14784 11211 14786
rect 10060 14728 11150 14784
rect 11206 14728 11211 14784
rect 10060 14726 11211 14728
rect 10060 14724 10066 14726
rect 11145 14723 11211 14726
rect 11329 14786 11395 14789
rect 13537 14786 13603 14789
rect 11329 14784 13603 14786
rect 11329 14728 11334 14784
rect 11390 14728 13542 14784
rect 13598 14728 13603 14784
rect 11329 14726 13603 14728
rect 11329 14723 11395 14726
rect 13537 14723 13603 14726
rect 15510 14724 15516 14788
rect 15580 14786 15586 14788
rect 20161 14786 20227 14789
rect 15580 14784 20227 14786
rect 15580 14728 20166 14784
rect 20222 14728 20227 14784
rect 15580 14726 20227 14728
rect 15580 14724 15586 14726
rect 20161 14723 20227 14726
rect 7808 14720 8128 14721
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 2681 14650 2747 14653
rect 6913 14650 6979 14653
rect 2681 14648 6979 14650
rect 2681 14592 2686 14648
rect 2742 14592 6918 14648
rect 6974 14592 6979 14648
rect 2681 14590 6979 14592
rect 2681 14587 2747 14590
rect 6913 14587 6979 14590
rect 12014 14588 12020 14652
rect 12084 14650 12090 14652
rect 14365 14650 14431 14653
rect 12084 14648 14431 14650
rect 12084 14592 14370 14648
rect 14426 14592 14431 14648
rect 12084 14590 14431 14592
rect 12084 14588 12090 14590
rect 14365 14587 14431 14590
rect 16982 14588 16988 14652
rect 17052 14650 17058 14652
rect 18045 14650 18111 14653
rect 17052 14648 18111 14650
rect 17052 14592 18050 14648
rect 18106 14592 18111 14648
rect 17052 14590 18111 14592
rect 17052 14588 17058 14590
rect 18045 14587 18111 14590
rect 0 14514 480 14544
rect 2773 14514 2839 14517
rect 0 14512 2839 14514
rect 0 14456 2778 14512
rect 2834 14456 2839 14512
rect 0 14454 2839 14456
rect 0 14424 480 14454
rect 2773 14451 2839 14454
rect 4613 14514 4679 14517
rect 5533 14514 5599 14517
rect 4613 14512 5599 14514
rect 4613 14456 4618 14512
rect 4674 14456 5538 14512
rect 5594 14456 5599 14512
rect 4613 14454 5599 14456
rect 4613 14451 4679 14454
rect 5533 14451 5599 14454
rect 5809 14514 5875 14517
rect 7557 14514 7623 14517
rect 5809 14512 7623 14514
rect 5809 14456 5814 14512
rect 5870 14456 7562 14512
rect 7618 14456 7623 14512
rect 5809 14454 7623 14456
rect 5809 14451 5875 14454
rect 7557 14451 7623 14454
rect 7833 14514 7899 14517
rect 18638 14514 18644 14516
rect 7833 14512 18644 14514
rect 7833 14456 7838 14512
rect 7894 14456 18644 14512
rect 7833 14454 18644 14456
rect 7833 14451 7899 14454
rect 18638 14452 18644 14454
rect 18708 14452 18714 14516
rect 19241 14514 19307 14517
rect 22320 14514 22800 14544
rect 19241 14512 22800 14514
rect 19241 14456 19246 14512
rect 19302 14456 22800 14512
rect 19241 14454 22800 14456
rect 19241 14451 19307 14454
rect 22320 14424 22800 14454
rect 6637 14378 6703 14381
rect 19609 14378 19675 14381
rect 6637 14376 19675 14378
rect 6637 14320 6642 14376
rect 6698 14320 19614 14376
rect 19670 14320 19675 14376
rect 6637 14318 19675 14320
rect 6637 14315 6703 14318
rect 19609 14315 19675 14318
rect 11789 14242 11855 14245
rect 12985 14242 13051 14245
rect 11789 14240 13051 14242
rect 11789 14184 11794 14240
rect 11850 14184 12990 14240
rect 13046 14184 13051 14240
rect 11789 14182 13051 14184
rect 11789 14179 11855 14182
rect 12985 14179 13051 14182
rect 13261 14242 13327 14245
rect 13721 14242 13787 14245
rect 13261 14240 13787 14242
rect 13261 14184 13266 14240
rect 13322 14184 13726 14240
rect 13782 14184 13787 14240
rect 13261 14182 13787 14184
rect 13261 14179 13327 14182
rect 13721 14179 13787 14182
rect 13854 14180 13860 14244
rect 13924 14242 13930 14244
rect 15326 14242 15332 14244
rect 13924 14182 15332 14242
rect 13924 14180 13930 14182
rect 15326 14180 15332 14182
rect 15396 14242 15402 14244
rect 15396 14182 18016 14242
rect 15396 14180 15402 14182
rect 4376 14176 4696 14177
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 9121 14106 9187 14109
rect 11697 14106 11763 14109
rect 13905 14106 13971 14109
rect 9121 14104 9322 14106
rect 9121 14048 9126 14104
rect 9182 14048 9322 14104
rect 9121 14046 9322 14048
rect 9121 14043 9187 14046
rect 0 13970 480 14000
rect 4061 13970 4127 13973
rect 0 13968 4127 13970
rect 0 13912 4066 13968
rect 4122 13912 4127 13968
rect 0 13910 4127 13912
rect 9262 13970 9322 14046
rect 11697 14104 13971 14106
rect 11697 14048 11702 14104
rect 11758 14048 13910 14104
rect 13966 14048 13971 14104
rect 11697 14046 13971 14048
rect 11697 14043 11763 14046
rect 13905 14043 13971 14046
rect 14181 14106 14247 14109
rect 15929 14106 15995 14109
rect 14181 14104 15995 14106
rect 14181 14048 14186 14104
rect 14242 14048 15934 14104
rect 15990 14048 15995 14104
rect 14181 14046 15995 14048
rect 14181 14043 14247 14046
rect 15929 14043 15995 14046
rect 14917 13970 14983 13973
rect 15469 13970 15535 13973
rect 17166 13970 17172 13972
rect 9262 13910 12864 13970
rect 0 13880 480 13910
rect 4061 13907 4127 13910
rect 3601 13834 3667 13837
rect 7465 13834 7531 13837
rect 3601 13832 7531 13834
rect 3601 13776 3606 13832
rect 3662 13776 7470 13832
rect 7526 13776 7531 13832
rect 3601 13774 7531 13776
rect 12804 13834 12864 13910
rect 14917 13968 17172 13970
rect 14917 13912 14922 13968
rect 14978 13912 15474 13968
rect 15530 13912 17172 13968
rect 14917 13910 17172 13912
rect 14917 13907 14983 13910
rect 15469 13907 15535 13910
rect 17166 13908 17172 13910
rect 17236 13908 17242 13972
rect 17956 13970 18016 14182
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 18413 13970 18479 13973
rect 17956 13968 18479 13970
rect 17956 13912 18418 13968
rect 18474 13912 18479 13968
rect 17956 13910 18479 13912
rect 18413 13907 18479 13910
rect 18781 13970 18847 13973
rect 19609 13970 19675 13973
rect 18781 13968 19675 13970
rect 18781 13912 18786 13968
rect 18842 13912 19614 13968
rect 19670 13912 19675 13968
rect 18781 13910 19675 13912
rect 18781 13907 18847 13910
rect 19609 13907 19675 13910
rect 21357 13970 21423 13973
rect 22320 13970 22800 14000
rect 21357 13968 22800 13970
rect 21357 13912 21362 13968
rect 21418 13912 22800 13968
rect 21357 13910 22800 13912
rect 21357 13907 21423 13910
rect 22320 13880 22800 13910
rect 14181 13834 14247 13837
rect 16941 13836 17007 13837
rect 12804 13832 14247 13834
rect 12804 13776 14186 13832
rect 14242 13776 14247 13832
rect 14598 13800 15210 13834
rect 12804 13774 14247 13776
rect 3601 13771 3667 13774
rect 7465 13771 7531 13774
rect 14181 13771 14247 13774
rect 14414 13774 15210 13800
rect 14414 13740 14658 13774
rect 12249 13698 12315 13701
rect 13854 13698 13860 13700
rect 12249 13696 13860 13698
rect 12249 13640 12254 13696
rect 12310 13640 13860 13696
rect 12249 13638 13860 13640
rect 12249 13635 12315 13638
rect 13854 13636 13860 13638
rect 13924 13636 13930 13700
rect 7808 13632 8128 13633
rect 0 13562 480 13592
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 3325 13562 3391 13565
rect 0 13560 3391 13562
rect 0 13504 3330 13560
rect 3386 13504 3391 13560
rect 0 13502 3391 13504
rect 0 13472 480 13502
rect 3325 13499 3391 13502
rect 11605 13562 11671 13565
rect 12382 13562 12388 13564
rect 11605 13560 12388 13562
rect 11605 13504 11610 13560
rect 11666 13504 12388 13560
rect 11605 13502 12388 13504
rect 11605 13499 11671 13502
rect 12382 13500 12388 13502
rect 12452 13562 12458 13564
rect 14414 13562 14474 13740
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 13567 14992 13568
rect 12452 13502 14474 13562
rect 15150 13562 15210 13774
rect 16941 13832 16988 13836
rect 17052 13834 17058 13836
rect 19425 13834 19491 13837
rect 19885 13834 19951 13837
rect 16941 13776 16946 13832
rect 16941 13772 16988 13776
rect 17052 13774 17098 13834
rect 19425 13832 19951 13834
rect 19425 13776 19430 13832
rect 19486 13776 19890 13832
rect 19946 13776 19951 13832
rect 19425 13774 19951 13776
rect 17052 13772 17058 13774
rect 16941 13771 17007 13772
rect 19425 13771 19491 13774
rect 19885 13771 19951 13774
rect 16757 13698 16823 13701
rect 19558 13698 19564 13700
rect 16757 13696 19564 13698
rect 16757 13640 16762 13696
rect 16818 13640 19564 13696
rect 16757 13638 19564 13640
rect 16757 13635 16823 13638
rect 19558 13636 19564 13638
rect 19628 13636 19634 13700
rect 19374 13562 19380 13564
rect 15150 13502 19380 13562
rect 12452 13500 12458 13502
rect 17174 13429 17234 13502
rect 19374 13500 19380 13502
rect 19444 13500 19450 13564
rect 20897 13562 20963 13565
rect 22320 13562 22800 13592
rect 20897 13560 22800 13562
rect 20897 13504 20902 13560
rect 20958 13504 22800 13560
rect 20897 13502 22800 13504
rect 20897 13499 20963 13502
rect 22320 13472 22800 13502
rect 5717 13426 5783 13429
rect 16757 13426 16823 13429
rect 5717 13424 16823 13426
rect 5717 13368 5722 13424
rect 5778 13368 16762 13424
rect 16818 13368 16823 13424
rect 5717 13366 16823 13368
rect 5717 13363 5826 13366
rect 16757 13363 16823 13366
rect 17125 13424 17234 13429
rect 17125 13368 17130 13424
rect 17186 13368 17234 13424
rect 17125 13366 17234 13368
rect 17125 13363 17191 13366
rect 4376 13088 4696 13089
rect 0 13018 480 13048
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 4245 13018 4311 13021
rect 0 13016 4311 13018
rect 0 12960 4250 13016
rect 4306 12960 4311 13016
rect 0 12958 4311 12960
rect 5766 13018 5826 13363
rect 13077 13292 13143 13293
rect 13353 13292 13419 13293
rect 13721 13292 13787 13293
rect 13077 13290 13124 13292
rect 6134 13230 11714 13290
rect 13032 13288 13124 13290
rect 13032 13232 13082 13288
rect 13032 13230 13124 13232
rect 5901 13018 5967 13021
rect 5766 13016 5967 13018
rect 5766 12960 5906 13016
rect 5962 12960 5967 13016
rect 5766 12958 5967 12960
rect 0 12928 480 12958
rect 4245 12955 4311 12958
rect 5901 12955 5967 12958
rect 5257 12882 5323 12885
rect 6134 12882 6194 13230
rect 8937 13154 9003 13157
rect 9581 13154 9647 13157
rect 8937 13152 9647 13154
rect 8937 13096 8942 13152
rect 8998 13096 9586 13152
rect 9642 13096 9647 13152
rect 8937 13094 9647 13096
rect 11654 13154 11714 13230
rect 13077 13228 13124 13230
rect 13188 13228 13194 13292
rect 13302 13290 13308 13292
rect 13262 13230 13308 13290
rect 13372 13288 13419 13292
rect 13670 13290 13676 13292
rect 13414 13232 13419 13288
rect 13302 13228 13308 13230
rect 13372 13228 13419 13232
rect 13630 13230 13676 13290
rect 13740 13288 13787 13292
rect 13905 13290 13971 13293
rect 13782 13232 13787 13288
rect 13670 13228 13676 13230
rect 13740 13228 13787 13232
rect 13077 13227 13143 13228
rect 13353 13227 13419 13228
rect 13721 13227 13787 13228
rect 13862 13288 13971 13290
rect 13862 13232 13910 13288
rect 13966 13232 13971 13288
rect 13862 13227 13971 13232
rect 16205 13290 16271 13293
rect 21173 13290 21239 13293
rect 16205 13288 21239 13290
rect 16205 13232 16210 13288
rect 16266 13232 21178 13288
rect 21234 13232 21239 13288
rect 16205 13230 21239 13232
rect 16205 13227 16271 13230
rect 21173 13227 21239 13230
rect 13862 13154 13922 13227
rect 11654 13094 13922 13154
rect 16941 13154 17007 13157
rect 17166 13154 17172 13156
rect 16941 13152 17172 13154
rect 16941 13096 16946 13152
rect 17002 13096 17172 13152
rect 16941 13094 17172 13096
rect 8937 13091 9003 13094
rect 9581 13091 9647 13094
rect 16941 13091 17007 13094
rect 17166 13092 17172 13094
rect 17236 13092 17242 13156
rect 18781 13154 18847 13157
rect 19885 13154 19951 13157
rect 18781 13152 19951 13154
rect 18781 13096 18786 13152
rect 18842 13096 19890 13152
rect 19946 13096 19951 13152
rect 18781 13094 19951 13096
rect 18781 13091 18847 13094
rect 19885 13091 19951 13094
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 7557 13018 7623 13021
rect 10317 13020 10383 13021
rect 8518 13018 8524 13020
rect 7557 13016 8524 13018
rect 7557 12960 7562 13016
rect 7618 12960 8524 13016
rect 7557 12958 8524 12960
rect 7557 12955 7623 12958
rect 8518 12956 8524 12958
rect 8588 12956 8594 13020
rect 10317 13018 10364 13020
rect 10272 13016 10364 13018
rect 10272 12960 10322 13016
rect 10272 12958 10364 12960
rect 10317 12956 10364 12958
rect 10428 12956 10434 13020
rect 12801 13018 12867 13021
rect 15142 13018 15148 13020
rect 12801 13016 15148 13018
rect 12801 12960 12806 13016
rect 12862 12960 15148 13016
rect 12801 12958 15148 12960
rect 10317 12955 10383 12956
rect 12801 12955 12867 12958
rect 15142 12956 15148 12958
rect 15212 13018 15218 13020
rect 17217 13018 17283 13021
rect 15212 13016 17283 13018
rect 15212 12960 17222 13016
rect 17278 12960 17283 13016
rect 15212 12958 17283 12960
rect 15212 12956 15218 12958
rect 17217 12955 17283 12958
rect 18873 13018 18939 13021
rect 19333 13020 19399 13021
rect 19006 13018 19012 13020
rect 18873 13016 19012 13018
rect 18873 12960 18878 13016
rect 18934 12960 19012 13016
rect 18873 12958 19012 12960
rect 18873 12955 18939 12958
rect 19006 12956 19012 12958
rect 19076 12956 19082 13020
rect 19333 13016 19380 13020
rect 19444 13018 19450 13020
rect 22320 13018 22800 13048
rect 19333 12960 19338 13016
rect 19333 12956 19380 12960
rect 19444 12958 19490 13018
rect 20118 12958 22800 13018
rect 19444 12956 19450 12958
rect 19333 12955 19399 12956
rect 5257 12880 6194 12882
rect 5257 12824 5262 12880
rect 5318 12824 6194 12880
rect 5257 12822 6194 12824
rect 10409 12882 10475 12885
rect 12249 12884 12315 12885
rect 13169 12884 13235 12885
rect 12198 12882 12204 12884
rect 10409 12880 12204 12882
rect 12268 12880 12315 12884
rect 10409 12824 10414 12880
rect 10470 12824 12204 12880
rect 12310 12824 12315 12880
rect 10409 12822 12204 12824
rect 5257 12819 5323 12822
rect 10409 12819 10475 12822
rect 12198 12820 12204 12822
rect 12268 12820 12315 12824
rect 13118 12820 13124 12884
rect 13188 12882 13235 12884
rect 19885 12882 19951 12885
rect 13188 12880 13280 12882
rect 13230 12824 13280 12880
rect 13188 12822 13280 12824
rect 13356 12880 19951 12882
rect 13356 12824 19890 12880
rect 19946 12824 19951 12880
rect 13356 12822 19951 12824
rect 13188 12820 13235 12822
rect 12249 12819 12315 12820
rect 13169 12819 13235 12820
rect 5441 12746 5507 12749
rect 4662 12744 5507 12746
rect 4662 12688 5446 12744
rect 5502 12688 5507 12744
rect 4662 12686 5507 12688
rect 0 12610 480 12640
rect 4662 12613 4722 12686
rect 5441 12683 5507 12686
rect 6361 12746 6427 12749
rect 9438 12746 9444 12748
rect 6361 12744 9444 12746
rect 6361 12688 6366 12744
rect 6422 12688 9444 12744
rect 6361 12686 9444 12688
rect 6361 12683 6427 12686
rect 9438 12684 9444 12686
rect 9508 12746 9514 12748
rect 10317 12746 10383 12749
rect 11697 12748 11763 12749
rect 9508 12744 10383 12746
rect 9508 12688 10322 12744
rect 10378 12688 10383 12744
rect 9508 12686 10383 12688
rect 9508 12684 9514 12686
rect 10317 12683 10383 12686
rect 11646 12684 11652 12748
rect 11716 12746 11763 12748
rect 11716 12744 11808 12746
rect 11758 12688 11808 12744
rect 11716 12686 11808 12688
rect 11716 12684 11763 12686
rect 11697 12683 11763 12684
rect 3969 12610 4035 12613
rect 0 12608 4035 12610
rect 0 12552 3974 12608
rect 4030 12552 4035 12608
rect 0 12550 4035 12552
rect 4662 12608 4771 12613
rect 4662 12552 4710 12608
rect 4766 12552 4771 12608
rect 4662 12550 4771 12552
rect 0 12520 480 12550
rect 3969 12547 4035 12550
rect 4705 12547 4771 12550
rect 4838 12548 4844 12612
rect 4908 12610 4914 12612
rect 5257 12610 5323 12613
rect 4908 12608 5323 12610
rect 4908 12552 5262 12608
rect 5318 12552 5323 12608
rect 4908 12550 5323 12552
rect 4908 12548 4914 12550
rect 5257 12547 5323 12550
rect 8293 12610 8359 12613
rect 11830 12610 11836 12612
rect 8293 12608 11836 12610
rect 8293 12552 8298 12608
rect 8354 12552 11836 12608
rect 8293 12550 11836 12552
rect 8293 12547 8359 12550
rect 11830 12548 11836 12550
rect 11900 12548 11906 12612
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 9213 12474 9279 12477
rect 9622 12474 9628 12476
rect 9213 12472 9628 12474
rect 9213 12416 9218 12472
rect 9274 12416 9628 12472
rect 9213 12414 9628 12416
rect 9213 12411 9279 12414
rect 9622 12412 9628 12414
rect 9692 12474 9698 12476
rect 13356 12474 13416 12822
rect 19885 12819 19951 12822
rect 13537 12746 13603 12749
rect 13670 12746 13676 12748
rect 13537 12744 13676 12746
rect 13537 12688 13542 12744
rect 13598 12688 13676 12744
rect 13537 12686 13676 12688
rect 13537 12683 13603 12686
rect 13670 12684 13676 12686
rect 13740 12684 13746 12748
rect 14181 12746 14247 12749
rect 14641 12746 14707 12749
rect 14181 12744 14707 12746
rect 14181 12688 14186 12744
rect 14242 12688 14646 12744
rect 14702 12688 14707 12744
rect 14181 12686 14707 12688
rect 14181 12683 14247 12686
rect 14641 12683 14707 12686
rect 14917 12746 14983 12749
rect 20118 12746 20178 12958
rect 22320 12928 22800 12958
rect 14917 12744 20178 12746
rect 14917 12688 14922 12744
rect 14978 12688 20178 12744
rect 14917 12686 20178 12688
rect 14917 12683 14983 12686
rect 15101 12612 15167 12613
rect 15101 12608 15148 12612
rect 15212 12610 15218 12612
rect 15101 12552 15106 12608
rect 15101 12548 15148 12552
rect 15212 12550 15258 12610
rect 15212 12548 15218 12550
rect 15101 12547 15167 12548
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 9692 12414 13416 12474
rect 15101 12474 15167 12477
rect 15334 12474 15394 12686
rect 17309 12612 17375 12613
rect 17585 12612 17651 12613
rect 17309 12610 17356 12612
rect 17264 12608 17356 12610
rect 17264 12552 17314 12608
rect 17264 12550 17356 12552
rect 17309 12548 17356 12550
rect 17420 12548 17426 12612
rect 17534 12610 17540 12612
rect 17494 12550 17540 12610
rect 17604 12608 17651 12612
rect 17769 12610 17835 12613
rect 17646 12552 17651 12608
rect 17534 12548 17540 12550
rect 17604 12548 17651 12552
rect 17309 12547 17375 12548
rect 17585 12547 17651 12548
rect 17726 12608 17835 12610
rect 17726 12552 17774 12608
rect 17830 12552 17835 12608
rect 17726 12547 17835 12552
rect 18689 12610 18755 12613
rect 19149 12610 19215 12613
rect 18689 12608 19215 12610
rect 18689 12552 18694 12608
rect 18750 12552 19154 12608
rect 19210 12552 19215 12608
rect 18689 12550 19215 12552
rect 18689 12547 18755 12550
rect 19149 12547 19215 12550
rect 19885 12610 19951 12613
rect 22320 12610 22800 12640
rect 19885 12608 22800 12610
rect 19885 12552 19890 12608
rect 19946 12552 22800 12608
rect 19885 12550 22800 12552
rect 19885 12547 19951 12550
rect 15101 12472 15394 12474
rect 15101 12416 15106 12472
rect 15162 12416 15394 12472
rect 15101 12414 15394 12416
rect 16941 12474 17007 12477
rect 17726 12474 17786 12547
rect 22320 12520 22800 12550
rect 16941 12472 17786 12474
rect 16941 12416 16946 12472
rect 17002 12416 17786 12472
rect 16941 12414 17786 12416
rect 18321 12474 18387 12477
rect 19149 12474 19215 12477
rect 18321 12472 19215 12474
rect 18321 12416 18326 12472
rect 18382 12416 19154 12472
rect 19210 12416 19215 12472
rect 18321 12414 19215 12416
rect 9692 12412 9698 12414
rect 15101 12411 15167 12414
rect 16941 12411 17007 12414
rect 18321 12411 18387 12414
rect 19149 12411 19215 12414
rect 8385 12338 8451 12341
rect 11513 12338 11579 12341
rect 8385 12336 11579 12338
rect 8385 12280 8390 12336
rect 8446 12280 11518 12336
rect 11574 12280 11579 12336
rect 8385 12278 11579 12280
rect 8385 12275 8451 12278
rect 11513 12275 11579 12278
rect 11646 12276 11652 12340
rect 11716 12338 11722 12340
rect 16614 12338 16620 12340
rect 11716 12278 16620 12338
rect 11716 12276 11722 12278
rect 16614 12276 16620 12278
rect 16684 12276 16690 12340
rect 17585 12338 17651 12341
rect 19190 12338 19196 12340
rect 17585 12336 19196 12338
rect 17585 12280 17590 12336
rect 17646 12280 19196 12336
rect 17585 12278 19196 12280
rect 17585 12275 17651 12278
rect 19190 12276 19196 12278
rect 19260 12276 19266 12340
rect 7925 12202 7991 12205
rect 4248 12200 7991 12202
rect 4248 12144 7930 12200
rect 7986 12144 7991 12200
rect 4248 12142 7991 12144
rect 0 12066 480 12096
rect 4248 12066 4308 12142
rect 7925 12139 7991 12142
rect 9305 12202 9371 12205
rect 11881 12204 11947 12205
rect 9305 12200 11760 12202
rect 9305 12144 9310 12200
rect 9366 12144 11760 12200
rect 9305 12142 11760 12144
rect 9305 12139 9371 12142
rect 0 12006 4308 12066
rect 0 11976 480 12006
rect 9254 12004 9260 12068
rect 9324 12066 9330 12068
rect 9673 12066 9739 12069
rect 9324 12064 9739 12066
rect 9324 12008 9678 12064
rect 9734 12008 9739 12064
rect 9324 12006 9739 12008
rect 9324 12004 9330 12006
rect 9673 12003 9739 12006
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 6126 11868 6132 11932
rect 6196 11930 6202 11932
rect 6545 11930 6611 11933
rect 10910 11930 10916 11932
rect 6196 11928 10916 11930
rect 6196 11872 6550 11928
rect 6606 11872 10916 11928
rect 6196 11870 10916 11872
rect 6196 11868 6202 11870
rect 6545 11867 6611 11870
rect 10910 11868 10916 11870
rect 10980 11868 10986 11932
rect 11700 11930 11760 12142
rect 11830 12140 11836 12204
rect 11900 12202 11947 12204
rect 12065 12202 12131 12205
rect 11900 12200 11992 12202
rect 11942 12144 11992 12200
rect 11900 12142 11992 12144
rect 12065 12200 18706 12202
rect 12065 12144 12070 12200
rect 12126 12144 18706 12200
rect 12065 12142 18706 12144
rect 11900 12140 11947 12142
rect 11881 12139 11947 12140
rect 12065 12139 12131 12142
rect 12709 12066 12775 12069
rect 13077 12066 13143 12069
rect 13445 12068 13511 12069
rect 13445 12066 13492 12068
rect 12709 12064 13143 12066
rect 12709 12008 12714 12064
rect 12770 12008 13082 12064
rect 13138 12008 13143 12064
rect 12709 12006 13143 12008
rect 13400 12064 13492 12066
rect 13400 12008 13450 12064
rect 13400 12006 13492 12008
rect 12709 12003 12775 12006
rect 13077 12003 13143 12006
rect 13445 12004 13492 12006
rect 13556 12004 13562 12068
rect 14181 12066 14247 12069
rect 14641 12066 14707 12069
rect 16205 12066 16271 12069
rect 14181 12064 16271 12066
rect 14181 12008 14186 12064
rect 14242 12008 14646 12064
rect 14702 12008 16210 12064
rect 16266 12008 16271 12064
rect 14181 12006 16271 12008
rect 18646 12066 18706 12142
rect 22320 12066 22800 12096
rect 18646 12006 22800 12066
rect 13445 12003 13511 12004
rect 14181 12003 14247 12006
rect 14641 12003 14707 12006
rect 16205 12003 16271 12006
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 22320 11976 22800 12006
rect 18104 11935 18424 11936
rect 11700 11870 17786 11930
rect 3509 11794 3575 11797
rect 8753 11794 8819 11797
rect 3509 11792 8819 11794
rect 3509 11736 3514 11792
rect 3570 11736 8758 11792
rect 8814 11736 8819 11792
rect 3509 11734 8819 11736
rect 3509 11731 3575 11734
rect 8753 11731 8819 11734
rect 11329 11794 11395 11797
rect 12065 11794 12131 11797
rect 11329 11792 12131 11794
rect 11329 11736 11334 11792
rect 11390 11736 12070 11792
rect 12126 11736 12131 11792
rect 11329 11734 12131 11736
rect 11329 11731 11395 11734
rect 12065 11731 12131 11734
rect 12249 11794 12315 11797
rect 15469 11794 15535 11797
rect 16849 11794 16915 11797
rect 17585 11796 17651 11797
rect 17534 11794 17540 11796
rect 12249 11792 15394 11794
rect 12249 11736 12254 11792
rect 12310 11736 15394 11792
rect 12249 11734 15394 11736
rect 12249 11731 12315 11734
rect 0 11658 480 11688
rect 12014 11658 12020 11660
rect 0 11598 12020 11658
rect 0 11568 480 11598
rect 12014 11596 12020 11598
rect 12084 11596 12090 11660
rect 13118 11596 13124 11660
rect 13188 11658 13194 11660
rect 15334 11658 15394 11734
rect 15469 11792 16915 11794
rect 15469 11736 15474 11792
rect 15530 11736 16854 11792
rect 16910 11736 16915 11792
rect 15469 11734 16915 11736
rect 17494 11734 17540 11794
rect 17604 11792 17651 11796
rect 17646 11736 17651 11792
rect 15469 11731 15535 11734
rect 16849 11731 16915 11734
rect 17534 11732 17540 11734
rect 17604 11732 17651 11736
rect 17726 11794 17786 11870
rect 19793 11794 19859 11797
rect 17726 11792 19859 11794
rect 17726 11736 19798 11792
rect 19854 11736 19859 11792
rect 17726 11734 19859 11736
rect 17585 11731 17651 11732
rect 19793 11731 19859 11734
rect 17677 11658 17743 11661
rect 22320 11658 22800 11688
rect 13188 11598 15164 11658
rect 15334 11656 17743 11658
rect 15334 11600 17682 11656
rect 17738 11600 17743 11656
rect 15334 11598 17743 11600
rect 13188 11596 13194 11598
rect 4102 11460 4108 11524
rect 4172 11522 4178 11524
rect 4245 11522 4311 11525
rect 4172 11520 4311 11522
rect 4172 11464 4250 11520
rect 4306 11464 4311 11520
rect 4172 11462 4311 11464
rect 4172 11460 4178 11462
rect 4245 11459 4311 11462
rect 8753 11522 8819 11525
rect 11646 11522 11652 11524
rect 8753 11520 11652 11522
rect 8753 11464 8758 11520
rect 8814 11464 11652 11520
rect 8753 11462 11652 11464
rect 8753 11459 8819 11462
rect 11646 11460 11652 11462
rect 11716 11460 11722 11524
rect 12934 11460 12940 11524
rect 13004 11522 13010 11524
rect 13261 11522 13327 11525
rect 13004 11520 13327 11522
rect 13004 11464 13266 11520
rect 13322 11464 13327 11520
rect 13004 11462 13327 11464
rect 15104 11522 15164 11598
rect 17677 11595 17743 11598
rect 20118 11598 22800 11658
rect 20118 11522 20178 11598
rect 22320 11568 22800 11598
rect 15104 11462 20178 11522
rect 13004 11460 13010 11462
rect 13261 11459 13327 11462
rect 7808 11456 8128 11457
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 3877 11386 3943 11389
rect 5390 11386 5396 11388
rect 3877 11384 5396 11386
rect 3877 11328 3882 11384
rect 3938 11328 5396 11384
rect 3877 11326 5396 11328
rect 3877 11323 3943 11326
rect 5390 11324 5396 11326
rect 5460 11324 5466 11388
rect 10358 11324 10364 11388
rect 10428 11386 10434 11388
rect 14181 11386 14247 11389
rect 10428 11384 14247 11386
rect 10428 11328 14186 11384
rect 14242 11328 14247 11384
rect 10428 11326 14247 11328
rect 10428 11324 10434 11326
rect 14181 11323 14247 11326
rect 15878 11324 15884 11388
rect 15948 11386 15954 11388
rect 16297 11386 16363 11389
rect 15948 11384 16363 11386
rect 15948 11328 16302 11384
rect 16358 11328 16363 11384
rect 15948 11326 16363 11328
rect 15948 11324 15954 11326
rect 16297 11323 16363 11326
rect 18781 11386 18847 11389
rect 21357 11386 21423 11389
rect 18781 11384 21423 11386
rect 18781 11328 18786 11384
rect 18842 11328 21362 11384
rect 21418 11328 21423 11384
rect 18781 11326 21423 11328
rect 18781 11323 18847 11326
rect 21357 11323 21423 11326
rect 5165 11250 5231 11253
rect 17677 11250 17743 11253
rect 4708 11248 17743 11250
rect 4708 11192 5170 11248
rect 5226 11192 17682 11248
rect 17738 11192 17743 11248
rect 4708 11190 17743 11192
rect 0 11114 480 11144
rect 4708 11114 4768 11190
rect 5165 11187 5231 11190
rect 17677 11187 17743 11190
rect 0 11054 4768 11114
rect 0 11024 480 11054
rect 10910 11052 10916 11116
rect 10980 11114 10986 11116
rect 15377 11114 15443 11117
rect 15510 11114 15516 11116
rect 10980 11054 13186 11114
rect 10980 11052 10986 11054
rect 4376 10912 4696 10913
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 5390 10780 5396 10844
rect 5460 10842 5466 10844
rect 9581 10842 9647 10845
rect 5460 10840 9647 10842
rect 5460 10784 9586 10840
rect 9642 10784 9647 10840
rect 5460 10782 9647 10784
rect 5460 10780 5466 10782
rect 9581 10779 9647 10782
rect 12617 10842 12683 10845
rect 12985 10842 13051 10845
rect 12617 10840 13051 10842
rect 12617 10784 12622 10840
rect 12678 10784 12990 10840
rect 13046 10784 13051 10840
rect 12617 10782 13051 10784
rect 13126 10842 13186 11054
rect 15377 11112 15516 11114
rect 15377 11056 15382 11112
rect 15438 11056 15516 11112
rect 15377 11054 15516 11056
rect 15377 11051 15443 11054
rect 15510 11052 15516 11054
rect 15580 11114 15586 11116
rect 17309 11114 17375 11117
rect 15580 11112 17375 11114
rect 15580 11056 17314 11112
rect 17370 11056 17375 11112
rect 15580 11054 17375 11056
rect 15580 11052 15586 11054
rect 17309 11051 17375 11054
rect 18822 11052 18828 11116
rect 18892 11114 18898 11116
rect 22320 11114 22800 11144
rect 18892 11054 22800 11114
rect 18892 11052 18898 11054
rect 22320 11024 22800 11054
rect 13302 10916 13308 10980
rect 13372 10978 13378 10980
rect 13997 10978 14063 10981
rect 13372 10976 14063 10978
rect 13372 10920 14002 10976
rect 14058 10920 14063 10976
rect 13372 10918 14063 10920
rect 13372 10916 13378 10918
rect 13997 10915 14063 10918
rect 14641 10978 14707 10981
rect 15745 10978 15811 10981
rect 14641 10976 15811 10978
rect 14641 10920 14646 10976
rect 14702 10920 15750 10976
rect 15806 10920 15811 10976
rect 14641 10918 15811 10920
rect 14641 10915 14707 10918
rect 15745 10915 15811 10918
rect 16481 10978 16547 10981
rect 17033 10978 17099 10981
rect 16481 10976 17099 10978
rect 16481 10920 16486 10976
rect 16542 10920 17038 10976
rect 17094 10920 17099 10976
rect 16481 10918 17099 10920
rect 16481 10915 16547 10918
rect 17033 10915 17099 10918
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 16021 10842 16087 10845
rect 13126 10840 16087 10842
rect 13126 10784 16026 10840
rect 16082 10784 16087 10840
rect 13126 10782 16087 10784
rect 12617 10779 12683 10782
rect 12985 10779 13051 10782
rect 16021 10779 16087 10782
rect 0 10706 480 10736
rect 6637 10706 6703 10709
rect 8845 10708 8911 10709
rect 8845 10706 8892 10708
rect 0 10704 6703 10706
rect 0 10648 6642 10704
rect 6698 10648 6703 10704
rect 0 10646 6703 10648
rect 8800 10704 8892 10706
rect 8800 10648 8850 10704
rect 8800 10646 8892 10648
rect 0 10616 480 10646
rect 6637 10643 6703 10646
rect 8845 10644 8892 10646
rect 8956 10644 8962 10708
rect 10409 10706 10475 10709
rect 11830 10706 11836 10708
rect 10409 10704 11836 10706
rect 10409 10648 10414 10704
rect 10470 10648 11836 10704
rect 10409 10646 11836 10648
rect 8845 10643 8911 10644
rect 10409 10643 10475 10646
rect 11830 10644 11836 10646
rect 11900 10644 11906 10708
rect 12985 10706 13051 10709
rect 13905 10706 13971 10709
rect 12985 10704 13971 10706
rect 12985 10648 12990 10704
rect 13046 10648 13910 10704
rect 13966 10648 13971 10704
rect 12985 10646 13971 10648
rect 12985 10643 13051 10646
rect 13905 10643 13971 10646
rect 14181 10706 14247 10709
rect 16982 10706 16988 10708
rect 14181 10704 16988 10706
rect 14181 10648 14186 10704
rect 14242 10648 16988 10704
rect 14181 10646 16988 10648
rect 14181 10643 14247 10646
rect 16982 10644 16988 10646
rect 17052 10644 17058 10708
rect 17217 10706 17283 10709
rect 22320 10706 22800 10736
rect 17217 10704 22800 10706
rect 17217 10648 17222 10704
rect 17278 10648 22800 10704
rect 17217 10646 22800 10648
rect 17217 10643 17283 10646
rect 22320 10616 22800 10646
rect 8109 10570 8175 10573
rect 9990 10570 9996 10572
rect 8109 10568 9996 10570
rect 8109 10512 8114 10568
rect 8170 10512 9996 10568
rect 8109 10510 9996 10512
rect 8109 10507 8175 10510
rect 9990 10508 9996 10510
rect 10060 10570 10066 10572
rect 13302 10570 13308 10572
rect 10060 10510 13308 10570
rect 10060 10508 10066 10510
rect 13302 10508 13308 10510
rect 13372 10508 13378 10572
rect 15009 10570 15075 10573
rect 16757 10570 16823 10573
rect 15009 10568 16823 10570
rect 15009 10512 15014 10568
rect 15070 10512 16762 10568
rect 16818 10512 16823 10568
rect 15009 10510 16823 10512
rect 15009 10507 15075 10510
rect 16757 10507 16823 10510
rect 18781 10568 18847 10573
rect 18781 10512 18786 10568
rect 18842 10512 18847 10568
rect 18781 10507 18847 10512
rect 9305 10434 9371 10437
rect 11053 10434 11119 10437
rect 9305 10432 11119 10434
rect 9305 10376 9310 10432
rect 9366 10376 11058 10432
rect 11114 10376 11119 10432
rect 9305 10374 11119 10376
rect 9305 10371 9371 10374
rect 11053 10371 11119 10374
rect 12249 10434 12315 10437
rect 12934 10434 12940 10436
rect 12249 10432 12940 10434
rect 12249 10376 12254 10432
rect 12310 10376 12940 10432
rect 12249 10374 12940 10376
rect 12249 10371 12315 10374
rect 12934 10372 12940 10374
rect 13004 10372 13010 10436
rect 15745 10434 15811 10437
rect 18784 10434 18844 10507
rect 15745 10432 18844 10434
rect 15745 10376 15750 10432
rect 15806 10376 18844 10432
rect 15745 10374 18844 10376
rect 15745 10371 15811 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 10303 14992 10304
rect 10174 10236 10180 10300
rect 10244 10298 10250 10300
rect 10685 10298 10751 10301
rect 10244 10296 10751 10298
rect 10244 10240 10690 10296
rect 10746 10240 10751 10296
rect 10244 10238 10751 10240
rect 10244 10236 10250 10238
rect 10685 10235 10751 10238
rect 10869 10298 10935 10301
rect 14181 10298 14247 10301
rect 10869 10296 14247 10298
rect 10869 10240 10874 10296
rect 10930 10240 14186 10296
rect 14242 10240 14247 10296
rect 10869 10238 14247 10240
rect 10869 10235 10935 10238
rect 14181 10235 14247 10238
rect 15193 10298 15259 10301
rect 17309 10298 17375 10301
rect 15193 10296 17375 10298
rect 15193 10240 15198 10296
rect 15254 10240 17314 10296
rect 17370 10240 17375 10296
rect 15193 10238 17375 10240
rect 15193 10235 15259 10238
rect 17309 10235 17375 10238
rect 0 10162 480 10192
rect 7414 10162 7420 10164
rect 0 10102 7420 10162
rect 0 10072 480 10102
rect 7414 10100 7420 10102
rect 7484 10162 7490 10164
rect 9765 10162 9831 10165
rect 10225 10162 10291 10165
rect 15837 10162 15903 10165
rect 22320 10162 22800 10192
rect 7484 10102 7712 10162
rect 7484 10100 7490 10102
rect 7652 10029 7712 10102
rect 9765 10160 18752 10162
rect 9765 10104 9770 10160
rect 9826 10104 10230 10160
rect 10286 10104 15842 10160
rect 15898 10104 18752 10160
rect 9765 10102 18752 10104
rect 9765 10099 9831 10102
rect 10225 10099 10291 10102
rect 15837 10099 15903 10102
rect 6085 10028 6151 10029
rect 6085 10026 6132 10028
rect 6040 10024 6132 10026
rect 6040 9968 6090 10024
rect 6040 9966 6132 9968
rect 6085 9964 6132 9966
rect 6196 9964 6202 10028
rect 7649 10024 7715 10029
rect 7649 9968 7654 10024
rect 7710 9968 7715 10024
rect 6085 9963 6151 9964
rect 7649 9963 7715 9968
rect 8569 10026 8635 10029
rect 16757 10026 16823 10029
rect 8569 10024 16823 10026
rect 8569 9968 8574 10024
rect 8630 9968 16762 10024
rect 16818 9968 16823 10024
rect 8569 9966 16823 9968
rect 8569 9963 8635 9966
rect 16070 9893 16130 9966
rect 16757 9963 16823 9966
rect 17309 10028 17375 10029
rect 17309 10024 17356 10028
rect 17420 10026 17426 10028
rect 18413 10026 18479 10029
rect 17309 9968 17314 10024
rect 17309 9964 17356 9968
rect 17420 9966 17466 10026
rect 17956 10024 18479 10026
rect 17956 9968 18418 10024
rect 18474 9968 18479 10024
rect 17956 9966 18479 9968
rect 17420 9964 17426 9966
rect 17309 9963 17375 9964
rect 12801 9892 12867 9893
rect 12750 9890 12756 9892
rect 11654 9830 12756 9890
rect 12820 9890 12867 9892
rect 12820 9888 12912 9890
rect 12862 9832 12912 9888
rect 4376 9824 4696 9825
rect 0 9754 480 9784
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 3877 9754 3943 9757
rect 0 9752 3943 9754
rect 0 9696 3882 9752
rect 3938 9696 3943 9752
rect 0 9694 3943 9696
rect 0 9664 480 9694
rect 3877 9691 3943 9694
rect 10409 9754 10475 9757
rect 10542 9754 10548 9756
rect 10409 9752 10548 9754
rect 10409 9696 10414 9752
rect 10470 9696 10548 9752
rect 10409 9694 10548 9696
rect 10409 9691 10475 9694
rect 10542 9692 10548 9694
rect 10612 9692 10618 9756
rect 10542 9556 10548 9620
rect 10612 9618 10618 9620
rect 11654 9618 11714 9830
rect 12750 9828 12756 9830
rect 12820 9830 12912 9832
rect 12820 9828 12867 9830
rect 15326 9828 15332 9892
rect 15396 9890 15402 9892
rect 15929 9890 15995 9893
rect 15396 9888 15995 9890
rect 15396 9832 15934 9888
rect 15990 9832 15995 9888
rect 15396 9830 15995 9832
rect 16070 9888 16179 9893
rect 16070 9832 16118 9888
rect 16174 9832 16179 9888
rect 16070 9830 16179 9832
rect 15396 9828 15402 9830
rect 12801 9827 12867 9828
rect 15929 9827 15995 9830
rect 16113 9827 16179 9830
rect 17166 9828 17172 9892
rect 17236 9890 17242 9892
rect 17401 9890 17467 9893
rect 17236 9888 17467 9890
rect 17236 9832 17406 9888
rect 17462 9832 17467 9888
rect 17236 9830 17467 9832
rect 17236 9828 17242 9830
rect 17401 9827 17467 9830
rect 11830 9692 11836 9756
rect 11900 9754 11906 9756
rect 12750 9754 12756 9756
rect 11900 9694 12756 9754
rect 11900 9692 11906 9694
rect 12750 9692 12756 9694
rect 12820 9692 12826 9756
rect 12934 9692 12940 9756
rect 13004 9754 13010 9756
rect 16389 9754 16455 9757
rect 17956 9754 18016 9966
rect 18413 9963 18479 9966
rect 18692 9890 18752 10102
rect 18876 10102 22800 10162
rect 18876 10029 18936 10102
rect 22320 10072 22800 10102
rect 18873 10024 18939 10029
rect 18873 9968 18878 10024
rect 18934 9968 18939 10024
rect 18873 9963 18939 9968
rect 19333 10028 19399 10029
rect 19333 10024 19380 10028
rect 19444 10026 19450 10028
rect 19333 9968 19338 10024
rect 19333 9964 19380 9968
rect 19444 9966 19490 10026
rect 19444 9964 19450 9966
rect 19333 9963 19399 9964
rect 18692 9830 19626 9890
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 13004 9752 18016 9754
rect 13004 9696 16394 9752
rect 16450 9696 18016 9752
rect 13004 9694 18016 9696
rect 19566 9754 19626 9830
rect 22320 9754 22800 9784
rect 19566 9694 22800 9754
rect 13004 9692 13010 9694
rect 16389 9691 16455 9694
rect 22320 9664 22800 9694
rect 10612 9558 11714 9618
rect 10612 9556 10618 9558
rect 12750 9556 12756 9620
rect 12820 9618 12826 9620
rect 18873 9618 18939 9621
rect 12820 9616 18939 9618
rect 12820 9560 18878 9616
rect 18934 9560 18939 9616
rect 12820 9558 18939 9560
rect 12820 9556 12826 9558
rect 18873 9555 18939 9558
rect 11053 9482 11119 9485
rect 15377 9482 15443 9485
rect 11053 9480 15443 9482
rect 11053 9424 11058 9480
rect 11114 9424 15382 9480
rect 15438 9424 15443 9480
rect 11053 9422 15443 9424
rect 11053 9419 11119 9422
rect 15377 9419 15443 9422
rect 18781 9482 18847 9485
rect 19190 9482 19196 9484
rect 18781 9480 19196 9482
rect 18781 9424 18786 9480
rect 18842 9424 19196 9480
rect 18781 9422 19196 9424
rect 18781 9419 18847 9422
rect 19190 9420 19196 9422
rect 19260 9420 19266 9484
rect 11237 9346 11303 9349
rect 12014 9346 12020 9348
rect 11237 9344 12020 9346
rect 11237 9288 11242 9344
rect 11298 9288 12020 9344
rect 11237 9286 12020 9288
rect 11237 9283 11303 9286
rect 12014 9284 12020 9286
rect 12084 9284 12090 9348
rect 15142 9284 15148 9348
rect 15212 9346 15218 9348
rect 19333 9346 19399 9349
rect 15212 9344 19399 9346
rect 15212 9288 19338 9344
rect 19394 9288 19399 9344
rect 15212 9286 19399 9288
rect 15212 9284 15218 9286
rect 19333 9283 19399 9286
rect 7808 9280 8128 9281
rect 0 9210 480 9240
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 14457 9210 14523 9213
rect 0 9150 4906 9210
rect 0 9120 480 9150
rect 4846 8938 4906 9150
rect 10964 9208 14523 9210
rect 10964 9152 14462 9208
rect 14518 9152 14523 9208
rect 10964 9150 14523 9152
rect 6361 9074 6427 9077
rect 10964 9074 11024 9150
rect 14457 9147 14523 9150
rect 17350 9148 17356 9212
rect 17420 9210 17426 9212
rect 17861 9210 17927 9213
rect 22320 9210 22800 9240
rect 17420 9208 17927 9210
rect 17420 9152 17866 9208
rect 17922 9152 17927 9208
rect 19382 9176 22800 9210
rect 17420 9150 17927 9152
rect 17420 9148 17426 9150
rect 17861 9147 17927 9150
rect 19198 9150 22800 9176
rect 19198 9116 19442 9150
rect 22320 9120 22800 9150
rect 6361 9072 11024 9074
rect 6361 9016 6366 9072
rect 6422 9016 11024 9072
rect 6361 9014 11024 9016
rect 12065 9074 12131 9077
rect 19198 9074 19258 9116
rect 12065 9072 19258 9074
rect 12065 9016 12070 9072
rect 12126 9016 19258 9072
rect 12065 9014 19258 9016
rect 6361 9011 6427 9014
rect 12065 9011 12131 9014
rect 9121 8938 9187 8941
rect 4846 8936 9187 8938
rect 4846 8880 9126 8936
rect 9182 8880 9187 8936
rect 4846 8878 9187 8880
rect 9121 8875 9187 8878
rect 10501 8938 10567 8941
rect 12249 8938 12315 8941
rect 12433 8938 12499 8941
rect 13862 8940 13922 9014
rect 10501 8936 12082 8938
rect 10501 8880 10506 8936
rect 10562 8880 12082 8936
rect 10501 8878 12082 8880
rect 10501 8875 10567 8878
rect 0 8802 480 8832
rect 4061 8802 4127 8805
rect 0 8800 4127 8802
rect 0 8744 4066 8800
rect 4122 8744 4127 8800
rect 0 8742 4127 8744
rect 0 8712 480 8742
rect 4061 8739 4127 8742
rect 6545 8802 6611 8805
rect 7465 8802 7531 8805
rect 8845 8802 8911 8805
rect 6545 8800 8911 8802
rect 6545 8744 6550 8800
rect 6606 8744 7470 8800
rect 7526 8744 8850 8800
rect 8906 8744 8911 8800
rect 6545 8742 8911 8744
rect 6545 8739 6611 8742
rect 7465 8739 7531 8742
rect 8845 8739 8911 8742
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 6361 8666 6427 8669
rect 9857 8666 9923 8669
rect 6361 8664 9923 8666
rect 6361 8608 6366 8664
rect 6422 8608 9862 8664
rect 9918 8608 9923 8664
rect 6361 8606 9923 8608
rect 12022 8666 12082 8878
rect 12249 8936 12499 8938
rect 12249 8880 12254 8936
rect 12310 8880 12438 8936
rect 12494 8880 12499 8936
rect 12249 8878 12499 8880
rect 12249 8875 12315 8878
rect 12433 8875 12499 8878
rect 13854 8876 13860 8940
rect 13924 8876 13930 8940
rect 14457 8938 14523 8941
rect 17309 8938 17375 8941
rect 19241 8938 19307 8941
rect 14457 8936 19307 8938
rect 14457 8880 14462 8936
rect 14518 8880 17314 8936
rect 17370 8880 19246 8936
rect 19302 8880 19307 8936
rect 14457 8878 19307 8880
rect 14457 8875 14523 8878
rect 17309 8875 17375 8878
rect 19241 8875 19307 8878
rect 12433 8802 12499 8805
rect 13118 8802 13124 8804
rect 12433 8800 13124 8802
rect 12433 8744 12438 8800
rect 12494 8744 13124 8800
rect 12433 8742 13124 8744
rect 12433 8739 12499 8742
rect 13118 8740 13124 8742
rect 13188 8740 13194 8804
rect 15745 8802 15811 8805
rect 16297 8804 16363 8805
rect 14782 8800 15811 8802
rect 14782 8744 15750 8800
rect 15806 8744 15811 8800
rect 14782 8742 15811 8744
rect 14782 8666 14842 8742
rect 15745 8739 15811 8742
rect 16246 8740 16252 8804
rect 16316 8802 16363 8804
rect 18965 8804 19031 8805
rect 18965 8802 19012 8804
rect 16316 8800 16408 8802
rect 16358 8744 16408 8800
rect 16316 8742 16408 8744
rect 18920 8800 19012 8802
rect 18920 8744 18970 8800
rect 18920 8742 19012 8744
rect 16316 8740 16363 8742
rect 16297 8739 16363 8740
rect 18965 8740 19012 8742
rect 19076 8740 19082 8804
rect 19333 8802 19399 8805
rect 22320 8802 22800 8832
rect 19333 8800 22800 8802
rect 19333 8744 19338 8800
rect 19394 8744 22800 8800
rect 19333 8742 22800 8744
rect 18965 8739 19031 8740
rect 19333 8739 19399 8742
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 22320 8712 22800 8742
rect 18104 8671 18424 8672
rect 12022 8606 14842 8666
rect 15009 8666 15075 8669
rect 16798 8666 16804 8668
rect 15009 8664 16804 8666
rect 15009 8608 15014 8664
rect 15070 8608 16804 8664
rect 15009 8606 16804 8608
rect 6361 8603 6427 8606
rect 9857 8603 9923 8606
rect 15009 8603 15075 8606
rect 16798 8604 16804 8606
rect 16868 8604 16874 8668
rect 5349 8532 5415 8533
rect 5349 8530 5396 8532
rect 5304 8528 5396 8530
rect 5304 8472 5354 8528
rect 5304 8470 5396 8472
rect 5349 8468 5396 8470
rect 5460 8468 5466 8532
rect 5993 8530 6059 8533
rect 6545 8530 6611 8533
rect 5993 8528 6611 8530
rect 5993 8472 5998 8528
rect 6054 8472 6550 8528
rect 6606 8472 6611 8528
rect 5993 8470 6611 8472
rect 5349 8467 5415 8468
rect 5993 8467 6059 8470
rect 6545 8467 6611 8470
rect 9857 8530 9923 8533
rect 15694 8530 15700 8532
rect 9857 8528 15700 8530
rect 9857 8472 9862 8528
rect 9918 8472 15700 8528
rect 9857 8470 15700 8472
rect 9857 8467 9923 8470
rect 15694 8468 15700 8470
rect 15764 8468 15770 8532
rect 18229 8530 18295 8533
rect 19425 8530 19491 8533
rect 18229 8528 19491 8530
rect 18229 8472 18234 8528
rect 18290 8472 19430 8528
rect 19486 8472 19491 8528
rect 18229 8470 19491 8472
rect 18229 8467 18295 8470
rect 19425 8467 19491 8470
rect 9857 8394 9923 8397
rect 10685 8394 10751 8397
rect 12014 8394 12020 8396
rect 9857 8392 12020 8394
rect 9857 8336 9862 8392
rect 9918 8336 10690 8392
rect 10746 8336 12020 8392
rect 9857 8334 12020 8336
rect 9857 8331 9923 8334
rect 10685 8331 10751 8334
rect 12014 8332 12020 8334
rect 12084 8332 12090 8396
rect 15009 8394 15075 8397
rect 15009 8392 19212 8394
rect 15009 8336 15014 8392
rect 15070 8336 19212 8392
rect 15009 8334 19212 8336
rect 15009 8331 15075 8334
rect 0 8258 480 8288
rect 4061 8258 4127 8261
rect 9857 8258 9923 8261
rect 0 8256 4127 8258
rect 0 8200 4066 8256
rect 4122 8200 4127 8256
rect 0 8198 4127 8200
rect 0 8168 480 8198
rect 4061 8195 4127 8198
rect 9078 8256 9923 8258
rect 9078 8200 9862 8256
rect 9918 8200 9923 8256
rect 9078 8198 9923 8200
rect 7808 8192 8128 8193
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 8661 8122 8727 8125
rect 9078 8122 9138 8198
rect 9857 8195 9923 8198
rect 10726 8196 10732 8260
rect 10796 8258 10802 8260
rect 13077 8258 13143 8261
rect 10796 8256 13143 8258
rect 10796 8200 13082 8256
rect 13138 8200 13143 8256
rect 10796 8198 13143 8200
rect 10796 8196 10802 8198
rect 13077 8195 13143 8198
rect 15377 8258 15443 8261
rect 18781 8258 18847 8261
rect 15377 8256 18847 8258
rect 15377 8200 15382 8256
rect 15438 8200 18786 8256
rect 18842 8200 18847 8256
rect 15377 8198 18847 8200
rect 19152 8258 19212 8334
rect 22320 8258 22800 8288
rect 19152 8198 22800 8258
rect 15377 8195 15443 8198
rect 18781 8195 18847 8198
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 22320 8168 22800 8198
rect 14672 8127 14992 8128
rect 8661 8120 9138 8122
rect 8661 8064 8666 8120
rect 8722 8064 9138 8120
rect 8661 8062 9138 8064
rect 9857 8122 9923 8125
rect 14457 8122 14523 8125
rect 9857 8120 14523 8122
rect 9857 8064 9862 8120
rect 9918 8064 14462 8120
rect 14518 8064 14523 8120
rect 9857 8062 14523 8064
rect 8661 8059 8727 8062
rect 9857 8059 9923 8062
rect 14457 8059 14523 8062
rect 10593 7986 10659 7989
rect 13629 7986 13695 7989
rect 18413 7986 18479 7989
rect 19006 7986 19012 7988
rect 10593 7984 19012 7986
rect 10593 7928 10598 7984
rect 10654 7928 13634 7984
rect 13690 7928 18418 7984
rect 18474 7928 19012 7984
rect 10593 7926 19012 7928
rect 10593 7923 10659 7926
rect 13629 7923 13695 7926
rect 18413 7923 18479 7926
rect 19006 7924 19012 7926
rect 19076 7924 19082 7988
rect 0 7850 480 7880
rect 3969 7850 4035 7853
rect 0 7848 4035 7850
rect 0 7792 3974 7848
rect 4030 7792 4035 7848
rect 0 7790 4035 7792
rect 0 7760 480 7790
rect 3969 7787 4035 7790
rect 10961 7850 11027 7853
rect 16297 7850 16363 7853
rect 10961 7848 16363 7850
rect 10961 7792 10966 7848
rect 11022 7792 16302 7848
rect 16358 7792 16363 7848
rect 10961 7790 16363 7792
rect 10961 7787 11027 7790
rect 16297 7787 16363 7790
rect 20713 7850 20779 7853
rect 22320 7850 22800 7880
rect 20713 7848 22800 7850
rect 20713 7792 20718 7848
rect 20774 7792 22800 7848
rect 20713 7790 22800 7792
rect 20713 7787 20779 7790
rect 22320 7760 22800 7790
rect 13353 7714 13419 7717
rect 13486 7714 13492 7716
rect 13353 7712 13492 7714
rect 13353 7656 13358 7712
rect 13414 7656 13492 7712
rect 13353 7654 13492 7656
rect 13353 7651 13419 7654
rect 13486 7652 13492 7654
rect 13556 7652 13562 7716
rect 14457 7714 14523 7717
rect 16021 7714 16087 7717
rect 14457 7712 16087 7714
rect 14457 7656 14462 7712
rect 14518 7656 16026 7712
rect 16082 7656 16087 7712
rect 14457 7654 16087 7656
rect 14457 7651 14523 7654
rect 16021 7651 16087 7654
rect 4376 7648 4696 7649
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 13353 7578 13419 7581
rect 14457 7578 14523 7581
rect 18689 7580 18755 7581
rect 13353 7576 14523 7578
rect 13353 7520 13358 7576
rect 13414 7520 14462 7576
rect 14518 7520 14523 7576
rect 13353 7518 14523 7520
rect 13353 7515 13419 7518
rect 14457 7515 14523 7518
rect 18638 7516 18644 7580
rect 18708 7578 18755 7580
rect 18708 7576 18800 7578
rect 18750 7520 18800 7576
rect 18708 7518 18800 7520
rect 18708 7516 18755 7518
rect 18689 7515 18755 7516
rect 2681 7442 2747 7445
rect 8385 7442 8451 7445
rect 2681 7440 15578 7442
rect 2681 7384 2686 7440
rect 2742 7384 8390 7440
rect 8446 7384 15578 7440
rect 2681 7382 15578 7384
rect 2681 7379 2747 7382
rect 8385 7379 8451 7382
rect 0 7306 480 7336
rect 4061 7306 4127 7309
rect 0 7304 4127 7306
rect 0 7248 4066 7304
rect 4122 7248 4127 7304
rect 0 7246 4127 7248
rect 0 7216 480 7246
rect 4061 7243 4127 7246
rect 4613 7306 4679 7309
rect 5073 7306 5139 7309
rect 15518 7306 15578 7382
rect 22320 7306 22800 7336
rect 4613 7304 15394 7306
rect 4613 7248 4618 7304
rect 4674 7248 5078 7304
rect 5134 7248 15394 7304
rect 4613 7246 15394 7248
rect 15518 7246 22800 7306
rect 4613 7243 4679 7246
rect 5073 7243 5139 7246
rect 12157 7170 12223 7173
rect 12566 7170 12572 7172
rect 12157 7168 12572 7170
rect 12157 7112 12162 7168
rect 12218 7112 12572 7168
rect 12157 7110 12572 7112
rect 12157 7107 12223 7110
rect 12566 7108 12572 7110
rect 12636 7108 12642 7172
rect 15334 7170 15394 7246
rect 22320 7216 22800 7246
rect 16757 7170 16823 7173
rect 15334 7168 16823 7170
rect 15334 7112 16762 7168
rect 16818 7112 16823 7168
rect 15334 7110 16823 7112
rect 16757 7107 16823 7110
rect 18822 7108 18828 7172
rect 18892 7170 18898 7172
rect 18965 7170 19031 7173
rect 18892 7168 19031 7170
rect 18892 7112 18970 7168
rect 19026 7112 19031 7168
rect 18892 7110 19031 7112
rect 18892 7108 18898 7110
rect 18965 7107 19031 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 7039 14992 7040
rect 4889 7034 4955 7037
rect 6085 7034 6151 7037
rect 4889 7032 6151 7034
rect 4889 6976 4894 7032
rect 4950 6976 6090 7032
rect 6146 6976 6151 7032
rect 4889 6974 6151 6976
rect 4889 6971 4955 6974
rect 6085 6971 6151 6974
rect 0 6898 480 6928
rect 9213 6898 9279 6901
rect 0 6896 9279 6898
rect 0 6840 9218 6896
rect 9274 6840 9279 6896
rect 0 6838 9279 6840
rect 0 6808 480 6838
rect 9213 6835 9279 6838
rect 9581 6898 9647 6901
rect 12985 6898 13051 6901
rect 9581 6896 13051 6898
rect 9581 6840 9586 6896
rect 9642 6840 12990 6896
rect 13046 6840 13051 6896
rect 9581 6838 13051 6840
rect 9581 6835 9647 6838
rect 12985 6835 13051 6838
rect 13169 6898 13235 6901
rect 15837 6898 15903 6901
rect 13169 6896 15903 6898
rect 13169 6840 13174 6896
rect 13230 6840 15842 6896
rect 15898 6840 15903 6896
rect 13169 6838 15903 6840
rect 13169 6835 13235 6838
rect 15837 6835 15903 6838
rect 18873 6898 18939 6901
rect 22320 6898 22800 6928
rect 18873 6896 22800 6898
rect 18873 6840 18878 6896
rect 18934 6840 22800 6896
rect 18873 6838 22800 6840
rect 18873 6835 18939 6838
rect 22320 6808 22800 6838
rect 6085 6762 6151 6765
rect 8753 6762 8819 6765
rect 10317 6764 10383 6765
rect 10317 6762 10364 6764
rect 6085 6760 8819 6762
rect 6085 6704 6090 6760
rect 6146 6704 8758 6760
rect 8814 6704 8819 6760
rect 6085 6702 8819 6704
rect 10272 6760 10364 6762
rect 10272 6704 10322 6760
rect 10272 6702 10364 6704
rect 6085 6699 6151 6702
rect 8753 6699 8819 6702
rect 10317 6700 10364 6702
rect 10428 6700 10434 6764
rect 10685 6762 10751 6765
rect 10685 6760 11714 6762
rect 10685 6704 10690 6760
rect 10746 6704 11714 6760
rect 10685 6702 11714 6704
rect 10317 6699 10383 6700
rect 10685 6699 10751 6702
rect 9857 6626 9923 6629
rect 10961 6626 11027 6629
rect 9857 6624 11027 6626
rect 9857 6568 9862 6624
rect 9918 6568 10966 6624
rect 11022 6568 11027 6624
rect 9857 6566 11027 6568
rect 11654 6626 11714 6702
rect 12014 6700 12020 6764
rect 12084 6762 12090 6764
rect 18321 6762 18387 6765
rect 12084 6760 18387 6762
rect 12084 6704 18326 6760
rect 18382 6704 18387 6760
rect 12084 6702 18387 6704
rect 12084 6700 12090 6702
rect 18321 6699 18387 6702
rect 17585 6626 17651 6629
rect 11654 6624 17651 6626
rect 11654 6568 17590 6624
rect 17646 6568 17651 6624
rect 11654 6566 17651 6568
rect 9857 6563 9923 6566
rect 10961 6563 11027 6566
rect 17585 6563 17651 6566
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 11789 6490 11855 6493
rect 13537 6490 13603 6493
rect 11789 6488 13603 6490
rect 11789 6432 11794 6488
rect 11850 6432 13542 6488
rect 13598 6432 13603 6488
rect 11789 6430 13603 6432
rect 11789 6427 11855 6430
rect 13537 6427 13603 6430
rect 14917 6490 14983 6493
rect 16665 6490 16731 6493
rect 14917 6488 16731 6490
rect 14917 6432 14922 6488
rect 14978 6432 16670 6488
rect 16726 6432 16731 6488
rect 14917 6430 16731 6432
rect 14917 6427 14983 6430
rect 16665 6427 16731 6430
rect 0 6354 480 6384
rect 6545 6354 6611 6357
rect 0 6352 6611 6354
rect 0 6296 6550 6352
rect 6606 6296 6611 6352
rect 0 6294 6611 6296
rect 0 6264 480 6294
rect 6545 6291 6611 6294
rect 11513 6354 11579 6357
rect 22320 6354 22800 6384
rect 11513 6352 22800 6354
rect 11513 6296 11518 6352
rect 11574 6296 22800 6352
rect 11513 6294 22800 6296
rect 11513 6291 11579 6294
rect 22320 6264 22800 6294
rect 12341 6218 12407 6221
rect 13169 6218 13235 6221
rect 15101 6218 15167 6221
rect 12341 6216 15167 6218
rect 12341 6160 12346 6216
rect 12402 6160 13174 6216
rect 13230 6160 15106 6216
rect 15162 6160 15167 6216
rect 12341 6158 15167 6160
rect 12341 6155 12407 6158
rect 13169 6155 13235 6158
rect 15101 6155 15167 6158
rect 10041 6082 10107 6085
rect 10961 6082 11027 6085
rect 10041 6080 11027 6082
rect 10041 6024 10046 6080
rect 10102 6024 10966 6080
rect 11022 6024 11027 6080
rect 10041 6022 11027 6024
rect 10041 6019 10107 6022
rect 10961 6019 11027 6022
rect 11145 6082 11211 6085
rect 12341 6082 12407 6085
rect 11145 6080 12407 6082
rect 11145 6024 11150 6080
rect 11206 6024 12346 6080
rect 12402 6024 12407 6080
rect 11145 6022 12407 6024
rect 11145 6019 11211 6022
rect 12341 6019 12407 6022
rect 15101 6082 15167 6085
rect 17585 6082 17651 6085
rect 15101 6080 17651 6082
rect 15101 6024 15106 6080
rect 15162 6024 17590 6080
rect 17646 6024 17651 6080
rect 15101 6022 17651 6024
rect 15101 6019 15167 6022
rect 17585 6019 17651 6022
rect 7808 6016 8128 6017
rect 0 5946 480 5976
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 4061 5946 4127 5949
rect 0 5944 4127 5946
rect 0 5888 4066 5944
rect 4122 5888 4127 5944
rect 0 5886 4127 5888
rect 0 5856 480 5886
rect 4061 5883 4127 5886
rect 10358 5884 10364 5948
rect 10428 5946 10434 5948
rect 13905 5946 13971 5949
rect 10428 5944 13971 5946
rect 10428 5888 13910 5944
rect 13966 5888 13971 5944
rect 10428 5886 13971 5888
rect 10428 5884 10434 5886
rect 13905 5883 13971 5886
rect 15101 5946 15167 5949
rect 22320 5946 22800 5976
rect 15101 5944 22800 5946
rect 15101 5888 15106 5944
rect 15162 5888 22800 5944
rect 15101 5886 22800 5888
rect 15101 5883 15167 5886
rect 22320 5856 22800 5886
rect 7189 5810 7255 5813
rect 8886 5810 8892 5812
rect 7189 5808 8892 5810
rect 7189 5752 7194 5808
rect 7250 5752 8892 5808
rect 7189 5750 8892 5752
rect 7189 5747 7255 5750
rect 8886 5748 8892 5750
rect 8956 5810 8962 5812
rect 11145 5810 11211 5813
rect 8956 5808 11211 5810
rect 8956 5752 11150 5808
rect 11206 5752 11211 5808
rect 8956 5750 11211 5752
rect 8956 5748 8962 5750
rect 11145 5747 11211 5750
rect 14457 5810 14523 5813
rect 17718 5810 17724 5812
rect 14457 5808 17724 5810
rect 14457 5752 14462 5808
rect 14518 5752 17724 5808
rect 14457 5750 17724 5752
rect 14457 5747 14523 5750
rect 17718 5748 17724 5750
rect 17788 5748 17794 5812
rect 18873 5810 18939 5813
rect 19006 5810 19012 5812
rect 18873 5808 19012 5810
rect 18873 5752 18878 5808
rect 18934 5752 19012 5808
rect 18873 5750 19012 5752
rect 18873 5747 18939 5750
rect 19006 5748 19012 5750
rect 19076 5748 19082 5812
rect 11053 5674 11119 5677
rect 11789 5674 11855 5677
rect 12382 5674 12388 5676
rect 11053 5672 11714 5674
rect 11053 5616 11058 5672
rect 11114 5616 11714 5672
rect 11053 5614 11714 5616
rect 11053 5611 11119 5614
rect 11654 5538 11714 5614
rect 11789 5672 12388 5674
rect 11789 5616 11794 5672
rect 11850 5616 12388 5672
rect 11789 5614 12388 5616
rect 11789 5611 11855 5614
rect 12382 5612 12388 5614
rect 12452 5612 12458 5676
rect 12525 5674 12591 5677
rect 14460 5674 14520 5747
rect 12525 5672 14520 5674
rect 12525 5616 12530 5672
rect 12586 5616 14520 5672
rect 12525 5614 14520 5616
rect 12525 5611 12591 5614
rect 16941 5538 17007 5541
rect 11654 5536 17007 5538
rect 11654 5480 16946 5536
rect 17002 5480 17007 5536
rect 11654 5478 17007 5480
rect 16941 5475 17007 5478
rect 4376 5472 4696 5473
rect 0 5402 480 5432
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 11697 5402 11763 5405
rect 17585 5402 17651 5405
rect 0 5342 4308 5402
rect 0 5312 480 5342
rect 4248 5266 4308 5342
rect 11697 5400 17651 5402
rect 11697 5344 11702 5400
rect 11758 5344 17590 5400
rect 17646 5344 17651 5400
rect 11697 5342 17651 5344
rect 11697 5339 11763 5342
rect 17585 5339 17651 5342
rect 18781 5402 18847 5405
rect 22320 5402 22800 5432
rect 18781 5400 22800 5402
rect 18781 5344 18786 5400
rect 18842 5344 22800 5400
rect 18781 5342 22800 5344
rect 18781 5339 18847 5342
rect 22320 5312 22800 5342
rect 12525 5266 12591 5269
rect 4248 5264 12591 5266
rect 4248 5208 12530 5264
rect 12586 5208 12591 5264
rect 4248 5206 12591 5208
rect 12525 5203 12591 5206
rect 13302 5204 13308 5268
rect 13372 5266 13378 5268
rect 15285 5266 15351 5269
rect 13372 5264 15351 5266
rect 13372 5208 15290 5264
rect 15346 5208 15351 5264
rect 13372 5206 15351 5208
rect 13372 5204 13378 5206
rect 13448 5133 13508 5206
rect 15285 5203 15351 5206
rect 8385 5130 8451 5133
rect 10869 5130 10935 5133
rect 11697 5130 11763 5133
rect 8385 5128 11763 5130
rect 8385 5072 8390 5128
rect 8446 5072 10874 5128
rect 10930 5072 11702 5128
rect 11758 5072 11763 5128
rect 8385 5070 11763 5072
rect 8385 5067 8451 5070
rect 10869 5067 10935 5070
rect 11697 5067 11763 5070
rect 12525 5130 12591 5133
rect 12985 5130 13051 5133
rect 12525 5128 13051 5130
rect 12525 5072 12530 5128
rect 12586 5072 12990 5128
rect 13046 5072 13051 5128
rect 12525 5070 13051 5072
rect 12525 5067 12591 5070
rect 12985 5067 13051 5070
rect 13445 5128 13511 5133
rect 16573 5130 16639 5133
rect 13445 5072 13450 5128
rect 13506 5072 13511 5128
rect 13445 5067 13511 5072
rect 14092 5128 16639 5130
rect 14092 5072 16578 5128
rect 16634 5072 16639 5128
rect 14092 5070 16639 5072
rect 0 4994 480 5024
rect 4061 4994 4127 4997
rect 0 4992 4127 4994
rect 0 4936 4066 4992
rect 4122 4936 4127 4992
rect 0 4934 4127 4936
rect 0 4904 480 4934
rect 4061 4931 4127 4934
rect 9857 4994 9923 4997
rect 14092 4994 14152 5070
rect 16573 5067 16639 5070
rect 9857 4992 14152 4994
rect 9857 4936 9862 4992
rect 9918 4936 14152 4992
rect 9857 4934 14152 4936
rect 16205 4994 16271 4997
rect 22320 4994 22800 5024
rect 16205 4992 22800 4994
rect 16205 4936 16210 4992
rect 16266 4936 22800 4992
rect 16205 4934 22800 4936
rect 9857 4931 9923 4934
rect 16205 4931 16271 4934
rect 7808 4928 8128 4929
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 22320 4904 22800 4934
rect 14672 4863 14992 4864
rect 8201 4858 8267 4861
rect 11973 4858 12039 4861
rect 8201 4856 12039 4858
rect 8201 4800 8206 4856
rect 8262 4800 11978 4856
rect 12034 4800 12039 4856
rect 8201 4798 12039 4800
rect 8201 4795 8267 4798
rect 11973 4795 12039 4798
rect 12341 4858 12407 4861
rect 13670 4858 13676 4860
rect 12341 4856 13676 4858
rect 12341 4800 12346 4856
rect 12402 4800 13676 4856
rect 12341 4798 13676 4800
rect 12341 4795 12407 4798
rect 13670 4796 13676 4798
rect 13740 4858 13746 4860
rect 14273 4858 14339 4861
rect 13740 4856 14339 4858
rect 13740 4800 14278 4856
rect 14334 4800 14339 4856
rect 13740 4798 14339 4800
rect 13740 4796 13746 4798
rect 14273 4795 14339 4798
rect 5441 4722 5507 4725
rect 13537 4722 13603 4725
rect 13854 4722 13860 4724
rect 5441 4720 13370 4722
rect 5441 4664 5446 4720
rect 5502 4664 13370 4720
rect 5441 4662 13370 4664
rect 5441 4659 5507 4662
rect 12893 4586 12959 4589
rect 3926 4584 12959 4586
rect 3926 4528 12898 4584
rect 12954 4528 12959 4584
rect 3926 4526 12959 4528
rect 13310 4586 13370 4662
rect 13537 4720 13860 4722
rect 13537 4664 13542 4720
rect 13598 4664 13860 4720
rect 13537 4662 13860 4664
rect 13537 4659 13603 4662
rect 13854 4660 13860 4662
rect 13924 4660 13930 4724
rect 13854 4586 13860 4588
rect 13310 4526 13860 4586
rect 0 4450 480 4480
rect 2773 4450 2839 4453
rect 3926 4450 3986 4526
rect 12893 4523 12959 4526
rect 13854 4524 13860 4526
rect 13924 4586 13930 4588
rect 15142 4586 15148 4588
rect 13924 4526 15148 4586
rect 13924 4524 13930 4526
rect 15142 4524 15148 4526
rect 15212 4524 15218 4588
rect 0 4448 3986 4450
rect 0 4392 2778 4448
rect 2834 4392 3986 4448
rect 0 4390 3986 4392
rect 10317 4450 10383 4453
rect 11053 4450 11119 4453
rect 10317 4448 11119 4450
rect 10317 4392 10322 4448
rect 10378 4392 11058 4448
rect 11114 4392 11119 4448
rect 10317 4390 11119 4392
rect 0 4360 480 4390
rect 2773 4387 2839 4390
rect 10317 4387 10383 4390
rect 11053 4387 11119 4390
rect 11973 4450 12039 4453
rect 13997 4450 14063 4453
rect 11973 4448 14063 4450
rect 11973 4392 11978 4448
rect 12034 4392 14002 4448
rect 14058 4392 14063 4448
rect 11973 4390 14063 4392
rect 11973 4387 12039 4390
rect 13997 4387 14063 4390
rect 20805 4450 20871 4453
rect 22320 4450 22800 4480
rect 20805 4448 22800 4450
rect 20805 4392 20810 4448
rect 20866 4392 22800 4448
rect 20805 4390 22800 4392
rect 20805 4387 20871 4390
rect 4376 4384 4696 4385
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 22320 4360 22800 4390
rect 18104 4319 18424 4320
rect 12341 4314 12407 4317
rect 12341 4312 13370 4314
rect 12341 4256 12346 4312
rect 12402 4256 13370 4312
rect 12341 4254 13370 4256
rect 12341 4251 12407 4254
rect 10501 4180 10567 4181
rect 10501 4178 10548 4180
rect 10456 4176 10548 4178
rect 10456 4120 10506 4176
rect 10456 4118 10548 4120
rect 10501 4116 10548 4118
rect 10612 4116 10618 4180
rect 12433 4178 12499 4181
rect 13169 4178 13235 4181
rect 12433 4176 13235 4178
rect 12433 4120 12438 4176
rect 12494 4120 13174 4176
rect 13230 4120 13235 4176
rect 12433 4118 13235 4120
rect 13310 4178 13370 4254
rect 13486 4252 13492 4316
rect 13556 4314 13562 4316
rect 17217 4314 17283 4317
rect 19609 4314 19675 4317
rect 13556 4312 17283 4314
rect 13556 4256 17222 4312
rect 17278 4256 17283 4312
rect 13556 4254 17283 4256
rect 13556 4252 13562 4254
rect 17217 4251 17283 4254
rect 18600 4312 19675 4314
rect 18600 4256 19614 4312
rect 19670 4256 19675 4312
rect 18600 4254 19675 4256
rect 18600 4212 18660 4254
rect 19609 4251 19675 4254
rect 17910 4178 18660 4212
rect 13310 4152 18660 4178
rect 13310 4118 17970 4152
rect 10501 4115 10567 4116
rect 12433 4115 12499 4118
rect 13169 4115 13235 4118
rect 0 4042 480 4072
rect 4061 4042 4127 4045
rect 10317 4042 10383 4045
rect 0 4040 4127 4042
rect 0 3984 4066 4040
rect 4122 3984 4127 4040
rect 0 3982 4127 3984
rect 0 3952 480 3982
rect 4061 3979 4127 3982
rect 4294 4040 10383 4042
rect 4294 3984 10322 4040
rect 10378 3984 10383 4040
rect 4294 3982 10383 3984
rect 3693 3906 3759 3909
rect 4294 3906 4354 3982
rect 10317 3979 10383 3982
rect 11145 4042 11211 4045
rect 18965 4042 19031 4045
rect 22320 4042 22800 4072
rect 11145 4040 19031 4042
rect 11145 3984 11150 4040
rect 11206 3984 18970 4040
rect 19026 3984 19031 4040
rect 11145 3982 19031 3984
rect 11145 3979 11211 3982
rect 18965 3979 19031 3982
rect 19566 3982 22800 4042
rect 3693 3904 4354 3906
rect 3693 3848 3698 3904
rect 3754 3848 4354 3904
rect 3693 3846 4354 3848
rect 10777 3906 10843 3909
rect 13997 3906 14063 3909
rect 16573 3908 16639 3909
rect 16573 3906 16620 3908
rect 10777 3904 14063 3906
rect 10777 3848 10782 3904
rect 10838 3848 14002 3904
rect 14058 3848 14063 3904
rect 10777 3846 14063 3848
rect 16528 3904 16620 3906
rect 16528 3848 16578 3904
rect 16528 3846 16620 3848
rect 3693 3843 3759 3846
rect 10777 3843 10843 3846
rect 13997 3843 14063 3846
rect 16573 3844 16620 3846
rect 16684 3844 16690 3908
rect 16573 3843 16639 3844
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 3775 14992 3776
rect 12525 3770 12591 3773
rect 14222 3770 14228 3772
rect 12525 3768 14228 3770
rect 12525 3712 12530 3768
rect 12586 3712 14228 3768
rect 12525 3710 14228 3712
rect 12525 3707 12591 3710
rect 14222 3708 14228 3710
rect 14292 3708 14298 3772
rect 17309 3770 17375 3773
rect 17902 3770 17908 3772
rect 17309 3768 17908 3770
rect 17309 3712 17314 3768
rect 17370 3712 17908 3768
rect 17309 3710 17908 3712
rect 17309 3707 17375 3710
rect 17902 3708 17908 3710
rect 17972 3708 17978 3772
rect 18873 3770 18939 3773
rect 19566 3770 19626 3982
rect 22320 3952 22800 3982
rect 18873 3768 19626 3770
rect 18873 3712 18878 3768
rect 18934 3712 19626 3768
rect 18873 3710 19626 3712
rect 18873 3707 18939 3710
rect 5901 3634 5967 3637
rect 9673 3634 9739 3637
rect 5901 3632 9739 3634
rect 5901 3576 5906 3632
rect 5962 3576 9678 3632
rect 9734 3576 9739 3632
rect 5901 3574 9739 3576
rect 5901 3571 5967 3574
rect 9673 3571 9739 3574
rect 11513 3634 11579 3637
rect 14406 3634 14412 3636
rect 11513 3632 14412 3634
rect 11513 3576 11518 3632
rect 11574 3576 14412 3632
rect 11513 3574 14412 3576
rect 11513 3571 11579 3574
rect 14406 3572 14412 3574
rect 14476 3572 14482 3636
rect 18781 3634 18847 3637
rect 19190 3634 19196 3636
rect 18781 3632 19196 3634
rect 18781 3576 18786 3632
rect 18842 3576 19196 3632
rect 18781 3574 19196 3576
rect 18781 3571 18847 3574
rect 19190 3572 19196 3574
rect 19260 3634 19266 3636
rect 19333 3634 19399 3637
rect 19260 3632 19399 3634
rect 19260 3576 19338 3632
rect 19394 3576 19399 3632
rect 19260 3574 19399 3576
rect 19260 3572 19266 3574
rect 19333 3571 19399 3574
rect 0 3498 480 3528
rect 3049 3498 3115 3501
rect 9213 3498 9279 3501
rect 10501 3498 10567 3501
rect 0 3496 3115 3498
rect 0 3440 3054 3496
rect 3110 3440 3115 3496
rect 0 3438 3115 3440
rect 0 3408 480 3438
rect 3049 3435 3115 3438
rect 4110 3496 10567 3498
rect 4110 3440 9218 3496
rect 9274 3440 10506 3496
rect 10562 3440 10567 3496
rect 4110 3438 10567 3440
rect 565 3362 631 3365
rect 4110 3362 4170 3438
rect 9213 3435 9279 3438
rect 10501 3435 10567 3438
rect 11102 3438 11714 3498
rect 565 3360 4170 3362
rect 565 3304 570 3360
rect 626 3304 4170 3360
rect 565 3302 4170 3304
rect 6729 3362 6795 3365
rect 7097 3362 7163 3365
rect 11102 3362 11162 3438
rect 6729 3360 11162 3362
rect 6729 3304 6734 3360
rect 6790 3304 7102 3360
rect 7158 3304 11162 3360
rect 6729 3302 11162 3304
rect 11654 3362 11714 3438
rect 12750 3436 12756 3500
rect 12820 3498 12826 3500
rect 12893 3498 12959 3501
rect 12820 3496 12959 3498
rect 12820 3440 12898 3496
rect 12954 3440 12959 3496
rect 12820 3438 12959 3440
rect 12820 3436 12826 3438
rect 12893 3435 12959 3438
rect 18045 3498 18111 3501
rect 19241 3498 19307 3501
rect 18045 3496 19307 3498
rect 18045 3440 18050 3496
rect 18106 3440 19246 3496
rect 19302 3440 19307 3496
rect 18045 3438 19307 3440
rect 18045 3435 18111 3438
rect 19241 3435 19307 3438
rect 20805 3498 20871 3501
rect 22320 3498 22800 3528
rect 20805 3496 22800 3498
rect 20805 3440 20810 3496
rect 20866 3440 22800 3496
rect 20805 3438 22800 3440
rect 20805 3435 20871 3438
rect 22320 3408 22800 3438
rect 13169 3362 13235 3365
rect 11654 3302 12634 3362
rect 565 3299 631 3302
rect 6729 3299 6795 3302
rect 7097 3299 7163 3302
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 12574 3226 12634 3302
rect 13169 3360 13508 3362
rect 13169 3304 13174 3360
rect 13230 3304 13508 3360
rect 13169 3302 13508 3304
rect 13169 3299 13235 3302
rect 13448 3226 13508 3302
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 13721 3226 13787 3229
rect 12574 3166 13370 3226
rect 13448 3224 13787 3226
rect 13448 3168 13726 3224
rect 13782 3168 13787 3224
rect 13448 3166 13787 3168
rect 0 3090 480 3120
rect 2313 3090 2379 3093
rect 0 3088 2379 3090
rect 0 3032 2318 3088
rect 2374 3032 2379 3088
rect 0 3030 2379 3032
rect 0 3000 480 3030
rect 2313 3027 2379 3030
rect 4061 3090 4127 3093
rect 9949 3090 10015 3093
rect 13169 3090 13235 3093
rect 4061 3088 13235 3090
rect 4061 3032 4066 3088
rect 4122 3032 9954 3088
rect 10010 3032 13174 3088
rect 13230 3032 13235 3088
rect 4061 3030 13235 3032
rect 13310 3090 13370 3166
rect 13721 3163 13787 3166
rect 13905 3226 13971 3229
rect 14641 3226 14707 3229
rect 17769 3226 17835 3229
rect 13905 3224 14707 3226
rect 13905 3168 13910 3224
rect 13966 3168 14646 3224
rect 14702 3168 14707 3224
rect 13905 3166 14707 3168
rect 13905 3163 13971 3166
rect 14641 3163 14707 3166
rect 14782 3224 17835 3226
rect 14782 3168 17774 3224
rect 17830 3168 17835 3224
rect 14782 3166 17835 3168
rect 14782 3090 14842 3166
rect 17769 3163 17835 3166
rect 18965 3226 19031 3229
rect 19609 3226 19675 3229
rect 18965 3224 19675 3226
rect 18965 3168 18970 3224
rect 19026 3168 19614 3224
rect 19670 3168 19675 3224
rect 18965 3166 19675 3168
rect 18965 3163 19031 3166
rect 19609 3163 19675 3166
rect 19742 3164 19748 3228
rect 19812 3226 19818 3228
rect 19885 3226 19951 3229
rect 19812 3224 19951 3226
rect 19812 3168 19890 3224
rect 19946 3168 19951 3224
rect 19812 3166 19951 3168
rect 19812 3164 19818 3166
rect 19885 3163 19951 3166
rect 13310 3030 14842 3090
rect 4061 3027 4127 3030
rect 9949 3027 10015 3030
rect 13169 3027 13235 3030
rect 16798 3028 16804 3092
rect 16868 3090 16874 3092
rect 17769 3090 17835 3093
rect 16868 3088 17835 3090
rect 16868 3032 17774 3088
rect 17830 3032 17835 3088
rect 16868 3030 17835 3032
rect 16868 3028 16874 3030
rect 17769 3027 17835 3030
rect 18321 3090 18387 3093
rect 18597 3090 18663 3093
rect 18321 3088 18663 3090
rect 18321 3032 18326 3088
rect 18382 3032 18602 3088
rect 18658 3032 18663 3088
rect 18321 3030 18663 3032
rect 18321 3027 18387 3030
rect 18597 3027 18663 3030
rect 19793 3090 19859 3093
rect 19926 3090 19932 3092
rect 19793 3088 19932 3090
rect 19793 3032 19798 3088
rect 19854 3032 19932 3088
rect 19793 3030 19932 3032
rect 19793 3027 19859 3030
rect 19926 3028 19932 3030
rect 19996 3028 20002 3092
rect 22320 3090 22800 3120
rect 20118 3030 22800 3090
rect 9029 2954 9095 2957
rect 12341 2954 12407 2957
rect 9029 2952 12407 2954
rect 9029 2896 9034 2952
rect 9090 2896 12346 2952
rect 12402 2896 12407 2952
rect 9029 2894 12407 2896
rect 9029 2891 9095 2894
rect 12341 2891 12407 2894
rect 12934 2892 12940 2956
rect 13004 2954 13010 2956
rect 13169 2954 13235 2957
rect 13004 2952 13235 2954
rect 13004 2896 13174 2952
rect 13230 2896 13235 2952
rect 13004 2894 13235 2896
rect 13004 2892 13010 2894
rect 13169 2891 13235 2894
rect 13537 2954 13603 2957
rect 14549 2954 14615 2957
rect 13537 2952 14615 2954
rect 13537 2896 13542 2952
rect 13598 2896 14554 2952
rect 14610 2896 14615 2952
rect 13537 2894 14615 2896
rect 13537 2891 13603 2894
rect 14549 2891 14615 2894
rect 17309 2954 17375 2957
rect 18638 2954 18644 2956
rect 17309 2952 18644 2954
rect 17309 2896 17314 2952
rect 17370 2896 18644 2952
rect 17309 2894 18644 2896
rect 17309 2891 17375 2894
rect 18638 2892 18644 2894
rect 18708 2954 18714 2956
rect 20118 2954 20178 3030
rect 22320 3000 22800 3030
rect 18708 2894 20178 2954
rect 18708 2892 18714 2894
rect 10225 2818 10291 2821
rect 10726 2818 10732 2820
rect 10225 2816 10732 2818
rect 10225 2760 10230 2816
rect 10286 2760 10732 2816
rect 10225 2758 10732 2760
rect 10225 2755 10291 2758
rect 10726 2756 10732 2758
rect 10796 2756 10802 2820
rect 12014 2756 12020 2820
rect 12084 2818 12090 2820
rect 13813 2818 13879 2821
rect 18873 2820 18939 2821
rect 12084 2816 13879 2818
rect 12084 2760 13818 2816
rect 13874 2760 13879 2816
rect 12084 2758 13879 2760
rect 12084 2756 12090 2758
rect 13813 2755 13879 2758
rect 18822 2756 18828 2820
rect 18892 2818 18939 2820
rect 18892 2816 18984 2818
rect 18934 2760 18984 2816
rect 18892 2758 18984 2760
rect 18892 2756 18939 2758
rect 18873 2755 18939 2756
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 10409 2684 10475 2685
rect 13905 2684 13971 2685
rect 10358 2682 10364 2684
rect 10318 2622 10364 2682
rect 10428 2680 10475 2684
rect 10470 2624 10475 2680
rect 10358 2620 10364 2622
rect 10428 2620 10475 2624
rect 13854 2620 13860 2684
rect 13924 2682 13971 2684
rect 15929 2682 15995 2685
rect 16062 2682 16068 2684
rect 13924 2680 14016 2682
rect 13966 2624 14016 2680
rect 13924 2622 14016 2624
rect 15929 2680 16068 2682
rect 15929 2624 15934 2680
rect 15990 2624 16068 2680
rect 15929 2622 16068 2624
rect 13924 2620 13971 2622
rect 10409 2619 10475 2620
rect 13905 2619 13971 2620
rect 15929 2619 15995 2622
rect 16062 2620 16068 2622
rect 16132 2620 16138 2684
rect 16430 2620 16436 2684
rect 16500 2682 16506 2684
rect 16941 2682 17007 2685
rect 20437 2684 20503 2685
rect 20437 2682 20484 2684
rect 16500 2680 17007 2682
rect 16500 2624 16946 2680
rect 17002 2624 17007 2680
rect 16500 2622 17007 2624
rect 20392 2680 20484 2682
rect 20392 2624 20442 2680
rect 20392 2622 20484 2624
rect 16500 2620 16506 2622
rect 16941 2619 17007 2622
rect 20437 2620 20484 2622
rect 20548 2620 20554 2684
rect 20437 2619 20503 2620
rect 0 2546 480 2576
rect 1853 2546 1919 2549
rect 0 2544 1919 2546
rect 0 2488 1858 2544
rect 1914 2488 1919 2544
rect 0 2486 1919 2488
rect 0 2456 480 2486
rect 1853 2483 1919 2486
rect 10133 2546 10199 2549
rect 10542 2546 10548 2548
rect 10133 2544 10548 2546
rect 10133 2488 10138 2544
rect 10194 2488 10548 2544
rect 10133 2486 10548 2488
rect 10133 2483 10199 2486
rect 10542 2484 10548 2486
rect 10612 2484 10618 2548
rect 12382 2484 12388 2548
rect 12452 2546 12458 2548
rect 13905 2546 13971 2549
rect 12452 2544 13971 2546
rect 12452 2488 13910 2544
rect 13966 2488 13971 2544
rect 12452 2486 13971 2488
rect 12452 2484 12458 2486
rect 13905 2483 13971 2486
rect 14038 2484 14044 2548
rect 14108 2546 14114 2548
rect 17217 2546 17283 2549
rect 14108 2544 17283 2546
rect 14108 2488 17222 2544
rect 17278 2488 17283 2544
rect 14108 2486 17283 2488
rect 14108 2484 14114 2486
rect 17217 2483 17283 2486
rect 19057 2546 19123 2549
rect 20294 2546 20300 2548
rect 19057 2544 20300 2546
rect 19057 2488 19062 2544
rect 19118 2488 20300 2544
rect 19057 2486 20300 2488
rect 19057 2483 19123 2486
rect 20294 2484 20300 2486
rect 20364 2484 20370 2548
rect 22320 2546 22800 2576
rect 20486 2486 22800 2546
rect 9673 2410 9739 2413
rect 15377 2410 15443 2413
rect 9673 2408 15443 2410
rect 9673 2352 9678 2408
rect 9734 2352 15382 2408
rect 15438 2352 15443 2408
rect 9673 2350 15443 2352
rect 9673 2347 9739 2350
rect 15377 2347 15443 2350
rect 18781 2410 18847 2413
rect 20486 2410 20546 2486
rect 22320 2456 22800 2486
rect 18781 2408 20546 2410
rect 18781 2352 18786 2408
rect 18842 2352 20546 2408
rect 18781 2350 20546 2352
rect 18781 2347 18847 2350
rect 4376 2208 4696 2209
rect 0 2138 480 2168
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 3233 2138 3299 2141
rect 22320 2138 22800 2168
rect 0 2136 3299 2138
rect 0 2080 3238 2136
rect 3294 2080 3299 2136
rect 0 2078 3299 2080
rect 0 2048 480 2078
rect 3233 2075 3299 2078
rect 18646 2078 22800 2138
rect 8477 2002 8543 2005
rect 14365 2002 14431 2005
rect 8477 2000 14431 2002
rect 8477 1944 8482 2000
rect 8538 1944 14370 2000
rect 14426 1944 14431 2000
rect 8477 1942 14431 1944
rect 8477 1939 8543 1942
rect 14365 1939 14431 1942
rect 16573 2002 16639 2005
rect 18646 2002 18706 2078
rect 22320 2048 22800 2078
rect 16573 2000 18706 2002
rect 16573 1944 16578 2000
rect 16634 1944 18706 2000
rect 16573 1942 18706 1944
rect 16573 1939 16639 1942
rect 17350 1804 17356 1868
rect 17420 1866 17426 1868
rect 18045 1866 18111 1869
rect 17420 1864 18111 1866
rect 17420 1808 18050 1864
rect 18106 1808 18111 1864
rect 17420 1806 18111 1808
rect 17420 1804 17426 1806
rect 18045 1803 18111 1806
rect 0 1594 480 1624
rect 5257 1594 5323 1597
rect 0 1592 5323 1594
rect 0 1536 5262 1592
rect 5318 1536 5323 1592
rect 0 1534 5323 1536
rect 0 1504 480 1534
rect 5257 1531 5323 1534
rect 17953 1594 18019 1597
rect 21265 1594 21331 1597
rect 22320 1594 22800 1624
rect 17953 1592 22800 1594
rect 17953 1536 17958 1592
rect 18014 1536 21270 1592
rect 21326 1536 22800 1592
rect 17953 1534 22800 1536
rect 17953 1531 18019 1534
rect 21265 1531 21331 1534
rect 22320 1504 22800 1534
rect 0 1186 480 1216
rect 4245 1186 4311 1189
rect 0 1184 4311 1186
rect 0 1128 4250 1184
rect 4306 1128 4311 1184
rect 0 1126 4311 1128
rect 0 1096 480 1126
rect 4245 1123 4311 1126
rect 17953 1186 18019 1189
rect 21357 1186 21423 1189
rect 22320 1186 22800 1216
rect 17953 1184 22800 1186
rect 17953 1128 17958 1184
rect 18014 1128 21362 1184
rect 21418 1128 22800 1184
rect 17953 1126 22800 1128
rect 17953 1123 18019 1126
rect 21357 1123 21423 1126
rect 22320 1096 22800 1126
rect 0 642 480 672
rect 3233 642 3299 645
rect 0 640 3299 642
rect 0 584 3238 640
rect 3294 584 3299 640
rect 0 582 3299 584
rect 0 552 480 582
rect 3233 579 3299 582
rect 19149 642 19215 645
rect 22320 642 22800 672
rect 19149 640 22800 642
rect 19149 584 19154 640
rect 19210 584 22800 640
rect 19149 582 22800 584
rect 19149 579 19215 582
rect 22320 552 22800 582
rect 0 234 480 264
rect 3969 234 4035 237
rect 0 232 4035 234
rect 0 176 3974 232
rect 4030 176 4035 232
rect 0 174 4035 176
rect 0 144 480 174
rect 3969 171 4035 174
rect 18873 234 18939 237
rect 22320 234 22800 264
rect 18873 232 22800 234
rect 18873 176 18878 232
rect 18934 176 22800 232
rect 18873 174 22800 176
rect 18873 171 18939 174
rect 22320 144 22800 174
<< via3 >>
rect 13860 20300 13924 20364
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 13676 19756 13740 19820
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 14228 19544 14292 19548
rect 14228 19488 14278 19544
rect 14278 19488 14292 19544
rect 14228 19484 14292 19488
rect 14412 19408 14476 19412
rect 14412 19352 14426 19408
rect 14426 19352 14476 19408
rect 14412 19348 14476 19352
rect 19932 19408 19996 19412
rect 19932 19352 19946 19408
rect 19946 19352 19996 19408
rect 19932 19348 19996 19352
rect 4108 19212 4172 19276
rect 12940 19272 13004 19276
rect 12940 19216 12990 19272
rect 12990 19216 13004 19272
rect 12940 19212 13004 19216
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4844 18668 4908 18732
rect 15148 18668 15212 18732
rect 15884 18668 15948 18732
rect 18828 18668 18892 18732
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 9260 18396 9324 18460
rect 19196 18456 19260 18460
rect 19196 18400 19246 18456
rect 19246 18400 19260 18456
rect 8524 18260 8588 18324
rect 19196 18396 19260 18400
rect 19380 18396 19444 18460
rect 15516 18260 15580 18324
rect 10180 18184 10244 18188
rect 10180 18128 10194 18184
rect 10194 18128 10244 18184
rect 10180 18124 10244 18128
rect 13492 18124 13556 18188
rect 14044 18124 14108 18188
rect 15332 18124 15396 18188
rect 17172 18124 17236 18188
rect 20484 18124 20548 18188
rect 7420 18048 7484 18052
rect 7420 17992 7470 18048
rect 7470 17992 7484 18048
rect 7420 17988 7484 17992
rect 13860 17988 13924 18052
rect 15700 18048 15764 18052
rect 15700 17992 15714 18048
rect 15714 17992 15764 18048
rect 15700 17988 15764 17992
rect 16068 18048 16132 18052
rect 16068 17992 16082 18048
rect 16082 17992 16132 18048
rect 16068 17988 16132 17992
rect 16436 17988 16500 18052
rect 16620 17988 16684 18052
rect 17908 17988 17972 18052
rect 19748 18048 19812 18052
rect 19748 17992 19762 18048
rect 19762 17992 19812 18048
rect 19748 17988 19812 17992
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 19564 17852 19628 17916
rect 12756 17716 12820 17780
rect 13124 17444 13188 17508
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 9444 17368 9508 17372
rect 9444 17312 9458 17368
rect 9458 17312 9508 17368
rect 9444 17308 9508 17312
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 11652 17172 11716 17236
rect 16988 17308 17052 17372
rect 12204 16900 12268 16964
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 15884 16628 15948 16692
rect 17724 16688 17788 16692
rect 17724 16632 17774 16688
rect 17774 16632 17788 16688
rect 17724 16628 17788 16632
rect 18644 16628 18708 16692
rect 12204 16492 12268 16556
rect 16804 16492 16868 16556
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 12572 15812 12636 15876
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 9628 15540 9692 15604
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 16252 15540 16316 15604
rect 12388 15404 12452 15468
rect 8524 15268 8588 15332
rect 20300 15328 20364 15332
rect 20300 15272 20350 15328
rect 20350 15272 20364 15328
rect 20300 15268 20364 15272
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 15332 14996 15396 15060
rect 15884 14996 15948 15060
rect 10548 14860 10612 14924
rect 11836 14860 11900 14924
rect 9996 14724 10060 14788
rect 15516 14724 15580 14788
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 12020 14588 12084 14652
rect 16988 14588 17052 14652
rect 18644 14452 18708 14516
rect 13860 14180 13924 14244
rect 15332 14180 15396 14244
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 17172 13908 17236 13972
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 13860 13636 13924 13700
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 12388 13500 12452 13564
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 16988 13832 17052 13836
rect 16988 13776 17002 13832
rect 17002 13776 17052 13832
rect 16988 13772 17052 13776
rect 19564 13636 19628 13700
rect 19380 13500 19444 13564
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 13124 13288 13188 13292
rect 13124 13232 13138 13288
rect 13138 13232 13188 13288
rect 13124 13228 13188 13232
rect 13308 13288 13372 13292
rect 13308 13232 13358 13288
rect 13358 13232 13372 13288
rect 13308 13228 13372 13232
rect 13676 13288 13740 13292
rect 13676 13232 13726 13288
rect 13726 13232 13740 13288
rect 13676 13228 13740 13232
rect 17172 13092 17236 13156
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 8524 12956 8588 13020
rect 10364 13016 10428 13020
rect 10364 12960 10378 13016
rect 10378 12960 10428 13016
rect 10364 12956 10428 12960
rect 15148 12956 15212 13020
rect 19012 12956 19076 13020
rect 19380 13016 19444 13020
rect 19380 12960 19394 13016
rect 19394 12960 19444 13016
rect 19380 12956 19444 12960
rect 12204 12880 12268 12884
rect 12204 12824 12254 12880
rect 12254 12824 12268 12880
rect 12204 12820 12268 12824
rect 13124 12880 13188 12884
rect 13124 12824 13174 12880
rect 13174 12824 13188 12880
rect 13124 12820 13188 12824
rect 9444 12684 9508 12748
rect 11652 12744 11716 12748
rect 11652 12688 11702 12744
rect 11702 12688 11716 12744
rect 11652 12684 11716 12688
rect 4844 12548 4908 12612
rect 11836 12548 11900 12612
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 9628 12412 9692 12476
rect 13676 12684 13740 12748
rect 15148 12608 15212 12612
rect 15148 12552 15162 12608
rect 15162 12552 15212 12608
rect 15148 12548 15212 12552
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 17356 12608 17420 12612
rect 17356 12552 17370 12608
rect 17370 12552 17420 12608
rect 17356 12548 17420 12552
rect 17540 12608 17604 12612
rect 17540 12552 17590 12608
rect 17590 12552 17604 12608
rect 17540 12548 17604 12552
rect 11652 12276 11716 12340
rect 16620 12276 16684 12340
rect 19196 12276 19260 12340
rect 9260 12004 9324 12068
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 6132 11868 6196 11932
rect 10916 11868 10980 11932
rect 11836 12200 11900 12204
rect 11836 12144 11886 12200
rect 11886 12144 11900 12200
rect 11836 12140 11900 12144
rect 13492 12064 13556 12068
rect 13492 12008 13506 12064
rect 13506 12008 13556 12064
rect 13492 12004 13556 12008
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 12020 11596 12084 11660
rect 13124 11596 13188 11660
rect 17540 11792 17604 11796
rect 17540 11736 17590 11792
rect 17590 11736 17604 11792
rect 17540 11732 17604 11736
rect 4108 11460 4172 11524
rect 11652 11460 11716 11524
rect 12940 11460 13004 11524
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 5396 11324 5460 11388
rect 10364 11324 10428 11388
rect 15884 11324 15948 11388
rect 10916 11052 10980 11116
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 5396 10780 5460 10844
rect 15516 11052 15580 11116
rect 18828 11052 18892 11116
rect 13308 10916 13372 10980
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 8892 10704 8956 10708
rect 8892 10648 8906 10704
rect 8906 10648 8956 10704
rect 8892 10644 8956 10648
rect 11836 10644 11900 10708
rect 16988 10644 17052 10708
rect 9996 10508 10060 10572
rect 13308 10508 13372 10572
rect 12940 10372 13004 10436
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 10180 10236 10244 10300
rect 7420 10100 7484 10164
rect 6132 10024 6196 10028
rect 6132 9968 6146 10024
rect 6146 9968 6196 10024
rect 6132 9964 6196 9968
rect 17356 10024 17420 10028
rect 17356 9968 17370 10024
rect 17370 9968 17420 10024
rect 17356 9964 17420 9968
rect 12756 9888 12820 9892
rect 12756 9832 12806 9888
rect 12806 9832 12820 9888
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 10548 9692 10612 9756
rect 10548 9556 10612 9620
rect 12756 9828 12820 9832
rect 15332 9828 15396 9892
rect 17172 9828 17236 9892
rect 11836 9692 11900 9756
rect 12756 9692 12820 9756
rect 12940 9692 13004 9756
rect 19380 10024 19444 10028
rect 19380 9968 19394 10024
rect 19394 9968 19444 10024
rect 19380 9964 19444 9968
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 12756 9556 12820 9620
rect 19196 9420 19260 9484
rect 12020 9284 12084 9348
rect 15148 9284 15212 9348
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 17356 9148 17420 9212
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 13860 8876 13924 8940
rect 13124 8740 13188 8804
rect 16252 8800 16316 8804
rect 16252 8744 16302 8800
rect 16302 8744 16316 8800
rect 16252 8740 16316 8744
rect 19012 8800 19076 8804
rect 19012 8744 19026 8800
rect 19026 8744 19076 8800
rect 19012 8740 19076 8744
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 16804 8604 16868 8668
rect 5396 8528 5460 8532
rect 5396 8472 5410 8528
rect 5410 8472 5460 8528
rect 5396 8468 5460 8472
rect 15700 8468 15764 8532
rect 12020 8332 12084 8396
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 10732 8196 10796 8260
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 19012 7924 19076 7988
rect 13492 7652 13556 7716
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 18644 7576 18708 7580
rect 18644 7520 18694 7576
rect 18694 7520 18708 7576
rect 18644 7516 18708 7520
rect 12572 7108 12636 7172
rect 18828 7108 18892 7172
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 10364 6760 10428 6764
rect 10364 6704 10378 6760
rect 10378 6704 10428 6760
rect 10364 6700 10428 6704
rect 12020 6700 12084 6764
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 10364 5884 10428 5948
rect 8892 5748 8956 5812
rect 17724 5748 17788 5812
rect 19012 5748 19076 5812
rect 12388 5612 12452 5676
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 13308 5204 13372 5268
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 13676 4796 13740 4860
rect 13860 4660 13924 4724
rect 13860 4524 13924 4588
rect 15148 4524 15212 4588
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 10548 4176 10612 4180
rect 10548 4120 10562 4176
rect 10562 4120 10612 4176
rect 10548 4116 10612 4120
rect 13492 4252 13556 4316
rect 16620 3904 16684 3908
rect 16620 3848 16634 3904
rect 16634 3848 16684 3904
rect 16620 3844 16684 3848
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 14228 3708 14292 3772
rect 17908 3708 17972 3772
rect 14412 3572 14476 3636
rect 19196 3572 19260 3636
rect 12756 3436 12820 3500
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 19748 3164 19812 3228
rect 16804 3028 16868 3092
rect 19932 3028 19996 3092
rect 12940 2892 13004 2956
rect 18644 2892 18708 2956
rect 10732 2756 10796 2820
rect 12020 2756 12084 2820
rect 18828 2816 18892 2820
rect 18828 2760 18878 2816
rect 18878 2760 18892 2816
rect 18828 2756 18892 2760
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 10364 2680 10428 2684
rect 10364 2624 10414 2680
rect 10414 2624 10428 2680
rect 10364 2620 10428 2624
rect 13860 2680 13924 2684
rect 13860 2624 13910 2680
rect 13910 2624 13924 2680
rect 13860 2620 13924 2624
rect 16068 2620 16132 2684
rect 16436 2620 16500 2684
rect 20484 2680 20548 2684
rect 20484 2624 20498 2680
rect 20498 2624 20548 2680
rect 20484 2620 20548 2624
rect 10548 2484 10612 2548
rect 12388 2484 12452 2548
rect 14044 2484 14108 2548
rect 20300 2484 20364 2548
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
rect 17356 1804 17420 1868
<< metal4 >>
rect 13859 20364 13925 20365
rect 13859 20300 13860 20364
rect 13924 20300 13925 20364
rect 13859 20299 13925 20300
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4107 19276 4173 19277
rect 4107 19212 4108 19276
rect 4172 19212 4173 19276
rect 4107 19211 4173 19212
rect 4110 11525 4170 19211
rect 4376 18528 4696 19552
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 4843 18732 4909 18733
rect 4843 18668 4844 18732
rect 4908 18668 4909 18732
rect 4843 18667 4909 18668
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4846 12613 4906 18667
rect 7419 18052 7485 18053
rect 7419 17988 7420 18052
rect 7484 17988 7485 18052
rect 7419 17987 7485 17988
rect 4843 12612 4909 12613
rect 4843 12548 4844 12612
rect 4908 12548 4909 12612
rect 4843 12547 4909 12548
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4107 11524 4173 11525
rect 4107 11460 4108 11524
rect 4172 11460 4173 11524
rect 4107 11459 4173 11460
rect 4376 10912 4696 11936
rect 6131 11932 6197 11933
rect 6131 11868 6132 11932
rect 6196 11868 6197 11932
rect 6131 11867 6197 11868
rect 5395 11388 5461 11389
rect 5395 11324 5396 11388
rect 5460 11324 5461 11388
rect 5395 11323 5461 11324
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 5398 10845 5458 11323
rect 5395 10844 5461 10845
rect 5395 10780 5396 10844
rect 5460 10780 5461 10844
rect 5395 10779 5461 10780
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 5398 8533 5458 10779
rect 6134 10029 6194 11867
rect 7422 10165 7482 17987
rect 7808 17984 8128 19008
rect 11240 19616 11560 20176
rect 13675 19820 13741 19821
rect 13675 19756 13676 19820
rect 13740 19756 13741 19820
rect 13675 19755 13741 19756
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 12939 19276 13005 19277
rect 12939 19212 12940 19276
rect 13004 19212 13005 19276
rect 12939 19211 13005 19212
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 9259 18460 9325 18461
rect 9259 18396 9260 18460
rect 9324 18396 9325 18460
rect 9259 18395 9325 18396
rect 8523 18324 8589 18325
rect 8523 18260 8524 18324
rect 8588 18260 8589 18324
rect 8523 18259 8589 18260
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 8526 15333 8586 18259
rect 8523 15332 8589 15333
rect 8523 15268 8524 15332
rect 8588 15268 8589 15332
rect 8523 15267 8589 15268
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 8526 13021 8586 15267
rect 8523 13020 8589 13021
rect 8523 12956 8524 13020
rect 8588 12956 8589 13020
rect 8523 12955 8589 12956
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 9262 12069 9322 18395
rect 10179 18188 10245 18189
rect 10179 18124 10180 18188
rect 10244 18124 10245 18188
rect 10179 18123 10245 18124
rect 9443 17372 9509 17373
rect 9443 17308 9444 17372
rect 9508 17308 9509 17372
rect 9443 17307 9509 17308
rect 9446 12749 9506 17307
rect 9627 15604 9693 15605
rect 9627 15540 9628 15604
rect 9692 15540 9693 15604
rect 9627 15539 9693 15540
rect 9443 12748 9509 12749
rect 9443 12684 9444 12748
rect 9508 12684 9509 12748
rect 9443 12683 9509 12684
rect 9630 12477 9690 15539
rect 9995 14788 10061 14789
rect 9995 14724 9996 14788
rect 10060 14724 10061 14788
rect 9995 14723 10061 14724
rect 9627 12476 9693 12477
rect 9627 12412 9628 12476
rect 9692 12412 9693 12476
rect 9627 12411 9693 12412
rect 9259 12068 9325 12069
rect 9259 12004 9260 12068
rect 9324 12004 9325 12068
rect 9259 12003 9325 12004
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 8891 10708 8957 10709
rect 8891 10644 8892 10708
rect 8956 10644 8957 10708
rect 8891 10643 8957 10644
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7419 10164 7485 10165
rect 7419 10100 7420 10164
rect 7484 10100 7485 10164
rect 7419 10099 7485 10100
rect 6131 10028 6197 10029
rect 6131 9964 6132 10028
rect 6196 9964 6197 10028
rect 6131 9963 6197 9964
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 5395 8532 5461 8533
rect 5395 8468 5396 8532
rect 5460 8468 5461 8532
rect 5395 8467 5461 8468
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 8894 5813 8954 10643
rect 9998 10573 10058 14723
rect 9995 10572 10061 10573
rect 9995 10508 9996 10572
rect 10060 10508 10061 10572
rect 9995 10507 10061 10508
rect 10182 10301 10242 18123
rect 11240 17440 11560 18464
rect 12755 17780 12821 17781
rect 12755 17716 12756 17780
rect 12820 17716 12821 17780
rect 12755 17715 12821 17716
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11651 17236 11717 17237
rect 11651 17172 11652 17236
rect 11716 17172 11717 17236
rect 11651 17171 11717 17172
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 10547 14924 10613 14925
rect 10547 14860 10548 14924
rect 10612 14860 10613 14924
rect 10547 14859 10613 14860
rect 10363 13020 10429 13021
rect 10363 12956 10364 13020
rect 10428 12956 10429 13020
rect 10363 12955 10429 12956
rect 10366 11389 10426 12955
rect 10363 11388 10429 11389
rect 10363 11324 10364 11388
rect 10428 11324 10429 11388
rect 10363 11323 10429 11324
rect 10179 10300 10245 10301
rect 10179 10236 10180 10300
rect 10244 10236 10245 10300
rect 10179 10235 10245 10236
rect 10550 9757 10610 14859
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11654 12749 11714 17171
rect 12203 16964 12269 16965
rect 12203 16900 12204 16964
rect 12268 16900 12269 16964
rect 12203 16899 12269 16900
rect 12206 16557 12266 16899
rect 12203 16556 12269 16557
rect 12203 16492 12204 16556
rect 12268 16492 12269 16556
rect 12203 16491 12269 16492
rect 11835 14924 11901 14925
rect 11835 14860 11836 14924
rect 11900 14860 11901 14924
rect 11835 14859 11901 14860
rect 11651 12748 11717 12749
rect 11651 12684 11652 12748
rect 11716 12684 11717 12748
rect 11651 12683 11717 12684
rect 11838 12613 11898 14859
rect 12019 14652 12085 14653
rect 12019 14588 12020 14652
rect 12084 14588 12085 14652
rect 12019 14587 12085 14588
rect 11835 12612 11901 12613
rect 11835 12548 11836 12612
rect 11900 12548 11901 12612
rect 11835 12547 11901 12548
rect 11651 12340 11717 12341
rect 11651 12276 11652 12340
rect 11716 12276 11717 12340
rect 11651 12275 11717 12276
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 10915 11932 10981 11933
rect 10915 11868 10916 11932
rect 10980 11868 10981 11932
rect 10915 11867 10981 11868
rect 10918 11117 10978 11867
rect 10915 11116 10981 11117
rect 10915 11052 10916 11116
rect 10980 11052 10981 11116
rect 10915 11051 10981 11052
rect 11240 10912 11560 11936
rect 11654 11525 11714 12275
rect 11838 12205 11898 12547
rect 11835 12204 11901 12205
rect 11835 12140 11836 12204
rect 11900 12140 11901 12204
rect 11835 12139 11901 12140
rect 12022 11661 12082 14587
rect 12206 12885 12266 16491
rect 12571 15876 12637 15877
rect 12571 15812 12572 15876
rect 12636 15812 12637 15876
rect 12571 15811 12637 15812
rect 12387 15468 12453 15469
rect 12387 15404 12388 15468
rect 12452 15404 12453 15468
rect 12387 15403 12453 15404
rect 12390 15330 12450 15403
rect 12574 15330 12634 15811
rect 12390 15270 12634 15330
rect 12387 13564 12453 13565
rect 12387 13500 12388 13564
rect 12452 13500 12453 13564
rect 12387 13499 12453 13500
rect 12203 12884 12269 12885
rect 12203 12820 12204 12884
rect 12268 12820 12269 12884
rect 12203 12819 12269 12820
rect 12019 11660 12085 11661
rect 12019 11596 12020 11660
rect 12084 11596 12085 11660
rect 12019 11595 12085 11596
rect 11651 11524 11717 11525
rect 11651 11460 11652 11524
rect 11716 11460 11717 11524
rect 11651 11459 11717 11460
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11835 10708 11901 10709
rect 11835 10644 11836 10708
rect 11900 10644 11901 10708
rect 11835 10643 11901 10644
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 10547 9756 10613 9757
rect 10547 9692 10548 9756
rect 10612 9692 10613 9756
rect 10547 9691 10613 9692
rect 10547 9620 10613 9621
rect 10547 9556 10548 9620
rect 10612 9556 10613 9620
rect 10547 9555 10613 9556
rect 10363 6764 10429 6765
rect 10363 6700 10364 6764
rect 10428 6700 10429 6764
rect 10363 6699 10429 6700
rect 10366 5949 10426 6699
rect 10363 5948 10429 5949
rect 10363 5884 10364 5948
rect 10428 5884 10429 5948
rect 10363 5883 10429 5884
rect 8891 5812 8957 5813
rect 8891 5748 8892 5812
rect 8956 5748 8957 5812
rect 8891 5747 8957 5748
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 10366 2685 10426 5883
rect 10550 4181 10610 9555
rect 11240 8736 11560 9760
rect 11838 9757 11898 10643
rect 11835 9756 11901 9757
rect 11835 9692 11836 9756
rect 11900 9692 11901 9756
rect 11835 9691 11901 9692
rect 12022 9349 12082 11595
rect 12019 9348 12085 9349
rect 12019 9284 12020 9348
rect 12084 9284 12085 9348
rect 12019 9283 12085 9284
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 10731 8260 10797 8261
rect 10731 8196 10732 8260
rect 10796 8196 10797 8260
rect 10731 8195 10797 8196
rect 10547 4180 10613 4181
rect 10547 4116 10548 4180
rect 10612 4116 10613 4180
rect 10547 4115 10613 4116
rect 10363 2684 10429 2685
rect 10363 2620 10364 2684
rect 10428 2620 10429 2684
rect 10363 2619 10429 2620
rect 10550 2549 10610 4115
rect 10734 2821 10794 8195
rect 11240 7648 11560 8672
rect 12019 8396 12085 8397
rect 12019 8332 12020 8396
rect 12084 8332 12085 8396
rect 12019 8331 12085 8332
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 12022 6765 12082 8331
rect 12390 7170 12450 13499
rect 12758 9893 12818 17715
rect 12942 11525 13002 19211
rect 13491 18188 13557 18189
rect 13491 18124 13492 18188
rect 13556 18124 13557 18188
rect 13491 18123 13557 18124
rect 13123 17508 13189 17509
rect 13123 17444 13124 17508
rect 13188 17444 13189 17508
rect 13123 17443 13189 17444
rect 13126 13293 13186 17443
rect 13123 13292 13189 13293
rect 13123 13228 13124 13292
rect 13188 13228 13189 13292
rect 13123 13227 13189 13228
rect 13307 13292 13373 13293
rect 13307 13228 13308 13292
rect 13372 13228 13373 13292
rect 13307 13227 13373 13228
rect 13123 12884 13189 12885
rect 13123 12820 13124 12884
rect 13188 12820 13189 12884
rect 13123 12819 13189 12820
rect 13126 11661 13186 12819
rect 13123 11660 13189 11661
rect 13123 11596 13124 11660
rect 13188 11596 13189 11660
rect 13123 11595 13189 11596
rect 12939 11524 13005 11525
rect 12939 11460 12940 11524
rect 13004 11460 13005 11524
rect 12939 11459 13005 11460
rect 12939 10436 13005 10437
rect 12939 10372 12940 10436
rect 13004 10372 13005 10436
rect 12939 10371 13005 10372
rect 12755 9892 12821 9893
rect 12755 9828 12756 9892
rect 12820 9828 12821 9892
rect 12755 9827 12821 9828
rect 12942 9757 13002 10371
rect 12755 9756 12821 9757
rect 12755 9692 12756 9756
rect 12820 9692 12821 9756
rect 12755 9691 12821 9692
rect 12939 9756 13005 9757
rect 12939 9692 12940 9756
rect 13004 9692 13005 9756
rect 12939 9691 13005 9692
rect 12758 9621 12818 9691
rect 12755 9620 12821 9621
rect 12755 9556 12756 9620
rect 12820 9556 12821 9620
rect 12755 9555 12821 9556
rect 12571 7172 12637 7173
rect 12571 7170 12572 7172
rect 12390 7110 12572 7170
rect 12571 7108 12572 7110
rect 12636 7108 12637 7172
rect 12571 7107 12637 7108
rect 12019 6764 12085 6765
rect 12019 6700 12020 6764
rect 12084 6700 12085 6764
rect 12019 6699 12085 6700
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 10731 2820 10797 2821
rect 10731 2756 10732 2820
rect 10796 2756 10797 2820
rect 10731 2755 10797 2756
rect 10547 2548 10613 2549
rect 10547 2484 10548 2548
rect 10612 2484 10613 2548
rect 10547 2483 10613 2484
rect 11240 2208 11560 3232
rect 12022 2821 12082 6699
rect 12387 5676 12453 5677
rect 12387 5612 12388 5676
rect 12452 5612 12453 5676
rect 12387 5611 12453 5612
rect 12019 2820 12085 2821
rect 12019 2756 12020 2820
rect 12084 2756 12085 2820
rect 12019 2755 12085 2756
rect 12390 2549 12450 5611
rect 12758 3501 12818 9555
rect 12755 3500 12821 3501
rect 12755 3436 12756 3500
rect 12820 3436 12821 3500
rect 12755 3435 12821 3436
rect 12942 2957 13002 9691
rect 13126 8805 13186 11595
rect 13310 10981 13370 13227
rect 13494 12069 13554 18123
rect 13678 13293 13738 19755
rect 13862 18053 13922 20299
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14227 19548 14293 19549
rect 14227 19484 14228 19548
rect 14292 19484 14293 19548
rect 14227 19483 14293 19484
rect 14043 18188 14109 18189
rect 14043 18124 14044 18188
rect 14108 18124 14109 18188
rect 14043 18123 14109 18124
rect 13859 18052 13925 18053
rect 13859 17988 13860 18052
rect 13924 17988 13925 18052
rect 13859 17987 13925 17988
rect 13859 14244 13925 14245
rect 13859 14180 13860 14244
rect 13924 14180 13925 14244
rect 13859 14179 13925 14180
rect 13862 13701 13922 14179
rect 13859 13700 13925 13701
rect 13859 13636 13860 13700
rect 13924 13636 13925 13700
rect 13859 13635 13925 13636
rect 13675 13292 13741 13293
rect 13675 13228 13676 13292
rect 13740 13228 13741 13292
rect 13675 13227 13741 13228
rect 13675 12748 13741 12749
rect 13675 12684 13676 12748
rect 13740 12684 13741 12748
rect 13675 12683 13741 12684
rect 13491 12068 13557 12069
rect 13491 12004 13492 12068
rect 13556 12004 13557 12068
rect 13491 12003 13557 12004
rect 13307 10980 13373 10981
rect 13307 10916 13308 10980
rect 13372 10916 13373 10980
rect 13307 10915 13373 10916
rect 13307 10572 13373 10573
rect 13307 10508 13308 10572
rect 13372 10508 13373 10572
rect 13307 10507 13373 10508
rect 13123 8804 13189 8805
rect 13123 8740 13124 8804
rect 13188 8740 13189 8804
rect 13123 8739 13189 8740
rect 13310 5269 13370 10507
rect 13491 7716 13557 7717
rect 13491 7652 13492 7716
rect 13556 7652 13557 7716
rect 13491 7651 13557 7652
rect 13307 5268 13373 5269
rect 13307 5204 13308 5268
rect 13372 5204 13373 5268
rect 13307 5203 13373 5204
rect 13494 4317 13554 7651
rect 13678 4861 13738 12683
rect 13859 8940 13925 8941
rect 13859 8876 13860 8940
rect 13924 8876 13925 8940
rect 13859 8875 13925 8876
rect 13675 4860 13741 4861
rect 13675 4796 13676 4860
rect 13740 4796 13741 4860
rect 13675 4795 13741 4796
rect 13862 4725 13922 8875
rect 13859 4724 13925 4725
rect 13859 4660 13860 4724
rect 13924 4660 13925 4724
rect 13859 4659 13925 4660
rect 13859 4588 13925 4589
rect 13859 4524 13860 4588
rect 13924 4524 13925 4588
rect 13859 4523 13925 4524
rect 13491 4316 13557 4317
rect 13491 4252 13492 4316
rect 13556 4252 13557 4316
rect 13491 4251 13557 4252
rect 12939 2956 13005 2957
rect 12939 2892 12940 2956
rect 13004 2892 13005 2956
rect 12939 2891 13005 2892
rect 13862 2685 13922 4523
rect 13859 2684 13925 2685
rect 13859 2620 13860 2684
rect 13924 2620 13925 2684
rect 13859 2619 13925 2620
rect 14046 2549 14106 18123
rect 14230 3773 14290 19483
rect 14411 19412 14477 19413
rect 14411 19348 14412 19412
rect 14476 19348 14477 19412
rect 14411 19347 14477 19348
rect 14227 3772 14293 3773
rect 14227 3708 14228 3772
rect 14292 3708 14293 3772
rect 14227 3707 14293 3708
rect 14414 3637 14474 19347
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 15147 18732 15213 18733
rect 15147 18668 15148 18732
rect 15212 18668 15213 18732
rect 15147 18667 15213 18668
rect 15883 18732 15949 18733
rect 15883 18668 15884 18732
rect 15948 18668 15949 18732
rect 15883 18667 15949 18668
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 15150 13021 15210 18667
rect 15515 18324 15581 18325
rect 15515 18260 15516 18324
rect 15580 18260 15581 18324
rect 15515 18259 15581 18260
rect 15331 18188 15397 18189
rect 15331 18124 15332 18188
rect 15396 18124 15397 18188
rect 15331 18123 15397 18124
rect 15334 15061 15394 18123
rect 15331 15060 15397 15061
rect 15331 14996 15332 15060
rect 15396 14996 15397 15060
rect 15331 14995 15397 14996
rect 15518 14789 15578 18259
rect 15699 18052 15765 18053
rect 15699 17988 15700 18052
rect 15764 17988 15765 18052
rect 15699 17987 15765 17988
rect 15515 14788 15581 14789
rect 15515 14724 15516 14788
rect 15580 14724 15581 14788
rect 15515 14723 15581 14724
rect 15331 14244 15397 14245
rect 15331 14180 15332 14244
rect 15396 14180 15397 14244
rect 15331 14179 15397 14180
rect 15147 13020 15213 13021
rect 15147 12956 15148 13020
rect 15212 12956 15213 13020
rect 15147 12955 15213 12956
rect 15147 12612 15213 12613
rect 15147 12548 15148 12612
rect 15212 12548 15213 12612
rect 15147 12547 15213 12548
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 15150 9349 15210 12547
rect 15334 9893 15394 14179
rect 15518 11117 15578 14723
rect 15515 11116 15581 11117
rect 15515 11052 15516 11116
rect 15580 11052 15581 11116
rect 15515 11051 15581 11052
rect 15331 9892 15397 9893
rect 15331 9828 15332 9892
rect 15396 9828 15397 9892
rect 15331 9827 15397 9828
rect 15147 9348 15213 9349
rect 15147 9284 15148 9348
rect 15212 9284 15213 9348
rect 15147 9283 15213 9284
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 15150 4589 15210 9283
rect 15702 8533 15762 17987
rect 15886 16693 15946 18667
rect 18104 18528 18424 19552
rect 19931 19412 19997 19413
rect 19931 19348 19932 19412
rect 19996 19348 19997 19412
rect 19931 19347 19997 19348
rect 18827 18732 18893 18733
rect 18827 18668 18828 18732
rect 18892 18668 18893 18732
rect 18827 18667 18893 18668
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 17171 18188 17237 18189
rect 17171 18124 17172 18188
rect 17236 18124 17237 18188
rect 17171 18123 17237 18124
rect 16067 18052 16133 18053
rect 16067 17988 16068 18052
rect 16132 17988 16133 18052
rect 16067 17987 16133 17988
rect 16435 18052 16501 18053
rect 16435 17988 16436 18052
rect 16500 17988 16501 18052
rect 16435 17987 16501 17988
rect 16619 18052 16685 18053
rect 16619 17988 16620 18052
rect 16684 17988 16685 18052
rect 16619 17987 16685 17988
rect 15883 16692 15949 16693
rect 15883 16628 15884 16692
rect 15948 16628 15949 16692
rect 15883 16627 15949 16628
rect 15883 15060 15949 15061
rect 15883 14996 15884 15060
rect 15948 14996 15949 15060
rect 15883 14995 15949 14996
rect 15886 11389 15946 14995
rect 15883 11388 15949 11389
rect 15883 11324 15884 11388
rect 15948 11324 15949 11388
rect 15883 11323 15949 11324
rect 15699 8532 15765 8533
rect 15699 8468 15700 8532
rect 15764 8468 15765 8532
rect 15699 8467 15765 8468
rect 15147 4588 15213 4589
rect 15147 4524 15148 4588
rect 15212 4524 15213 4588
rect 15147 4523 15213 4524
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14411 3636 14477 3637
rect 14411 3572 14412 3636
rect 14476 3572 14477 3636
rect 14411 3571 14477 3572
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 12387 2548 12453 2549
rect 12387 2484 12388 2548
rect 12452 2484 12453 2548
rect 12387 2483 12453 2484
rect 14043 2548 14109 2549
rect 14043 2484 14044 2548
rect 14108 2484 14109 2548
rect 14043 2483 14109 2484
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 2128 14992 2688
rect 16070 2685 16130 17987
rect 16251 15604 16317 15605
rect 16251 15540 16252 15604
rect 16316 15540 16317 15604
rect 16251 15539 16317 15540
rect 16254 8805 16314 15539
rect 16251 8804 16317 8805
rect 16251 8740 16252 8804
rect 16316 8740 16317 8804
rect 16251 8739 16317 8740
rect 16438 2685 16498 17987
rect 16622 12341 16682 17987
rect 16987 17372 17053 17373
rect 16987 17308 16988 17372
rect 17052 17308 17053 17372
rect 16987 17307 17053 17308
rect 16803 16556 16869 16557
rect 16803 16492 16804 16556
rect 16868 16492 16869 16556
rect 16803 16491 16869 16492
rect 16619 12340 16685 12341
rect 16619 12276 16620 12340
rect 16684 12276 16685 12340
rect 16619 12275 16685 12276
rect 16806 11250 16866 16491
rect 16990 14653 17050 17307
rect 16987 14652 17053 14653
rect 16987 14588 16988 14652
rect 17052 14588 17053 14652
rect 16987 14587 17053 14588
rect 17174 13973 17234 18123
rect 17907 18052 17973 18053
rect 17907 17988 17908 18052
rect 17972 17988 17973 18052
rect 17907 17987 17973 17988
rect 17723 16692 17789 16693
rect 17723 16628 17724 16692
rect 17788 16628 17789 16692
rect 17723 16627 17789 16628
rect 17171 13972 17237 13973
rect 17171 13908 17172 13972
rect 17236 13908 17237 13972
rect 17171 13907 17237 13908
rect 16987 13836 17053 13837
rect 16987 13772 16988 13836
rect 17052 13772 17053 13836
rect 16987 13771 17053 13772
rect 16622 11190 16866 11250
rect 16622 3909 16682 11190
rect 16990 10709 17050 13771
rect 17171 13156 17237 13157
rect 17171 13092 17172 13156
rect 17236 13092 17237 13156
rect 17171 13091 17237 13092
rect 16987 10708 17053 10709
rect 16987 10644 16988 10708
rect 17052 10644 17053 10708
rect 16987 10643 17053 10644
rect 17174 9893 17234 13091
rect 17355 12612 17421 12613
rect 17355 12548 17356 12612
rect 17420 12548 17421 12612
rect 17355 12547 17421 12548
rect 17539 12612 17605 12613
rect 17539 12548 17540 12612
rect 17604 12548 17605 12612
rect 17539 12547 17605 12548
rect 17358 10029 17418 12547
rect 17542 11797 17602 12547
rect 17539 11796 17605 11797
rect 17539 11732 17540 11796
rect 17604 11732 17605 11796
rect 17539 11731 17605 11732
rect 17355 10028 17421 10029
rect 17355 9964 17356 10028
rect 17420 9964 17421 10028
rect 17355 9963 17421 9964
rect 17171 9892 17237 9893
rect 17171 9828 17172 9892
rect 17236 9828 17237 9892
rect 17171 9827 17237 9828
rect 17355 9212 17421 9213
rect 17355 9148 17356 9212
rect 17420 9148 17421 9212
rect 17355 9147 17421 9148
rect 16803 8668 16869 8669
rect 16803 8604 16804 8668
rect 16868 8604 16869 8668
rect 16803 8603 16869 8604
rect 16619 3908 16685 3909
rect 16619 3844 16620 3908
rect 16684 3844 16685 3908
rect 16619 3843 16685 3844
rect 16806 3093 16866 8603
rect 16803 3092 16869 3093
rect 16803 3028 16804 3092
rect 16868 3028 16869 3092
rect 16803 3027 16869 3028
rect 16067 2684 16133 2685
rect 16067 2620 16068 2684
rect 16132 2620 16133 2684
rect 16067 2619 16133 2620
rect 16435 2684 16501 2685
rect 16435 2620 16436 2684
rect 16500 2620 16501 2684
rect 16435 2619 16501 2620
rect 17358 1869 17418 9147
rect 17726 5813 17786 16627
rect 17723 5812 17789 5813
rect 17723 5748 17724 5812
rect 17788 5748 17789 5812
rect 17723 5747 17789 5748
rect 17910 3773 17970 17987
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18643 16692 18709 16693
rect 18643 16628 18644 16692
rect 18708 16628 18709 16692
rect 18643 16627 18709 16628
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18646 14517 18706 16627
rect 18643 14516 18709 14517
rect 18643 14452 18644 14516
rect 18708 14452 18709 14516
rect 18643 14451 18709 14452
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18830 11117 18890 18667
rect 19195 18460 19261 18461
rect 19195 18396 19196 18460
rect 19260 18396 19261 18460
rect 19195 18395 19261 18396
rect 19379 18460 19445 18461
rect 19379 18396 19380 18460
rect 19444 18396 19445 18460
rect 19379 18395 19445 18396
rect 19011 13020 19077 13021
rect 19011 12956 19012 13020
rect 19076 12956 19077 13020
rect 19011 12955 19077 12956
rect 18827 11116 18893 11117
rect 18827 11052 18828 11116
rect 18892 11052 18893 11116
rect 18827 11051 18893 11052
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 19014 8805 19074 12955
rect 19198 12341 19258 18395
rect 19382 13565 19442 18395
rect 19747 18052 19813 18053
rect 19747 17988 19748 18052
rect 19812 17988 19813 18052
rect 19747 17987 19813 17988
rect 19563 17916 19629 17917
rect 19563 17852 19564 17916
rect 19628 17852 19629 17916
rect 19563 17851 19629 17852
rect 19566 13701 19626 17851
rect 19563 13700 19629 13701
rect 19563 13636 19564 13700
rect 19628 13636 19629 13700
rect 19563 13635 19629 13636
rect 19379 13564 19445 13565
rect 19379 13500 19380 13564
rect 19444 13500 19445 13564
rect 19379 13499 19445 13500
rect 19379 13020 19445 13021
rect 19379 12956 19380 13020
rect 19444 12956 19445 13020
rect 19379 12955 19445 12956
rect 19195 12340 19261 12341
rect 19195 12276 19196 12340
rect 19260 12276 19261 12340
rect 19195 12275 19261 12276
rect 19382 10029 19442 12955
rect 19379 10028 19445 10029
rect 19379 9964 19380 10028
rect 19444 9964 19445 10028
rect 19379 9963 19445 9964
rect 19195 9484 19261 9485
rect 19195 9420 19196 9484
rect 19260 9420 19261 9484
rect 19195 9419 19261 9420
rect 19011 8804 19077 8805
rect 19011 8740 19012 8804
rect 19076 8740 19077 8804
rect 19011 8739 19077 8740
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 19011 7988 19077 7989
rect 19011 7924 19012 7988
rect 19076 7924 19077 7988
rect 19011 7923 19077 7924
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18643 7580 18709 7581
rect 18643 7516 18644 7580
rect 18708 7516 18709 7580
rect 18643 7515 18709 7516
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 17907 3772 17973 3773
rect 17907 3708 17908 3772
rect 17972 3708 17973 3772
rect 17907 3707 17973 3708
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18646 2957 18706 7515
rect 18827 7172 18893 7173
rect 18827 7108 18828 7172
rect 18892 7108 18893 7172
rect 18827 7107 18893 7108
rect 18643 2956 18709 2957
rect 18643 2892 18644 2956
rect 18708 2892 18709 2956
rect 18643 2891 18709 2892
rect 18830 2821 18890 7107
rect 19014 5813 19074 7923
rect 19011 5812 19077 5813
rect 19011 5748 19012 5812
rect 19076 5748 19077 5812
rect 19011 5747 19077 5748
rect 19198 3637 19258 9419
rect 19195 3636 19261 3637
rect 19195 3572 19196 3636
rect 19260 3572 19261 3636
rect 19195 3571 19261 3572
rect 19750 3229 19810 17987
rect 19747 3228 19813 3229
rect 19747 3164 19748 3228
rect 19812 3164 19813 3228
rect 19747 3163 19813 3164
rect 19934 3093 19994 19347
rect 20483 18188 20549 18189
rect 20483 18124 20484 18188
rect 20548 18124 20549 18188
rect 20483 18123 20549 18124
rect 20299 15332 20365 15333
rect 20299 15268 20300 15332
rect 20364 15268 20365 15332
rect 20299 15267 20365 15268
rect 19931 3092 19997 3093
rect 19931 3028 19932 3092
rect 19996 3028 19997 3092
rect 19931 3027 19997 3028
rect 18827 2820 18893 2821
rect 18827 2756 18828 2820
rect 18892 2756 18893 2820
rect 18827 2755 18893 2756
rect 20302 2549 20362 15267
rect 20486 2685 20546 18123
rect 20483 2684 20549 2685
rect 20483 2620 20484 2684
rect 20548 2620 20549 2684
rect 20483 2619 20549 2620
rect 20299 2548 20365 2549
rect 20299 2484 20300 2548
rect 20364 2484 20365 2548
rect 20299 2483 20365 2484
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
rect 17355 1868 17421 1869
rect 17355 1804 17356 1868
rect 17420 1804 17421 1868
rect 17355 1803 17421 1804
use sky130_fd_sc_hd__decap_8  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1605641404
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1748 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2576 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 2760 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1605641404
transform 1 0 2116 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_20
timestamp 1605641404
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_4_
timestamp 1605641404
transform 1 0 2944 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3128 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4784 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4600 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1605641404
transform 1 0 4416 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1605641404
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32
timestamp 1605641404
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_38
timestamp 1605641404
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 6808 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_5_
timestamp 1605641404
transform 1 0 5796 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1605641404
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1605641404
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47
timestamp 1605641404
transform 1 0 5428 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1605641404
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_56
timestamp 1605641404
transform 1 0 6256 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 8740 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_4_
timestamp 1605641404
transform 1 0 7912 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_2_
timestamp 1605641404
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72
timestamp 1605641404
transform 1 0 7728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83
timestamp 1605641404
transform 1 0 8740 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_78
timestamp 1605641404
transform 1 0 8280 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_82
timestamp 1605641404
transform 1 0 8648 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _109_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 9108 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 10396 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1605641404
transform 1 0 9844 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1605641404
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_91
timestamp 1605641404
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94
timestamp 1605641404
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_104
timestamp 1605641404
transform 1 0 10672 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_99
timestamp 1605641404
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 10856 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1605641404
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1605641404
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1605641404
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1605641404
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_125
timestamp 1605641404
transform 1 0 12604 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_117
timestamp 1605641404
transform 1 0 11868 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1605641404
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1605641404
transform 1 0 12696 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13432 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13708 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1605641404
transform 1 0 14444 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_135
timestamp 1605641404
transform 1 0 13524 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1605641404
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_143
timestamp 1605641404
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1605641404
transform 1 0 14812 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1605641404
transform 1 0 15456 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1605641404
transform 1 0 15456 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1605641404
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_146
timestamp 1605641404
transform 1 0 14536 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1605641404
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_165
timestamp 1605641404
transform 1 0 16284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_154
timestamp 1605641404
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_165 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 16284 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_171
timestamp 1605641404
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_176
timestamp 1605641404
transform 1 0 17296 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1605641404
transform 1 0 16928 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 16468 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_184
timestamp 1605641404
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1605641404
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1605641404
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1605641404
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1605641404
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 17480 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_187
timestamp 1605641404
transform 1 0 18308 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1605641404
transform 1 0 18492 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1605641404
transform 1 0 20056 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_3_
timestamp 1605641404
transform 1 0 19412 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1605641404
transform 1 0 19044 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_1_
timestamp 1605641404
transform 1 0 18400 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_0_193
timestamp 1605641404
transform 1 0 18860 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_204
timestamp 1605641404
transform 1 0 19872 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_197
timestamp 1605641404
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_208
timestamp 1605641404
transform 1 0 20240 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1605641404
transform 1 0 20516 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1605641404
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1605641404
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1605641404
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1605641404
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1605641404
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1605641404
transform 1 0 20884 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_219
timestamp 1605641404
transform 1 0 21252 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_3_
timestamp 1605641404
transform 1 0 1932 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1605641404
transform 1 0 2944 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1605641404
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1605641404
transform 1 0 1380 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_18
timestamp 1605641404
transform 1 0 2760 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1605641404
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1605641404
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_41
timestamp 1605641404
transform 1 0 4876 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 5704 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_2_49
timestamp 1605641404
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1605641404
transform 1 0 8556 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1605641404
transform 1 0 7360 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1605641404
transform 1 0 8372 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_66
timestamp 1605641404
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_77
timestamp 1605641404
transform 1 0 8188 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1605641404
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1605641404
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1605641404
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_90
timestamp 1605641404
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_104
timestamp 1605641404
transform 1 0 10672 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1605641404
transform 1 0 11500 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1605641404
transform 1 0 12512 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 10764 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_111
timestamp 1605641404
transform 1 0 11316 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_122
timestamp 1605641404
transform 1 0 12328 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1605641404
transform 1 0 13524 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_133
timestamp 1605641404
transform 1 0 13340 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_144
timestamp 1605641404
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 16376 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1605641404
transform 1 0 14536 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_3_
timestamp 1605641404
transform 1 0 15364 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1605641404
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_150
timestamp 1605641404
transform 1 0 14904 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_154
timestamp 1605641404
transform 1 0 15272 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_164
timestamp 1605641404
transform 1 0 16192 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1605641404
transform 1 0 17848 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_2_
timestamp 1605641404
transform 1 0 16836 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_169
timestamp 1605641404
transform 1 0 16652 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_180
timestamp 1605641404
transform 1 0 17664 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 18860 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1605641404
transform 1 0 19596 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_191
timestamp 1605641404
transform 1 0 18676 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_199
timestamp 1605641404
transform 1 0 19412 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1605641404
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1605641404
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_210
timestamp 1605641404
transform 1 0 20424 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1605641404
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1605641404
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 2024 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1605641404
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1605641404
transform 1 0 1380 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_9
timestamp 1605641404
transform 1 0 1932 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_4_
timestamp 1605641404
transform 1 0 4048 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1605641404
transform 1 0 4876 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_3_26
timestamp 1605641404
transform 1 0 3496 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_1_
timestamp 1605641404
transform 1 0 5704 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1605641404
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1605641404
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_62
timestamp 1605641404
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8464 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1605641404
transform 1 0 6992 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_3_73
timestamp 1605641404
transform 1 0 7820 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_79
timestamp 1605641404
transform 1 0 8372 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1605641404
transform 1 0 10120 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_96
timestamp 1605641404
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12420 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1605641404
transform 1 0 11132 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1605641404
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_107
timestamp 1605641404
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_118
timestamp 1605641404
transform 1 0 11960 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14076 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_139
timestamp 1605641404
transform 1 0 13892 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1605641404
transform 1 0 16284 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1605641404
transform 1 0 15272 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_3_150
timestamp 1605641404
transform 1 0 14904 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_163
timestamp 1605641404
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1605641404
transform 1 0 17388 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1605641404
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1605641404
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_174
timestamp 1605641404
transform 1 0 17112 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1605641404
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 18952 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1605641404
transform 1 0 19872 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1605641404
transform 1 0 19688 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_193
timestamp 1605641404
transform 1 0 18860 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_200
timestamp 1605641404
transform 1 0 19504 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1605641404
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_213
timestamp 1605641404
transform 1 0 20700 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_219
timestamp 1605641404
transform 1 0 21252 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1605641404
transform 1 0 2852 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1605641404
transform 1 0 2024 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1605641404
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp 1605641404
transform 1 0 1380 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_9
timestamp 1605641404
transform 1 0 1932 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1605641404
transform 1 0 3128 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1605641404
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1605641404
transform 1 0 4876 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_32
timestamp 1605641404
transform 1 0 4048 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_40
timestamp 1605641404
transform 1 0 4784 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1605641404
transform 1 0 6256 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1605641404
transform 1 0 5060 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_52
timestamp 1605641404
transform 1 0 5888 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1605641404
transform 1 0 7912 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_72
timestamp 1605641404
transform 1 0 7728 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_83
timestamp 1605641404
transform 1 0 8740 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1605641404
transform 1 0 10672 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1605641404
transform 1 0 9016 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1605641404
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1605641404
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1605641404
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_102
timestamp 1605641404
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1605641404
transform 1 0 11040 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1605641404
transform 1 0 12236 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1605641404
transform 1 0 12052 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_117
timestamp 1605641404
transform 1 0 11868 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13248 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_4_
timestamp 1605641404
transform 1 0 14168 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_130
timestamp 1605641404
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_138
timestamp 1605641404
transform 1 0 13800 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15272 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1605641404
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1605641404
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 17388 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_4_170
timestamp 1605641404
transform 1 0 16744 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_176
timestamp 1605641404
transform 1 0 17296 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1605641404
transform 1 0 19044 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1605641404
transform 1 0 19596 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_193
timestamp 1605641404
transform 1 0 18860 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_199
timestamp 1605641404
transform 1 0 19412 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1605641404
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1605641404
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1605641404
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_210
timestamp 1605641404
transform 1 0 20424 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_218
timestamp 1605641404
transform 1 0 21160 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1605641404
transform 1 0 2024 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1605641404
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1605641404
transform 1 0 1380 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_9
timestamp 1605641404
transform 1 0 1932 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_19
timestamp 1605641404
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4324 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1605641404
transform 1 0 3036 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_30
timestamp 1605641404
transform 1 0 3864 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_34
timestamp 1605641404
transform 1 0 4232 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l5_in_0_
timestamp 1605641404
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1605641404
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1605641404
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1605641404
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8096 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_71
timestamp 1605641404
transform 1 0 7636 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_75
timestamp 1605641404
transform 1 0 8004 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1605641404
transform 1 0 10580 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1605641404
transform 1 0 9568 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_85
timestamp 1605641404
transform 1 0 8924 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_91
timestamp 1605641404
transform 1 0 9476 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_101
timestamp 1605641404
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 11592 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1605641404
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_112
timestamp 1605641404
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1605641404
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 13432 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1605641404
transform 1 0 14260 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_132
timestamp 1605641404
transform 1 0 13248 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_140
timestamp 1605641404
transform 1 0 13984 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1605641404
transform 1 0 16376 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1605641404
transform 1 0 15272 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_152
timestamp 1605641404
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_163
timestamp 1605641404
transform 1 0 16100 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_4_
timestamp 1605641404
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1605641404
transform 1 0 16928 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1605641404
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_170
timestamp 1605641404
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1605641404
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 19320 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_193
timestamp 1605641404
transform 1 0 18860 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_197
timestamp 1605641404
transform 1 0 19228 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1605641404
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_214
timestamp 1605641404
transform 1 0 20792 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 1748 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 1472 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1605641404
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1605641404
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1605641404
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1605641404
transform 1 0 1380 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_20
timestamp 1605641404
transform 1 0 2944 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1605641404
transform 1 0 3404 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4048 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4600 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1605641404
transform 1 0 3496 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1605641404
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_23
timestamp 1605641404
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_28
timestamp 1605641404
transform 1 0 3680 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_35
timestamp 1605641404
transform 1 0 4324 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_3_
timestamp 1605641404
transform 1 0 6256 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1605641404
transform 1 0 5612 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1605641404
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_48
timestamp 1605641404
transform 1 0 5520 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_47
timestamp 1605641404
transform 1 0 5428 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_58
timestamp 1605641404
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_62
timestamp 1605641404
transform 1 0 6808 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7268 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_7_
timestamp 1605641404
transform 1 0 6900 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1605641404
transform 1 0 8004 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_65
timestamp 1605641404
transform 1 0 7084 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_83
timestamp 1605641404
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_72
timestamp 1605641404
transform 1 0 7728 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1605641404
transform 1 0 8924 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9660 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9016 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1605641404
transform 1 0 10672 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1605641404
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_88
timestamp 1605641404
transform 1 0 9200 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_84
timestamp 1605641404
transform 1 0 8832 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_102
timestamp 1605641404
transform 1 0 10488 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1605641404
transform 1 0 11776 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 12420 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12328 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1605641404
transform 1 0 11316 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1605641404
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_109
timestamp 1605641404
transform 1 0 11132 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_120
timestamp 1605641404
transform 1 0 12144 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_113
timestamp 1605641404
transform 1 0 11500 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1605641404
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_4_
timestamp 1605641404
transform 1 0 14168 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1605641404
transform 1 0 14168 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1605641404
transform 1 0 13984 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1605641404
transform 1 0 13800 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_139
timestamp 1605641404
transform 1 0 13892 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 15272 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 15180 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1605641404
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1605641404
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_151
timestamp 1605641404
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1605641404
transform 1 0 16836 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1605641404
transform 1 0 16928 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1605641404
transform 1 0 17940 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1605641404
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_170
timestamp 1605641404
transform 1 0 16744 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_181
timestamp 1605641404
transform 1 0 17756 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1605641404
transform 1 0 16652 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_180
timestamp 1605641404
transform 1 0 17664 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_184
timestamp 1605641404
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1605641404
transform 1 0 18952 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1605641404
transform 1 0 18400 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 18952 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1605641404
transform 1 0 19504 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_192
timestamp 1605641404
transform 1 0 18768 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_198
timestamp 1605641404
transform 1 0 19320 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_192
timestamp 1605641404
transform 1 0 18768 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_210
timestamp 1605641404
transform 1 0 20424 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1605641404
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1605641404
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_209
timestamp 1605641404
transform 1 0 20332 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1605641404
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 20608 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_218
timestamp 1605641404
transform 1 0 21160 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1605641404
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1605641404
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1605641404
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1605641404
transform 1 0 2024 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1605641404
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1605641404
transform 1 0 1380 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1605641404
transform 1 0 1932 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_19
timestamp 1605641404
transform 1 0 2852 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4508 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 3036 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1605641404
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1605641404
transform 1 0 4324 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1605641404
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_8_32
timestamp 1605641404
transform 1 0 4048 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1605641404
transform 1 0 5520 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_46
timestamp 1605641404
transform 1 0 5336 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_57
timestamp 1605641404
transform 1 0 6348 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1605641404
transform 1 0 7912 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_6_
timestamp 1605641404
transform 1 0 6900 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_72
timestamp 1605641404
transform 1 0 7728 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_83
timestamp 1605641404
transform 1 0 8740 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_4_
timestamp 1605641404
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1605641404
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1605641404
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_102
timestamp 1605641404
transform 1 0 10488 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1605641404
transform 1 0 10856 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 11316 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_109
timestamp 1605641404
transform 1 0 11132 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1605641404
transform 1 0 12972 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14168 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_127
timestamp 1605641404
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_138
timestamp 1605641404
transform 1 0 13800 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1605641404
transform 1 0 15364 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1605641404
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1605641404
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_154
timestamp 1605641404
transform 1 0 15272 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_164
timestamp 1605641404
transform 1 0 16192 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 16560 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_184
timestamp 1605641404
transform 1 0 18032 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1605641404
transform 1 0 18492 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 19136 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_188
timestamp 1605641404
transform 1 0 18400 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_193
timestamp 1605641404
transform 1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1605641404
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1605641404
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1605641404
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1605641404
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1605641404
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2484 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1605641404
transform 1 0 1472 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1605641404
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1605641404
transform 1 0 1380 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_13
timestamp 1605641404
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_4_
timestamp 1605641404
transform 1 0 4140 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_31
timestamp 1605641404
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1605641404
transform 1 0 5704 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1605641404
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_42
timestamp 1605641404
transform 1 0 4968 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1605641404
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_62
timestamp 1605641404
transform 1 0 6808 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7360 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1605641404
transform 1 0 8832 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_3_
timestamp 1605641404
transform 1 0 10488 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1605641404
transform 1 0 9476 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1605641404
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_87
timestamp 1605641404
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_100
timestamp 1605641404
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1605641404
transform 1 0 11776 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1605641404
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_111
timestamp 1605641404
transform 1 0 11316 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_115
timestamp 1605641404
transform 1 0 11684 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1605641404
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1605641404
transform 1 0 13800 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 14352 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 13432 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1605641404
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_137
timestamp 1605641404
transform 1 0 13708 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_142
timestamp 1605641404
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1605641404
transform 1 0 16192 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1605641404
transform 1 0 15364 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_153
timestamp 1605641404
transform 1 0 15180 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16928 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1605641404
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1605641404
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1605641404
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_168
timestamp 1605641404
transform 1 0 16560 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1605641404
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 19320 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_193
timestamp 1605641404
transform 1 0 18860 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_197
timestamp 1605641404
transform 1 0 19228 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1605641404
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_214
timestamp 1605641404
transform 1 0 20792 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1605641404
transform 1 0 1472 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1605641404
transform 1 0 2484 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1605641404
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1605641404
transform 1 0 1380 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_13
timestamp 1605641404
transform 1 0 2300 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1605641404
transform 1 0 3496 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4324 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1605641404
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_24
timestamp 1605641404
transform 1 0 3312 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1605641404
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_32
timestamp 1605641404
transform 1 0 4048 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1605641404
transform 1 0 5980 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_51
timestamp 1605641404
transform 1 0 5796 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_62
timestamp 1605641404
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8556 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1605641404
transform 1 0 6992 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1605641404
transform 1 0 8188 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_73
timestamp 1605641404
transform 1 0 7820 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_80
timestamp 1605641404
transform 1 0 8464 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1605641404
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1605641404
transform 1 0 10672 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1605641404
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1605641404
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_102
timestamp 1605641404
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1605641404
transform 1 0 11684 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_113
timestamp 1605641404
transform 1 0 11500 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_124
timestamp 1605641404
transform 1 0 12512 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1605641404
transform 1 0 13708 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1605641404
transform 1 0 12696 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_135
timestamp 1605641404
transform 1 0 13524 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1605641404
transform 1 0 14720 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1605641404
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1605641404
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_146
timestamp 1605641404
transform 1 0 14536 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1605641404
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_163
timestamp 1605641404
transform 1 0 16100 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1605641404
transform 1 0 16468 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 17020 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_171
timestamp 1605641404
transform 1 0 16836 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1605641404
transform 1 0 19688 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1605641404
transform 1 0 18676 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_189
timestamp 1605641404
transform 1 0 18492 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_200
timestamp 1605641404
transform 1 0 19504 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1605641404
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1605641404
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1605641404
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_211
timestamp 1605641404
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_218
timestamp 1605641404
transform 1 0 21160 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 1380 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1605641404
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_19
timestamp 1605641404
transform 1 0 2852 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 3680 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_27
timestamp 1605641404
transform 1 0 3588 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1605641404
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1605641404
transform 1 0 5336 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1605641404
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1605641404
transform 1 0 6348 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_44
timestamp 1605641404
transform 1 0 5152 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_55
timestamp 1605641404
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1605641404
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8280 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_11_71
timestamp 1605641404
transform 1 0 7636 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_77
timestamp 1605641404
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1605641404
transform 1 0 10120 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1605641404
transform 1 0 9936 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_94
timestamp 1605641404
transform 1 0 9752 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12420 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1605641404
transform 1 0 11132 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1605641404
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_107
timestamp 1605641404
transform 1 0 10948 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_118
timestamp 1605641404
transform 1 0 11960 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1605641404
transform 1 0 14076 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_139
timestamp 1605641404
transform 1 0 13892 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_3_
timestamp 1605641404
transform 1 0 16100 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1605641404
transform 1 0 15088 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_150
timestamp 1605641404
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_161
timestamp 1605641404
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1605641404
transform 1 0 17112 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1605641404
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1605641404
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1605641404
transform 1 0 17664 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_172
timestamp 1605641404
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_178
timestamp 1605641404
transform 1 0 17480 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1605641404
transform 1 0 19044 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1605641404
transform 1 0 20056 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_193
timestamp 1605641404
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_204
timestamp 1605641404
transform 1 0 19872 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1605641404
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_215
timestamp 1605641404
transform 1 0 20884 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_219
timestamp 1605641404
transform 1 0 21252 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2300 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1605641404
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_3
timestamp 1605641404
transform 1 0 1380 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_11
timestamp 1605641404
transform 1 0 2116 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4876 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1605641404
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1605641404
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_32
timestamp 1605641404
transform 1 0 4048 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_40
timestamp 1605641404
transform 1 0 4784 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1605641404
transform 1 0 5888 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_50
timestamp 1605641404
transform 1 0 5704 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_61
timestamp 1605641404
transform 1 0 6716 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6900 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1605641404
transform 1 0 7912 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_72
timestamp 1605641404
transform 1 0 7728 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_83
timestamp 1605641404
transform 1 0 8740 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1605641404
transform 1 0 9752 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1605641404
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1605641404
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_93
timestamp 1605641404
transform 1 0 9660 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_103
timestamp 1605641404
transform 1 0 10580 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l4_in_0_
timestamp 1605641404
transform 1 0 11776 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1605641404
transform 1 0 10764 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_114
timestamp 1605641404
transform 1 0 11592 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_125
timestamp 1605641404
transform 1 0 12604 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 13340 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15272 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1605641404
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1605641404
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1605641404
transform 1 0 17940 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1605641404
transform 1 0 16928 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_170
timestamp 1605641404
transform 1 0 16744 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_181
timestamp 1605641404
transform 1 0 17756 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_2_
timestamp 1605641404
transform 1 0 18952 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 19964 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_192
timestamp 1605641404
transform 1 0 18768 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_203
timestamp 1605641404
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1605641404
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1605641404
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_211
timestamp 1605641404
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1605641404
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1605641404
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1605641404
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_6
timestamp 1605641404
transform 1 0 1656 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1605641404
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1605641404
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_3_
timestamp 1605641404
transform 1 0 1748 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_2_
timestamp 1605641404
transform 1 0 1840 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1605641404
transform 1 0 1380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_16
timestamp 1605641404
transform 1 0 2576 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_17
timestamp 1605641404
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_7_
timestamp 1605641404
transform 1 0 2852 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 4232 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4048 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1605641404
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_28
timestamp 1605641404
transform 1 0 3680 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1605641404
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1605641404
transform 1 0 5888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 6808 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_1_
timestamp 1605641404
transform 1 0 5704 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1605641404
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_50
timestamp 1605641404
transform 1 0 5704 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_55
timestamp 1605641404
transform 1 0 6164 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_48
timestamp 1605641404
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_59
timestamp 1605641404
transform 1 0 6532 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7360 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1605641404
transform 1 0 7084 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_78
timestamp 1605641404
transform 1 0 8280 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9108 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1605641404
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_86
timestamp 1605641404
transform 1 0 9016 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_103
timestamp 1605641404
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_84
timestamp 1605641404
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_109
timestamp 1605641404
transform 1 0 11132 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_114
timestamp 1605641404
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1605641404
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1605641404
transform 1 0 11316 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_120
timestamp 1605641404
transform 1 0 12144 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_119
timestamp 1605641404
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1605641404
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1605641404
transform 1 0 12328 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1605641404
transform 1 0 11776 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12420 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1605641404
transform 1 0 14168 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_1_
timestamp 1605641404
transform 1 0 13340 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1605641404
transform 1 0 14352 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_139
timestamp 1605641404
transform 1 0 13892 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_145
timestamp 1605641404
transform 1 0 14444 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_131
timestamp 1605641404
transform 1 0 13156 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_142
timestamp 1605641404
transform 1 0 14168 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1605641404
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_147
timestamp 1605641404
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1605641404
transform 1 0 14812 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1605641404
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_163
timestamp 1605641404
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_163
timestamp 1605641404
transform 1 0 16100 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1605641404
transform 1 0 16284 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16284 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 14628 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1605641404
transform 1 0 17388 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 18032 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l4_in_0_
timestamp 1605641404
transform 1 0 17296 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1605641404
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_174
timestamp 1605641404
transform 1 0 17112 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1605641404
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_174
timestamp 1605641404
transform 1 0 17112 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_185
timestamp 1605641404
transform 1 0 18124 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1605641404
transform 1 0 18400 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1605641404
transform 1 0 18952 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1605641404
transform 1 0 19688 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_200
timestamp 1605641404
transform 1 0 19504 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_192
timestamp 1605641404
transform 1 0 18768 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1605641404
transform 1 0 20700 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1605641404
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1605641404
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1605641404
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_211
timestamp 1605641404
transform 1 0 20516 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_217
timestamp 1605641404
transform 1 0 21068 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_210
timestamp 1605641404
transform 1 0 20424 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1605641404
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1605641404
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_1_
timestamp 1605641404
transform 1 0 1656 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1605641404
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1605641404
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_15
timestamp 1605641404
transform 1 0 2484 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l4_in_0_
timestamp 1605641404
transform 1 0 4784 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1605641404
transform 1 0 3588 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1605641404
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_23
timestamp 1605641404
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_36
timestamp 1605641404
transform 1 0 4416 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1605641404
transform 1 0 5888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_2_
timestamp 1605641404
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1605641404
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_49
timestamp 1605641404
transform 1 0 5612 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_55
timestamp 1605641404
transform 1 0 6164 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1605641404
transform 1 0 7820 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_71
timestamp 1605641404
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_82
timestamp 1605641404
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 9844 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8832 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_93
timestamp 1605641404
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 12420 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_2_
timestamp 1605641404
transform 1 0 11500 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1605641404
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_111
timestamp 1605641404
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1605641404
transform 1 0 14076 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_139
timestamp 1605641404
transform 1 0 13892 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 15180 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_15_150
timestamp 1605641404
transform 1 0 14904 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_1_
timestamp 1605641404
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1605641404
transform 1 0 16836 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1605641404
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1605641404
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_180
timestamp 1605641404
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 19504 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_15_193
timestamp 1605641404
transform 1 0 18860 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_199
timestamp 1605641404
transform 1 0 19412 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1605641404
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_216
timestamp 1605641404
transform 1 0 20976 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1605641404
transform 1 0 1748 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 2300 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1605641404
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1605641404
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_11
timestamp 1605641404
transform 1 0 2116 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_3_
timestamp 1605641404
transform 1 0 4416 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1605641404
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1605641404
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_32
timestamp 1605641404
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6716 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_3_
timestamp 1605641404
transform 1 0 5428 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1605641404
transform 1 0 6440 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_45
timestamp 1605641404
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_56
timestamp 1605641404
transform 1 0 6256 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1605641404
transform 1 0 8372 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_77
timestamp 1605641404
transform 1 0 8188 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1605641404
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 10488 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_16_88
timestamp 1605641404
transform 1 0 9200 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_93
timestamp 1605641404
transform 1 0 9660 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_101
timestamp 1605641404
transform 1 0 10396 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_122
timestamp 1605641404
transform 1 0 12328 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12696 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_3_
timestamp 1605641404
transform 1 0 13708 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_135
timestamp 1605641404
transform 1 0 13524 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1605641404
transform 1 0 14720 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1605641404
transform 1 0 16284 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1605641404
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1605641404
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_146
timestamp 1605641404
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1605641404
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_163
timestamp 1605641404
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_2_
timestamp 1605641404
transform 1 0 17296 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_174
timestamp 1605641404
transform 1 0 17112 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_185
timestamp 1605641404
transform 1 0 18124 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1605641404
transform 1 0 18584 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 19136 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_16_189
timestamp 1605641404
transform 1 0 18492 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1605641404
transform 1 0 18952 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1605641404
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1605641404
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1605641404
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1605641404
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_218
timestamp 1605641404
transform 1 0 21160 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 1564 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1605641404
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1605641404
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1605641404
transform 1 0 4232 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_1_
timestamp 1605641404
transform 1 0 4692 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1605641404
transform 1 0 3220 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_21
timestamp 1605641404
transform 1 0 3036 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_32
timestamp 1605641404
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_37
timestamp 1605641404
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l4_in_0_
timestamp 1605641404
transform 1 0 5704 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1605641404
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_48
timestamp 1605641404
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1605641404
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1605641404
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1605641404
transform 1 0 8004 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1605641404
transform 1 0 6992 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1605641404
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9936 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1605641404
transform 1 0 9108 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_17_84
timestamp 1605641404
transform 1 0 8832 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12420 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1605641404
transform 1 0 11408 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1605641404
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1605641404
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1605641404
transform 1 0 14168 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_17_139
timestamp 1605641404
transform 1 0 13892 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1605641404
transform 1 0 16192 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l4_in_0_
timestamp 1605641404
transform 1 0 15180 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_151
timestamp 1605641404
transform 1 0 14996 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_162
timestamp 1605641404
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1605641404
transform 1 0 17388 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1605641404
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_173
timestamp 1605641404
transform 1 0 17020 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1605641404
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1605641404
transform 1 0 19688 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1605641404
transform 1 0 19504 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_196
timestamp 1605641404
transform 1 0 19136 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1605641404
transform 1 0 20700 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1605641404
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_211
timestamp 1605641404
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_217
timestamp 1605641404
transform 1 0 21068 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1605641404
transform 1 0 1472 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1605641404
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1605641404
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_20
timestamp 1605641404
transform 1 0 2944 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1605641404
transform 1 0 3128 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1605641404
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1605641404
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_26
timestamp 1605641404
transform 1 0 3496 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1605641404
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_41
timestamp 1605641404
transform 1 0 4876 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 5520 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_18_47
timestamp 1605641404
transform 1 0 5428 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 7176 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_64
timestamp 1605641404
transform 1 0 6992 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_82
timestamp 1605641404
transform 1 0 8648 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1605641404
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1605641404
transform 1 0 10672 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1605641404
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1605641404
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1605641404
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1605641404
transform 1 0 11500 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1605641404
transform 1 0 11776 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_125
timestamp 1605641404
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_3_
timestamp 1605641404
transform 1 0 14168 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1605641404
transform 1 0 12972 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1605641404
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_138
timestamp 1605641404
transform 1 0 13800 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 15272 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1605641404
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1605641404
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1605641404
transform 1 0 16836 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 18032 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1605641404
transform 1 0 17204 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_170
timestamp 1605641404
transform 1 0 16744 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1605641404
transform 1 0 19504 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_203
timestamp 1605641404
transform 1 0 19780 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1605641404
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1605641404
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_211
timestamp 1605641404
transform 1 0 20516 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1605641404
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1605641404
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_10
timestamp 1605641404
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1605641404
transform 1 0 1380 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1605641404
transform 1 0 1748 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1605641404
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1605641404
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1605641404
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l5_in_0_
timestamp 1605641404
transform 1 0 1840 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1472 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_17
timestamp 1605641404
transform 1 0 2668 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2208 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1605641404
transform 1 0 3036 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1605641404
transform 1 0 4048 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1605641404
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1605641404
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_30
timestamp 1605641404
transform 1 0 3864 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_41
timestamp 1605641404
transform 1 0 4876 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_28
timestamp 1605641404
transform 1 0 3680 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_41
timestamp 1605641404
transform 1 0 4876 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1605641404
transform 1 0 6072 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1605641404
transform 1 0 6072 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1605641404
transform 1 0 5060 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1605641404
transform 1 0 5060 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1605641404
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_52
timestamp 1605641404
transform 1 0 5888 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_58
timestamp 1605641404
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_62
timestamp 1605641404
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_52
timestamp 1605641404
transform 1 0 5888 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 7544 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1605641404
transform 1 0 7820 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1605641404
transform 1 0 7176 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1605641404
transform 1 0 7084 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_69
timestamp 1605641404
transform 1 0 7452 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_63
timestamp 1605641404
transform 1 0 6900 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_68
timestamp 1605641404
transform 1 0 7360 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_72
timestamp 1605641404
transform 1 0 7728 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_82
timestamp 1605641404
transform 1 0 8648 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_93
timestamp 1605641404
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1605641404
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_86
timestamp 1605641404
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1605641404
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1605641404
transform 1 0 9200 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _135_
timestamp 1605641404
transform 1 0 9016 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_101
timestamp 1605641404
transform 1 0 10396 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_97
timestamp 1605641404
transform 1 0 10028 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1605641404
transform 1 0 10488 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9752 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _132_
timestamp 1605641404
transform 1 0 11776 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 11592 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12512 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1605641404
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_111
timestamp 1605641404
transform 1 0 11316 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_115
timestamp 1605641404
transform 1 0 11684 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1605641404
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_123
timestamp 1605641404
transform 1 0 12420 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_110
timestamp 1605641404
transform 1 0 11224 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1605641404
transform 1 0 13156 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1605641404
transform 1 0 13892 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1605641404
transform 1 0 14168 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1605641404
transform 1 0 13708 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_140
timestamp 1605641404
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_145
timestamp 1605641404
transform 1 0 14444 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_130
timestamp 1605641404
transform 1 0 13064 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_135
timestamp 1605641404
transform 1 0 13524 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 14536 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_2_
timestamp 1605641404
transform 1 0 16192 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_1_
timestamp 1605641404
transform 1 0 15456 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1605641404
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_162
timestamp 1605641404
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_148
timestamp 1605641404
transform 1 0 14720 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1605641404
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_154
timestamp 1605641404
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_165
timestamp 1605641404
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_174
timestamp 1605641404
transform 1 0 17112 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_173
timestamp 1605641404
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1605641404
transform 1 0 16468 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 17204 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1605641404
transform 1 0 17296 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1605641404
transform 1 0 16744 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1605641404
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1605641404
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1605641404
transform 1 0 18124 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 18032 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 19504 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_3_
timestamp 1605641404
transform 1 0 19320 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1605641404
transform 1 0 19136 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1605641404
transform 1 0 18952 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_207
timestamp 1605641404
transform 1 0 20148 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1605641404
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1605641404
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1605641404
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_216
timestamp 1605641404
transform 1 0 20976 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1605641404
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1605641404
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1605641404
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 2852 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_6_
timestamp 1605641404
transform 1 0 1840 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1605641404
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1605641404
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1605641404
transform 1 0 1748 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_17
timestamp 1605641404
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 4508 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_35
timestamp 1605641404
transform 1 0 4324 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1605641404
transform 1 0 6164 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6808 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1605641404
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_53
timestamp 1605641404
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1605641404
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8464 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_78
timestamp 1605641404
transform 1 0 8280 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _133_
timestamp 1605641404
transform 1 0 9844 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 10396 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1605641404
transform 1 0 9476 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_89
timestamp 1605641404
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_94
timestamp 1605641404
transform 1 0 9752 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_99
timestamp 1605641404
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1605641404
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_117
timestamp 1605641404
transform 1 0 11868 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1605641404
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1605641404
transform 1 0 13432 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1605641404
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_143
timestamp 1605641404
transform 1 0 14260 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1605641404
transform 1 0 14720 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15272 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_147
timestamp 1605641404
transform 1 0 14628 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_152
timestamp 1605641404
transform 1 0 15088 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 18032 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16928 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1605641404
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_170
timestamp 1605641404
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1605641404
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1605641404
transform 1 0 19688 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_200
timestamp 1605641404
transform 1 0 19504 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1605641404
transform 1 0 20700 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1605641404
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_211
timestamp 1605641404
transform 1 0 20516 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_217
timestamp 1605641404
transform 1 0 21068 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_5_
timestamp 1605641404
transform 1 0 2208 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1472 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1605641404
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1605641404
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_10
timestamp 1605641404
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 4048 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 3220 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1605641404
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_21
timestamp 1605641404
transform 1 0 3036 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1605641404
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5704 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1605641404
transform 1 0 6716 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_48
timestamp 1605641404
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_59
timestamp 1605641404
transform 1 0 6532 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7912 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_2_
timestamp 1605641404
transform 1 0 6900 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1605641404
transform 1 0 7728 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_83
timestamp 1605641404
transform 1 0 8740 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _134_
timestamp 1605641404
transform 1 0 9016 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_3_
timestamp 1605641404
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1605641404
transform 1 0 10672 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1605641404
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1605641404
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_102
timestamp 1605641404
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1605641404
transform 1 0 11960 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12512 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_113
timestamp 1605641404
transform 1 0 11500 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_117
timestamp 1605641404
transform 1 0 11868 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_122
timestamp 1605641404
transform 1 0 12328 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1605641404
transform 1 0 14168 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_140
timestamp 1605641404
transform 1 0 13984 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 15272 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1605641404
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1605641404
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 17112 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_170
timestamp 1605641404
transform 1 0 16744 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_3_
timestamp 1605641404
transform 1 0 19780 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1605641404
transform 1 0 18584 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1605641404
transform 1 0 19596 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_199
timestamp 1605641404
transform 1 0 19412 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1605641404
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1605641404
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1605641404
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1605641404
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_218
timestamp 1605641404
transform 1 0 21160 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 1472 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_4_
timestamp 1605641404
transform 1 0 2208 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1605641404
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_3
timestamp 1605641404
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_10
timestamp 1605641404
transform 1 0 2024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1605641404
transform 1 0 3220 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1605641404
transform 1 0 3956 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_21
timestamp 1605641404
transform 1 0 3036 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_27
timestamp 1605641404
transform 1 0 3588 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_40
timestamp 1605641404
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1605641404
transform 1 0 6164 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1605641404
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1605641404
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1605641404
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1605641404
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1605641404
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1605641404
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1605641404
transform 1 0 7636 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1605641404
transform 1 0 8648 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_80
timestamp 1605641404
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1605641404
transform 1 0 8832 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1605641404
transform 1 0 9844 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_93
timestamp 1605641404
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_104
timestamp 1605641404
transform 1 0 10672 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1605641404
transform 1 0 11868 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1605641404
transform 1 0 10856 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1605641404
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_115
timestamp 1605641404
transform 1 0 11684 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1605641404
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_123
timestamp 1605641404
transform 1 0 12420 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1605641404
transform 1 0 12788 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 13340 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_131
timestamp 1605641404
transform 1 0 13156 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1605641404
transform 1 0 14996 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 15548 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_149
timestamp 1605641404
transform 1 0 14812 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_155
timestamp 1605641404
transform 1 0 15364 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l4_in_0_
timestamp 1605641404
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 17204 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1605641404
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_173
timestamp 1605641404
transform 1 0 17020 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1605641404
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_2_
timestamp 1605641404
transform 1 0 20056 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_3_
timestamp 1605641404
transform 1 0 19044 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_193
timestamp 1605641404
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_204
timestamp 1605641404
transform 1 0 19872 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1605641404
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1605641404
transform 1 0 20884 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_219
timestamp 1605641404
transform 1 0 21252 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1605641404
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_4_
timestamp 1605641404
transform 1 0 1932 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_6_
timestamp 1605641404
transform 1 0 2944 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1605641404
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1605641404
transform 1 0 1748 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_18
timestamp 1605641404
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_7_
timestamp 1605641404
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1605641404
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1605641404
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_41
timestamp 1605641404
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1605641404
transform 1 0 5060 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 5612 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_47
timestamp 1605641404
transform 1 0 5428 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 7268 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_65
timestamp 1605641404
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_83
timestamp 1605641404
transform 1 0 8740 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _127_
timestamp 1605641404
transform 1 0 9016 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9660 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1605641404
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1605641404
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1605641404
transform 1 0 11316 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1605641404
transform 1 0 11776 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_109
timestamp 1605641404
transform 1 0 11132 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_114
timestamp 1605641404
transform 1 0 11592 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_125
timestamp 1605641404
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12788 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1605641404
transform 1 0 13800 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_136
timestamp 1605641404
transform 1 0 13616 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_1_
timestamp 1605641404
transform 1 0 15548 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1605641404
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1605641404
transform 1 0 14812 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_147
timestamp 1605641404
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1605641404
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_154
timestamp 1605641404
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_166
timestamp 1605641404
transform 1 0 16376 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 16836 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_24_170
timestamp 1605641404
transform 1 0 16744 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_187
timestamp 1605641404
transform 1 0 18308 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1605641404
transform 1 0 18768 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_1_
timestamp 1605641404
transform 1 0 19596 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_24_191
timestamp 1605641404
transform 1 0 18676 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1605641404
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1605641404
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_210
timestamp 1605641404
transform 1 0 20424 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1605641404
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1605641404
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1605641404
transform 1 0 1472 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_5_
timestamp 1605641404
transform 1 0 2024 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1605641404
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1605641404
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_8
timestamp 1605641404
transform 1 0 1840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_19
timestamp 1605641404
transform 1 0 2852 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 3036 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_2_
timestamp 1605641404
transform 1 0 4692 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_37
timestamp 1605641404
transform 1 0 4508 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5704 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1605641404
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_48
timestamp 1605641404
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1605641404
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_62
timestamp 1605641404
transform 1 0 6808 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _130_
timestamp 1605641404
transform 1 0 6900 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 7452 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_67
timestamp 1605641404
transform 1 0 7268 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1605641404
transform 1 0 9384 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9936 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_85
timestamp 1605641404
transform 1 0 8924 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_89
timestamp 1605641404
transform 1 0 9292 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_94
timestamp 1605641404
transform 1 0 9752 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1605641404
transform 1 0 11776 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1605641404
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1605641404
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_112
timestamp 1605641404
transform 1 0 11408 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_120
timestamp 1605641404
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13432 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_132
timestamp 1605641404
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_143
timestamp 1605641404
transform 1 0 14260 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1605641404
transform 1 0 14628 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1605641404
transform 1 0 15640 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_156
timestamp 1605641404
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_3_
timestamp 1605641404
transform 1 0 16652 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1605641404
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_167
timestamp 1605641404
transform 1 0 16468 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_178
timestamp 1605641404
transform 1 0 17480 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1605641404
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_184
timestamp 1605641404
transform 1 0 18032 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l5_in_0_
timestamp 1605641404
transform 1 0 19872 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1605641404
transform 1 0 19044 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1605641404
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_192
timestamp 1605641404
transform 1 0 18768 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1605641404
transform 1 0 20884 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1605641404
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_213
timestamp 1605641404
transform 1 0 20700 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_218
timestamp 1605641404
transform 1 0 21160 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1605641404
transform 1 0 1380 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_7
timestamp 1605641404
transform 1 0 1748 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1605641404
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1605641404
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1605641404
transform 1 0 1472 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 1932 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1605641404
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_13
timestamp 1605641404
transform 1 0 2300 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_18
timestamp 1605641404
transform 1 0 2760 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_1_
timestamp 1605641404
transform 1 0 2944 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 2484 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1605641404
transform 1 0 4140 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_3_
timestamp 1605641404
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1605641404
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1605641404
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_41
timestamp 1605641404
transform 1 0 4876 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_31
timestamp 1605641404
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _128_
timestamp 1605641404
transform 1 0 6164 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1605641404
transform 1 0 6440 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1605641404
transform 1 0 5428 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1605641404
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_56
timestamp 1605641404
transform 1 0 6256 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_49
timestamp 1605641404
transform 1 0 5612 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1605641404
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_62
timestamp 1605641404
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1605641404
transform 1 0 7452 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7912 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1605641404
transform 1 0 7084 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_4_
timestamp 1605641404
transform 1 0 7912 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_67
timestamp 1605641404
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_72
timestamp 1605641404
transform 1 0 7728 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_83
timestamp 1605641404
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_93
timestamp 1605641404
transform 1 0 9660 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1605641404
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1605641404
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1605641404
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1605641404
transform 1 0 9108 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_96
timestamp 1605641404
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_98
timestamp 1605641404
transform 1 0 10120 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1605641404
transform 1 0 10120 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1605641404
transform 1 0 9752 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 10304 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1605641404
transform 1 0 12512 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1605641404
transform 1 0 12052 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_2_
timestamp 1605641404
transform 1 0 11132 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1605641404
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_116
timestamp 1605641404
transform 1 0 11776 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_107
timestamp 1605641404
transform 1 0 10948 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_118
timestamp 1605641404
transform 1 0 11960 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp 1605641404
transform 1 0 12420 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13432 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 14260 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1605641404
transform 1 0 13064 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_26_128
timestamp 1605641404
transform 1 0 12880 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_128
timestamp 1605641404
transform 1 0 12880 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_139
timestamp 1605641404
transform 1 0 13892 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 15272 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 16192 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1605641404
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_150
timestamp 1605641404
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_159
timestamp 1605641404
transform 1 0 15732 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_163
timestamp 1605641404
transform 1 0 16100 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1605641404
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_2_
timestamp 1605641404
transform 1 0 18124 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_2_
timestamp 1605641404
transform 1 0 17112 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1605641404
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1605641404
transform 1 0 16928 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_170
timestamp 1605641404
transform 1 0 16744 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_183
timestamp 1605641404
transform 1 0 17940 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_180
timestamp 1605641404
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1605641404
transform 1 0 19136 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1605641404
transform 1 0 19964 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1605641404
transform 1 0 19872 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1605641404
transform 1 0 18860 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1605641404
transform 1 0 18952 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_202
timestamp 1605641404
transform 1 0 19688 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1605641404
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 20700 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1605641404
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1605641404
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1605641404
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1605641404
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_219
timestamp 1605641404
transform 1 0 21252 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1605641404
transform 1 0 1472 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2024 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1605641404
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 1605641404
transform 1 0 1380 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_8
timestamp 1605641404
transform 1 0 1840 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_16
timestamp 1605641404
transform 1 0 2576 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1605641404
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1605641404
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1605641404
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_41
timestamp 1605641404
transform 1 0 4876 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1605641404
transform 1 0 5060 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5428 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_28_46
timestamp 1605641404
transform 1 0 5336 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1605641404
transform 1 0 8464 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1605641404
transform 1 0 7268 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1605641404
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_63
timestamp 1605641404
transform 1 0 6900 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_76
timestamp 1605641404
transform 1 0 8096 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1605641404
transform 1 0 10672 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1605641404
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1605641404
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_89
timestamp 1605641404
transform 1 0 9292 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_102
timestamp 1605641404
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 11132 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_107
timestamp 1605641404
transform 1 0 10948 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_125
timestamp 1605641404
transform 1 0 12604 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1605641404
transform 1 0 12788 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1605641404
transform 1 0 13984 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1605641404
transform 1 0 13616 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l4_in_0_
timestamp 1605641404
transform 1 0 16284 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1605641404
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_149
timestamp 1605641404
transform 1 0 14812 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_163
timestamp 1605641404
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1605641404
transform 1 0 17296 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1605641404
transform 1 0 18308 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_174
timestamp 1605641404
transform 1 0 17112 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_185
timestamp 1605641404
transform 1 0 18124 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1605641404
transform 1 0 19504 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_196
timestamp 1605641404
transform 1 0 19136 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1605641404
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1605641404
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1605641404
transform 1 0 20332 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1605641404
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1605641404
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1605641404
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1605641404
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1605641404
transform 1 0 2300 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1605641404
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1605641404
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_11
timestamp 1605641404
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_17
timestamp 1605641404
transform 1 0 2668 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1605641404
transform 1 0 3128 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1605641404
transform 1 0 4140 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_29_21
timestamp 1605641404
transform 1 0 3036 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_31
timestamp 1605641404
transform 1 0 3956 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1605641404
transform 1 0 6808 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 6164 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l5_in_0_
timestamp 1605641404
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1605641404
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_42
timestamp 1605641404
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1605641404
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1605641404
transform 1 0 7636 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1605641404
transform 1 0 7452 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_66
timestamp 1605641404
transform 1 0 7176 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_80
timestamp 1605641404
transform 1 0 8464 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1605641404
transform 1 0 9936 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1605641404
transform 1 0 8924 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_29_84
timestamp 1605641404
transform 1 0 8832 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_94
timestamp 1605641404
transform 1 0 9752 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1605641404
transform 1 0 11316 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1605641404
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1605641404
transform 1 0 10764 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1605641404
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13800 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_29_132
timestamp 1605641404
transform 1 0 13248 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1605641404
transform 1 0 14812 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15824 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_147
timestamp 1605641404
transform 1 0 14628 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_158
timestamp 1605641404
transform 1 0 15640 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_4_
timestamp 1605641404
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_5_
timestamp 1605641404
transform 1 0 16836 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1605641404
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1605641404
transform 1 0 16652 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_180
timestamp 1605641404
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1605641404
transform 1 0 19412 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_29_193
timestamp 1605641404
transform 1 0 18860 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_208
timestamp 1605641404
transform 1 0 20240 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 20424 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1605641404
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_216
timestamp 1605641404
transform 1 0 20976 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1605641404
transform 1 0 1564 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 2116 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1605641404
transform 1 0 2944 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1605641404
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1605641404
transform 1 0 1380 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_9
timestamp 1605641404
transform 1 0 1932 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_17
timestamp 1605641404
transform 1 0 2668 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1605641404
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4692 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1605641404
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1605641404
transform 1 0 4416 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1605641404
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_38
timestamp 1605641404
transform 1 0 4600 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 6716 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1605641404
transform 1 0 5704 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_48
timestamp 1605641404
transform 1 0 5520 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_59
timestamp 1605641404
transform 1 0 6532 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8556 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_77
timestamp 1605641404
transform 1 0 8188 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10028 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1605641404
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1605641404
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_93
timestamp 1605641404
transform 1 0 9660 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_1_
timestamp 1605641404
transform 1 0 11684 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_113
timestamp 1605641404
transform 1 0 11500 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_124
timestamp 1605641404
transform 1 0 12512 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 13524 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 12788 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_133
timestamp 1605641404
transform 1 0 13340 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16284 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1605641404
transform 1 0 15272 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1605641404
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_151
timestamp 1605641404
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_163
timestamp 1605641404
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1605641404
transform 1 0 17388 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_30_174
timestamp 1605641404
transform 1 0 17112 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_186
timestamp 1605641404
transform 1 0 18216 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1605641404
transform 1 0 19228 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1605641404
transform 1 0 18400 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1605641404
transform 1 0 19780 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1605641404
transform 1 0 18768 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_196
timestamp 1605641404
transform 1 0 19136 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_201
timestamp 1605641404
transform 1 0 19596 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1605641404
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1605641404
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1605641404
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1605641404
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1605641404
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1605641404
transform 1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1605641404
transform 1 0 2300 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1605641404
transform 1 0 2852 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1605641404
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1605641404
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1605641404
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_17
timestamp 1605641404
transform 1 0 2668 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4692 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1605641404
transform 1 0 3680 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_31_23
timestamp 1605641404
transform 1 0 3220 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_27
timestamp 1605641404
transform 1 0 3588 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_37
timestamp 1605641404
transform 1 0 4508 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 6808 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1605641404
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_55
timestamp 1605641404
transform 1 0 6164 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8464 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_78
timestamp 1605641404
transform 1 0 8280 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _126_
timestamp 1605641404
transform 1 0 10120 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 10672 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_96
timestamp 1605641404
transform 1 0 9936 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_102
timestamp 1605641404
transform 1 0 10488 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 12420 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1605641404
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1605641404
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_3_
timestamp 1605641404
transform 1 0 14076 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1605641404
transform 1 0 13892 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1605641404
transform 1 0 15088 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 16100 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_150
timestamp 1605641404
transform 1 0 14904 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_161
timestamp 1605641404
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1605641404
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 17020 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1605641404
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_169
timestamp 1605641404
transform 1 0 16652 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_179
timestamp 1605641404
transform 1 0 17572 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1605641404
transform 1 0 18400 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1605641404
transform 1 0 19136 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_6_
timestamp 1605641404
transform 1 0 19688 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1605641404
transform 1 0 18952 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_192
timestamp 1605641404
transform 1 0 18768 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_200
timestamp 1605641404
transform 1 0 19504 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1605641404
transform 1 0 20700 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1605641404
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_211
timestamp 1605641404
transform 1 0 20516 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_217
timestamp 1605641404
transform 1 0 21068 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1605641404
transform 1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1605641404
transform 1 0 2300 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _131_
timestamp 1605641404
transform 1 0 2852 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1605641404
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1605641404
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_11
timestamp 1605641404
transform 1 0 2116 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_17
timestamp 1605641404
transform 1 0 2668 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _129_
timestamp 1605641404
transform 1 0 3404 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4416 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1605641404
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_23
timestamp 1605641404
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1605641404
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_32
timestamp 1605641404
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 6072 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1605641404
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_52
timestamp 1605641404
transform 1 0 5888 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_60
timestamp 1605641404
transform 1 0 6624 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1605641404
transform 1 0 6900 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8464 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1605641404
transform 1 0 7452 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_32_67
timestamp 1605641404
transform 1 0 7268 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_78
timestamp 1605641404
transform 1 0 8280 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1605641404
transform 1 0 9752 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1605641404
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_89
timestamp 1605641404
transform 1 0 9292 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_103
timestamp 1605641404
transform 1 0 10580 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1605641404
transform 1 0 12604 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 10764 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1605641404
transform 1 0 11500 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1605641404
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_111
timestamp 1605641404
transform 1 0 11316 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_122
timestamp 1605641404
transform 1 0 12328 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1605641404
transform 1 0 14076 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l4_in_0_
timestamp 1605641404
transform 1 0 13064 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_32_128
timestamp 1605641404
transform 1 0 12880 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_139
timestamp 1605641404
transform 1 0 13892 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1605641404
transform 1 0 15456 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 16008 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1605641404
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_150
timestamp 1605641404
transform 1 0 14904 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_154
timestamp 1605641404
transform 1 0 15272 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_160
timestamp 1605641404
transform 1 0 15824 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1605641404
transform 1 0 17664 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1605641404
transform 1 0 16744 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1605641404
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_168
timestamp 1605641404
transform 1 0 16560 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_176
timestamp 1605641404
transform 1 0 17296 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_184
timestamp 1605641404
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_187
timestamp 1605641404
transform 1 0 18308 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1605641404
transform 1 0 18768 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1605641404
transform 1 0 19320 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_7_
timestamp 1605641404
transform 1 0 19872 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_32_191
timestamp 1605641404
transform 1 0 18676 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_196
timestamp 1605641404
transform 1 0 19136 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_202
timestamp 1605641404
transform 1 0 19688 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1605641404
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1605641404
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_213
timestamp 1605641404
transform 1 0 20700 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1605641404
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_42_
port 0 nsew default input
rlabel metal2 s 570 0 626 480 6 bottom_left_grid_pin_43_
port 1 nsew default input
rlabel metal2 s 1030 0 1086 480 6 bottom_left_grid_pin_44_
port 2 nsew default input
rlabel metal2 s 1490 0 1546 480 6 bottom_left_grid_pin_45_
port 3 nsew default input
rlabel metal2 s 1950 0 2006 480 6 bottom_left_grid_pin_46_
port 4 nsew default input
rlabel metal2 s 2410 0 2466 480 6 bottom_left_grid_pin_47_
port 5 nsew default input
rlabel metal2 s 2870 0 2926 480 6 bottom_left_grid_pin_48_
port 6 nsew default input
rlabel metal2 s 3330 0 3386 480 6 bottom_left_grid_pin_49_
port 7 nsew default input
rlabel metal2 s 4158 0 4214 480 6 ccff_head
port 8 nsew default input
rlabel metal2 s 4618 0 4674 480 6 ccff_tail
port 9 nsew default tristate
rlabel metal3 s 0 3952 480 4072 6 chanx_left_in[0]
port 10 nsew default input
rlabel metal3 s 0 8712 480 8832 6 chanx_left_in[10]
port 11 nsew default input
rlabel metal3 s 0 9120 480 9240 6 chanx_left_in[11]
port 12 nsew default input
rlabel metal3 s 0 9664 480 9784 6 chanx_left_in[12]
port 13 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[13]
port 14 nsew default input
rlabel metal3 s 0 10616 480 10736 6 chanx_left_in[14]
port 15 nsew default input
rlabel metal3 s 0 11024 480 11144 6 chanx_left_in[15]
port 16 nsew default input
rlabel metal3 s 0 11568 480 11688 6 chanx_left_in[16]
port 17 nsew default input
rlabel metal3 s 0 11976 480 12096 6 chanx_left_in[17]
port 18 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[18]
port 19 nsew default input
rlabel metal3 s 0 12928 480 13048 6 chanx_left_in[19]
port 20 nsew default input
rlabel metal3 s 0 4360 480 4480 6 chanx_left_in[1]
port 21 nsew default input
rlabel metal3 s 0 4904 480 5024 6 chanx_left_in[2]
port 22 nsew default input
rlabel metal3 s 0 5312 480 5432 6 chanx_left_in[3]
port 23 nsew default input
rlabel metal3 s 0 5856 480 5976 6 chanx_left_in[4]
port 24 nsew default input
rlabel metal3 s 0 6264 480 6384 6 chanx_left_in[5]
port 25 nsew default input
rlabel metal3 s 0 6808 480 6928 6 chanx_left_in[6]
port 26 nsew default input
rlabel metal3 s 0 7216 480 7336 6 chanx_left_in[7]
port 27 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[8]
port 28 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[9]
port 29 nsew default input
rlabel metal3 s 0 13472 480 13592 6 chanx_left_out[0]
port 30 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chanx_left_out[10]
port 31 nsew default tristate
rlabel metal3 s 0 18640 480 18760 6 chanx_left_out[11]
port 32 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chanx_left_out[12]
port 33 nsew default tristate
rlabel metal3 s 0 19592 480 19712 6 chanx_left_out[13]
port 34 nsew default tristate
rlabel metal3 s 0 20136 480 20256 6 chanx_left_out[14]
port 35 nsew default tristate
rlabel metal3 s 0 20544 480 20664 6 chanx_left_out[15]
port 36 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[16]
port 37 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[17]
port 38 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[18]
port 39 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[19]
port 40 nsew default tristate
rlabel metal3 s 0 13880 480 14000 6 chanx_left_out[1]
port 41 nsew default tristate
rlabel metal3 s 0 14424 480 14544 6 chanx_left_out[2]
port 42 nsew default tristate
rlabel metal3 s 0 14832 480 14952 6 chanx_left_out[3]
port 43 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 chanx_left_out[4]
port 44 nsew default tristate
rlabel metal3 s 0 15784 480 15904 6 chanx_left_out[5]
port 45 nsew default tristate
rlabel metal3 s 0 16328 480 16448 6 chanx_left_out[6]
port 46 nsew default tristate
rlabel metal3 s 0 16736 480 16856 6 chanx_left_out[7]
port 47 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[8]
port 48 nsew default tristate
rlabel metal3 s 0 17688 480 17808 6 chanx_left_out[9]
port 49 nsew default tristate
rlabel metal3 s 22320 3952 22800 4072 6 chanx_right_in[0]
port 50 nsew default input
rlabel metal3 s 22320 8712 22800 8832 6 chanx_right_in[10]
port 51 nsew default input
rlabel metal3 s 22320 9120 22800 9240 6 chanx_right_in[11]
port 52 nsew default input
rlabel metal3 s 22320 9664 22800 9784 6 chanx_right_in[12]
port 53 nsew default input
rlabel metal3 s 22320 10072 22800 10192 6 chanx_right_in[13]
port 54 nsew default input
rlabel metal3 s 22320 10616 22800 10736 6 chanx_right_in[14]
port 55 nsew default input
rlabel metal3 s 22320 11024 22800 11144 6 chanx_right_in[15]
port 56 nsew default input
rlabel metal3 s 22320 11568 22800 11688 6 chanx_right_in[16]
port 57 nsew default input
rlabel metal3 s 22320 11976 22800 12096 6 chanx_right_in[17]
port 58 nsew default input
rlabel metal3 s 22320 12520 22800 12640 6 chanx_right_in[18]
port 59 nsew default input
rlabel metal3 s 22320 12928 22800 13048 6 chanx_right_in[19]
port 60 nsew default input
rlabel metal3 s 22320 4360 22800 4480 6 chanx_right_in[1]
port 61 nsew default input
rlabel metal3 s 22320 4904 22800 5024 6 chanx_right_in[2]
port 62 nsew default input
rlabel metal3 s 22320 5312 22800 5432 6 chanx_right_in[3]
port 63 nsew default input
rlabel metal3 s 22320 5856 22800 5976 6 chanx_right_in[4]
port 64 nsew default input
rlabel metal3 s 22320 6264 22800 6384 6 chanx_right_in[5]
port 65 nsew default input
rlabel metal3 s 22320 6808 22800 6928 6 chanx_right_in[6]
port 66 nsew default input
rlabel metal3 s 22320 7216 22800 7336 6 chanx_right_in[7]
port 67 nsew default input
rlabel metal3 s 22320 7760 22800 7880 6 chanx_right_in[8]
port 68 nsew default input
rlabel metal3 s 22320 8168 22800 8288 6 chanx_right_in[9]
port 69 nsew default input
rlabel metal3 s 22320 13472 22800 13592 6 chanx_right_out[0]
port 70 nsew default tristate
rlabel metal3 s 22320 18232 22800 18352 6 chanx_right_out[10]
port 71 nsew default tristate
rlabel metal3 s 22320 18640 22800 18760 6 chanx_right_out[11]
port 72 nsew default tristate
rlabel metal3 s 22320 19184 22800 19304 6 chanx_right_out[12]
port 73 nsew default tristate
rlabel metal3 s 22320 19592 22800 19712 6 chanx_right_out[13]
port 74 nsew default tristate
rlabel metal3 s 22320 20136 22800 20256 6 chanx_right_out[14]
port 75 nsew default tristate
rlabel metal3 s 22320 20544 22800 20664 6 chanx_right_out[15]
port 76 nsew default tristate
rlabel metal3 s 22320 21088 22800 21208 6 chanx_right_out[16]
port 77 nsew default tristate
rlabel metal3 s 22320 21496 22800 21616 6 chanx_right_out[17]
port 78 nsew default tristate
rlabel metal3 s 22320 22040 22800 22160 6 chanx_right_out[18]
port 79 nsew default tristate
rlabel metal3 s 22320 22448 22800 22568 6 chanx_right_out[19]
port 80 nsew default tristate
rlabel metal3 s 22320 13880 22800 14000 6 chanx_right_out[1]
port 81 nsew default tristate
rlabel metal3 s 22320 14424 22800 14544 6 chanx_right_out[2]
port 82 nsew default tristate
rlabel metal3 s 22320 14832 22800 14952 6 chanx_right_out[3]
port 83 nsew default tristate
rlabel metal3 s 22320 15376 22800 15496 6 chanx_right_out[4]
port 84 nsew default tristate
rlabel metal3 s 22320 15784 22800 15904 6 chanx_right_out[5]
port 85 nsew default tristate
rlabel metal3 s 22320 16328 22800 16448 6 chanx_right_out[6]
port 86 nsew default tristate
rlabel metal3 s 22320 16736 22800 16856 6 chanx_right_out[7]
port 87 nsew default tristate
rlabel metal3 s 22320 17280 22800 17400 6 chanx_right_out[8]
port 88 nsew default tristate
rlabel metal3 s 22320 17688 22800 17808 6 chanx_right_out[9]
port 89 nsew default tristate
rlabel metal2 s 5078 0 5134 480 6 chany_bottom_in[0]
port 90 nsew default input
rlabel metal2 s 9586 0 9642 480 6 chany_bottom_in[10]
port 91 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[11]
port 92 nsew default input
rlabel metal2 s 10414 0 10470 480 6 chany_bottom_in[12]
port 93 nsew default input
rlabel metal2 s 10874 0 10930 480 6 chany_bottom_in[13]
port 94 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[14]
port 95 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_in[15]
port 96 nsew default input
rlabel metal2 s 12254 0 12310 480 6 chany_bottom_in[16]
port 97 nsew default input
rlabel metal2 s 12714 0 12770 480 6 chany_bottom_in[17]
port 98 nsew default input
rlabel metal2 s 13174 0 13230 480 6 chany_bottom_in[18]
port 99 nsew default input
rlabel metal2 s 13542 0 13598 480 6 chany_bottom_in[19]
port 100 nsew default input
rlabel metal2 s 5538 0 5594 480 6 chany_bottom_in[1]
port 101 nsew default input
rlabel metal2 s 5998 0 6054 480 6 chany_bottom_in[2]
port 102 nsew default input
rlabel metal2 s 6458 0 6514 480 6 chany_bottom_in[3]
port 103 nsew default input
rlabel metal2 s 6826 0 6882 480 6 chany_bottom_in[4]
port 104 nsew default input
rlabel metal2 s 7286 0 7342 480 6 chany_bottom_in[5]
port 105 nsew default input
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_in[6]
port 106 nsew default input
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[7]
port 107 nsew default input
rlabel metal2 s 8666 0 8722 480 6 chany_bottom_in[8]
port 108 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[9]
port 109 nsew default input
rlabel metal2 s 14002 0 14058 480 6 chany_bottom_out[0]
port 110 nsew default tristate
rlabel metal2 s 18510 0 18566 480 6 chany_bottom_out[10]
port 111 nsew default tristate
rlabel metal2 s 18970 0 19026 480 6 chany_bottom_out[11]
port 112 nsew default tristate
rlabel metal2 s 19430 0 19486 480 6 chany_bottom_out[12]
port 113 nsew default tristate
rlabel metal2 s 19798 0 19854 480 6 chany_bottom_out[13]
port 114 nsew default tristate
rlabel metal2 s 20258 0 20314 480 6 chany_bottom_out[14]
port 115 nsew default tristate
rlabel metal2 s 20718 0 20774 480 6 chany_bottom_out[15]
port 116 nsew default tristate
rlabel metal2 s 21178 0 21234 480 6 chany_bottom_out[16]
port 117 nsew default tristate
rlabel metal2 s 21638 0 21694 480 6 chany_bottom_out[17]
port 118 nsew default tristate
rlabel metal2 s 22098 0 22154 480 6 chany_bottom_out[18]
port 119 nsew default tristate
rlabel metal2 s 22558 0 22614 480 6 chany_bottom_out[19]
port 120 nsew default tristate
rlabel metal2 s 14462 0 14518 480 6 chany_bottom_out[1]
port 121 nsew default tristate
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_out[2]
port 122 nsew default tristate
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_out[3]
port 123 nsew default tristate
rlabel metal2 s 15842 0 15898 480 6 chany_bottom_out[4]
port 124 nsew default tristate
rlabel metal2 s 16302 0 16358 480 6 chany_bottom_out[5]
port 125 nsew default tristate
rlabel metal2 s 16670 0 16726 480 6 chany_bottom_out[6]
port 126 nsew default tristate
rlabel metal2 s 17130 0 17186 480 6 chany_bottom_out[7]
port 127 nsew default tristate
rlabel metal2 s 17590 0 17646 480 6 chany_bottom_out[8]
port 128 nsew default tristate
rlabel metal2 s 18050 0 18106 480 6 chany_bottom_out[9]
port 129 nsew default tristate
rlabel metal2 s 3974 22320 4030 22800 6 chany_top_in[0]
port 130 nsew default input
rlabel metal2 s 8758 22320 8814 22800 6 chany_top_in[10]
port 131 nsew default input
rlabel metal2 s 9218 22320 9274 22800 6 chany_top_in[11]
port 132 nsew default input
rlabel metal2 s 9678 22320 9734 22800 6 chany_top_in[12]
port 133 nsew default input
rlabel metal2 s 10138 22320 10194 22800 6 chany_top_in[13]
port 134 nsew default input
rlabel metal2 s 10598 22320 10654 22800 6 chany_top_in[14]
port 135 nsew default input
rlabel metal2 s 11058 22320 11114 22800 6 chany_top_in[15]
port 136 nsew default input
rlabel metal2 s 11610 22320 11666 22800 6 chany_top_in[16]
port 137 nsew default input
rlabel metal2 s 12070 22320 12126 22800 6 chany_top_in[17]
port 138 nsew default input
rlabel metal2 s 12530 22320 12586 22800 6 chany_top_in[18]
port 139 nsew default input
rlabel metal2 s 12990 22320 13046 22800 6 chany_top_in[19]
port 140 nsew default input
rlabel metal2 s 4434 22320 4490 22800 6 chany_top_in[1]
port 141 nsew default input
rlabel metal2 s 4894 22320 4950 22800 6 chany_top_in[2]
port 142 nsew default input
rlabel metal2 s 5354 22320 5410 22800 6 chany_top_in[3]
port 143 nsew default input
rlabel metal2 s 5906 22320 5962 22800 6 chany_top_in[4]
port 144 nsew default input
rlabel metal2 s 6366 22320 6422 22800 6 chany_top_in[5]
port 145 nsew default input
rlabel metal2 s 6826 22320 6882 22800 6 chany_top_in[6]
port 146 nsew default input
rlabel metal2 s 7286 22320 7342 22800 6 chany_top_in[7]
port 147 nsew default input
rlabel metal2 s 7746 22320 7802 22800 6 chany_top_in[8]
port 148 nsew default input
rlabel metal2 s 8206 22320 8262 22800 6 chany_top_in[9]
port 149 nsew default input
rlabel metal2 s 13450 22320 13506 22800 6 chany_top_out[0]
port 150 nsew default tristate
rlabel metal2 s 18234 22320 18290 22800 6 chany_top_out[10]
port 151 nsew default tristate
rlabel metal2 s 18694 22320 18750 22800 6 chany_top_out[11]
port 152 nsew default tristate
rlabel metal2 s 19154 22320 19210 22800 6 chany_top_out[12]
port 153 nsew default tristate
rlabel metal2 s 19614 22320 19670 22800 6 chany_top_out[13]
port 154 nsew default tristate
rlabel metal2 s 20166 22320 20222 22800 6 chany_top_out[14]
port 155 nsew default tristate
rlabel metal2 s 20626 22320 20682 22800 6 chany_top_out[15]
port 156 nsew default tristate
rlabel metal2 s 21086 22320 21142 22800 6 chany_top_out[16]
port 157 nsew default tristate
rlabel metal2 s 21546 22320 21602 22800 6 chany_top_out[17]
port 158 nsew default tristate
rlabel metal2 s 22006 22320 22062 22800 6 chany_top_out[18]
port 159 nsew default tristate
rlabel metal2 s 22466 22320 22522 22800 6 chany_top_out[19]
port 160 nsew default tristate
rlabel metal2 s 13910 22320 13966 22800 6 chany_top_out[1]
port 161 nsew default tristate
rlabel metal2 s 14462 22320 14518 22800 6 chany_top_out[2]
port 162 nsew default tristate
rlabel metal2 s 14922 22320 14978 22800 6 chany_top_out[3]
port 163 nsew default tristate
rlabel metal2 s 15382 22320 15438 22800 6 chany_top_out[4]
port 164 nsew default tristate
rlabel metal2 s 15842 22320 15898 22800 6 chany_top_out[5]
port 165 nsew default tristate
rlabel metal2 s 16302 22320 16358 22800 6 chany_top_out[6]
port 166 nsew default tristate
rlabel metal2 s 16762 22320 16818 22800 6 chany_top_out[7]
port 167 nsew default tristate
rlabel metal2 s 17314 22320 17370 22800 6 chany_top_out[8]
port 168 nsew default tristate
rlabel metal2 s 17774 22320 17830 22800 6 chany_top_out[9]
port 169 nsew default tristate
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_34_
port 170 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_35_
port 171 nsew default input
rlabel metal3 s 0 1096 480 1216 6 left_bottom_grid_pin_36_
port 172 nsew default input
rlabel metal3 s 0 1504 480 1624 6 left_bottom_grid_pin_37_
port 173 nsew default input
rlabel metal3 s 0 2048 480 2168 6 left_bottom_grid_pin_38_
port 174 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_39_
port 175 nsew default input
rlabel metal3 s 0 3000 480 3120 6 left_bottom_grid_pin_40_
port 176 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_bottom_grid_pin_41_
port 177 nsew default input
rlabel metal2 s 3698 0 3754 480 6 prog_clk
port 178 nsew default input
rlabel metal3 s 22320 144 22800 264 6 right_bottom_grid_pin_34_
port 179 nsew default input
rlabel metal3 s 22320 552 22800 672 6 right_bottom_grid_pin_35_
port 180 nsew default input
rlabel metal3 s 22320 1096 22800 1216 6 right_bottom_grid_pin_36_
port 181 nsew default input
rlabel metal3 s 22320 1504 22800 1624 6 right_bottom_grid_pin_37_
port 182 nsew default input
rlabel metal3 s 22320 2048 22800 2168 6 right_bottom_grid_pin_38_
port 183 nsew default input
rlabel metal3 s 22320 2456 22800 2576 6 right_bottom_grid_pin_39_
port 184 nsew default input
rlabel metal3 s 22320 3000 22800 3120 6 right_bottom_grid_pin_40_
port 185 nsew default input
rlabel metal3 s 22320 3408 22800 3528 6 right_bottom_grid_pin_41_
port 186 nsew default input
rlabel metal2 s 202 22320 258 22800 6 top_left_grid_pin_42_
port 187 nsew default input
rlabel metal2 s 662 22320 718 22800 6 top_left_grid_pin_43_
port 188 nsew default input
rlabel metal2 s 1122 22320 1178 22800 6 top_left_grid_pin_44_
port 189 nsew default input
rlabel metal2 s 1582 22320 1638 22800 6 top_left_grid_pin_45_
port 190 nsew default input
rlabel metal2 s 2042 22320 2098 22800 6 top_left_grid_pin_46_
port 191 nsew default input
rlabel metal2 s 2502 22320 2558 22800 6 top_left_grid_pin_47_
port 192 nsew default input
rlabel metal2 s 3054 22320 3110 22800 6 top_left_grid_pin_48_
port 193 nsew default input
rlabel metal2 s 3514 22320 3570 22800 6 top_left_grid_pin_49_
port 194 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 195 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 196 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22800
<< end >>
