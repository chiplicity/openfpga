magic
tech sky130A
magscale 1 2
timestamp 1606931724
<< locali >>
rect 2789 16983 2823 17085
rect 9689 9979 9723 10149
rect 9689 6409 9788 6443
rect 9689 6375 9723 6409
rect 9723 6069 9781 6103
rect 12081 5695 12115 5865
rect 12173 5083 12207 5253
rect 12265 4675 12299 4777
rect 4997 3927 5031 4097
rect 9781 2839 9815 3077
rect 14105 2975 14139 3077
rect 17417 2975 17451 3145
<< viali >>
rect 1961 20009 1995 20043
rect 1777 19873 1811 19907
rect 7021 19465 7055 19499
rect 1777 19261 1811 19295
rect 2329 19261 2363 19295
rect 6837 19261 6871 19295
rect 1961 19125 1995 19159
rect 2513 19125 2547 19159
rect 8033 18921 8067 18955
rect 3157 18853 3191 18887
rect 7389 18853 7423 18887
rect 2145 18785 2179 18819
rect 2881 18785 2915 18819
rect 7113 18785 7147 18819
rect 7849 18785 7883 18819
rect 2329 18717 2363 18751
rect 2513 18377 2547 18411
rect 3065 18377 3099 18411
rect 3617 18377 3651 18411
rect 1777 18173 1811 18207
rect 2329 18173 2363 18207
rect 2881 18173 2915 18207
rect 3433 18173 3467 18207
rect 1961 18037 1995 18071
rect 1869 17833 1903 17867
rect 2513 17765 2547 17799
rect 8217 17765 8251 17799
rect 10425 17765 10459 17799
rect 1685 17697 1719 17731
rect 2237 17697 2271 17731
rect 7941 17697 7975 17731
rect 10149 17697 10183 17731
rect 3801 17289 3835 17323
rect 10793 17289 10827 17323
rect 5549 17221 5583 17255
rect 3065 17153 3099 17187
rect 6193 17153 6227 17187
rect 8677 17153 8711 17187
rect 9873 17153 9907 17187
rect 11437 17153 11471 17187
rect 1593 17085 1627 17119
rect 2145 17085 2179 17119
rect 2421 17085 2455 17119
rect 2789 17085 2823 17119
rect 2881 17085 2915 17119
rect 3617 17085 3651 17119
rect 8493 17085 8527 17119
rect 11161 17017 11195 17051
rect 11805 17017 11839 17051
rect 1777 16949 1811 16983
rect 2789 16949 2823 16983
rect 4169 16949 4203 16983
rect 5917 16949 5951 16983
rect 6009 16949 6043 16983
rect 9229 16949 9263 16983
rect 9597 16949 9631 16983
rect 9689 16949 9723 16983
rect 11253 16949 11287 16983
rect 5825 16745 5859 16779
rect 7481 16745 7515 16779
rect 9137 16745 9171 16779
rect 11069 16745 11103 16779
rect 12725 16745 12759 16779
rect 1961 16677 1995 16711
rect 6346 16677 6380 16711
rect 1685 16609 1719 16643
rect 2421 16609 2455 16643
rect 2697 16609 2731 16643
rect 3157 16609 3191 16643
rect 4445 16609 4479 16643
rect 4712 16609 4746 16643
rect 9689 16609 9723 16643
rect 9956 16609 9990 16643
rect 11345 16609 11379 16643
rect 11612 16609 11646 16643
rect 6101 16541 6135 16575
rect 8125 16541 8159 16575
rect 3341 16473 3375 16507
rect 4997 16201 5031 16235
rect 5733 16201 5767 16235
rect 7297 16201 7331 16235
rect 11621 16201 11655 16235
rect 2329 16065 2363 16099
rect 3617 16065 3651 16099
rect 5273 16065 5307 16099
rect 6285 16065 6319 16099
rect 7941 16065 7975 16099
rect 1501 15997 1535 16031
rect 2053 15997 2087 16031
rect 2789 15997 2823 16031
rect 7665 15997 7699 16031
rect 8309 15997 8343 16031
rect 10241 15997 10275 16031
rect 10508 15997 10542 16031
rect 3884 15929 3918 15963
rect 6193 15929 6227 15963
rect 8576 15929 8610 15963
rect 1685 15861 1719 15895
rect 2973 15861 3007 15895
rect 6101 15861 6135 15895
rect 7757 15861 7791 15895
rect 9689 15861 9723 15895
rect 2881 15657 2915 15691
rect 4077 15657 4111 15691
rect 4445 15657 4479 15691
rect 9137 15657 9171 15691
rect 9689 15657 9723 15691
rect 11069 15657 11103 15691
rect 2421 15589 2455 15623
rect 3249 15589 3283 15623
rect 5089 15589 5123 15623
rect 6184 15589 6218 15623
rect 10057 15589 10091 15623
rect 10149 15589 10183 15623
rect 10609 15589 10643 15623
rect 1593 15521 1627 15555
rect 2145 15521 2179 15555
rect 4537 15521 4571 15555
rect 5917 15521 5951 15555
rect 7757 15521 7791 15555
rect 8024 15521 8058 15555
rect 11437 15521 11471 15555
rect 11529 15521 11563 15555
rect 3341 15453 3375 15487
rect 3525 15453 3559 15487
rect 4629 15453 4663 15487
rect 10241 15453 10275 15487
rect 10977 15453 11011 15487
rect 11621 15453 11655 15487
rect 1777 15317 1811 15351
rect 7297 15317 7331 15351
rect 4169 15113 4203 15147
rect 4629 15113 4663 15147
rect 5733 15113 5767 15147
rect 8217 15113 8251 15147
rect 10609 15113 10643 15147
rect 2329 14977 2363 15011
rect 5181 14977 5215 15011
rect 6377 14977 6411 15011
rect 7573 14977 7607 15011
rect 8861 14977 8895 15011
rect 1501 14909 1535 14943
rect 2053 14909 2087 14943
rect 2789 14909 2823 14943
rect 8585 14909 8619 14943
rect 9229 14909 9263 14943
rect 3056 14841 3090 14875
rect 4537 14841 4571 14875
rect 5089 14841 5123 14875
rect 9474 14841 9508 14875
rect 1685 14773 1719 14807
rect 4997 14773 5031 14807
rect 6101 14773 6135 14807
rect 6193 14773 6227 14807
rect 7021 14773 7055 14807
rect 7389 14773 7423 14807
rect 7481 14773 7515 14807
rect 7849 14773 7883 14807
rect 8677 14773 8711 14807
rect 9137 14773 9171 14807
rect 3525 14569 3559 14603
rect 4445 14569 4479 14603
rect 5825 14569 5859 14603
rect 7665 14569 7699 14603
rect 8585 14569 8619 14603
rect 1685 14501 1719 14535
rect 6552 14501 6586 14535
rect 9045 14501 9079 14535
rect 1409 14433 1443 14467
rect 2412 14433 2446 14467
rect 4813 14433 4847 14467
rect 6285 14433 6319 14467
rect 8953 14433 8987 14467
rect 9956 14433 9990 14467
rect 2145 14365 2179 14399
rect 4905 14365 4939 14399
rect 5089 14365 5123 14399
rect 9229 14365 9263 14399
rect 9689 14365 9723 14399
rect 11069 14229 11103 14263
rect 3157 14025 3191 14059
rect 5549 14025 5583 14059
rect 9965 14025 9999 14059
rect 3065 13957 3099 13991
rect 1961 13889 1995 13923
rect 3801 13889 3835 13923
rect 10241 13889 10275 13923
rect 1685 13821 1719 13855
rect 2237 13821 2271 13855
rect 2513 13821 2547 13855
rect 3617 13821 3651 13855
rect 4169 13821 4203 13855
rect 6837 13821 6871 13855
rect 7104 13821 7138 13855
rect 8585 13821 8619 13855
rect 4436 13753 4470 13787
rect 5825 13753 5859 13787
rect 8852 13753 8886 13787
rect 3525 13685 3559 13719
rect 8217 13685 8251 13719
rect 3617 13481 3651 13515
rect 5457 13481 5491 13515
rect 5733 13481 5767 13515
rect 7113 13481 7147 13515
rect 7573 13481 7607 13515
rect 9689 13481 9723 13515
rect 4344 13413 4378 13447
rect 1685 13345 1719 13379
rect 2789 13345 2823 13379
rect 3433 13345 3467 13379
rect 4077 13345 4111 13379
rect 6101 13345 6135 13379
rect 7297 13345 7331 13379
rect 7941 13345 7975 13379
rect 8033 13345 8067 13379
rect 10057 13345 10091 13379
rect 1869 13277 1903 13311
rect 2881 13277 2915 13311
rect 2973 13277 3007 13311
rect 6193 13277 6227 13311
rect 6377 13277 6411 13311
rect 8217 13277 8251 13311
rect 10149 13277 10183 13311
rect 10241 13277 10275 13311
rect 2421 13141 2455 13175
rect 6377 12937 6411 12971
rect 9045 12937 9079 12971
rect 10057 12937 10091 12971
rect 4261 12869 4295 12903
rect 2053 12801 2087 12835
rect 4537 12801 4571 12835
rect 7205 12801 7239 12835
rect 7665 12801 7699 12835
rect 1869 12733 1903 12767
rect 2881 12733 2915 12767
rect 4997 12733 5031 12767
rect 5264 12733 5298 12767
rect 10241 12733 10275 12767
rect 3148 12665 3182 12699
rect 7932 12665 7966 12699
rect 1685 12393 1719 12427
rect 2053 12393 2087 12427
rect 2421 12393 2455 12427
rect 3249 12393 3283 12427
rect 4261 12393 4295 12427
rect 4537 12393 4571 12427
rect 6929 12393 6963 12427
rect 9689 12393 9723 12427
rect 1501 12257 1535 12291
rect 3065 12257 3099 12291
rect 4445 12257 4479 12291
rect 4905 12257 4939 12291
rect 4997 12257 5031 12291
rect 5549 12257 5583 12291
rect 5816 12257 5850 12291
rect 7564 12257 7598 12291
rect 10057 12257 10091 12291
rect 19533 12257 19567 12291
rect 2513 12189 2547 12223
rect 2697 12189 2731 12223
rect 5181 12189 5215 12223
rect 7297 12189 7331 12223
rect 10149 12189 10183 12223
rect 10241 12189 10275 12223
rect 8677 12121 8711 12155
rect 19717 12053 19751 12087
rect 3801 11849 3835 11883
rect 6377 11849 6411 11883
rect 7021 11849 7055 11883
rect 7757 11849 7791 11883
rect 10701 11849 10735 11883
rect 3525 11781 3559 11815
rect 4261 11713 4295 11747
rect 4353 11713 4387 11747
rect 8401 11713 8435 11747
rect 2145 11645 2179 11679
rect 2412 11645 2446 11679
rect 4997 11645 5031 11679
rect 7205 11645 7239 11679
rect 9321 11645 9355 11679
rect 19073 11645 19107 11679
rect 4169 11577 4203 11611
rect 5264 11577 5298 11611
rect 8125 11577 8159 11611
rect 8769 11577 8803 11611
rect 9588 11577 9622 11611
rect 8217 11509 8251 11543
rect 19257 11509 19291 11543
rect 2329 11305 2363 11339
rect 2789 11305 2823 11339
rect 3341 11305 3375 11339
rect 4537 11305 4571 11339
rect 5549 11305 5583 11339
rect 6929 11305 6963 11339
rect 8585 11305 8619 11339
rect 5917 11237 5951 11271
rect 8953 11237 8987 11271
rect 2697 11169 2731 11203
rect 4077 11169 4111 11203
rect 4905 11169 4939 11203
rect 7297 11169 7331 11203
rect 9689 11169 9723 11203
rect 9956 11169 9990 11203
rect 18613 11169 18647 11203
rect 2973 11101 3007 11135
rect 4997 11101 5031 11135
rect 5181 11101 5215 11135
rect 6009 11101 6043 11135
rect 6193 11101 6227 11135
rect 7389 11101 7423 11135
rect 7573 11101 7607 11135
rect 9045 11101 9079 11135
rect 9229 11101 9263 11135
rect 11069 11033 11103 11067
rect 18797 11033 18831 11067
rect 2973 10761 3007 10795
rect 3709 10761 3743 10795
rect 6377 10761 6411 10795
rect 10517 10761 10551 10795
rect 9045 10693 9079 10727
rect 9689 10693 9723 10727
rect 1593 10625 1627 10659
rect 4353 10625 4387 10659
rect 4997 10625 5031 10659
rect 10241 10625 10275 10659
rect 10977 10625 11011 10659
rect 11069 10625 11103 10659
rect 1860 10557 1894 10591
rect 7389 10557 7423 10591
rect 7665 10557 7699 10591
rect 7921 10557 7955 10591
rect 10149 10557 10183 10591
rect 18245 10557 18279 10591
rect 4077 10489 4111 10523
rect 5264 10489 5298 10523
rect 9413 10489 9447 10523
rect 10885 10489 10919 10523
rect 4169 10421 4203 10455
rect 7205 10421 7239 10455
rect 10057 10421 10091 10455
rect 18429 10421 18463 10455
rect 3065 10217 3099 10251
rect 3157 10217 3191 10251
rect 5641 10217 5675 10251
rect 8217 10217 8251 10251
rect 8493 10217 8527 10251
rect 11161 10217 11195 10251
rect 6193 10149 6227 10183
rect 9689 10149 9723 10183
rect 4528 10081 4562 10115
rect 5917 10081 5951 10115
rect 6837 10081 6871 10115
rect 7104 10081 7138 10115
rect 8861 10081 8895 10115
rect 3249 10013 3283 10047
rect 4261 10013 4295 10047
rect 8953 10013 8987 10047
rect 9045 10013 9079 10047
rect 9873 10081 9907 10115
rect 2697 9945 2731 9979
rect 9689 9945 9723 9979
rect 2973 9673 3007 9707
rect 4905 9673 4939 9707
rect 10149 9673 10183 9707
rect 5181 9605 5215 9639
rect 6837 9605 6871 9639
rect 10425 9605 10459 9639
rect 5733 9537 5767 9571
rect 7389 9537 7423 9571
rect 7849 9537 7883 9571
rect 1593 9469 1627 9503
rect 3525 9469 3559 9503
rect 3792 9469 3826 9503
rect 5641 9469 5675 9503
rect 8769 9469 8803 9503
rect 9036 9469 9070 9503
rect 10609 9469 10643 9503
rect 1860 9401 1894 9435
rect 7297 9401 7331 9435
rect 5549 9333 5583 9367
rect 6193 9333 6227 9367
rect 7205 9333 7239 9367
rect 2789 9129 2823 9163
rect 4445 9129 4479 9163
rect 4537 9129 4571 9163
rect 5089 9129 5123 9163
rect 5457 9129 5491 9163
rect 8585 9129 8619 9163
rect 8953 9129 8987 9163
rect 1676 8993 1710 9027
rect 6745 8993 6779 9027
rect 6837 8993 6871 9027
rect 7941 8993 7975 9027
rect 8033 8993 8067 9027
rect 10324 8993 10358 9027
rect 1409 8925 1443 8959
rect 4721 8925 4755 8959
rect 5549 8925 5583 8959
rect 5641 8925 5675 8959
rect 6929 8925 6963 8959
rect 8125 8925 8159 8959
rect 9045 8925 9079 8959
rect 9229 8925 9263 8959
rect 10057 8925 10091 8959
rect 4077 8789 4111 8823
rect 6377 8789 6411 8823
rect 7573 8789 7607 8823
rect 11437 8789 11471 8823
rect 1777 8585 1811 8619
rect 8769 8585 8803 8619
rect 11069 8585 11103 8619
rect 11805 8585 11839 8619
rect 4445 8517 4479 8551
rect 9229 8517 9263 8551
rect 2329 8449 2363 8483
rect 4997 8449 5031 8483
rect 6009 8449 6043 8483
rect 6837 8449 6871 8483
rect 7389 8449 7423 8483
rect 9689 8449 9723 8483
rect 2789 8381 2823 8415
rect 4813 8381 4847 8415
rect 5825 8381 5859 8415
rect 6653 8381 6687 8415
rect 9413 8381 9447 8415
rect 9956 8381 9990 8415
rect 11989 8381 12023 8415
rect 3056 8313 3090 8347
rect 5917 8313 5951 8347
rect 7656 8313 7690 8347
rect 2145 8245 2179 8279
rect 2237 8245 2271 8279
rect 4169 8245 4203 8279
rect 4905 8245 4939 8279
rect 5457 8245 5491 8279
rect 6469 8245 6503 8279
rect 11345 8245 11379 8279
rect 2237 8041 2271 8075
rect 2697 8041 2731 8075
rect 4077 8041 4111 8075
rect 7021 8041 7055 8075
rect 7481 8041 7515 8075
rect 8217 8041 8251 8075
rect 10701 8041 10735 8075
rect 11253 8041 11287 8075
rect 16681 8041 16715 8075
rect 5448 7973 5482 8007
rect 10609 7973 10643 8007
rect 15568 7973 15602 8007
rect 2605 7905 2639 7939
rect 3249 7905 3283 7939
rect 3893 7905 3927 7939
rect 4445 7905 4479 7939
rect 4537 7905 4571 7939
rect 7389 7905 7423 7939
rect 8585 7905 8619 7939
rect 11621 7905 11655 7939
rect 2789 7837 2823 7871
rect 4629 7837 4663 7871
rect 5181 7837 5215 7871
rect 7665 7837 7699 7871
rect 8677 7837 8711 7871
rect 8861 7837 8895 7871
rect 10885 7837 10919 7871
rect 11713 7837 11747 7871
rect 11805 7837 11839 7871
rect 15301 7837 15335 7871
rect 3709 7769 3743 7803
rect 10241 7769 10275 7803
rect 6561 7701 6595 7735
rect 1961 7497 1995 7531
rect 6837 7497 6871 7531
rect 8125 7497 8159 7531
rect 14289 7429 14323 7463
rect 2513 7361 2547 7395
rect 3617 7361 3651 7395
rect 4445 7361 4479 7395
rect 7297 7361 7331 7395
rect 7389 7361 7423 7395
rect 8769 7361 8803 7395
rect 10333 7361 10367 7395
rect 14933 7361 14967 7395
rect 4712 7293 4746 7327
rect 8493 7293 8527 7327
rect 12173 7293 12207 7327
rect 16957 7293 16991 7327
rect 2329 7225 2363 7259
rect 3433 7225 3467 7259
rect 6285 7225 6319 7259
rect 7205 7225 7239 7259
rect 10600 7225 10634 7259
rect 14749 7225 14783 7259
rect 17233 7225 17267 7259
rect 2421 7157 2455 7191
rect 3065 7157 3099 7191
rect 3525 7157 3559 7191
rect 5825 7157 5859 7191
rect 8585 7157 8619 7191
rect 11713 7157 11747 7191
rect 11989 7157 12023 7191
rect 12449 7157 12483 7191
rect 13645 7157 13679 7191
rect 14657 7157 14691 7191
rect 15577 7157 15611 7191
rect 4077 6953 4111 6987
rect 10517 6953 10551 6987
rect 12449 6953 12483 6987
rect 4445 6885 4479 6919
rect 10425 6885 10459 6919
rect 11336 6885 11370 6919
rect 2228 6817 2262 6851
rect 4537 6817 4571 6851
rect 5273 6817 5307 6851
rect 5632 6817 5666 6851
rect 7277 6817 7311 6851
rect 13093 6817 13127 6851
rect 13360 6817 13394 6851
rect 15568 6817 15602 6851
rect 16957 6817 16991 6851
rect 1961 6749 1995 6783
rect 4721 6749 4755 6783
rect 5372 6749 5406 6783
rect 7021 6749 7055 6783
rect 10701 6749 10735 6783
rect 11069 6749 11103 6783
rect 15301 6749 15335 6783
rect 17233 6749 17267 6783
rect 3341 6681 3375 6715
rect 6745 6681 6779 6715
rect 5089 6613 5123 6647
rect 8401 6613 8435 6647
rect 10057 6613 10091 6647
rect 14473 6613 14507 6647
rect 16681 6613 16715 6647
rect 2789 6409 2823 6443
rect 9788 6409 9822 6443
rect 13921 6409 13955 6443
rect 15209 6409 15243 6443
rect 9689 6341 9723 6375
rect 9873 6341 9907 6375
rect 6285 6273 6319 6307
rect 7389 6273 7423 6307
rect 10425 6273 10459 6307
rect 11713 6273 11747 6307
rect 14749 6273 14783 6307
rect 15761 6273 15795 6307
rect 1409 6205 1443 6239
rect 3709 6205 3743 6239
rect 3976 6205 4010 6239
rect 6009 6205 6043 6239
rect 7205 6205 7239 6239
rect 8217 6205 8251 6239
rect 8484 6205 8518 6239
rect 10241 6205 10275 6239
rect 11529 6205 11563 6239
rect 12541 6205 12575 6239
rect 14565 6205 14599 6239
rect 15577 6205 15611 6239
rect 15669 6205 15703 6239
rect 16313 6205 16347 6239
rect 1676 6137 1710 6171
rect 7297 6137 7331 6171
rect 12808 6137 12842 6171
rect 14657 6137 14691 6171
rect 16580 6137 16614 6171
rect 3065 6069 3099 6103
rect 5089 6069 5123 6103
rect 5641 6069 5675 6103
rect 6101 6069 6135 6103
rect 6837 6069 6871 6103
rect 9597 6069 9631 6103
rect 9689 6069 9723 6103
rect 9781 6069 9815 6103
rect 10333 6069 10367 6103
rect 11161 6069 11195 6103
rect 11621 6069 11655 6103
rect 14197 6069 14231 6103
rect 17693 6069 17727 6103
rect 1593 5865 1627 5899
rect 1961 5865 1995 5899
rect 4077 5865 4111 5899
rect 9045 5865 9079 5899
rect 10241 5865 10275 5899
rect 12081 5865 12115 5899
rect 14289 5865 14323 5899
rect 17417 5865 17451 5899
rect 2973 5729 3007 5763
rect 4445 5729 4479 5763
rect 5549 5729 5583 5763
rect 5816 5729 5850 5763
rect 7573 5729 7607 5763
rect 8953 5729 8987 5763
rect 9689 5729 9723 5763
rect 10425 5729 10459 5763
rect 10784 5729 10818 5763
rect 14197 5797 14231 5831
rect 16304 5797 16338 5831
rect 12440 5729 12474 5763
rect 15025 5729 15059 5763
rect 15301 5729 15335 5763
rect 17693 5729 17727 5763
rect 2053 5661 2087 5695
rect 2237 5661 2271 5695
rect 3065 5661 3099 5695
rect 3249 5661 3283 5695
rect 4537 5661 4571 5695
rect 4721 5661 4755 5695
rect 7665 5661 7699 5695
rect 7849 5661 7883 5695
rect 9229 5661 9263 5695
rect 10517 5661 10551 5695
rect 12081 5661 12115 5695
rect 12173 5661 12207 5695
rect 14381 5661 14415 5695
rect 15485 5661 15519 5695
rect 16037 5661 16071 5695
rect 11897 5593 11931 5627
rect 2605 5525 2639 5559
rect 6929 5525 6963 5559
rect 7205 5525 7239 5559
rect 8585 5525 8619 5559
rect 13553 5525 13587 5559
rect 13829 5525 13863 5559
rect 14841 5525 14875 5559
rect 17877 5525 17911 5559
rect 5733 5321 5767 5355
rect 8309 5321 8343 5355
rect 10149 5253 10183 5287
rect 10425 5253 10459 5287
rect 12173 5253 12207 5287
rect 2421 5185 2455 5219
rect 3341 5185 3375 5219
rect 4721 5185 4755 5219
rect 6377 5185 6411 5219
rect 10977 5185 11011 5219
rect 3157 5117 3191 5151
rect 4537 5117 4571 5151
rect 6193 5117 6227 5151
rect 6929 5117 6963 5151
rect 8769 5117 8803 5151
rect 9025 5117 9059 5151
rect 11621 5117 11655 5151
rect 13001 5185 13035 5219
rect 15761 5185 15795 5219
rect 15945 5185 15979 5219
rect 16957 5185 16991 5219
rect 12909 5117 12943 5151
rect 13645 5117 13679 5151
rect 14381 5117 14415 5151
rect 15669 5117 15703 5151
rect 17325 5117 17359 5151
rect 7196 5049 7230 5083
rect 10793 5049 10827 5083
rect 11897 5049 11931 5083
rect 12173 5049 12207 5083
rect 13921 5049 13955 5083
rect 14657 5049 14691 5083
rect 16681 5049 16715 5083
rect 1777 4981 1811 5015
rect 2145 4981 2179 5015
rect 2237 4981 2271 5015
rect 2789 4981 2823 5015
rect 3249 4981 3283 5015
rect 4169 4981 4203 5015
rect 4629 4981 4663 5015
rect 6101 4981 6135 5015
rect 10885 4981 10919 5015
rect 12449 4981 12483 5015
rect 12817 4981 12851 5015
rect 15301 4981 15335 5015
rect 16313 4981 16347 5015
rect 16773 4981 16807 5015
rect 3433 4777 3467 4811
rect 4997 4777 5031 4811
rect 5549 4777 5583 4811
rect 5917 4777 5951 4811
rect 6561 4777 6595 4811
rect 12265 4777 12299 4811
rect 14105 4777 14139 4811
rect 2044 4709 2078 4743
rect 8217 4709 8251 4743
rect 9934 4709 9968 4743
rect 14197 4709 14231 4743
rect 18236 4709 18270 4743
rect 1777 4641 1811 4675
rect 4905 4641 4939 4675
rect 6009 4641 6043 4675
rect 6929 4641 6963 4675
rect 11713 4641 11747 4675
rect 12265 4641 12299 4675
rect 12449 4641 12483 4675
rect 15660 4641 15694 4675
rect 17049 4641 17083 4675
rect 17969 4641 18003 4675
rect 5181 4573 5215 4607
rect 6193 4573 6227 4607
rect 7021 4573 7055 4607
rect 7205 4573 7239 4607
rect 8309 4573 8343 4607
rect 8493 4573 8527 4607
rect 9689 4573 9723 4607
rect 11989 4573 12023 4607
rect 12725 4573 12759 4607
rect 14381 4573 14415 4607
rect 15393 4573 15427 4607
rect 17233 4573 17267 4607
rect 3157 4437 3191 4471
rect 4537 4437 4571 4471
rect 7849 4437 7883 4471
rect 11069 4437 11103 4471
rect 13737 4437 13771 4471
rect 16773 4437 16807 4471
rect 19349 4437 19383 4471
rect 6469 4233 6503 4267
rect 14657 4233 14691 4267
rect 16313 4233 16347 4267
rect 16589 4233 16623 4267
rect 2605 4097 2639 4131
rect 4997 4097 5031 4131
rect 6929 4097 6963 4131
rect 8217 4097 8251 4131
rect 8309 4097 8343 4131
rect 9413 4097 9447 4131
rect 12449 4097 12483 4131
rect 14933 4097 14967 4131
rect 17141 4097 17175 4131
rect 2329 4029 2363 4063
rect 2973 4029 3007 4063
rect 3240 4029 3274 4063
rect 5089 4029 5123 4063
rect 9229 4029 9263 4063
rect 9781 4029 9815 4063
rect 10048 4029 10082 4063
rect 11437 4029 11471 4063
rect 13277 4029 13311 4063
rect 15189 4029 15223 4063
rect 5334 3961 5368 3995
rect 11713 3961 11747 3995
rect 13544 3961 13578 3995
rect 1961 3893 1995 3927
rect 2421 3893 2455 3927
rect 4353 3893 4387 3927
rect 4997 3893 5031 3927
rect 7757 3893 7791 3927
rect 8125 3893 8159 3927
rect 8769 3893 8803 3927
rect 9137 3893 9171 3927
rect 11161 3893 11195 3927
rect 16957 3893 16991 3927
rect 17049 3893 17083 3927
rect 4077 3689 4111 3723
rect 6377 3689 6411 3723
rect 6837 3689 6871 3723
rect 10241 3689 10275 3723
rect 12173 3689 12207 3723
rect 13829 3689 13863 3723
rect 15853 3689 15887 3723
rect 11060 3621 11094 3655
rect 12694 3621 12728 3655
rect 1593 3553 1627 3587
rect 1860 3553 1894 3587
rect 4537 3553 4571 3587
rect 4804 3553 4838 3587
rect 6745 3553 6779 3587
rect 8013 3553 8047 3587
rect 10149 3553 10183 3587
rect 14473 3553 14507 3587
rect 15761 3553 15795 3587
rect 16405 3553 16439 3587
rect 17233 3553 17267 3587
rect 17785 3553 17819 3587
rect 19993 3553 20027 3587
rect 6929 3485 6963 3519
rect 7757 3485 7791 3519
rect 10425 3485 10459 3519
rect 10793 3485 10827 3519
rect 12449 3485 12483 3519
rect 14565 3485 14599 3519
rect 14657 3485 14691 3519
rect 15945 3485 15979 3519
rect 16681 3485 16715 3519
rect 15393 3417 15427 3451
rect 2973 3349 3007 3383
rect 5917 3349 5951 3383
rect 9137 3349 9171 3383
rect 9781 3349 9815 3383
rect 14105 3349 14139 3383
rect 17417 3349 17451 3383
rect 17969 3349 18003 3383
rect 20177 3349 20211 3383
rect 11345 3145 11379 3179
rect 17417 3145 17451 3179
rect 3525 3077 3559 3111
rect 5273 3077 5307 3111
rect 9781 3077 9815 3111
rect 2145 3009 2179 3043
rect 3893 3009 3927 3043
rect 6285 3009 6319 3043
rect 9505 3009 9539 3043
rect 2412 2941 2446 2975
rect 4160 2941 4194 2975
rect 7297 2941 7331 2975
rect 7564 2941 7598 2975
rect 9321 2873 9355 2907
rect 14105 3077 14139 3111
rect 16589 3077 16623 3111
rect 10425 3009 10459 3043
rect 10609 3009 10643 3043
rect 11989 3009 12023 3043
rect 18429 3009 18463 3043
rect 10333 2941 10367 2975
rect 11805 2941 11839 2975
rect 12449 2941 12483 2975
rect 12725 2941 12759 2975
rect 13185 2941 13219 2975
rect 13737 2941 13771 2975
rect 14105 2941 14139 2975
rect 14289 2941 14323 2975
rect 14933 2941 14967 2975
rect 15669 2941 15703 2975
rect 16405 2941 16439 2975
rect 16957 2941 16991 2975
rect 17417 2941 17451 2975
rect 17509 2941 17543 2975
rect 18245 2941 18279 2975
rect 20545 2941 20579 2975
rect 15209 2873 15243 2907
rect 15945 2873 15979 2907
rect 5733 2805 5767 2839
rect 6101 2805 6135 2839
rect 6193 2805 6227 2839
rect 8677 2805 8711 2839
rect 8953 2805 8987 2839
rect 9413 2805 9447 2839
rect 9781 2805 9815 2839
rect 9965 2805 9999 2839
rect 11713 2805 11747 2839
rect 13369 2805 13403 2839
rect 13921 2805 13955 2839
rect 14473 2805 14507 2839
rect 17141 2805 17175 2839
rect 20729 2805 20763 2839
rect 1961 2601 1995 2635
rect 2421 2601 2455 2635
rect 2973 2601 3007 2635
rect 3433 2601 3467 2635
rect 5365 2601 5399 2635
rect 5457 2601 5491 2635
rect 6929 2601 6963 2635
rect 7389 2601 7423 2635
rect 8401 2601 8435 2635
rect 8493 2601 8527 2635
rect 9781 2601 9815 2635
rect 10241 2601 10275 2635
rect 12081 2601 12115 2635
rect 13737 2601 13771 2635
rect 2329 2533 2363 2567
rect 7297 2533 7331 2567
rect 9045 2533 9079 2567
rect 3341 2465 3375 2499
rect 10149 2465 10183 2499
rect 10793 2465 10827 2499
rect 11069 2465 11103 2499
rect 11529 2465 11563 2499
rect 12633 2465 12667 2499
rect 14197 2465 14231 2499
rect 14749 2465 14783 2499
rect 15485 2465 15519 2499
rect 16037 2465 16071 2499
rect 16681 2465 16715 2499
rect 2605 2397 2639 2431
rect 3617 2397 3651 2431
rect 5549 2397 5583 2431
rect 7481 2397 7515 2431
rect 8677 2397 8711 2431
rect 10425 2397 10459 2431
rect 4997 2329 5031 2363
rect 8033 2329 8067 2363
rect 11713 2261 11747 2295
rect 12817 2261 12851 2295
rect 14381 2261 14415 2295
rect 14933 2261 14967 2295
rect 15669 2261 15703 2295
rect 16221 2261 16255 2295
rect 16865 2261 16899 2295
<< metal1 >>
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 1946 20040 1952 20052
rect 1907 20012 1952 20040
rect 1946 20000 1952 20012
rect 2004 20000 2010 20052
rect 1765 19907 1823 19913
rect 1765 19873 1777 19907
rect 1811 19904 1823 19907
rect 2222 19904 2228 19916
rect 1811 19876 2228 19904
rect 1811 19873 1823 19876
rect 1765 19867 1823 19873
rect 2222 19864 2228 19876
rect 2280 19864 2286 19916
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 3694 19456 3700 19508
rect 3752 19496 3758 19508
rect 7009 19499 7067 19505
rect 7009 19496 7021 19499
rect 3752 19468 7021 19496
rect 3752 19456 3758 19468
rect 7009 19465 7021 19468
rect 7055 19465 7067 19499
rect 7009 19459 7067 19465
rect 1765 19295 1823 19301
rect 1765 19261 1777 19295
rect 1811 19292 1823 19295
rect 2038 19292 2044 19304
rect 1811 19264 2044 19292
rect 1811 19261 1823 19264
rect 1765 19255 1823 19261
rect 2038 19252 2044 19264
rect 2096 19252 2102 19304
rect 2314 19292 2320 19304
rect 2275 19264 2320 19292
rect 2314 19252 2320 19264
rect 2372 19252 2378 19304
rect 6822 19292 6828 19304
rect 6783 19264 6828 19292
rect 6822 19252 6828 19264
rect 6880 19252 6886 19304
rect 2866 19224 2872 19236
rect 1964 19196 2872 19224
rect 1964 19165 1992 19196
rect 2866 19184 2872 19196
rect 2924 19184 2930 19236
rect 1949 19159 2007 19165
rect 1949 19125 1961 19159
rect 1995 19125 2007 19159
rect 1949 19119 2007 19125
rect 2501 19159 2559 19165
rect 2501 19125 2513 19159
rect 2547 19156 2559 19159
rect 2774 19156 2780 19168
rect 2547 19128 2780 19156
rect 2547 19125 2559 19128
rect 2501 19119 2559 19125
rect 2774 19116 2780 19128
rect 2832 19116 2838 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 4062 18912 4068 18964
rect 4120 18952 4126 18964
rect 8021 18955 8079 18961
rect 8021 18952 8033 18955
rect 4120 18924 8033 18952
rect 4120 18912 4126 18924
rect 8021 18921 8033 18924
rect 8067 18921 8079 18955
rect 8021 18915 8079 18921
rect 2314 18844 2320 18896
rect 2372 18884 2378 18896
rect 3145 18887 3203 18893
rect 3145 18884 3157 18887
rect 2372 18856 3157 18884
rect 2372 18844 2378 18856
rect 3145 18853 3157 18856
rect 3191 18853 3203 18887
rect 3145 18847 3203 18853
rect 6822 18844 6828 18896
rect 6880 18884 6886 18896
rect 7377 18887 7435 18893
rect 7377 18884 7389 18887
rect 6880 18856 7389 18884
rect 6880 18844 6886 18856
rect 7377 18853 7389 18856
rect 7423 18853 7435 18887
rect 7377 18847 7435 18853
rect 2133 18819 2191 18825
rect 2133 18785 2145 18819
rect 2179 18785 2191 18819
rect 2133 18779 2191 18785
rect 2869 18819 2927 18825
rect 2869 18785 2881 18819
rect 2915 18785 2927 18819
rect 2869 18779 2927 18785
rect 7101 18819 7159 18825
rect 7101 18785 7113 18819
rect 7147 18816 7159 18819
rect 7650 18816 7656 18828
rect 7147 18788 7656 18816
rect 7147 18785 7159 18788
rect 7101 18779 7159 18785
rect 2148 18680 2176 18779
rect 2222 18708 2228 18760
rect 2280 18748 2286 18760
rect 2317 18751 2375 18757
rect 2317 18748 2329 18751
rect 2280 18720 2329 18748
rect 2280 18708 2286 18720
rect 2317 18717 2329 18720
rect 2363 18717 2375 18751
rect 2884 18748 2912 18779
rect 7650 18776 7656 18788
rect 7708 18776 7714 18828
rect 7837 18819 7895 18825
rect 7837 18785 7849 18819
rect 7883 18816 7895 18819
rect 8202 18816 8208 18828
rect 7883 18788 8208 18816
rect 7883 18785 7895 18788
rect 7837 18779 7895 18785
rect 8202 18776 8208 18788
rect 8260 18776 8266 18828
rect 8570 18748 8576 18760
rect 2884 18720 8576 18748
rect 2317 18711 2375 18717
rect 8570 18708 8576 18720
rect 8628 18708 8634 18760
rect 7190 18680 7196 18692
rect 2148 18652 7196 18680
rect 7190 18640 7196 18652
rect 7248 18640 7254 18692
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 2501 18411 2559 18417
rect 2501 18377 2513 18411
rect 2547 18408 2559 18411
rect 2774 18408 2780 18420
rect 2547 18380 2780 18408
rect 2547 18377 2559 18380
rect 2501 18371 2559 18377
rect 2774 18368 2780 18380
rect 2832 18368 2838 18420
rect 3050 18408 3056 18420
rect 3011 18380 3056 18408
rect 3050 18368 3056 18380
rect 3108 18368 3114 18420
rect 3602 18408 3608 18420
rect 3563 18380 3608 18408
rect 3602 18368 3608 18380
rect 3660 18368 3666 18420
rect 1765 18207 1823 18213
rect 1765 18173 1777 18207
rect 1811 18173 1823 18207
rect 2314 18204 2320 18216
rect 2275 18176 2320 18204
rect 1765 18167 1823 18173
rect 1780 18136 1808 18167
rect 2314 18164 2320 18176
rect 2372 18164 2378 18216
rect 2869 18207 2927 18213
rect 2869 18173 2881 18207
rect 2915 18173 2927 18207
rect 2869 18167 2927 18173
rect 3421 18207 3479 18213
rect 3421 18173 3433 18207
rect 3467 18204 3479 18207
rect 8662 18204 8668 18216
rect 3467 18176 8668 18204
rect 3467 18173 3479 18176
rect 3421 18167 3479 18173
rect 2406 18136 2412 18148
rect 1780 18108 2412 18136
rect 2406 18096 2412 18108
rect 2464 18096 2470 18148
rect 2884 18136 2912 18167
rect 8662 18164 8668 18176
rect 8720 18164 8726 18216
rect 10410 18136 10416 18148
rect 2884 18108 10416 18136
rect 10410 18096 10416 18108
rect 10468 18096 10474 18148
rect 1946 18068 1952 18080
rect 1907 18040 1952 18068
rect 1946 18028 1952 18040
rect 2004 18028 2010 18080
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 1854 17864 1860 17876
rect 1815 17836 1860 17864
rect 1854 17824 1860 17836
rect 1912 17824 1918 17876
rect 2314 17756 2320 17808
rect 2372 17796 2378 17808
rect 2501 17799 2559 17805
rect 2501 17796 2513 17799
rect 2372 17768 2513 17796
rect 2372 17756 2378 17768
rect 2501 17765 2513 17768
rect 2547 17765 2559 17799
rect 8202 17796 8208 17808
rect 8163 17768 8208 17796
rect 2501 17759 2559 17765
rect 8202 17756 8208 17768
rect 8260 17756 8266 17808
rect 10410 17796 10416 17808
rect 10371 17768 10416 17796
rect 10410 17756 10416 17768
rect 10468 17756 10474 17808
rect 1673 17731 1731 17737
rect 1673 17697 1685 17731
rect 1719 17697 1731 17731
rect 1673 17691 1731 17697
rect 2225 17731 2283 17737
rect 2225 17697 2237 17731
rect 2271 17728 2283 17731
rect 7006 17728 7012 17740
rect 2271 17700 7012 17728
rect 2271 17697 2283 17700
rect 2225 17691 2283 17697
rect 1688 17660 1716 17691
rect 7006 17688 7012 17700
rect 7064 17688 7070 17740
rect 7929 17731 7987 17737
rect 7929 17697 7941 17731
rect 7975 17697 7987 17731
rect 7929 17691 7987 17697
rect 10137 17731 10195 17737
rect 10137 17697 10149 17731
rect 10183 17728 10195 17731
rect 10778 17728 10784 17740
rect 10183 17700 10784 17728
rect 10183 17697 10195 17700
rect 10137 17691 10195 17697
rect 3050 17660 3056 17672
rect 1688 17632 3056 17660
rect 3050 17620 3056 17632
rect 3108 17620 3114 17672
rect 7944 17660 7972 17691
rect 10778 17688 10784 17700
rect 10836 17688 10842 17740
rect 10410 17660 10416 17672
rect 7944 17632 10416 17660
rect 10410 17620 10416 17632
rect 10468 17620 10474 17672
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 3786 17320 3792 17332
rect 3747 17292 3792 17320
rect 3786 17280 3792 17292
rect 3844 17280 3850 17332
rect 10778 17320 10784 17332
rect 10739 17292 10784 17320
rect 10778 17280 10784 17292
rect 10836 17280 10842 17332
rect 5537 17255 5595 17261
rect 5537 17252 5549 17255
rect 2884 17224 5549 17252
rect 2884 17184 2912 17224
rect 5537 17221 5549 17224
rect 5583 17221 5595 17255
rect 5537 17215 5595 17221
rect 3050 17184 3056 17196
rect 2148 17156 2912 17184
rect 3011 17156 3056 17184
rect 1581 17119 1639 17125
rect 1581 17085 1593 17119
rect 1627 17116 1639 17119
rect 1946 17116 1952 17128
rect 1627 17088 1952 17116
rect 1627 17085 1639 17088
rect 1581 17079 1639 17085
rect 1946 17076 1952 17088
rect 2004 17076 2010 17128
rect 2148 17125 2176 17156
rect 3050 17144 3056 17156
rect 3108 17144 3114 17196
rect 6178 17184 6184 17196
rect 6139 17156 6184 17184
rect 6178 17144 6184 17156
rect 6236 17144 6242 17196
rect 8662 17184 8668 17196
rect 8623 17156 8668 17184
rect 8662 17144 8668 17156
rect 8720 17144 8726 17196
rect 9858 17184 9864 17196
rect 9819 17156 9864 17184
rect 9858 17144 9864 17156
rect 9916 17144 9922 17196
rect 11422 17184 11428 17196
rect 11383 17156 11428 17184
rect 11422 17144 11428 17156
rect 11480 17144 11486 17196
rect 2133 17119 2191 17125
rect 2133 17085 2145 17119
rect 2179 17085 2191 17119
rect 2406 17116 2412 17128
rect 2367 17088 2412 17116
rect 2133 17079 2191 17085
rect 2406 17076 2412 17088
rect 2464 17076 2470 17128
rect 2777 17119 2835 17125
rect 2777 17085 2789 17119
rect 2823 17116 2835 17119
rect 2869 17119 2927 17125
rect 2869 17116 2881 17119
rect 2823 17088 2881 17116
rect 2823 17085 2835 17088
rect 2777 17079 2835 17085
rect 2869 17085 2881 17088
rect 2915 17085 2927 17119
rect 3605 17119 3663 17125
rect 3605 17116 3617 17119
rect 2869 17079 2927 17085
rect 3068 17088 3617 17116
rect 2682 17008 2688 17060
rect 2740 17048 2746 17060
rect 3068 17048 3096 17088
rect 3605 17085 3617 17088
rect 3651 17085 3663 17119
rect 3605 17079 3663 17085
rect 8481 17119 8539 17125
rect 8481 17085 8493 17119
rect 8527 17116 8539 17119
rect 8527 17088 9260 17116
rect 8527 17085 8539 17088
rect 8481 17079 8539 17085
rect 5718 17048 5724 17060
rect 2740 17020 3096 17048
rect 3988 17020 5724 17048
rect 2740 17008 2746 17020
rect 1762 16980 1768 16992
rect 1723 16952 1768 16980
rect 1762 16940 1768 16952
rect 1820 16940 1826 16992
rect 2777 16983 2835 16989
rect 2777 16949 2789 16983
rect 2823 16980 2835 16983
rect 3988 16980 4016 17020
rect 5718 17008 5724 17020
rect 5776 17008 5782 17060
rect 4154 16980 4160 16992
rect 2823 16952 4016 16980
rect 4115 16952 4160 16980
rect 2823 16949 2835 16952
rect 2777 16943 2835 16949
rect 4154 16940 4160 16952
rect 4212 16940 4218 16992
rect 5902 16980 5908 16992
rect 5863 16952 5908 16980
rect 5902 16940 5908 16952
rect 5960 16940 5966 16992
rect 5994 16940 6000 16992
rect 6052 16980 6058 16992
rect 9232 16989 9260 17088
rect 11149 17051 11207 17057
rect 11149 17017 11161 17051
rect 11195 17048 11207 17051
rect 11793 17051 11851 17057
rect 11793 17048 11805 17051
rect 11195 17020 11805 17048
rect 11195 17017 11207 17020
rect 11149 17011 11207 17017
rect 11793 17017 11805 17020
rect 11839 17017 11851 17051
rect 11793 17011 11851 17017
rect 9217 16983 9275 16989
rect 6052 16952 6097 16980
rect 6052 16940 6058 16952
rect 9217 16949 9229 16983
rect 9263 16949 9275 16983
rect 9582 16980 9588 16992
rect 9543 16952 9588 16980
rect 9217 16943 9275 16949
rect 9582 16940 9588 16952
rect 9640 16940 9646 16992
rect 9674 16940 9680 16992
rect 9732 16980 9738 16992
rect 9732 16952 9777 16980
rect 9732 16940 9738 16952
rect 11054 16940 11060 16992
rect 11112 16980 11118 16992
rect 11241 16983 11299 16989
rect 11241 16980 11253 16983
rect 11112 16952 11253 16980
rect 11112 16940 11118 16952
rect 11241 16949 11253 16952
rect 11287 16949 11299 16983
rect 11241 16943 11299 16949
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 5813 16779 5871 16785
rect 1688 16748 5120 16776
rect 1688 16649 1716 16748
rect 1949 16711 2007 16717
rect 1949 16677 1961 16711
rect 1995 16708 2007 16711
rect 2038 16708 2044 16720
rect 1995 16680 2044 16708
rect 1995 16677 2007 16680
rect 1949 16671 2007 16677
rect 2038 16668 2044 16680
rect 2096 16668 2102 16720
rect 4062 16708 4068 16720
rect 2424 16680 4068 16708
rect 2424 16649 2452 16680
rect 4062 16668 4068 16680
rect 4120 16668 4126 16720
rect 1673 16643 1731 16649
rect 1673 16609 1685 16643
rect 1719 16609 1731 16643
rect 1673 16603 1731 16609
rect 2409 16643 2467 16649
rect 2409 16609 2421 16643
rect 2455 16609 2467 16643
rect 2682 16640 2688 16652
rect 2643 16612 2688 16640
rect 2409 16603 2467 16609
rect 2682 16600 2688 16612
rect 2740 16600 2746 16652
rect 3142 16640 3148 16652
rect 3103 16612 3148 16640
rect 3142 16600 3148 16612
rect 3200 16600 3206 16652
rect 3602 16600 3608 16652
rect 3660 16640 3666 16652
rect 4433 16643 4491 16649
rect 4433 16640 4445 16643
rect 3660 16612 4445 16640
rect 3660 16600 3666 16612
rect 4433 16609 4445 16612
rect 4479 16609 4491 16643
rect 4433 16603 4491 16609
rect 4700 16643 4758 16649
rect 4700 16609 4712 16643
rect 4746 16640 4758 16643
rect 4982 16640 4988 16652
rect 4746 16612 4988 16640
rect 4746 16609 4758 16612
rect 4700 16603 4758 16609
rect 4982 16600 4988 16612
rect 5040 16600 5046 16652
rect 5092 16640 5120 16748
rect 5813 16745 5825 16779
rect 5859 16745 5871 16779
rect 5813 16739 5871 16745
rect 5828 16708 5856 16739
rect 6178 16736 6184 16788
rect 6236 16776 6242 16788
rect 7469 16779 7527 16785
rect 7469 16776 7481 16779
rect 6236 16748 7481 16776
rect 6236 16736 6242 16748
rect 7469 16745 7481 16748
rect 7515 16745 7527 16779
rect 7469 16739 7527 16745
rect 9125 16779 9183 16785
rect 9125 16745 9137 16779
rect 9171 16776 9183 16779
rect 9582 16776 9588 16788
rect 9171 16748 9588 16776
rect 9171 16745 9183 16748
rect 9125 16739 9183 16745
rect 9582 16736 9588 16748
rect 9640 16736 9646 16788
rect 9858 16736 9864 16788
rect 9916 16776 9922 16788
rect 10502 16776 10508 16788
rect 9916 16748 10508 16776
rect 9916 16736 9922 16748
rect 10502 16736 10508 16748
rect 10560 16776 10566 16788
rect 11057 16779 11115 16785
rect 11057 16776 11069 16779
rect 10560 16748 11069 16776
rect 10560 16736 10566 16748
rect 11057 16745 11069 16748
rect 11103 16745 11115 16779
rect 11057 16739 11115 16745
rect 11422 16736 11428 16788
rect 11480 16776 11486 16788
rect 12713 16779 12771 16785
rect 12713 16776 12725 16779
rect 11480 16748 12725 16776
rect 11480 16736 11486 16748
rect 12713 16745 12725 16748
rect 12759 16776 12771 16779
rect 17954 16776 17960 16788
rect 12759 16748 17960 16776
rect 12759 16745 12771 16748
rect 12713 16739 12771 16745
rect 17954 16736 17960 16748
rect 18012 16736 18018 16788
rect 6270 16708 6276 16720
rect 5828 16680 6276 16708
rect 6270 16668 6276 16680
rect 6328 16717 6334 16720
rect 6328 16711 6392 16717
rect 6328 16677 6346 16711
rect 6380 16677 6392 16711
rect 6328 16671 6392 16677
rect 9692 16680 10364 16708
rect 6328 16668 6334 16671
rect 7282 16640 7288 16652
rect 5092 16612 7288 16640
rect 7282 16600 7288 16612
rect 7340 16600 7346 16652
rect 9692 16649 9720 16680
rect 10336 16652 10364 16680
rect 9677 16643 9735 16649
rect 9677 16609 9689 16643
rect 9723 16609 9735 16643
rect 9677 16603 9735 16609
rect 9944 16643 10002 16649
rect 9944 16609 9956 16643
rect 9990 16640 10002 16643
rect 10226 16640 10232 16652
rect 9990 16612 10232 16640
rect 9990 16609 10002 16612
rect 9944 16603 10002 16609
rect 10226 16600 10232 16612
rect 10284 16600 10290 16652
rect 10318 16600 10324 16652
rect 10376 16640 10382 16652
rect 11606 16649 11612 16652
rect 11333 16643 11391 16649
rect 11333 16640 11345 16643
rect 10376 16612 11345 16640
rect 10376 16600 10382 16612
rect 11333 16609 11345 16612
rect 11379 16609 11391 16643
rect 11333 16603 11391 16609
rect 11600 16603 11612 16649
rect 11664 16640 11670 16652
rect 11664 16612 11700 16640
rect 11606 16600 11612 16603
rect 11664 16600 11670 16612
rect 6086 16572 6092 16584
rect 6047 16544 6092 16572
rect 6086 16532 6092 16544
rect 6144 16532 6150 16584
rect 8110 16572 8116 16584
rect 8071 16544 8116 16572
rect 8110 16532 8116 16544
rect 8168 16532 8174 16584
rect 3326 16504 3332 16516
rect 3287 16476 3332 16504
rect 3326 16464 3332 16476
rect 3384 16464 3390 16516
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 4982 16232 4988 16244
rect 4943 16204 4988 16232
rect 4982 16192 4988 16204
rect 5040 16192 5046 16244
rect 5721 16235 5779 16241
rect 5721 16201 5733 16235
rect 5767 16232 5779 16235
rect 5994 16232 6000 16244
rect 5767 16204 6000 16232
rect 5767 16201 5779 16204
rect 5721 16195 5779 16201
rect 5994 16192 6000 16204
rect 6052 16192 6058 16244
rect 7282 16232 7288 16244
rect 7243 16204 7288 16232
rect 7282 16192 7288 16204
rect 7340 16192 7346 16244
rect 11606 16232 11612 16244
rect 11567 16204 11612 16232
rect 11606 16192 11612 16204
rect 11664 16192 11670 16244
rect 2866 16124 2872 16176
rect 2924 16164 2930 16176
rect 2924 16136 3648 16164
rect 2924 16124 2930 16136
rect 3620 16108 3648 16136
rect 2317 16099 2375 16105
rect 2317 16065 2329 16099
rect 2363 16096 2375 16099
rect 3142 16096 3148 16108
rect 2363 16068 3148 16096
rect 2363 16065 2375 16068
rect 2317 16059 2375 16065
rect 3142 16056 3148 16068
rect 3200 16056 3206 16108
rect 3602 16096 3608 16108
rect 3563 16068 3608 16096
rect 3602 16056 3608 16068
rect 3660 16056 3666 16108
rect 5261 16099 5319 16105
rect 5261 16065 5273 16099
rect 5307 16096 5319 16099
rect 5902 16096 5908 16108
rect 5307 16068 5908 16096
rect 5307 16065 5319 16068
rect 5261 16059 5319 16065
rect 5902 16056 5908 16068
rect 5960 16056 5966 16108
rect 6270 16096 6276 16108
rect 6231 16068 6276 16096
rect 6270 16056 6276 16068
rect 6328 16056 6334 16108
rect 7929 16099 7987 16105
rect 7929 16065 7941 16099
rect 7975 16096 7987 16099
rect 7975 16068 8432 16096
rect 7975 16065 7987 16068
rect 7929 16059 7987 16065
rect 1486 16028 1492 16040
rect 1447 16000 1492 16028
rect 1486 15988 1492 16000
rect 1544 15988 1550 16040
rect 2041 16031 2099 16037
rect 2041 15997 2053 16031
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 2056 15960 2084 15991
rect 2774 15988 2780 16040
rect 2832 16028 2838 16040
rect 7653 16031 7711 16037
rect 2832 16000 2877 16028
rect 2832 15988 2838 16000
rect 7653 15997 7665 16031
rect 7699 16028 7711 16031
rect 8110 16028 8116 16040
rect 7699 16000 8116 16028
rect 7699 15997 7711 16000
rect 7653 15991 7711 15997
rect 8110 15988 8116 16000
rect 8168 15988 8174 16040
rect 8202 15988 8208 16040
rect 8260 16028 8266 16040
rect 8297 16031 8355 16037
rect 8297 16028 8309 16031
rect 8260 16000 8309 16028
rect 8260 15988 8266 16000
rect 8297 15997 8309 16000
rect 8343 15997 8355 16031
rect 8297 15991 8355 15997
rect 3872 15963 3930 15969
rect 2056 15932 3648 15960
rect 1670 15892 1676 15904
rect 1631 15864 1676 15892
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 2958 15892 2964 15904
rect 2919 15864 2964 15892
rect 2958 15852 2964 15864
rect 3016 15852 3022 15904
rect 3620 15892 3648 15932
rect 3872 15929 3884 15963
rect 3918 15960 3930 15963
rect 4246 15960 4252 15972
rect 3918 15932 4252 15960
rect 3918 15929 3930 15932
rect 3872 15923 3930 15929
rect 4246 15920 4252 15932
rect 4304 15920 4310 15972
rect 6181 15963 6239 15969
rect 6181 15929 6193 15963
rect 6227 15960 6239 15963
rect 6822 15960 6828 15972
rect 6227 15932 6828 15960
rect 6227 15929 6239 15932
rect 6181 15923 6239 15929
rect 6822 15920 6828 15932
rect 6880 15920 6886 15972
rect 8404 15960 8432 16068
rect 10229 16031 10287 16037
rect 10229 15997 10241 16031
rect 10275 16028 10287 16031
rect 10318 16028 10324 16040
rect 10275 16000 10324 16028
rect 10275 15997 10287 16000
rect 10229 15991 10287 15997
rect 10318 15988 10324 16000
rect 10376 15988 10382 16040
rect 10502 16037 10508 16040
rect 10496 16028 10508 16037
rect 10463 16000 10508 16028
rect 10496 15991 10508 16000
rect 10502 15988 10508 15991
rect 10560 15988 10566 16040
rect 8564 15963 8622 15969
rect 8564 15960 8576 15963
rect 8404 15932 8576 15960
rect 8564 15929 8576 15932
rect 8610 15960 8622 15963
rect 9122 15960 9128 15972
rect 8610 15932 9128 15960
rect 8610 15929 8622 15932
rect 8564 15923 8622 15929
rect 9122 15920 9128 15932
rect 9180 15920 9186 15972
rect 4798 15892 4804 15904
rect 3620 15864 4804 15892
rect 4798 15852 4804 15864
rect 4856 15852 4862 15904
rect 6089 15895 6147 15901
rect 6089 15861 6101 15895
rect 6135 15892 6147 15895
rect 6270 15892 6276 15904
rect 6135 15864 6276 15892
rect 6135 15861 6147 15864
rect 6089 15855 6147 15861
rect 6270 15852 6276 15864
rect 6328 15852 6334 15904
rect 7742 15892 7748 15904
rect 7703 15864 7748 15892
rect 7742 15852 7748 15864
rect 7800 15852 7806 15904
rect 9677 15895 9735 15901
rect 9677 15861 9689 15895
rect 9723 15892 9735 15895
rect 10226 15892 10232 15904
rect 9723 15864 10232 15892
rect 9723 15861 9735 15864
rect 9677 15855 9735 15861
rect 10226 15852 10232 15864
rect 10284 15852 10290 15904
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 2869 15691 2927 15697
rect 2869 15657 2881 15691
rect 2915 15657 2927 15691
rect 4062 15688 4068 15700
rect 4023 15660 4068 15688
rect 2869 15651 2927 15657
rect 1946 15580 1952 15632
rect 2004 15620 2010 15632
rect 2409 15623 2467 15629
rect 2409 15620 2421 15623
rect 2004 15592 2421 15620
rect 2004 15580 2010 15592
rect 2409 15589 2421 15592
rect 2455 15589 2467 15623
rect 2409 15583 2467 15589
rect 1581 15555 1639 15561
rect 1581 15521 1593 15555
rect 1627 15521 1639 15555
rect 1581 15515 1639 15521
rect 2133 15555 2191 15561
rect 2133 15521 2145 15555
rect 2179 15552 2191 15555
rect 2884 15552 2912 15651
rect 4062 15648 4068 15660
rect 4120 15648 4126 15700
rect 4154 15648 4160 15700
rect 4212 15688 4218 15700
rect 4433 15691 4491 15697
rect 4433 15688 4445 15691
rect 4212 15660 4445 15688
rect 4212 15648 4218 15660
rect 4433 15657 4445 15660
rect 4479 15657 4491 15691
rect 4433 15651 4491 15657
rect 6270 15648 6276 15700
rect 6328 15688 6334 15700
rect 6546 15688 6552 15700
rect 6328 15660 6552 15688
rect 6328 15648 6334 15660
rect 6546 15648 6552 15660
rect 6604 15688 6610 15700
rect 9122 15688 9128 15700
rect 6604 15660 8340 15688
rect 9083 15660 9128 15688
rect 6604 15648 6610 15660
rect 6178 15629 6184 15632
rect 3237 15623 3295 15629
rect 3237 15589 3249 15623
rect 3283 15620 3295 15623
rect 5077 15623 5135 15629
rect 5077 15620 5089 15623
rect 3283 15592 5089 15620
rect 3283 15589 3295 15592
rect 3237 15583 3295 15589
rect 5077 15589 5089 15592
rect 5123 15589 5135 15623
rect 6172 15620 6184 15629
rect 6139 15592 6184 15620
rect 5077 15583 5135 15589
rect 6172 15583 6184 15592
rect 6178 15580 6184 15583
rect 6236 15580 6242 15632
rect 8202 15620 8208 15632
rect 7760 15592 8208 15620
rect 2179 15524 2912 15552
rect 4525 15555 4583 15561
rect 2179 15521 2191 15524
rect 2133 15515 2191 15521
rect 4525 15521 4537 15555
rect 4571 15552 4583 15555
rect 4706 15552 4712 15564
rect 4571 15524 4712 15552
rect 4571 15521 4583 15524
rect 4525 15515 4583 15521
rect 1596 15484 1624 15515
rect 4706 15512 4712 15524
rect 4764 15512 4770 15564
rect 5905 15555 5963 15561
rect 5905 15521 5917 15555
rect 5951 15552 5963 15555
rect 5994 15552 6000 15564
rect 5951 15524 6000 15552
rect 5951 15521 5963 15524
rect 5905 15515 5963 15521
rect 5994 15512 6000 15524
rect 6052 15552 6058 15564
rect 7760 15561 7788 15592
rect 8202 15580 8208 15592
rect 8260 15580 8266 15632
rect 8312 15620 8340 15660
rect 9122 15648 9128 15660
rect 9180 15648 9186 15700
rect 9674 15688 9680 15700
rect 9635 15660 9680 15688
rect 9674 15648 9680 15660
rect 9732 15648 9738 15700
rect 11054 15688 11060 15700
rect 11015 15660 11060 15688
rect 11054 15648 11060 15660
rect 11112 15648 11118 15700
rect 10045 15623 10103 15629
rect 10045 15620 10057 15623
rect 8312 15592 10057 15620
rect 10045 15589 10057 15592
rect 10091 15589 10103 15623
rect 10045 15583 10103 15589
rect 10137 15623 10195 15629
rect 10137 15589 10149 15623
rect 10183 15620 10195 15623
rect 10597 15623 10655 15629
rect 10597 15620 10609 15623
rect 10183 15592 10609 15620
rect 10183 15589 10195 15592
rect 10137 15583 10195 15589
rect 10597 15589 10609 15592
rect 10643 15620 10655 15623
rect 11698 15620 11704 15632
rect 10643 15592 11704 15620
rect 10643 15589 10655 15592
rect 10597 15583 10655 15589
rect 11698 15580 11704 15592
rect 11756 15580 11762 15632
rect 7745 15555 7803 15561
rect 7745 15552 7757 15555
rect 6052 15524 7757 15552
rect 6052 15512 6058 15524
rect 7745 15521 7757 15524
rect 7791 15521 7803 15555
rect 7745 15515 7803 15521
rect 8012 15555 8070 15561
rect 8012 15521 8024 15555
rect 8058 15552 8070 15555
rect 8846 15552 8852 15564
rect 8058 15524 8852 15552
rect 8058 15521 8070 15524
rect 8012 15515 8070 15521
rect 8846 15512 8852 15524
rect 8904 15512 8910 15564
rect 11054 15512 11060 15564
rect 11112 15552 11118 15564
rect 11425 15555 11483 15561
rect 11425 15552 11437 15555
rect 11112 15524 11437 15552
rect 11112 15512 11118 15524
rect 11425 15521 11437 15524
rect 11471 15521 11483 15555
rect 11425 15515 11483 15521
rect 11517 15555 11575 15561
rect 11517 15521 11529 15555
rect 11563 15552 11575 15555
rect 12066 15552 12072 15564
rect 11563 15524 12072 15552
rect 11563 15521 11575 15524
rect 11517 15515 11575 15521
rect 2498 15484 2504 15496
rect 1596 15456 2504 15484
rect 2498 15444 2504 15456
rect 2556 15444 2562 15496
rect 3326 15484 3332 15496
rect 3287 15456 3332 15484
rect 3326 15444 3332 15456
rect 3384 15444 3390 15496
rect 3510 15484 3516 15496
rect 3471 15456 3516 15484
rect 3510 15444 3516 15456
rect 3568 15444 3574 15496
rect 4617 15487 4675 15493
rect 4617 15453 4629 15487
rect 4663 15484 4675 15487
rect 4982 15484 4988 15496
rect 4663 15456 4988 15484
rect 4663 15453 4675 15456
rect 4617 15447 4675 15453
rect 4982 15444 4988 15456
rect 5040 15444 5046 15496
rect 10226 15444 10232 15496
rect 10284 15484 10290 15496
rect 10965 15487 11023 15493
rect 10284 15456 10329 15484
rect 10284 15444 10290 15456
rect 10965 15453 10977 15487
rect 11011 15484 11023 15487
rect 11532 15484 11560 15515
rect 12066 15512 12072 15524
rect 12124 15512 12130 15564
rect 11011 15456 11560 15484
rect 11011 15453 11023 15456
rect 10965 15447 11023 15453
rect 11606 15444 11612 15496
rect 11664 15484 11670 15496
rect 11664 15456 11709 15484
rect 11664 15444 11670 15456
rect 1762 15348 1768 15360
rect 1723 15320 1768 15348
rect 1762 15308 1768 15320
rect 1820 15308 1826 15360
rect 7285 15351 7343 15357
rect 7285 15317 7297 15351
rect 7331 15348 7343 15351
rect 7558 15348 7564 15360
rect 7331 15320 7564 15348
rect 7331 15317 7343 15320
rect 7285 15311 7343 15317
rect 7558 15308 7564 15320
rect 7616 15308 7622 15360
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 4157 15147 4215 15153
rect 4157 15113 4169 15147
rect 4203 15144 4215 15147
rect 4246 15144 4252 15156
rect 4203 15116 4252 15144
rect 4203 15113 4215 15116
rect 4157 15107 4215 15113
rect 4246 15104 4252 15116
rect 4304 15104 4310 15156
rect 4617 15147 4675 15153
rect 4617 15113 4629 15147
rect 4663 15144 4675 15147
rect 4706 15144 4712 15156
rect 4663 15116 4712 15144
rect 4663 15113 4675 15116
rect 4617 15107 4675 15113
rect 4706 15104 4712 15116
rect 4764 15104 4770 15156
rect 5718 15144 5724 15156
rect 5679 15116 5724 15144
rect 5718 15104 5724 15116
rect 5776 15104 5782 15156
rect 7742 15104 7748 15156
rect 7800 15144 7806 15156
rect 8205 15147 8263 15153
rect 8205 15144 8217 15147
rect 7800 15116 8217 15144
rect 7800 15104 7806 15116
rect 8205 15113 8217 15116
rect 8251 15113 8263 15147
rect 8846 15144 8852 15156
rect 8759 15116 8852 15144
rect 8205 15107 8263 15113
rect 8846 15104 8852 15116
rect 8904 15144 8910 15156
rect 10597 15147 10655 15153
rect 10597 15144 10609 15147
rect 8904 15116 10609 15144
rect 8904 15104 8910 15116
rect 10597 15113 10609 15116
rect 10643 15113 10655 15147
rect 10597 15107 10655 15113
rect 2774 15076 2780 15088
rect 2332 15048 2780 15076
rect 2332 15017 2360 15048
rect 2774 15036 2780 15048
rect 2832 15036 2838 15088
rect 2317 15011 2375 15017
rect 2317 14977 2329 15011
rect 2363 14977 2375 15011
rect 4264 15008 4292 15104
rect 5169 15011 5227 15017
rect 5169 15008 5181 15011
rect 4264 14980 5181 15008
rect 2317 14971 2375 14977
rect 5169 14977 5181 14980
rect 5215 14977 5227 15011
rect 5169 14971 5227 14977
rect 5258 14968 5264 15020
rect 5316 15008 5322 15020
rect 6362 15008 6368 15020
rect 5316 14980 6224 15008
rect 6323 14980 6368 15008
rect 5316 14968 5322 14980
rect 1489 14943 1547 14949
rect 1489 14909 1501 14943
rect 1535 14940 1547 14943
rect 1946 14940 1952 14952
rect 1535 14912 1952 14940
rect 1535 14909 1547 14912
rect 1489 14903 1547 14909
rect 1946 14900 1952 14912
rect 2004 14900 2010 14952
rect 2041 14943 2099 14949
rect 2041 14909 2053 14943
rect 2087 14909 2099 14943
rect 2041 14903 2099 14909
rect 2777 14943 2835 14949
rect 2777 14909 2789 14943
rect 2823 14940 2835 14943
rect 2866 14940 2872 14952
rect 2823 14912 2872 14940
rect 2823 14909 2835 14912
rect 2777 14903 2835 14909
rect 2056 14872 2084 14903
rect 2866 14900 2872 14912
rect 2924 14900 2930 14952
rect 5718 14940 5724 14952
rect 2976 14912 5724 14940
rect 2976 14872 3004 14912
rect 5718 14900 5724 14912
rect 5776 14900 5782 14952
rect 6196 14940 6224 14980
rect 6362 14968 6368 14980
rect 6420 14968 6426 15020
rect 7558 15008 7564 15020
rect 7519 14980 7564 15008
rect 7558 14968 7564 14980
rect 7616 14968 7622 15020
rect 8202 14968 8208 15020
rect 8260 15008 8266 15020
rect 8864 15017 8892 15104
rect 8849 15011 8907 15017
rect 8260 14980 8708 15008
rect 8260 14968 8266 14980
rect 8573 14943 8631 14949
rect 8573 14940 8585 14943
rect 6196 14912 8585 14940
rect 8573 14909 8585 14912
rect 8619 14909 8631 14943
rect 8680 14940 8708 14980
rect 8849 14977 8861 15011
rect 8895 14977 8907 15011
rect 8849 14971 8907 14977
rect 9217 14943 9275 14949
rect 9217 14940 9229 14943
rect 8680 14912 9229 14940
rect 8573 14903 8631 14909
rect 9217 14909 9229 14912
rect 9263 14909 9275 14943
rect 9217 14903 9275 14909
rect 2056 14844 3004 14872
rect 3044 14875 3102 14881
rect 3044 14841 3056 14875
rect 3090 14872 3102 14875
rect 3510 14872 3516 14884
rect 3090 14844 3516 14872
rect 3090 14841 3102 14844
rect 3044 14835 3102 14841
rect 3510 14832 3516 14844
rect 3568 14832 3574 14884
rect 4525 14875 4583 14881
rect 4525 14841 4537 14875
rect 4571 14872 4583 14875
rect 5077 14875 5135 14881
rect 5077 14872 5089 14875
rect 4571 14844 5089 14872
rect 4571 14841 4583 14844
rect 4525 14835 4583 14841
rect 5077 14841 5089 14844
rect 5123 14872 5135 14875
rect 7742 14872 7748 14884
rect 5123 14844 7748 14872
rect 5123 14841 5135 14844
rect 5077 14835 5135 14841
rect 7742 14832 7748 14844
rect 7800 14832 7806 14884
rect 9398 14832 9404 14884
rect 9456 14881 9462 14884
rect 9456 14875 9520 14881
rect 9456 14841 9474 14875
rect 9508 14841 9520 14875
rect 9456 14835 9520 14841
rect 9456 14832 9462 14835
rect 1670 14804 1676 14816
rect 1631 14776 1676 14804
rect 1670 14764 1676 14776
rect 1728 14764 1734 14816
rect 4985 14807 5043 14813
rect 4985 14773 4997 14807
rect 5031 14804 5043 14807
rect 5258 14804 5264 14816
rect 5031 14776 5264 14804
rect 5031 14773 5043 14776
rect 4985 14767 5043 14773
rect 5258 14764 5264 14776
rect 5316 14764 5322 14816
rect 5810 14764 5816 14816
rect 5868 14804 5874 14816
rect 6089 14807 6147 14813
rect 6089 14804 6101 14807
rect 5868 14776 6101 14804
rect 5868 14764 5874 14776
rect 6089 14773 6101 14776
rect 6135 14773 6147 14807
rect 6089 14767 6147 14773
rect 6181 14807 6239 14813
rect 6181 14773 6193 14807
rect 6227 14804 6239 14807
rect 7009 14807 7067 14813
rect 7009 14804 7021 14807
rect 6227 14776 7021 14804
rect 6227 14773 6239 14776
rect 6181 14767 6239 14773
rect 7009 14773 7021 14776
rect 7055 14773 7067 14807
rect 7374 14804 7380 14816
rect 7335 14776 7380 14804
rect 7009 14767 7067 14773
rect 7374 14764 7380 14776
rect 7432 14764 7438 14816
rect 7466 14764 7472 14816
rect 7524 14804 7530 14816
rect 7837 14807 7895 14813
rect 7837 14804 7849 14807
rect 7524 14776 7849 14804
rect 7524 14764 7530 14776
rect 7837 14773 7849 14776
rect 7883 14773 7895 14807
rect 7837 14767 7895 14773
rect 8665 14807 8723 14813
rect 8665 14773 8677 14807
rect 8711 14804 8723 14807
rect 9125 14807 9183 14813
rect 9125 14804 9137 14807
rect 8711 14776 9137 14804
rect 8711 14773 8723 14776
rect 8665 14767 8723 14773
rect 9125 14773 9137 14776
rect 9171 14804 9183 14807
rect 10686 14804 10692 14816
rect 9171 14776 10692 14804
rect 9171 14773 9183 14776
rect 9125 14767 9183 14773
rect 10686 14764 10692 14776
rect 10744 14764 10750 14816
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 3510 14600 3516 14612
rect 3471 14572 3516 14600
rect 3510 14560 3516 14572
rect 3568 14560 3574 14612
rect 4433 14603 4491 14609
rect 4433 14569 4445 14603
rect 4479 14600 4491 14603
rect 4798 14600 4804 14612
rect 4479 14572 4804 14600
rect 4479 14569 4491 14572
rect 4433 14563 4491 14569
rect 4798 14560 4804 14572
rect 4856 14560 4862 14612
rect 5810 14600 5816 14612
rect 5771 14572 5816 14600
rect 5810 14560 5816 14572
rect 5868 14560 5874 14612
rect 6362 14560 6368 14612
rect 6420 14600 6426 14612
rect 7098 14600 7104 14612
rect 6420 14572 7104 14600
rect 6420 14560 6426 14572
rect 7098 14560 7104 14572
rect 7156 14600 7162 14612
rect 7653 14603 7711 14609
rect 7653 14600 7665 14603
rect 7156 14572 7665 14600
rect 7156 14560 7162 14572
rect 7653 14569 7665 14572
rect 7699 14569 7711 14603
rect 8570 14600 8576 14612
rect 8531 14572 8576 14600
rect 7653 14563 7711 14569
rect 8570 14560 8576 14572
rect 8628 14560 8634 14612
rect 11054 14600 11060 14612
rect 8680 14572 11060 14600
rect 1486 14492 1492 14544
rect 1544 14532 1550 14544
rect 1673 14535 1731 14541
rect 1673 14532 1685 14535
rect 1544 14504 1685 14532
rect 1544 14492 1550 14504
rect 1673 14501 1685 14504
rect 1719 14501 1731 14535
rect 4246 14532 4252 14544
rect 1673 14495 1731 14501
rect 2332 14504 4252 14532
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14464 1455 14467
rect 2332 14464 2360 14504
rect 4246 14492 4252 14504
rect 4304 14492 4310 14544
rect 6540 14535 6598 14541
rect 6540 14501 6552 14535
rect 6586 14532 6598 14535
rect 7558 14532 7564 14544
rect 6586 14504 7564 14532
rect 6586 14501 6598 14504
rect 6540 14495 6598 14501
rect 7558 14492 7564 14504
rect 7616 14492 7622 14544
rect 1443 14436 2360 14464
rect 2400 14467 2458 14473
rect 1443 14433 1455 14436
rect 1397 14427 1455 14433
rect 2400 14433 2412 14467
rect 2446 14464 2458 14467
rect 3970 14464 3976 14476
rect 2446 14436 3976 14464
rect 2446 14433 2458 14436
rect 2400 14427 2458 14433
rect 3970 14424 3976 14436
rect 4028 14424 4034 14476
rect 4801 14467 4859 14473
rect 4801 14433 4813 14467
rect 4847 14464 4859 14467
rect 5810 14464 5816 14476
rect 4847 14436 5816 14464
rect 4847 14433 4859 14436
rect 4801 14427 4859 14433
rect 5810 14424 5816 14436
rect 5868 14424 5874 14476
rect 6086 14424 6092 14476
rect 6144 14464 6150 14476
rect 6273 14467 6331 14473
rect 6273 14464 6285 14467
rect 6144 14436 6285 14464
rect 6144 14424 6150 14436
rect 6273 14433 6285 14436
rect 6319 14464 6331 14467
rect 6914 14464 6920 14476
rect 6319 14436 6920 14464
rect 6319 14433 6331 14436
rect 6273 14427 6331 14433
rect 6914 14424 6920 14436
rect 6972 14424 6978 14476
rect 7374 14424 7380 14476
rect 7432 14464 7438 14476
rect 8680 14464 8708 14572
rect 11054 14560 11060 14572
rect 11112 14560 11118 14612
rect 9033 14535 9091 14541
rect 9033 14501 9045 14535
rect 9079 14532 9091 14535
rect 9674 14532 9680 14544
rect 9079 14504 9680 14532
rect 9079 14501 9091 14504
rect 9033 14495 9091 14501
rect 9674 14492 9680 14504
rect 9732 14492 9738 14544
rect 10318 14532 10324 14544
rect 9784 14504 10324 14532
rect 7432 14436 8708 14464
rect 8941 14467 8999 14473
rect 7432 14424 7438 14436
rect 8941 14433 8953 14467
rect 8987 14464 8999 14467
rect 9582 14464 9588 14476
rect 8987 14436 9588 14464
rect 8987 14433 8999 14436
rect 8941 14427 8999 14433
rect 9582 14424 9588 14436
rect 9640 14424 9646 14476
rect 2133 14399 2191 14405
rect 2133 14365 2145 14399
rect 2179 14365 2191 14399
rect 4890 14396 4896 14408
rect 4851 14368 4896 14396
rect 2133 14359 2191 14365
rect 2148 14260 2176 14359
rect 4890 14356 4896 14368
rect 4948 14356 4954 14408
rect 5074 14396 5080 14408
rect 5035 14368 5080 14396
rect 5074 14356 5080 14368
rect 5132 14356 5138 14408
rect 9217 14399 9275 14405
rect 9217 14365 9229 14399
rect 9263 14396 9275 14399
rect 9398 14396 9404 14408
rect 9263 14368 9404 14396
rect 9263 14365 9275 14368
rect 9217 14359 9275 14365
rect 9398 14356 9404 14368
rect 9456 14356 9462 14408
rect 9677 14399 9735 14405
rect 9677 14365 9689 14399
rect 9723 14396 9735 14399
rect 9784 14396 9812 14504
rect 10318 14492 10324 14504
rect 10376 14492 10382 14544
rect 9950 14473 9956 14476
rect 9944 14427 9956 14473
rect 10008 14464 10014 14476
rect 10008 14436 10044 14464
rect 9950 14424 9956 14427
rect 10008 14424 10014 14436
rect 9723 14368 9812 14396
rect 9723 14365 9735 14368
rect 9677 14359 9735 14365
rect 2866 14260 2872 14272
rect 2148 14232 2872 14260
rect 2866 14220 2872 14232
rect 2924 14220 2930 14272
rect 9416 14260 9444 14356
rect 11057 14263 11115 14269
rect 11057 14260 11069 14263
rect 9416 14232 11069 14260
rect 11057 14229 11069 14232
rect 11103 14229 11115 14263
rect 11057 14223 11115 14229
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 3145 14059 3203 14065
rect 3145 14025 3157 14059
rect 3191 14056 3203 14059
rect 3326 14056 3332 14068
rect 3191 14028 3332 14056
rect 3191 14025 3203 14028
rect 3145 14019 3203 14025
rect 3326 14016 3332 14028
rect 3384 14016 3390 14068
rect 3970 14056 3976 14068
rect 3883 14028 3976 14056
rect 3970 14016 3976 14028
rect 4028 14056 4034 14068
rect 5537 14059 5595 14065
rect 5537 14056 5549 14059
rect 4028 14028 5549 14056
rect 4028 14016 4034 14028
rect 5537 14025 5549 14028
rect 5583 14025 5595 14059
rect 9950 14056 9956 14068
rect 9911 14028 9956 14056
rect 5537 14019 5595 14025
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 3053 13991 3111 13997
rect 3053 13957 3065 13991
rect 3099 13988 3111 13991
rect 3099 13960 3648 13988
rect 3099 13957 3111 13960
rect 3053 13951 3111 13957
rect 1949 13923 2007 13929
rect 1949 13889 1961 13923
rect 1995 13920 2007 13923
rect 3418 13920 3424 13932
rect 1995 13892 3424 13920
rect 1995 13889 2007 13892
rect 1949 13883 2007 13889
rect 3418 13880 3424 13892
rect 3476 13880 3482 13932
rect 1673 13855 1731 13861
rect 1673 13821 1685 13855
rect 1719 13852 1731 13855
rect 1762 13852 1768 13864
rect 1719 13824 1768 13852
rect 1719 13821 1731 13824
rect 1673 13815 1731 13821
rect 1762 13812 1768 13824
rect 1820 13812 1826 13864
rect 2225 13855 2283 13861
rect 2225 13821 2237 13855
rect 2271 13852 2283 13855
rect 2498 13852 2504 13864
rect 2271 13824 2360 13852
rect 2459 13824 2504 13852
rect 2271 13821 2283 13824
rect 2225 13815 2283 13821
rect 2332 13784 2360 13824
rect 2498 13812 2504 13824
rect 2556 13812 2562 13864
rect 3326 13852 3332 13864
rect 2608 13824 3332 13852
rect 2608 13784 2636 13824
rect 3326 13812 3332 13824
rect 3384 13812 3390 13864
rect 3620 13861 3648 13960
rect 3789 13923 3847 13929
rect 3789 13889 3801 13923
rect 3835 13920 3847 13923
rect 3988 13920 4016 14016
rect 3835 13892 4016 13920
rect 3835 13889 3847 13892
rect 3789 13883 3847 13889
rect 9582 13880 9588 13932
rect 9640 13920 9646 13932
rect 10229 13923 10287 13929
rect 10229 13920 10241 13923
rect 9640 13892 10241 13920
rect 9640 13880 9646 13892
rect 10229 13889 10241 13892
rect 10275 13889 10287 13923
rect 10229 13883 10287 13889
rect 3605 13855 3663 13861
rect 3605 13821 3617 13855
rect 3651 13852 3663 13855
rect 3694 13852 3700 13864
rect 3651 13824 3700 13852
rect 3651 13821 3663 13824
rect 3605 13815 3663 13821
rect 3694 13812 3700 13824
rect 3752 13812 3758 13864
rect 4157 13855 4215 13861
rect 4157 13821 4169 13855
rect 4203 13821 4215 13855
rect 4157 13815 4215 13821
rect 6825 13855 6883 13861
rect 6825 13821 6837 13855
rect 6871 13852 6883 13855
rect 6914 13852 6920 13864
rect 6871 13824 6920 13852
rect 6871 13821 6883 13824
rect 6825 13815 6883 13821
rect 2332 13756 2636 13784
rect 2866 13744 2872 13796
rect 2924 13784 2930 13796
rect 4062 13784 4068 13796
rect 2924 13756 4068 13784
rect 2924 13744 2930 13756
rect 4062 13744 4068 13756
rect 4120 13784 4126 13796
rect 4172 13784 4200 13815
rect 6914 13812 6920 13824
rect 6972 13812 6978 13864
rect 7098 13861 7104 13864
rect 7092 13852 7104 13861
rect 7059 13824 7104 13852
rect 7092 13815 7104 13824
rect 7098 13812 7104 13815
rect 7156 13812 7162 13864
rect 7558 13852 7564 13864
rect 7300 13824 7564 13852
rect 4120 13756 4200 13784
rect 4424 13787 4482 13793
rect 4120 13744 4126 13756
rect 4424 13753 4436 13787
rect 4470 13784 4482 13787
rect 5074 13784 5080 13796
rect 4470 13756 5080 13784
rect 4470 13753 4482 13756
rect 4424 13747 4482 13753
rect 5074 13744 5080 13756
rect 5132 13744 5138 13796
rect 5810 13784 5816 13796
rect 5771 13756 5816 13784
rect 5810 13744 5816 13756
rect 5868 13744 5874 13796
rect 6932 13784 6960 13812
rect 7300 13784 7328 13824
rect 7558 13812 7564 13824
rect 7616 13852 7622 13864
rect 8573 13855 8631 13861
rect 8573 13852 8585 13855
rect 7616 13824 8585 13852
rect 7616 13812 7622 13824
rect 8573 13821 8585 13824
rect 8619 13821 8631 13855
rect 8573 13815 8631 13821
rect 6932 13756 7328 13784
rect 8840 13787 8898 13793
rect 8840 13753 8852 13787
rect 8886 13784 8898 13787
rect 9030 13784 9036 13796
rect 8886 13756 9036 13784
rect 8886 13753 8898 13756
rect 8840 13747 8898 13753
rect 9030 13744 9036 13756
rect 9088 13744 9094 13796
rect 3513 13719 3571 13725
rect 3513 13685 3525 13719
rect 3559 13716 3571 13719
rect 5350 13716 5356 13728
rect 3559 13688 5356 13716
rect 3559 13685 3571 13688
rect 3513 13679 3571 13685
rect 5350 13676 5356 13688
rect 5408 13676 5414 13728
rect 8202 13716 8208 13728
rect 8163 13688 8208 13716
rect 8202 13676 8208 13688
rect 8260 13676 8266 13728
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 3602 13512 3608 13524
rect 3563 13484 3608 13512
rect 3602 13472 3608 13484
rect 3660 13472 3666 13524
rect 5074 13472 5080 13524
rect 5132 13512 5138 13524
rect 5445 13515 5503 13521
rect 5445 13512 5457 13515
rect 5132 13484 5457 13512
rect 5132 13472 5138 13484
rect 5445 13481 5457 13484
rect 5491 13481 5503 13515
rect 5718 13512 5724 13524
rect 5679 13484 5724 13512
rect 5445 13475 5503 13481
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 6914 13472 6920 13524
rect 6972 13512 6978 13524
rect 7101 13515 7159 13521
rect 7101 13512 7113 13515
rect 6972 13484 7113 13512
rect 6972 13472 6978 13484
rect 7101 13481 7113 13484
rect 7147 13481 7159 13515
rect 7101 13475 7159 13481
rect 7190 13472 7196 13524
rect 7248 13512 7254 13524
rect 7561 13515 7619 13521
rect 7561 13512 7573 13515
rect 7248 13484 7573 13512
rect 7248 13472 7254 13484
rect 7561 13481 7573 13484
rect 7607 13481 7619 13515
rect 9674 13512 9680 13524
rect 9635 13484 9680 13512
rect 7561 13475 7619 13481
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 4332 13447 4390 13453
rect 4332 13413 4344 13447
rect 4378 13444 4390 13447
rect 5166 13444 5172 13456
rect 4378 13416 5172 13444
rect 4378 13413 4390 13416
rect 4332 13407 4390 13413
rect 5166 13404 5172 13416
rect 5224 13404 5230 13456
rect 5350 13404 5356 13456
rect 5408 13444 5414 13456
rect 5408 13416 9352 13444
rect 5408 13404 5414 13416
rect 1670 13376 1676 13388
rect 1631 13348 1676 13376
rect 1670 13336 1676 13348
rect 1728 13336 1734 13388
rect 2774 13336 2780 13388
rect 2832 13376 2838 13388
rect 3418 13376 3424 13388
rect 2832 13348 2877 13376
rect 3379 13348 3424 13376
rect 2832 13336 2838 13348
rect 3418 13336 3424 13348
rect 3476 13336 3482 13388
rect 4062 13376 4068 13388
rect 4023 13348 4068 13376
rect 4062 13336 4068 13348
rect 4120 13336 4126 13388
rect 4798 13336 4804 13388
rect 4856 13376 4862 13388
rect 6089 13379 6147 13385
rect 6089 13376 6101 13379
rect 4856 13348 6101 13376
rect 4856 13336 4862 13348
rect 6089 13345 6101 13348
rect 6135 13345 6147 13379
rect 6089 13339 6147 13345
rect 7098 13336 7104 13388
rect 7156 13376 7162 13388
rect 7285 13379 7343 13385
rect 7285 13376 7297 13379
rect 7156 13348 7297 13376
rect 7156 13336 7162 13348
rect 7285 13345 7297 13348
rect 7331 13345 7343 13379
rect 7285 13339 7343 13345
rect 7929 13379 7987 13385
rect 7929 13345 7941 13379
rect 7975 13345 7987 13379
rect 7929 13339 7987 13345
rect 8021 13379 8079 13385
rect 8021 13345 8033 13379
rect 8067 13376 8079 13379
rect 9214 13376 9220 13388
rect 8067 13348 9220 13376
rect 8067 13345 8079 13348
rect 8021 13339 8079 13345
rect 1486 13268 1492 13320
rect 1544 13308 1550 13320
rect 1857 13311 1915 13317
rect 1857 13308 1869 13311
rect 1544 13280 1869 13308
rect 1544 13268 1550 13280
rect 1857 13277 1869 13280
rect 1903 13277 1915 13311
rect 1857 13271 1915 13277
rect 2869 13311 2927 13317
rect 2869 13277 2881 13311
rect 2915 13277 2927 13311
rect 2869 13271 2927 13277
rect 2884 13240 2912 13271
rect 2958 13268 2964 13320
rect 3016 13308 3022 13320
rect 6178 13308 6184 13320
rect 3016 13280 3061 13308
rect 6139 13280 6184 13308
rect 3016 13268 3022 13280
rect 6178 13268 6184 13280
rect 6236 13268 6242 13320
rect 6362 13308 6368 13320
rect 6323 13280 6368 13308
rect 6362 13268 6368 13280
rect 6420 13268 6426 13320
rect 7190 13268 7196 13320
rect 7248 13308 7254 13320
rect 7944 13308 7972 13339
rect 9214 13336 9220 13348
rect 9272 13336 9278 13388
rect 9324 13376 9352 13416
rect 9950 13404 9956 13456
rect 10008 13444 10014 13456
rect 10008 13416 10272 13444
rect 10008 13404 10014 13416
rect 10045 13379 10103 13385
rect 10045 13376 10057 13379
rect 9324 13348 10057 13376
rect 10045 13345 10057 13348
rect 10091 13345 10103 13379
rect 10045 13339 10103 13345
rect 7248 13280 7972 13308
rect 8205 13311 8263 13317
rect 7248 13268 7254 13280
rect 8205 13277 8217 13311
rect 8251 13308 8263 13311
rect 9030 13308 9036 13320
rect 8251 13280 9036 13308
rect 8251 13277 8263 13280
rect 8205 13271 8263 13277
rect 9030 13268 9036 13280
rect 9088 13268 9094 13320
rect 10244 13317 10272 13416
rect 10137 13311 10195 13317
rect 10137 13308 10149 13311
rect 10060 13280 10149 13308
rect 10060 13252 10088 13280
rect 10137 13277 10149 13280
rect 10183 13277 10195 13311
rect 10137 13271 10195 13277
rect 10229 13311 10287 13317
rect 10229 13277 10241 13311
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 2884 13212 3004 13240
rect 2406 13172 2412 13184
rect 2367 13144 2412 13172
rect 2406 13132 2412 13144
rect 2464 13132 2470 13184
rect 2976 13172 3004 13212
rect 10042 13200 10048 13252
rect 10100 13200 10106 13252
rect 3142 13172 3148 13184
rect 2976 13144 3148 13172
rect 3142 13132 3148 13144
rect 3200 13172 3206 13184
rect 7374 13172 7380 13184
rect 3200 13144 7380 13172
rect 3200 13132 3206 13144
rect 7374 13132 7380 13144
rect 7432 13132 7438 13184
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 5166 12928 5172 12980
rect 5224 12968 5230 12980
rect 6365 12971 6423 12977
rect 6365 12968 6377 12971
rect 5224 12940 6377 12968
rect 5224 12928 5230 12940
rect 6365 12937 6377 12940
rect 6411 12937 6423 12971
rect 9030 12968 9036 12980
rect 8991 12940 9036 12968
rect 6365 12931 6423 12937
rect 9030 12928 9036 12940
rect 9088 12928 9094 12980
rect 10045 12971 10103 12977
rect 10045 12937 10057 12971
rect 10091 12968 10103 12971
rect 10318 12968 10324 12980
rect 10091 12940 10324 12968
rect 10091 12937 10103 12940
rect 10045 12931 10103 12937
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 4249 12903 4307 12909
rect 4249 12869 4261 12903
rect 4295 12900 4307 12903
rect 4706 12900 4712 12912
rect 4295 12872 4712 12900
rect 4295 12869 4307 12872
rect 4249 12863 4307 12869
rect 4706 12860 4712 12872
rect 4764 12860 4770 12912
rect 1946 12792 1952 12844
rect 2004 12832 2010 12844
rect 2041 12835 2099 12841
rect 2041 12832 2053 12835
rect 2004 12804 2053 12832
rect 2004 12792 2010 12804
rect 2041 12801 2053 12804
rect 2087 12801 2099 12835
rect 2041 12795 2099 12801
rect 4525 12835 4583 12841
rect 4525 12801 4537 12835
rect 4571 12832 4583 12835
rect 4798 12832 4804 12844
rect 4571 12804 4804 12832
rect 4571 12801 4583 12804
rect 4525 12795 4583 12801
rect 4798 12792 4804 12804
rect 4856 12792 4862 12844
rect 7190 12832 7196 12844
rect 7151 12804 7196 12832
rect 7190 12792 7196 12804
rect 7248 12792 7254 12844
rect 7558 12792 7564 12844
rect 7616 12832 7622 12844
rect 7653 12835 7711 12841
rect 7653 12832 7665 12835
rect 7616 12804 7665 12832
rect 7616 12792 7622 12804
rect 7653 12801 7665 12804
rect 7699 12801 7711 12835
rect 7653 12795 7711 12801
rect 1854 12764 1860 12776
rect 1815 12736 1860 12764
rect 1854 12724 1860 12736
rect 1912 12724 1918 12776
rect 2682 12724 2688 12776
rect 2740 12764 2746 12776
rect 2866 12764 2872 12776
rect 2740 12736 2872 12764
rect 2740 12724 2746 12736
rect 2866 12724 2872 12736
rect 2924 12724 2930 12776
rect 4982 12764 4988 12776
rect 4943 12736 4988 12764
rect 4982 12724 4988 12736
rect 5040 12724 5046 12776
rect 5252 12767 5310 12773
rect 5252 12733 5264 12767
rect 5298 12764 5310 12767
rect 6362 12764 6368 12776
rect 5298 12736 6368 12764
rect 5298 12733 5310 12736
rect 5252 12727 5310 12733
rect 6362 12724 6368 12736
rect 6420 12724 6426 12776
rect 10229 12767 10287 12773
rect 10229 12733 10241 12767
rect 10275 12764 10287 12767
rect 10410 12764 10416 12776
rect 10275 12736 10416 12764
rect 10275 12733 10287 12736
rect 10229 12727 10287 12733
rect 10410 12724 10416 12736
rect 10468 12724 10474 12776
rect 3136 12699 3194 12705
rect 3136 12665 3148 12699
rect 3182 12696 3194 12699
rect 3510 12696 3516 12708
rect 3182 12668 3516 12696
rect 3182 12665 3194 12668
rect 3136 12659 3194 12665
rect 3510 12656 3516 12668
rect 3568 12656 3574 12708
rect 4798 12656 4804 12708
rect 4856 12696 4862 12708
rect 5350 12696 5356 12708
rect 4856 12668 5356 12696
rect 4856 12656 4862 12668
rect 5350 12656 5356 12668
rect 5408 12656 5414 12708
rect 7920 12699 7978 12705
rect 7920 12665 7932 12699
rect 7966 12696 7978 12699
rect 8662 12696 8668 12708
rect 7966 12668 8668 12696
rect 7966 12665 7978 12668
rect 7920 12659 7978 12665
rect 8662 12656 8668 12668
rect 8720 12656 8726 12708
rect 4154 12588 4160 12640
rect 4212 12628 4218 12640
rect 4982 12628 4988 12640
rect 4212 12600 4988 12628
rect 4212 12588 4218 12600
rect 4982 12588 4988 12600
rect 5040 12588 5046 12640
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 1578 12384 1584 12436
rect 1636 12424 1642 12436
rect 1673 12427 1731 12433
rect 1673 12424 1685 12427
rect 1636 12396 1685 12424
rect 1636 12384 1642 12396
rect 1673 12393 1685 12396
rect 1719 12393 1731 12427
rect 1673 12387 1731 12393
rect 1854 12384 1860 12436
rect 1912 12424 1918 12436
rect 2041 12427 2099 12433
rect 2041 12424 2053 12427
rect 1912 12396 2053 12424
rect 1912 12384 1918 12396
rect 2041 12393 2053 12396
rect 2087 12393 2099 12427
rect 2406 12424 2412 12436
rect 2367 12396 2412 12424
rect 2041 12387 2099 12393
rect 2406 12384 2412 12396
rect 2464 12384 2470 12436
rect 3234 12424 3240 12436
rect 3195 12396 3240 12424
rect 3234 12384 3240 12396
rect 3292 12384 3298 12436
rect 4154 12384 4160 12436
rect 4212 12424 4218 12436
rect 4249 12427 4307 12433
rect 4249 12424 4261 12427
rect 4212 12396 4261 12424
rect 4212 12384 4218 12396
rect 4249 12393 4261 12396
rect 4295 12393 4307 12427
rect 4249 12387 4307 12393
rect 4525 12427 4583 12433
rect 4525 12393 4537 12427
rect 4571 12424 4583 12427
rect 4890 12424 4896 12436
rect 4571 12396 4896 12424
rect 4571 12393 4583 12396
rect 4525 12387 4583 12393
rect 4890 12384 4896 12396
rect 4948 12384 4954 12436
rect 5000 12396 5764 12424
rect 3418 12316 3424 12368
rect 3476 12356 3482 12368
rect 5000 12356 5028 12396
rect 3476 12328 5028 12356
rect 3476 12316 3482 12328
rect 5074 12316 5080 12368
rect 5132 12356 5138 12368
rect 5736 12356 5764 12396
rect 6362 12384 6368 12436
rect 6420 12424 6426 12436
rect 6917 12427 6975 12433
rect 6917 12424 6929 12427
rect 6420 12396 6929 12424
rect 6420 12384 6426 12396
rect 6917 12393 6929 12396
rect 6963 12393 6975 12427
rect 6917 12387 6975 12393
rect 9214 12384 9220 12436
rect 9272 12424 9278 12436
rect 9677 12427 9735 12433
rect 9677 12424 9689 12427
rect 9272 12396 9689 12424
rect 9272 12384 9278 12396
rect 9677 12393 9689 12396
rect 9723 12393 9735 12427
rect 9677 12387 9735 12393
rect 5132 12328 5580 12356
rect 5736 12328 19564 12356
rect 5132 12316 5138 12328
rect 1486 12288 1492 12300
rect 1447 12260 1492 12288
rect 1486 12248 1492 12260
rect 1544 12248 1550 12300
rect 3053 12291 3111 12297
rect 3053 12257 3065 12291
rect 3099 12288 3111 12291
rect 3602 12288 3608 12300
rect 3099 12260 3608 12288
rect 3099 12257 3111 12260
rect 3053 12251 3111 12257
rect 3602 12248 3608 12260
rect 3660 12248 3666 12300
rect 4433 12291 4491 12297
rect 4433 12257 4445 12291
rect 4479 12257 4491 12291
rect 4890 12288 4896 12300
rect 4851 12260 4896 12288
rect 4433 12251 4491 12257
rect 2498 12220 2504 12232
rect 2459 12192 2504 12220
rect 2498 12180 2504 12192
rect 2556 12180 2562 12232
rect 2685 12223 2743 12229
rect 2685 12189 2697 12223
rect 2731 12220 2743 12223
rect 3510 12220 3516 12232
rect 2731 12192 3516 12220
rect 2731 12189 2743 12192
rect 2685 12183 2743 12189
rect 3510 12180 3516 12192
rect 3568 12180 3574 12232
rect 4448 12152 4476 12251
rect 4890 12248 4896 12260
rect 4948 12248 4954 12300
rect 5552 12297 5580 12328
rect 4985 12291 5043 12297
rect 4985 12257 4997 12291
rect 5031 12288 5043 12291
rect 5537 12291 5595 12297
rect 5031 12260 5488 12288
rect 5031 12257 5043 12260
rect 4985 12251 5043 12257
rect 5166 12220 5172 12232
rect 5127 12192 5172 12220
rect 5166 12180 5172 12192
rect 5224 12180 5230 12232
rect 5460 12220 5488 12260
rect 5537 12257 5549 12291
rect 5583 12257 5595 12291
rect 5537 12251 5595 12257
rect 5626 12248 5632 12300
rect 5684 12248 5690 12300
rect 5804 12291 5862 12297
rect 5804 12257 5816 12291
rect 5850 12288 5862 12291
rect 6362 12288 6368 12300
rect 5850 12260 6368 12288
rect 5850 12257 5862 12260
rect 5804 12251 5862 12257
rect 6362 12248 6368 12260
rect 6420 12248 6426 12300
rect 6822 12248 6828 12300
rect 6880 12288 6886 12300
rect 7374 12288 7380 12300
rect 6880 12260 7380 12288
rect 6880 12248 6886 12260
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 7552 12291 7610 12297
rect 7552 12257 7564 12291
rect 7598 12288 7610 12291
rect 8386 12288 8392 12300
rect 7598 12260 8392 12288
rect 7598 12257 7610 12260
rect 7552 12251 7610 12257
rect 8386 12248 8392 12260
rect 8444 12248 8450 12300
rect 8478 12248 8484 12300
rect 8536 12288 8542 12300
rect 19536 12297 19564 12328
rect 10045 12291 10103 12297
rect 10045 12288 10057 12291
rect 8536 12260 10057 12288
rect 8536 12248 8542 12260
rect 10045 12257 10057 12260
rect 10091 12257 10103 12291
rect 10045 12251 10103 12257
rect 19521 12291 19579 12297
rect 19521 12257 19533 12291
rect 19567 12257 19579 12291
rect 19521 12251 19579 12257
rect 5644 12220 5672 12248
rect 5460 12192 5672 12220
rect 6914 12180 6920 12232
rect 6972 12220 6978 12232
rect 7285 12223 7343 12229
rect 7285 12220 7297 12223
rect 6972 12192 7297 12220
rect 6972 12180 6978 12192
rect 7285 12189 7297 12192
rect 7331 12189 7343 12223
rect 7285 12183 7343 12189
rect 9950 12180 9956 12232
rect 10008 12220 10014 12232
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 10008 12192 10149 12220
rect 10008 12180 10014 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 8662 12152 8668 12164
rect 4448 12124 5028 12152
rect 8575 12124 8668 12152
rect 2866 12044 2872 12096
rect 2924 12084 2930 12096
rect 4890 12084 4896 12096
rect 2924 12056 4896 12084
rect 2924 12044 2930 12056
rect 4890 12044 4896 12056
rect 4948 12044 4954 12096
rect 5000 12084 5028 12124
rect 8662 12112 8668 12124
rect 8720 12152 8726 12164
rect 10244 12152 10272 12183
rect 8720 12124 10272 12152
rect 8720 12112 8726 12124
rect 7098 12084 7104 12096
rect 5000 12056 7104 12084
rect 7098 12044 7104 12056
rect 7156 12044 7162 12096
rect 19705 12087 19763 12093
rect 19705 12053 19717 12087
rect 19751 12084 19763 12087
rect 20346 12084 20352 12096
rect 19751 12056 20352 12084
rect 19751 12053 19763 12056
rect 19705 12047 19763 12053
rect 20346 12044 20352 12056
rect 20404 12044 20410 12096
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 2498 11840 2504 11892
rect 2556 11880 2562 11892
rect 3789 11883 3847 11889
rect 3789 11880 3801 11883
rect 2556 11852 3801 11880
rect 2556 11840 2562 11852
rect 3789 11849 3801 11852
rect 3835 11849 3847 11883
rect 3789 11843 3847 11849
rect 4062 11840 4068 11892
rect 4120 11880 4126 11892
rect 6362 11880 6368 11892
rect 4120 11852 5948 11880
rect 6323 11852 6368 11880
rect 4120 11840 4126 11852
rect 3510 11812 3516 11824
rect 3471 11784 3516 11812
rect 3510 11772 3516 11784
rect 3568 11772 3574 11824
rect 5920 11812 5948 11852
rect 6362 11840 6368 11852
rect 6420 11840 6426 11892
rect 7009 11883 7067 11889
rect 7009 11849 7021 11883
rect 7055 11880 7067 11883
rect 7098 11880 7104 11892
rect 7055 11852 7104 11880
rect 7055 11849 7067 11852
rect 7009 11843 7067 11849
rect 7098 11840 7104 11852
rect 7156 11840 7162 11892
rect 7650 11840 7656 11892
rect 7708 11880 7714 11892
rect 7745 11883 7803 11889
rect 7745 11880 7757 11883
rect 7708 11852 7757 11880
rect 7708 11840 7714 11852
rect 7745 11849 7757 11852
rect 7791 11849 7803 11883
rect 10689 11883 10747 11889
rect 10689 11880 10701 11883
rect 7745 11843 7803 11849
rect 8864 11852 10701 11880
rect 5920 11784 7328 11812
rect 3418 11704 3424 11756
rect 3476 11744 3482 11756
rect 4249 11747 4307 11753
rect 4249 11744 4261 11747
rect 3476 11716 4261 11744
rect 3476 11704 3482 11716
rect 4249 11713 4261 11716
rect 4295 11713 4307 11747
rect 4249 11707 4307 11713
rect 4341 11747 4399 11753
rect 4341 11713 4353 11747
rect 4387 11713 4399 11747
rect 4341 11707 4399 11713
rect 1578 11636 1584 11688
rect 1636 11676 1642 11688
rect 2133 11679 2191 11685
rect 2133 11676 2145 11679
rect 1636 11648 2145 11676
rect 1636 11636 1642 11648
rect 2133 11645 2145 11648
rect 2179 11645 2191 11679
rect 2133 11639 2191 11645
rect 2400 11679 2458 11685
rect 2400 11645 2412 11679
rect 2446 11676 2458 11679
rect 2958 11676 2964 11688
rect 2446 11648 2964 11676
rect 2446 11645 2458 11648
rect 2400 11639 2458 11645
rect 2148 11608 2176 11639
rect 2958 11636 2964 11648
rect 3016 11676 3022 11688
rect 4356 11676 4384 11707
rect 3016 11648 4384 11676
rect 3016 11636 3022 11648
rect 4890 11636 4896 11688
rect 4948 11676 4954 11688
rect 4985 11679 5043 11685
rect 4985 11676 4997 11679
rect 4948 11648 4997 11676
rect 4948 11636 4954 11648
rect 4985 11645 4997 11648
rect 5031 11645 5043 11679
rect 4985 11639 5043 11645
rect 7098 11636 7104 11688
rect 7156 11676 7162 11688
rect 7193 11679 7251 11685
rect 7193 11676 7205 11679
rect 7156 11648 7205 11676
rect 7156 11636 7162 11648
rect 7193 11645 7205 11648
rect 7239 11645 7251 11679
rect 7300 11676 7328 11784
rect 8386 11744 8392 11756
rect 8299 11716 8392 11744
rect 8386 11704 8392 11716
rect 8444 11744 8450 11756
rect 8864 11744 8892 11852
rect 10689 11849 10701 11852
rect 10735 11849 10747 11883
rect 10689 11843 10747 11849
rect 8444 11716 8892 11744
rect 8444 11704 8450 11716
rect 9309 11679 9367 11685
rect 7300 11648 8892 11676
rect 7193 11639 7251 11645
rect 2682 11608 2688 11620
rect 2148 11580 2688 11608
rect 2682 11568 2688 11580
rect 2740 11568 2746 11620
rect 2774 11568 2780 11620
rect 2832 11608 2838 11620
rect 3234 11608 3240 11620
rect 2832 11580 3240 11608
rect 2832 11568 2838 11580
rect 3234 11568 3240 11580
rect 3292 11568 3298 11620
rect 4157 11611 4215 11617
rect 4157 11608 4169 11611
rect 3436 11580 4169 11608
rect 2314 11500 2320 11552
rect 2372 11540 2378 11552
rect 3436 11540 3464 11580
rect 4157 11577 4169 11580
rect 4203 11577 4215 11611
rect 4157 11571 4215 11577
rect 5252 11611 5310 11617
rect 5252 11577 5264 11611
rect 5298 11608 5310 11611
rect 5626 11608 5632 11620
rect 5298 11580 5632 11608
rect 5298 11577 5310 11580
rect 5252 11571 5310 11577
rect 5626 11568 5632 11580
rect 5684 11568 5690 11620
rect 8113 11611 8171 11617
rect 8113 11577 8125 11611
rect 8159 11608 8171 11611
rect 8757 11611 8815 11617
rect 8757 11608 8769 11611
rect 8159 11580 8769 11608
rect 8159 11577 8171 11580
rect 8113 11571 8171 11577
rect 8757 11577 8769 11580
rect 8803 11577 8815 11611
rect 8757 11571 8815 11577
rect 2372 11512 3464 11540
rect 2372 11500 2378 11512
rect 3602 11500 3608 11552
rect 3660 11540 3666 11552
rect 5534 11540 5540 11552
rect 3660 11512 5540 11540
rect 3660 11500 3666 11512
rect 5534 11500 5540 11512
rect 5592 11500 5598 11552
rect 5718 11500 5724 11552
rect 5776 11540 5782 11552
rect 6270 11540 6276 11552
rect 5776 11512 6276 11540
rect 5776 11500 5782 11512
rect 6270 11500 6276 11512
rect 6328 11500 6334 11552
rect 8205 11543 8263 11549
rect 8205 11509 8217 11543
rect 8251 11540 8263 11543
rect 8570 11540 8576 11552
rect 8251 11512 8576 11540
rect 8251 11509 8263 11512
rect 8205 11503 8263 11509
rect 8570 11500 8576 11512
rect 8628 11500 8634 11552
rect 8864 11540 8892 11648
rect 9309 11645 9321 11679
rect 9355 11676 9367 11679
rect 10318 11676 10324 11688
rect 9355 11648 10324 11676
rect 9355 11645 9367 11648
rect 9309 11639 9367 11645
rect 9692 11620 9720 11648
rect 10318 11636 10324 11648
rect 10376 11636 10382 11688
rect 19058 11676 19064 11688
rect 19019 11648 19064 11676
rect 19058 11636 19064 11648
rect 19116 11636 19122 11688
rect 9582 11617 9588 11620
rect 9576 11608 9588 11617
rect 9543 11580 9588 11608
rect 9576 11571 9588 11580
rect 9582 11568 9588 11571
rect 9640 11568 9646 11620
rect 9674 11568 9680 11620
rect 9732 11568 9738 11620
rect 11146 11540 11152 11552
rect 8864 11512 11152 11540
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 19245 11543 19303 11549
rect 19245 11509 19257 11543
rect 19291 11540 19303 11543
rect 19886 11540 19892 11552
rect 19291 11512 19892 11540
rect 19291 11509 19303 11512
rect 19245 11503 19303 11509
rect 19886 11500 19892 11512
rect 19944 11500 19950 11552
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 2314 11336 2320 11348
rect 2275 11308 2320 11336
rect 2314 11296 2320 11308
rect 2372 11296 2378 11348
rect 2777 11339 2835 11345
rect 2777 11305 2789 11339
rect 2823 11336 2835 11339
rect 2866 11336 2872 11348
rect 2823 11308 2872 11336
rect 2823 11305 2835 11308
rect 2777 11299 2835 11305
rect 2866 11296 2872 11308
rect 2924 11296 2930 11348
rect 3234 11296 3240 11348
rect 3292 11336 3298 11348
rect 3329 11339 3387 11345
rect 3329 11336 3341 11339
rect 3292 11308 3341 11336
rect 3292 11296 3298 11308
rect 3329 11305 3341 11308
rect 3375 11305 3387 11339
rect 3329 11299 3387 11305
rect 4246 11296 4252 11348
rect 4304 11336 4310 11348
rect 4525 11339 4583 11345
rect 4525 11336 4537 11339
rect 4304 11308 4537 11336
rect 4304 11296 4310 11308
rect 4525 11305 4537 11308
rect 4571 11305 4583 11339
rect 4525 11299 4583 11305
rect 5537 11339 5595 11345
rect 5537 11305 5549 11339
rect 5583 11336 5595 11339
rect 6178 11336 6184 11348
rect 5583 11308 6184 11336
rect 5583 11305 5595 11308
rect 5537 11299 5595 11305
rect 6178 11296 6184 11308
rect 6236 11296 6242 11348
rect 6917 11339 6975 11345
rect 6917 11305 6929 11339
rect 6963 11336 6975 11339
rect 7006 11336 7012 11348
rect 6963 11308 7012 11336
rect 6963 11305 6975 11308
rect 6917 11299 6975 11305
rect 7006 11296 7012 11308
rect 7064 11296 7070 11348
rect 8570 11336 8576 11348
rect 7107 11308 7328 11336
rect 8531 11308 8576 11336
rect 5905 11271 5963 11277
rect 5905 11237 5917 11271
rect 5951 11268 5963 11271
rect 6086 11268 6092 11280
rect 5951 11240 6092 11268
rect 5951 11237 5963 11240
rect 5905 11231 5963 11237
rect 6086 11228 6092 11240
rect 6144 11268 6150 11280
rect 7107 11268 7135 11308
rect 6144 11240 7135 11268
rect 7300 11268 7328 11308
rect 8570 11296 8576 11308
rect 8628 11296 8634 11348
rect 8662 11296 8668 11348
rect 8720 11336 8726 11348
rect 8720 11308 11100 11336
rect 8720 11296 8726 11308
rect 8941 11271 8999 11277
rect 8941 11268 8953 11271
rect 7300 11240 8953 11268
rect 6144 11228 6150 11240
rect 8941 11237 8953 11240
rect 8987 11237 8999 11271
rect 9582 11268 9588 11280
rect 8941 11231 8999 11237
rect 9232 11240 9588 11268
rect 2685 11203 2743 11209
rect 2685 11169 2697 11203
rect 2731 11200 2743 11203
rect 3234 11200 3240 11212
rect 2731 11172 3240 11200
rect 2731 11169 2743 11172
rect 2685 11163 2743 11169
rect 3234 11160 3240 11172
rect 3292 11160 3298 11212
rect 4065 11203 4123 11209
rect 4065 11169 4077 11203
rect 4111 11200 4123 11203
rect 4893 11203 4951 11209
rect 4893 11200 4905 11203
rect 4111 11172 4905 11200
rect 4111 11169 4123 11172
rect 4065 11163 4123 11169
rect 4893 11169 4905 11172
rect 4939 11169 4951 11203
rect 4893 11163 4951 11169
rect 7285 11203 7343 11209
rect 7285 11169 7297 11203
rect 7331 11200 7343 11203
rect 8478 11200 8484 11212
rect 7331 11172 8484 11200
rect 7331 11169 7343 11172
rect 7285 11163 7343 11169
rect 8478 11160 8484 11172
rect 8536 11160 8542 11212
rect 2961 11135 3019 11141
rect 2961 11101 2973 11135
rect 3007 11101 3019 11135
rect 4982 11132 4988 11144
rect 4943 11104 4988 11132
rect 2961 11095 3019 11101
rect 2682 11024 2688 11076
rect 2740 11064 2746 11076
rect 2976 11064 3004 11095
rect 4982 11092 4988 11104
rect 5040 11092 5046 11144
rect 5169 11135 5227 11141
rect 5169 11101 5181 11135
rect 5215 11132 5227 11135
rect 5626 11132 5632 11144
rect 5215 11104 5632 11132
rect 5215 11101 5227 11104
rect 5169 11095 5227 11101
rect 5626 11092 5632 11104
rect 5684 11092 5690 11144
rect 5997 11135 6055 11141
rect 5997 11132 6009 11135
rect 5920 11104 6009 11132
rect 5920 11076 5948 11104
rect 5997 11101 6009 11104
rect 6043 11101 6055 11135
rect 5997 11095 6055 11101
rect 6181 11135 6239 11141
rect 6181 11101 6193 11135
rect 6227 11132 6239 11135
rect 6362 11132 6368 11144
rect 6227 11104 6368 11132
rect 6227 11101 6239 11104
rect 6181 11095 6239 11101
rect 6362 11092 6368 11104
rect 6420 11092 6426 11144
rect 7377 11135 7435 11141
rect 7377 11101 7389 11135
rect 7423 11101 7435 11135
rect 7377 11095 7435 11101
rect 7561 11135 7619 11141
rect 7561 11101 7573 11135
rect 7607 11132 7619 11135
rect 7742 11132 7748 11144
rect 7607 11104 7748 11132
rect 7607 11101 7619 11104
rect 7561 11095 7619 11101
rect 2740 11036 3004 11064
rect 2740 11024 2746 11036
rect 3234 11024 3240 11076
rect 3292 11064 3298 11076
rect 5258 11064 5264 11076
rect 3292 11036 5264 11064
rect 3292 11024 3298 11036
rect 5258 11024 5264 11036
rect 5316 11024 5322 11076
rect 5902 11024 5908 11076
rect 5960 11024 5966 11076
rect 7392 11064 7420 11095
rect 7742 11092 7748 11104
rect 7800 11092 7806 11144
rect 9232 11141 9260 11240
rect 9582 11228 9588 11240
rect 9640 11268 9646 11280
rect 11072 11268 11100 11308
rect 11146 11296 11152 11348
rect 11204 11336 11210 11348
rect 19058 11336 19064 11348
rect 11204 11308 19064 11336
rect 11204 11296 11210 11308
rect 19058 11296 19064 11308
rect 19116 11296 19122 11348
rect 9640 11240 10916 11268
rect 11072 11240 18644 11268
rect 9640 11228 9646 11240
rect 9674 11200 9680 11212
rect 9635 11172 9680 11200
rect 9674 11160 9680 11172
rect 9732 11160 9738 11212
rect 9944 11203 10002 11209
rect 9944 11169 9956 11203
rect 9990 11200 10002 11203
rect 10778 11200 10784 11212
rect 9990 11172 10784 11200
rect 9990 11169 10002 11172
rect 9944 11163 10002 11169
rect 10778 11160 10784 11172
rect 10836 11160 10842 11212
rect 9033 11135 9091 11141
rect 9033 11101 9045 11135
rect 9079 11101 9091 11135
rect 9033 11095 9091 11101
rect 9217 11135 9275 11141
rect 9217 11101 9229 11135
rect 9263 11101 9275 11135
rect 10888 11132 10916 11240
rect 18616 11209 18644 11240
rect 18601 11203 18659 11209
rect 18601 11169 18613 11203
rect 18647 11169 18659 11203
rect 18601 11163 18659 11169
rect 10888 11104 11100 11132
rect 9217 11095 9275 11101
rect 8570 11064 8576 11076
rect 7392 11036 8576 11064
rect 8570 11024 8576 11036
rect 8628 11024 8634 11076
rect 9048 11064 9076 11095
rect 9398 11064 9404 11076
rect 9048 11036 9404 11064
rect 9398 11024 9404 11036
rect 9456 11024 9462 11076
rect 11072 11073 11100 11104
rect 11057 11067 11115 11073
rect 11057 11033 11069 11067
rect 11103 11033 11115 11067
rect 11057 11027 11115 11033
rect 18785 11067 18843 11073
rect 18785 11033 18797 11067
rect 18831 11064 18843 11067
rect 19426 11064 19432 11076
rect 18831 11036 19432 11064
rect 18831 11033 18843 11036
rect 18785 11027 18843 11033
rect 19426 11024 19432 11036
rect 19484 11024 19490 11076
rect 4062 10956 4068 11008
rect 4120 10996 4126 11008
rect 9674 10996 9680 11008
rect 4120 10968 9680 10996
rect 4120 10956 4126 10968
rect 9674 10956 9680 10968
rect 9732 10956 9738 11008
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 2958 10792 2964 10804
rect 2919 10764 2964 10792
rect 2958 10752 2964 10764
rect 3016 10752 3022 10804
rect 3326 10752 3332 10804
rect 3384 10792 3390 10804
rect 3697 10795 3755 10801
rect 3697 10792 3709 10795
rect 3384 10764 3709 10792
rect 3384 10752 3390 10764
rect 3697 10761 3709 10764
rect 3743 10761 3755 10795
rect 3697 10755 3755 10761
rect 5626 10752 5632 10804
rect 5684 10792 5690 10804
rect 6365 10795 6423 10801
rect 6365 10792 6377 10795
rect 5684 10764 6377 10792
rect 5684 10752 5690 10764
rect 6365 10761 6377 10764
rect 6411 10761 6423 10795
rect 9490 10792 9496 10804
rect 6365 10755 6423 10761
rect 7392 10764 9496 10792
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 4338 10656 4344 10668
rect 4299 10628 4344 10656
rect 4338 10616 4344 10628
rect 4396 10616 4402 10668
rect 4890 10616 4896 10668
rect 4948 10656 4954 10668
rect 4985 10659 5043 10665
rect 4985 10656 4997 10659
rect 4948 10628 4997 10656
rect 4948 10616 4954 10628
rect 4985 10625 4997 10628
rect 5031 10625 5043 10659
rect 4985 10619 5043 10625
rect 1848 10591 1906 10597
rect 1848 10557 1860 10591
rect 1894 10588 1906 10591
rect 2682 10588 2688 10600
rect 1894 10560 2688 10588
rect 1894 10557 1906 10560
rect 1848 10551 1906 10557
rect 2682 10548 2688 10560
rect 2740 10548 2746 10600
rect 3050 10548 3056 10600
rect 3108 10588 3114 10600
rect 7392 10597 7420 10764
rect 9490 10752 9496 10764
rect 9548 10752 9554 10804
rect 10502 10792 10508 10804
rect 10463 10764 10508 10792
rect 10502 10752 10508 10764
rect 10560 10752 10566 10804
rect 9030 10724 9036 10736
rect 8991 10696 9036 10724
rect 9030 10684 9036 10696
rect 9088 10724 9094 10736
rect 9677 10727 9735 10733
rect 9088 10696 9260 10724
rect 9088 10684 9094 10696
rect 9232 10656 9260 10696
rect 9677 10693 9689 10727
rect 9723 10724 9735 10727
rect 9723 10696 11008 10724
rect 9723 10693 9735 10696
rect 9677 10687 9735 10693
rect 10980 10665 11008 10696
rect 10229 10659 10287 10665
rect 10229 10656 10241 10659
rect 9232 10628 10241 10656
rect 10229 10625 10241 10628
rect 10275 10625 10287 10659
rect 10229 10619 10287 10625
rect 10965 10659 11023 10665
rect 10965 10625 10977 10659
rect 11011 10625 11023 10659
rect 10965 10619 11023 10625
rect 11057 10659 11115 10665
rect 11057 10625 11069 10659
rect 11103 10625 11115 10659
rect 11057 10619 11115 10625
rect 7377 10591 7435 10597
rect 3108 10560 5764 10588
rect 3108 10548 3114 10560
rect 5736 10532 5764 10560
rect 7377 10557 7389 10591
rect 7423 10557 7435 10591
rect 7650 10588 7656 10600
rect 7611 10560 7656 10588
rect 7377 10551 7435 10557
rect 7650 10548 7656 10560
rect 7708 10548 7714 10600
rect 7742 10548 7748 10600
rect 7800 10588 7806 10600
rect 7909 10591 7967 10597
rect 7909 10588 7921 10591
rect 7800 10560 7921 10588
rect 7800 10548 7806 10560
rect 7909 10557 7921 10560
rect 7955 10557 7967 10591
rect 7909 10551 7967 10557
rect 9122 10548 9128 10600
rect 9180 10588 9186 10600
rect 10137 10591 10195 10597
rect 10137 10588 10149 10591
rect 9180 10560 10149 10588
rect 9180 10548 9186 10560
rect 10137 10557 10149 10560
rect 10183 10557 10195 10591
rect 10137 10551 10195 10557
rect 10778 10548 10784 10600
rect 10836 10588 10842 10600
rect 11072 10588 11100 10619
rect 18230 10588 18236 10600
rect 10836 10560 11100 10588
rect 18191 10560 18236 10588
rect 10836 10548 10842 10560
rect 18230 10548 18236 10560
rect 18288 10548 18294 10600
rect 4065 10523 4123 10529
rect 4065 10489 4077 10523
rect 4111 10520 4123 10523
rect 5074 10520 5080 10532
rect 4111 10492 5080 10520
rect 4111 10489 4123 10492
rect 4065 10483 4123 10489
rect 5074 10480 5080 10492
rect 5132 10480 5138 10532
rect 5252 10523 5310 10529
rect 5252 10489 5264 10523
rect 5298 10520 5310 10523
rect 5442 10520 5448 10532
rect 5298 10492 5448 10520
rect 5298 10489 5310 10492
rect 5252 10483 5310 10489
rect 5442 10480 5448 10492
rect 5500 10480 5506 10532
rect 5718 10480 5724 10532
rect 5776 10520 5782 10532
rect 9401 10523 9459 10529
rect 5776 10492 7328 10520
rect 5776 10480 5782 10492
rect 2774 10412 2780 10464
rect 2832 10452 2838 10464
rect 3418 10452 3424 10464
rect 2832 10424 3424 10452
rect 2832 10412 2838 10424
rect 3418 10412 3424 10424
rect 3476 10412 3482 10464
rect 4157 10455 4215 10461
rect 4157 10421 4169 10455
rect 4203 10452 4215 10455
rect 6822 10452 6828 10464
rect 4203 10424 6828 10452
rect 4203 10421 4215 10424
rect 4157 10415 4215 10421
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 7098 10412 7104 10464
rect 7156 10452 7162 10464
rect 7193 10455 7251 10461
rect 7193 10452 7205 10455
rect 7156 10424 7205 10452
rect 7156 10412 7162 10424
rect 7193 10421 7205 10424
rect 7239 10421 7251 10455
rect 7300 10452 7328 10492
rect 9401 10489 9413 10523
rect 9447 10520 9459 10523
rect 10873 10523 10931 10529
rect 10873 10520 10885 10523
rect 9447 10492 10885 10520
rect 9447 10489 9459 10492
rect 9401 10483 9459 10489
rect 10873 10489 10885 10492
rect 10919 10489 10931 10523
rect 10873 10483 10931 10489
rect 10045 10455 10103 10461
rect 10045 10452 10057 10455
rect 7300 10424 10057 10452
rect 7193 10415 7251 10421
rect 10045 10421 10057 10424
rect 10091 10421 10103 10455
rect 10045 10415 10103 10421
rect 18417 10455 18475 10461
rect 18417 10421 18429 10455
rect 18463 10452 18475 10455
rect 18690 10452 18696 10464
rect 18463 10424 18696 10452
rect 18463 10421 18475 10424
rect 18417 10415 18475 10421
rect 18690 10412 18696 10424
rect 18748 10412 18754 10464
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 3050 10248 3056 10260
rect 3011 10220 3056 10248
rect 3050 10208 3056 10220
rect 3108 10208 3114 10260
rect 3145 10251 3203 10257
rect 3145 10217 3157 10251
rect 3191 10248 3203 10251
rect 4246 10248 4252 10260
rect 3191 10220 4252 10248
rect 3191 10217 3203 10220
rect 3145 10211 3203 10217
rect 4246 10208 4252 10220
rect 4304 10208 4310 10260
rect 5442 10208 5448 10260
rect 5500 10248 5506 10260
rect 5629 10251 5687 10257
rect 5629 10248 5641 10251
rect 5500 10220 5641 10248
rect 5500 10208 5506 10220
rect 5629 10217 5641 10220
rect 5675 10217 5687 10251
rect 5629 10211 5687 10217
rect 7742 10208 7748 10260
rect 7800 10248 7806 10260
rect 8205 10251 8263 10257
rect 8205 10248 8217 10251
rect 7800 10220 8217 10248
rect 7800 10208 7806 10220
rect 8205 10217 8217 10220
rect 8251 10217 8263 10251
rect 8478 10248 8484 10260
rect 8439 10220 8484 10248
rect 8205 10211 8263 10217
rect 8478 10208 8484 10220
rect 8536 10208 8542 10260
rect 9582 10208 9588 10260
rect 9640 10248 9646 10260
rect 11149 10251 11207 10257
rect 11149 10248 11161 10251
rect 9640 10220 11161 10248
rect 9640 10208 9646 10220
rect 11149 10217 11161 10220
rect 11195 10248 11207 10251
rect 11974 10248 11980 10260
rect 11195 10220 11980 10248
rect 11195 10217 11207 10220
rect 11149 10211 11207 10217
rect 11974 10208 11980 10220
rect 12032 10208 12038 10260
rect 2682 10140 2688 10192
rect 2740 10180 2746 10192
rect 2740 10152 3280 10180
rect 2740 10140 2746 10152
rect 2774 10044 2780 10056
rect 2700 10016 2780 10044
rect 2700 9985 2728 10016
rect 2774 10004 2780 10016
rect 2832 10004 2838 10056
rect 3252 10053 3280 10152
rect 3694 10140 3700 10192
rect 3752 10180 3758 10192
rect 3752 10152 5295 10180
rect 3752 10140 3758 10152
rect 4338 10072 4344 10124
rect 4396 10112 4402 10124
rect 4516 10115 4574 10121
rect 4516 10112 4528 10115
rect 4396 10084 4528 10112
rect 4396 10072 4402 10084
rect 4516 10081 4528 10084
rect 4562 10112 4574 10115
rect 4890 10112 4896 10124
rect 4562 10084 4896 10112
rect 4562 10081 4574 10084
rect 4516 10075 4574 10081
rect 4890 10072 4896 10084
rect 4948 10072 4954 10124
rect 3237 10047 3295 10053
rect 3237 10013 3249 10047
rect 3283 10013 3295 10047
rect 3237 10007 3295 10013
rect 3510 10004 3516 10056
rect 3568 10044 3574 10056
rect 4249 10047 4307 10053
rect 4249 10044 4261 10047
rect 3568 10016 4261 10044
rect 3568 10004 3574 10016
rect 4249 10013 4261 10016
rect 4295 10013 4307 10047
rect 5267 10044 5295 10152
rect 5534 10140 5540 10192
rect 5592 10180 5598 10192
rect 6181 10183 6239 10189
rect 6181 10180 6193 10183
rect 5592 10152 6193 10180
rect 5592 10140 5598 10152
rect 6181 10149 6193 10152
rect 6227 10149 6239 10183
rect 6181 10143 6239 10149
rect 6638 10140 6644 10192
rect 6696 10180 6702 10192
rect 9677 10183 9735 10189
rect 9677 10180 9689 10183
rect 6696 10152 9689 10180
rect 6696 10140 6702 10152
rect 9677 10149 9689 10152
rect 9723 10149 9735 10183
rect 9677 10143 9735 10149
rect 5905 10115 5963 10121
rect 5905 10081 5917 10115
rect 5951 10112 5963 10115
rect 6454 10112 6460 10124
rect 5951 10084 6460 10112
rect 5951 10081 5963 10084
rect 5905 10075 5963 10081
rect 6454 10072 6460 10084
rect 6512 10072 6518 10124
rect 6825 10115 6883 10121
rect 6825 10081 6837 10115
rect 6871 10112 6883 10115
rect 6914 10112 6920 10124
rect 6871 10084 6920 10112
rect 6871 10081 6883 10084
rect 6825 10075 6883 10081
rect 6914 10072 6920 10084
rect 6972 10072 6978 10124
rect 7092 10115 7150 10121
rect 7092 10081 7104 10115
rect 7138 10112 7150 10115
rect 8202 10112 8208 10124
rect 7138 10084 8208 10112
rect 7138 10081 7150 10084
rect 7092 10075 7150 10081
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 8294 10072 8300 10124
rect 8352 10112 8358 10124
rect 8849 10115 8907 10121
rect 8849 10112 8861 10115
rect 8352 10084 8861 10112
rect 8352 10072 8358 10084
rect 8849 10081 8861 10084
rect 8895 10081 8907 10115
rect 8849 10075 8907 10081
rect 9861 10115 9919 10121
rect 9861 10081 9873 10115
rect 9907 10112 9919 10115
rect 10318 10112 10324 10124
rect 9907 10084 10324 10112
rect 9907 10081 9919 10084
rect 9861 10075 9919 10081
rect 10318 10072 10324 10084
rect 10376 10072 10382 10124
rect 6546 10044 6552 10056
rect 5267 10016 6552 10044
rect 4249 10007 4307 10013
rect 6546 10004 6552 10016
rect 6604 10004 6610 10056
rect 8662 10004 8668 10056
rect 8720 10044 8726 10056
rect 8941 10047 8999 10053
rect 8941 10044 8953 10047
rect 8720 10016 8953 10044
rect 8720 10004 8726 10016
rect 8941 10013 8953 10016
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 9033 10047 9091 10053
rect 9033 10013 9045 10047
rect 9079 10013 9091 10047
rect 9033 10007 9091 10013
rect 2685 9979 2743 9985
rect 2685 9945 2697 9979
rect 2731 9945 2743 9979
rect 2685 9939 2743 9945
rect 8202 9936 8208 9988
rect 8260 9976 8266 9988
rect 9048 9976 9076 10007
rect 9214 9976 9220 9988
rect 8260 9948 9220 9976
rect 8260 9936 8266 9948
rect 9214 9936 9220 9948
rect 9272 9936 9278 9988
rect 9677 9979 9735 9985
rect 9677 9945 9689 9979
rect 9723 9976 9735 9979
rect 18230 9976 18236 9988
rect 9723 9948 18236 9976
rect 9723 9945 9735 9948
rect 9677 9939 9735 9945
rect 18230 9936 18236 9948
rect 18288 9936 18294 9988
rect 4062 9868 4068 9920
rect 4120 9908 4126 9920
rect 10870 9908 10876 9920
rect 4120 9880 10876 9908
rect 4120 9868 4126 9880
rect 10870 9868 10876 9880
rect 10928 9868 10934 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 2682 9664 2688 9716
rect 2740 9704 2746 9716
rect 2961 9707 3019 9713
rect 2961 9704 2973 9707
rect 2740 9676 2973 9704
rect 2740 9664 2746 9676
rect 2961 9673 2973 9676
rect 3007 9673 3019 9707
rect 2961 9667 3019 9673
rect 3786 9664 3792 9716
rect 3844 9704 3850 9716
rect 3878 9704 3884 9716
rect 3844 9676 3884 9704
rect 3844 9664 3850 9676
rect 3878 9664 3884 9676
rect 3936 9664 3942 9716
rect 4890 9704 4896 9716
rect 4851 9676 4896 9704
rect 4890 9664 4896 9676
rect 4948 9664 4954 9716
rect 10137 9707 10195 9713
rect 10137 9673 10149 9707
rect 10183 9704 10195 9707
rect 10778 9704 10784 9716
rect 10183 9676 10784 9704
rect 10183 9673 10195 9676
rect 10137 9667 10195 9673
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 10870 9664 10876 9716
rect 10928 9704 10934 9716
rect 14366 9704 14372 9716
rect 10928 9676 14372 9704
rect 10928 9664 10934 9676
rect 14366 9664 14372 9676
rect 14424 9664 14430 9716
rect 4982 9596 4988 9648
rect 5040 9636 5046 9648
rect 5169 9639 5227 9645
rect 5169 9636 5181 9639
rect 5040 9608 5181 9636
rect 5040 9596 5046 9608
rect 5169 9605 5181 9608
rect 5215 9605 5227 9639
rect 6822 9636 6828 9648
rect 6783 9608 6828 9636
rect 5169 9599 5227 9605
rect 6822 9596 6828 9608
rect 6880 9596 6886 9648
rect 10410 9636 10416 9648
rect 10371 9608 10416 9636
rect 10410 9596 10416 9608
rect 10468 9596 10474 9648
rect 5442 9528 5448 9580
rect 5500 9568 5506 9580
rect 5721 9571 5779 9577
rect 5721 9568 5733 9571
rect 5500 9540 5733 9568
rect 5500 9528 5506 9540
rect 5721 9537 5733 9540
rect 5767 9537 5779 9571
rect 7377 9571 7435 9577
rect 7377 9568 7389 9571
rect 5721 9531 5779 9537
rect 5828 9540 7389 9568
rect 1578 9500 1584 9512
rect 1539 9472 1584 9500
rect 1578 9460 1584 9472
rect 1636 9500 1642 9512
rect 3510 9500 3516 9512
rect 1636 9472 3516 9500
rect 1636 9460 1642 9472
rect 3510 9460 3516 9472
rect 3568 9460 3574 9512
rect 3780 9503 3838 9509
rect 3780 9469 3792 9503
rect 3826 9500 3838 9503
rect 4706 9500 4712 9512
rect 3826 9472 4712 9500
rect 3826 9469 3838 9472
rect 3780 9463 3838 9469
rect 4706 9460 4712 9472
rect 4764 9460 4770 9512
rect 5534 9460 5540 9512
rect 5592 9500 5598 9512
rect 5629 9503 5687 9509
rect 5629 9500 5641 9503
rect 5592 9472 5641 9500
rect 5592 9460 5598 9472
rect 5629 9469 5641 9472
rect 5675 9469 5687 9503
rect 5629 9463 5687 9469
rect 1848 9435 1906 9441
rect 1848 9401 1860 9435
rect 1894 9432 1906 9435
rect 2314 9432 2320 9444
rect 1894 9404 2320 9432
rect 1894 9401 1906 9404
rect 1848 9395 1906 9401
rect 2314 9392 2320 9404
rect 2372 9432 2378 9444
rect 2774 9432 2780 9444
rect 2372 9404 2780 9432
rect 2372 9392 2378 9404
rect 2774 9392 2780 9404
rect 2832 9392 2838 9444
rect 4724 9432 4752 9460
rect 5828 9432 5856 9540
rect 7377 9537 7389 9540
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 7837 9571 7895 9577
rect 7837 9537 7849 9571
rect 7883 9568 7895 9571
rect 8294 9568 8300 9580
rect 7883 9540 8300 9568
rect 7883 9537 7895 9540
rect 7837 9531 7895 9537
rect 8294 9528 8300 9540
rect 8352 9528 8358 9580
rect 7650 9460 7656 9512
rect 7708 9500 7714 9512
rect 9030 9509 9036 9512
rect 8757 9503 8815 9509
rect 8757 9500 8769 9503
rect 7708 9472 8769 9500
rect 7708 9460 7714 9472
rect 8757 9469 8769 9472
rect 8803 9469 8815 9503
rect 9024 9500 9036 9509
rect 8991 9472 9036 9500
rect 8757 9463 8815 9469
rect 9024 9463 9036 9472
rect 9030 9460 9036 9463
rect 9088 9460 9094 9512
rect 10597 9503 10655 9509
rect 10597 9469 10609 9503
rect 10643 9500 10655 9503
rect 11790 9500 11796 9512
rect 10643 9472 11796 9500
rect 10643 9469 10655 9472
rect 10597 9463 10655 9469
rect 11790 9460 11796 9472
rect 11848 9460 11854 9512
rect 4724 9404 5856 9432
rect 6914 9392 6920 9444
rect 6972 9432 6978 9444
rect 7285 9435 7343 9441
rect 7285 9432 7297 9435
rect 6972 9404 7297 9432
rect 6972 9392 6978 9404
rect 7285 9401 7297 9404
rect 7331 9401 7343 9435
rect 7285 9395 7343 9401
rect 9674 9392 9680 9444
rect 9732 9432 9738 9444
rect 11146 9432 11152 9444
rect 9732 9404 11152 9432
rect 9732 9392 9738 9404
rect 11146 9392 11152 9404
rect 11204 9392 11210 9444
rect 4430 9324 4436 9376
rect 4488 9364 4494 9376
rect 4798 9364 4804 9376
rect 4488 9336 4804 9364
rect 4488 9324 4494 9336
rect 4798 9324 4804 9336
rect 4856 9364 4862 9376
rect 4982 9364 4988 9376
rect 4856 9336 4988 9364
rect 4856 9324 4862 9336
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 5537 9367 5595 9373
rect 5537 9333 5549 9367
rect 5583 9364 5595 9367
rect 5718 9364 5724 9376
rect 5583 9336 5724 9364
rect 5583 9333 5595 9336
rect 5537 9327 5595 9333
rect 5718 9324 5724 9336
rect 5776 9324 5782 9376
rect 6178 9364 6184 9376
rect 6139 9336 6184 9364
rect 6178 9324 6184 9336
rect 6236 9324 6242 9376
rect 6822 9324 6828 9376
rect 6880 9364 6886 9376
rect 7193 9367 7251 9373
rect 7193 9364 7205 9367
rect 6880 9336 7205 9364
rect 6880 9324 6886 9336
rect 7193 9333 7205 9336
rect 7239 9364 7251 9367
rect 8938 9364 8944 9376
rect 7239 9336 8944 9364
rect 7239 9333 7251 9336
rect 7193 9327 7251 9333
rect 8938 9324 8944 9336
rect 8996 9324 9002 9376
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 2774 9160 2780 9172
rect 2735 9132 2780 9160
rect 2774 9120 2780 9132
rect 2832 9120 2838 9172
rect 4430 9160 4436 9172
rect 4391 9132 4436 9160
rect 4430 9120 4436 9132
rect 4488 9120 4494 9172
rect 4525 9163 4583 9169
rect 4525 9129 4537 9163
rect 4571 9160 4583 9163
rect 5074 9160 5080 9172
rect 4571 9132 4936 9160
rect 5035 9132 5080 9160
rect 4571 9129 4583 9132
rect 4525 9123 4583 9129
rect 4706 9052 4712 9104
rect 4764 9052 4770 9104
rect 4908 9092 4936 9132
rect 5074 9120 5080 9132
rect 5132 9120 5138 9172
rect 5445 9163 5503 9169
rect 5445 9129 5457 9163
rect 5491 9160 5503 9163
rect 6178 9160 6184 9172
rect 5491 9132 6184 9160
rect 5491 9129 5503 9132
rect 5445 9123 5503 9129
rect 6178 9120 6184 9132
rect 6236 9120 6242 9172
rect 8570 9160 8576 9172
rect 8531 9132 8576 9160
rect 8570 9120 8576 9132
rect 8628 9120 8634 9172
rect 8938 9160 8944 9172
rect 8899 9132 8944 9160
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 4908 9064 5764 9092
rect 1664 9027 1722 9033
rect 1664 8993 1676 9027
rect 1710 9024 1722 9027
rect 2498 9024 2504 9036
rect 1710 8996 2504 9024
rect 1710 8993 1722 8996
rect 1664 8987 1722 8993
rect 2498 8984 2504 8996
rect 2556 8984 2562 9036
rect 4724 9024 4752 9052
rect 5736 9024 5764 9064
rect 5810 9052 5816 9104
rect 5868 9092 5874 9104
rect 12250 9092 12256 9104
rect 5868 9064 12256 9092
rect 5868 9052 5874 9064
rect 12250 9052 12256 9064
rect 12308 9052 12314 9104
rect 6178 9024 6184 9036
rect 4724 8996 5672 9024
rect 5736 8996 6184 9024
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8925 1455 8959
rect 4706 8956 4712 8968
rect 4667 8928 4712 8956
rect 1397 8919 1455 8925
rect 1412 8820 1440 8919
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 5258 8916 5264 8968
rect 5316 8956 5322 8968
rect 5644 8965 5672 8996
rect 6178 8984 6184 8996
rect 6236 8984 6242 9036
rect 6730 9024 6736 9036
rect 6691 8996 6736 9024
rect 6730 8984 6736 8996
rect 6788 8984 6794 9036
rect 6825 9027 6883 9033
rect 6825 8993 6837 9027
rect 6871 9024 6883 9027
rect 7006 9024 7012 9036
rect 6871 8996 7012 9024
rect 6871 8993 6883 8996
rect 6825 8987 6883 8993
rect 7006 8984 7012 8996
rect 7064 8984 7070 9036
rect 7742 8984 7748 9036
rect 7800 9024 7806 9036
rect 7929 9027 7987 9033
rect 7929 9024 7941 9027
rect 7800 8996 7941 9024
rect 7800 8984 7806 8996
rect 7929 8993 7941 8996
rect 7975 8993 7987 9027
rect 7929 8987 7987 8993
rect 8021 9027 8079 9033
rect 8021 8993 8033 9027
rect 8067 9024 8079 9027
rect 8202 9024 8208 9036
rect 8067 8996 8208 9024
rect 8067 8993 8079 8996
rect 8021 8987 8079 8993
rect 8202 8984 8208 8996
rect 8260 8984 8266 9036
rect 10312 9027 10370 9033
rect 10312 8993 10324 9027
rect 10358 9024 10370 9027
rect 10870 9024 10876 9036
rect 10358 8996 10876 9024
rect 10358 8993 10370 8996
rect 10312 8987 10370 8993
rect 10870 8984 10876 8996
rect 10928 8984 10934 9036
rect 5537 8959 5595 8965
rect 5537 8956 5549 8959
rect 5316 8928 5549 8956
rect 5316 8916 5322 8928
rect 5537 8925 5549 8928
rect 5583 8925 5595 8959
rect 5537 8919 5595 8925
rect 5629 8959 5687 8965
rect 5629 8925 5641 8959
rect 5675 8925 5687 8959
rect 5629 8919 5687 8925
rect 6546 8916 6552 8968
rect 6604 8956 6610 8968
rect 6917 8959 6975 8965
rect 6917 8956 6929 8959
rect 6604 8928 6929 8956
rect 6604 8916 6610 8928
rect 6917 8925 6929 8928
rect 6963 8956 6975 8959
rect 8110 8956 8116 8968
rect 6963 8928 8116 8956
rect 6963 8925 6975 8928
rect 6917 8919 6975 8925
rect 8110 8916 8116 8928
rect 8168 8916 8174 8968
rect 8570 8916 8576 8968
rect 8628 8956 8634 8968
rect 9033 8959 9091 8965
rect 9033 8956 9045 8959
rect 8628 8928 9045 8956
rect 8628 8916 8634 8928
rect 9033 8925 9045 8928
rect 9079 8925 9091 8959
rect 9214 8956 9220 8968
rect 9175 8928 9220 8956
rect 9033 8919 9091 8925
rect 9214 8916 9220 8928
rect 9272 8916 9278 8968
rect 9674 8916 9680 8968
rect 9732 8956 9738 8968
rect 10045 8959 10103 8965
rect 10045 8956 10057 8959
rect 9732 8928 10057 8956
rect 9732 8916 9738 8928
rect 10045 8925 10057 8928
rect 10091 8925 10103 8959
rect 10045 8919 10103 8925
rect 3970 8848 3976 8900
rect 4028 8888 4034 8900
rect 9306 8888 9312 8900
rect 4028 8860 9312 8888
rect 4028 8848 4034 8860
rect 9306 8848 9312 8860
rect 9364 8848 9370 8900
rect 1578 8820 1584 8832
rect 1412 8792 1584 8820
rect 1578 8780 1584 8792
rect 1636 8820 1642 8832
rect 2590 8820 2596 8832
rect 1636 8792 2596 8820
rect 1636 8780 1642 8792
rect 2590 8780 2596 8792
rect 2648 8780 2654 8832
rect 4065 8823 4123 8829
rect 4065 8789 4077 8823
rect 4111 8820 4123 8823
rect 4798 8820 4804 8832
rect 4111 8792 4804 8820
rect 4111 8789 4123 8792
rect 4065 8783 4123 8789
rect 4798 8780 4804 8792
rect 4856 8780 4862 8832
rect 6365 8823 6423 8829
rect 6365 8789 6377 8823
rect 6411 8820 6423 8823
rect 7190 8820 7196 8832
rect 6411 8792 7196 8820
rect 6411 8789 6423 8792
rect 6365 8783 6423 8789
rect 7190 8780 7196 8792
rect 7248 8780 7254 8832
rect 7282 8780 7288 8832
rect 7340 8820 7346 8832
rect 7561 8823 7619 8829
rect 7561 8820 7573 8823
rect 7340 8792 7573 8820
rect 7340 8780 7346 8792
rect 7561 8789 7573 8792
rect 7607 8789 7619 8823
rect 7561 8783 7619 8789
rect 8846 8780 8852 8832
rect 8904 8820 8910 8832
rect 11425 8823 11483 8829
rect 11425 8820 11437 8823
rect 8904 8792 11437 8820
rect 8904 8780 8910 8792
rect 11425 8789 11437 8792
rect 11471 8789 11483 8823
rect 11425 8783 11483 8789
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 1670 8576 1676 8628
rect 1728 8616 1734 8628
rect 1765 8619 1823 8625
rect 1765 8616 1777 8619
rect 1728 8588 1777 8616
rect 1728 8576 1734 8588
rect 1765 8585 1777 8588
rect 1811 8585 1823 8619
rect 7650 8616 7656 8628
rect 1765 8579 1823 8585
rect 7392 8588 7656 8616
rect 4430 8548 4436 8560
rect 4391 8520 4436 8548
rect 4430 8508 4436 8520
rect 4488 8508 4494 8560
rect 4706 8508 4712 8560
rect 4764 8548 4770 8560
rect 4764 8520 6040 8548
rect 4764 8508 4770 8520
rect 2314 8480 2320 8492
rect 2275 8452 2320 8480
rect 2314 8440 2320 8452
rect 2372 8440 2378 8492
rect 4890 8440 4896 8492
rect 4948 8480 4954 8492
rect 6012 8489 6040 8520
rect 4985 8483 5043 8489
rect 4985 8480 4997 8483
rect 4948 8452 4997 8480
rect 4948 8440 4954 8452
rect 4985 8449 4997 8452
rect 5031 8449 5043 8483
rect 4985 8443 5043 8449
rect 5997 8483 6055 8489
rect 5997 8449 6009 8483
rect 6043 8449 6055 8483
rect 5997 8443 6055 8449
rect 6730 8440 6736 8492
rect 6788 8480 6794 8492
rect 7392 8489 7420 8588
rect 7650 8576 7656 8588
rect 7708 8576 7714 8628
rect 8110 8576 8116 8628
rect 8168 8616 8174 8628
rect 8757 8619 8815 8625
rect 8757 8616 8769 8619
rect 8168 8588 8769 8616
rect 8168 8576 8174 8588
rect 8757 8585 8769 8588
rect 8803 8585 8815 8619
rect 8757 8579 8815 8585
rect 10870 8576 10876 8628
rect 10928 8616 10934 8628
rect 11057 8619 11115 8625
rect 11057 8616 11069 8619
rect 10928 8588 11069 8616
rect 10928 8576 10934 8588
rect 11057 8585 11069 8588
rect 11103 8585 11115 8619
rect 11790 8616 11796 8628
rect 11751 8588 11796 8616
rect 11057 8579 11115 8585
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 9217 8551 9275 8557
rect 9217 8548 9229 8551
rect 9140 8520 9229 8548
rect 6825 8483 6883 8489
rect 6825 8480 6837 8483
rect 6788 8452 6837 8480
rect 6788 8440 6794 8452
rect 6825 8449 6837 8452
rect 6871 8449 6883 8483
rect 6825 8443 6883 8449
rect 7377 8483 7435 8489
rect 7377 8449 7389 8483
rect 7423 8449 7435 8483
rect 7377 8443 7435 8449
rect 9140 8480 9168 8520
rect 9217 8517 9229 8520
rect 9263 8517 9275 8551
rect 9217 8511 9275 8517
rect 9674 8480 9680 8492
rect 9140 8452 9680 8480
rect 2774 8372 2780 8424
rect 2832 8412 2838 8424
rect 2832 8384 2877 8412
rect 2832 8372 2838 8384
rect 3786 8372 3792 8424
rect 3844 8412 3850 8424
rect 4798 8412 4804 8424
rect 3844 8384 4660 8412
rect 4759 8384 4804 8412
rect 3844 8372 3850 8384
rect 3044 8347 3102 8353
rect 3044 8313 3056 8347
rect 3090 8344 3102 8347
rect 4632 8344 4660 8384
rect 4798 8372 4804 8384
rect 4856 8372 4862 8424
rect 5813 8415 5871 8421
rect 5813 8412 5825 8415
rect 5092 8384 5825 8412
rect 5092 8344 5120 8384
rect 5813 8381 5825 8384
rect 5859 8412 5871 8415
rect 6641 8415 6699 8421
rect 5859 8384 6592 8412
rect 5859 8381 5871 8384
rect 5813 8375 5871 8381
rect 3090 8316 4292 8344
rect 4632 8316 5120 8344
rect 3090 8313 3102 8316
rect 3044 8307 3102 8313
rect 2130 8276 2136 8288
rect 2091 8248 2136 8276
rect 2130 8236 2136 8248
rect 2188 8236 2194 8288
rect 2222 8236 2228 8288
rect 2280 8276 2286 8288
rect 2280 8248 2325 8276
rect 2280 8236 2286 8248
rect 2774 8236 2780 8288
rect 2832 8276 2838 8288
rect 4154 8276 4160 8288
rect 2832 8248 4160 8276
rect 2832 8236 2838 8248
rect 4154 8236 4160 8248
rect 4212 8236 4218 8288
rect 4264 8276 4292 8316
rect 5166 8304 5172 8356
rect 5224 8344 5230 8356
rect 5905 8347 5963 8353
rect 5224 8316 5580 8344
rect 5224 8304 5230 8316
rect 4798 8276 4804 8288
rect 4264 8248 4804 8276
rect 4798 8236 4804 8248
rect 4856 8236 4862 8288
rect 4893 8279 4951 8285
rect 4893 8245 4905 8279
rect 4939 8276 4951 8279
rect 5445 8279 5503 8285
rect 5445 8276 5457 8279
rect 4939 8248 5457 8276
rect 4939 8245 4951 8248
rect 4893 8239 4951 8245
rect 5445 8245 5457 8248
rect 5491 8245 5503 8279
rect 5552 8276 5580 8316
rect 5905 8313 5917 8347
rect 5951 8344 5963 8347
rect 6086 8344 6092 8356
rect 5951 8316 6092 8344
rect 5951 8313 5963 8316
rect 5905 8307 5963 8313
rect 6086 8304 6092 8316
rect 6144 8304 6150 8356
rect 6564 8344 6592 8384
rect 6641 8381 6653 8415
rect 6687 8412 6699 8415
rect 7098 8412 7104 8424
rect 6687 8384 7104 8412
rect 6687 8381 6699 8384
rect 6641 8375 6699 8381
rect 7098 8372 7104 8384
rect 7156 8372 7162 8424
rect 7392 8412 7420 8443
rect 9140 8412 9168 8452
rect 9674 8440 9680 8452
rect 9732 8440 9738 8492
rect 7392 8384 9168 8412
rect 9401 8415 9459 8421
rect 9401 8381 9413 8415
rect 9447 8381 9459 8415
rect 9401 8375 9459 8381
rect 9944 8415 10002 8421
rect 9944 8381 9956 8415
rect 9990 8412 10002 8415
rect 11698 8412 11704 8424
rect 9990 8384 11704 8412
rect 9990 8381 10002 8384
rect 9944 8375 10002 8381
rect 6822 8344 6828 8356
rect 6564 8316 6828 8344
rect 6822 8304 6828 8316
rect 6880 8304 6886 8356
rect 7650 8353 7656 8356
rect 7644 8344 7656 8353
rect 7611 8316 7656 8344
rect 7644 8307 7656 8316
rect 7650 8304 7656 8307
rect 7708 8304 7714 8356
rect 9416 8344 9444 8375
rect 11698 8372 11704 8384
rect 11756 8372 11762 8424
rect 11974 8412 11980 8424
rect 11935 8384 11980 8412
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 10410 8344 10416 8356
rect 9416 8316 10416 8344
rect 10410 8304 10416 8316
rect 10468 8304 10474 8356
rect 6457 8279 6515 8285
rect 6457 8276 6469 8279
rect 5552 8248 6469 8276
rect 5445 8239 5503 8245
rect 6457 8245 6469 8248
rect 6503 8245 6515 8279
rect 11330 8276 11336 8288
rect 11291 8248 11336 8276
rect 6457 8239 6515 8245
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 2130 8032 2136 8084
rect 2188 8072 2194 8084
rect 2225 8075 2283 8081
rect 2225 8072 2237 8075
rect 2188 8044 2237 8072
rect 2188 8032 2194 8044
rect 2225 8041 2237 8044
rect 2271 8041 2283 8075
rect 2225 8035 2283 8041
rect 2685 8075 2743 8081
rect 2685 8041 2697 8075
rect 2731 8072 2743 8075
rect 4065 8075 4123 8081
rect 4065 8072 4077 8075
rect 2731 8044 4077 8072
rect 2731 8041 2743 8044
rect 2685 8035 2743 8041
rect 4065 8041 4077 8044
rect 4111 8041 4123 8075
rect 5166 8072 5172 8084
rect 4065 8035 4123 8041
rect 4356 8044 5172 8072
rect 2593 7939 2651 7945
rect 2593 7905 2605 7939
rect 2639 7936 2651 7939
rect 3237 7939 3295 7945
rect 3237 7936 3249 7939
rect 2639 7908 3249 7936
rect 2639 7905 2651 7908
rect 2593 7899 2651 7905
rect 3237 7905 3249 7908
rect 3283 7905 3295 7939
rect 3237 7899 3295 7905
rect 3881 7939 3939 7945
rect 3881 7905 3893 7939
rect 3927 7936 3939 7939
rect 4356 7936 4384 8044
rect 5166 8032 5172 8044
rect 5224 8032 5230 8084
rect 7006 8072 7012 8084
rect 6967 8044 7012 8072
rect 7006 8032 7012 8044
rect 7064 8032 7070 8084
rect 7469 8075 7527 8081
rect 7469 8072 7481 8075
rect 7208 8044 7481 8072
rect 5258 8004 5264 8016
rect 4448 7976 5264 8004
rect 4448 7945 4476 7976
rect 5258 7964 5264 7976
rect 5316 7964 5322 8016
rect 5436 8007 5494 8013
rect 5436 7973 5448 8007
rect 5482 8004 5494 8007
rect 6546 8004 6552 8016
rect 5482 7976 6552 8004
rect 5482 7973 5494 7976
rect 5436 7967 5494 7973
rect 6546 7964 6552 7976
rect 6604 7964 6610 8016
rect 3927 7908 4384 7936
rect 4433 7939 4491 7945
rect 3927 7905 3939 7908
rect 3881 7899 3939 7905
rect 4433 7905 4445 7939
rect 4479 7905 4491 7939
rect 4433 7899 4491 7905
rect 4525 7939 4583 7945
rect 4525 7905 4537 7939
rect 4571 7936 4583 7939
rect 4890 7936 4896 7948
rect 4571 7908 4896 7936
rect 4571 7905 4583 7908
rect 4525 7899 4583 7905
rect 2498 7828 2504 7880
rect 2556 7868 2562 7880
rect 2774 7868 2780 7880
rect 2556 7840 2780 7868
rect 2556 7828 2562 7840
rect 2774 7828 2780 7840
rect 2832 7828 2838 7880
rect 4154 7828 4160 7880
rect 4212 7868 4218 7880
rect 4448 7868 4476 7899
rect 4890 7896 4896 7908
rect 4948 7936 4954 7948
rect 6362 7936 6368 7948
rect 4948 7908 6368 7936
rect 4948 7896 4954 7908
rect 6362 7896 6368 7908
rect 6420 7936 6426 7948
rect 7208 7936 7236 8044
rect 7469 8041 7481 8044
rect 7515 8041 7527 8075
rect 7469 8035 7527 8041
rect 7742 8032 7748 8084
rect 7800 8072 7806 8084
rect 8205 8075 8263 8081
rect 8205 8072 8217 8075
rect 7800 8044 8217 8072
rect 7800 8032 7806 8044
rect 8205 8041 8217 8044
rect 8251 8041 8263 8075
rect 8205 8035 8263 8041
rect 10689 8075 10747 8081
rect 10689 8041 10701 8075
rect 10735 8072 10747 8075
rect 11241 8075 11299 8081
rect 11241 8072 11253 8075
rect 10735 8044 11253 8072
rect 10735 8041 10747 8044
rect 10689 8035 10747 8041
rect 11241 8041 11253 8044
rect 11287 8041 11299 8075
rect 11241 8035 11299 8041
rect 16669 8075 16727 8081
rect 16669 8041 16681 8075
rect 16715 8041 16727 8075
rect 16669 8035 16727 8041
rect 10597 8007 10655 8013
rect 10597 7973 10609 8007
rect 10643 8004 10655 8007
rect 11330 8004 11336 8016
rect 10643 7976 11336 8004
rect 10643 7973 10655 7976
rect 10597 7967 10655 7973
rect 11330 7964 11336 7976
rect 11388 7964 11394 8016
rect 11698 7964 11704 8016
rect 11756 7964 11762 8016
rect 15556 8007 15614 8013
rect 15556 7973 15568 8007
rect 15602 8004 15614 8007
rect 15746 8004 15752 8016
rect 15602 7976 15752 8004
rect 15602 7973 15614 7976
rect 15556 7967 15614 7973
rect 15746 7964 15752 7976
rect 15804 7964 15810 8016
rect 6420 7908 7236 7936
rect 7377 7939 7435 7945
rect 6420 7896 6426 7908
rect 7377 7905 7389 7939
rect 7423 7905 7435 7939
rect 8573 7939 8631 7945
rect 8573 7936 8585 7939
rect 7377 7899 7435 7905
rect 7484 7908 8585 7936
rect 4212 7840 4476 7868
rect 4617 7871 4675 7877
rect 4212 7828 4218 7840
rect 4617 7837 4629 7871
rect 4663 7868 4675 7871
rect 4798 7868 4804 7880
rect 4663 7840 4804 7868
rect 4663 7837 4675 7840
rect 4617 7831 4675 7837
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 2682 7760 2688 7812
rect 2740 7800 2746 7812
rect 3694 7800 3700 7812
rect 2740 7772 3700 7800
rect 2740 7760 2746 7772
rect 3694 7760 3700 7772
rect 3752 7800 3758 7812
rect 5184 7800 5212 7831
rect 7098 7828 7104 7880
rect 7156 7868 7162 7880
rect 7392 7868 7420 7899
rect 7156 7840 7420 7868
rect 7156 7828 7162 7840
rect 7484 7800 7512 7908
rect 8573 7905 8585 7908
rect 8619 7905 8631 7939
rect 8573 7899 8631 7905
rect 11146 7896 11152 7948
rect 11204 7936 11210 7948
rect 11609 7939 11667 7945
rect 11609 7936 11621 7939
rect 11204 7908 11621 7936
rect 11204 7896 11210 7908
rect 11609 7905 11621 7908
rect 11655 7905 11667 7939
rect 11716 7936 11744 7964
rect 16684 7936 16712 8035
rect 11716 7908 16712 7936
rect 11609 7899 11667 7905
rect 7650 7868 7656 7880
rect 7563 7840 7656 7868
rect 7650 7828 7656 7840
rect 7708 7828 7714 7880
rect 8478 7828 8484 7880
rect 8536 7868 8542 7880
rect 8665 7871 8723 7877
rect 8665 7868 8677 7871
rect 8536 7840 8677 7868
rect 8536 7828 8542 7840
rect 8665 7837 8677 7840
rect 8711 7837 8723 7871
rect 8846 7868 8852 7880
rect 8807 7840 8852 7868
rect 8665 7831 8723 7837
rect 8846 7828 8852 7840
rect 8904 7828 8910 7880
rect 10870 7868 10876 7880
rect 10831 7840 10876 7868
rect 10870 7828 10876 7840
rect 10928 7828 10934 7880
rect 10962 7828 10968 7880
rect 11020 7868 11026 7880
rect 11808 7877 11836 7908
rect 11701 7871 11759 7877
rect 11701 7868 11713 7871
rect 11020 7840 11713 7868
rect 11020 7828 11026 7840
rect 11701 7837 11713 7840
rect 11747 7837 11759 7871
rect 11701 7831 11759 7837
rect 11793 7871 11851 7877
rect 11793 7837 11805 7871
rect 11839 7837 11851 7871
rect 11793 7831 11851 7837
rect 15010 7828 15016 7880
rect 15068 7868 15074 7880
rect 15289 7871 15347 7877
rect 15289 7868 15301 7871
rect 15068 7840 15301 7868
rect 15068 7828 15074 7840
rect 15289 7837 15301 7840
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 3752 7772 5212 7800
rect 6380 7772 7512 7800
rect 7668 7800 7696 7828
rect 8864 7800 8892 7828
rect 7668 7772 8892 7800
rect 10229 7803 10287 7809
rect 3752 7760 3758 7772
rect 4982 7692 4988 7744
rect 5040 7732 5046 7744
rect 6380 7732 6408 7772
rect 10229 7769 10241 7803
rect 10275 7800 10287 7803
rect 14642 7800 14648 7812
rect 10275 7772 14648 7800
rect 10275 7769 10287 7772
rect 10229 7763 10287 7769
rect 14642 7760 14648 7772
rect 14700 7760 14706 7812
rect 6546 7732 6552 7744
rect 5040 7704 6408 7732
rect 6507 7704 6552 7732
rect 5040 7692 5046 7704
rect 6546 7692 6552 7704
rect 6604 7692 6610 7744
rect 7006 7692 7012 7744
rect 7064 7732 7070 7744
rect 7558 7732 7564 7744
rect 7064 7704 7564 7732
rect 7064 7692 7070 7704
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 1762 7488 1768 7540
rect 1820 7528 1826 7540
rect 1949 7531 2007 7537
rect 1949 7528 1961 7531
rect 1820 7500 1961 7528
rect 1820 7488 1826 7500
rect 1949 7497 1961 7500
rect 1995 7497 2007 7531
rect 1949 7491 2007 7497
rect 4062 7488 4068 7540
rect 4120 7528 4126 7540
rect 5718 7528 5724 7540
rect 4120 7500 5724 7528
rect 4120 7488 4126 7500
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 6454 7488 6460 7540
rect 6512 7528 6518 7540
rect 6825 7531 6883 7537
rect 6825 7528 6837 7531
rect 6512 7500 6837 7528
rect 6512 7488 6518 7500
rect 6825 7497 6837 7500
rect 6871 7497 6883 7531
rect 6825 7491 6883 7497
rect 8113 7531 8171 7537
rect 8113 7497 8125 7531
rect 8159 7528 8171 7531
rect 8202 7528 8208 7540
rect 8159 7500 8208 7528
rect 8159 7497 8171 7500
rect 8113 7491 8171 7497
rect 8202 7488 8208 7500
rect 8260 7488 8266 7540
rect 5442 7420 5448 7472
rect 5500 7460 5506 7472
rect 7098 7460 7104 7472
rect 5500 7432 7104 7460
rect 5500 7420 5506 7432
rect 7098 7420 7104 7432
rect 7156 7460 7162 7472
rect 8662 7460 8668 7472
rect 7156 7432 8668 7460
rect 7156 7420 7162 7432
rect 8662 7420 8668 7432
rect 8720 7420 8726 7472
rect 14277 7463 14335 7469
rect 14277 7429 14289 7463
rect 14323 7460 14335 7463
rect 15654 7460 15660 7472
rect 14323 7432 15660 7460
rect 14323 7429 14335 7432
rect 14277 7423 14335 7429
rect 15654 7420 15660 7432
rect 15712 7420 15718 7472
rect 2498 7392 2504 7404
rect 2459 7364 2504 7392
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 3602 7392 3608 7404
rect 3563 7364 3608 7392
rect 3602 7352 3608 7364
rect 3660 7352 3666 7404
rect 3694 7352 3700 7404
rect 3752 7392 3758 7404
rect 4433 7395 4491 7401
rect 4433 7392 4445 7395
rect 3752 7364 4445 7392
rect 3752 7352 3758 7364
rect 4433 7361 4445 7364
rect 4479 7361 4491 7395
rect 7282 7392 7288 7404
rect 7243 7364 7288 7392
rect 4433 7355 4491 7361
rect 7282 7352 7288 7364
rect 7340 7352 7346 7404
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 8757 7395 8815 7401
rect 8757 7361 8769 7395
rect 8803 7392 8815 7395
rect 8846 7392 8852 7404
rect 8803 7364 8852 7392
rect 8803 7361 8815 7364
rect 8757 7355 8815 7361
rect 4700 7327 4758 7333
rect 4700 7293 4712 7327
rect 4746 7324 4758 7327
rect 6546 7324 6552 7336
rect 4746 7296 6552 7324
rect 4746 7293 4758 7296
rect 4700 7287 4758 7293
rect 6546 7284 6552 7296
rect 6604 7324 6610 7336
rect 7392 7324 7420 7355
rect 8846 7352 8852 7364
rect 8904 7352 8910 7404
rect 9674 7352 9680 7404
rect 9732 7392 9738 7404
rect 10321 7395 10379 7401
rect 10321 7392 10333 7395
rect 9732 7364 10333 7392
rect 9732 7352 9738 7364
rect 10321 7361 10333 7364
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 14921 7395 14979 7401
rect 14921 7361 14933 7395
rect 14967 7392 14979 7395
rect 15194 7392 15200 7404
rect 14967 7364 15200 7392
rect 14967 7361 14979 7364
rect 14921 7355 14979 7361
rect 6604 7296 7420 7324
rect 8481 7327 8539 7333
rect 6604 7284 6610 7296
rect 8481 7293 8493 7327
rect 8527 7324 8539 7327
rect 8938 7324 8944 7336
rect 8527 7296 8944 7324
rect 8527 7293 8539 7296
rect 8481 7287 8539 7293
rect 8938 7284 8944 7296
rect 8996 7284 9002 7336
rect 10336 7324 10364 7355
rect 15194 7352 15200 7364
rect 15252 7352 15258 7404
rect 10962 7324 10968 7336
rect 10336 7296 10968 7324
rect 10962 7284 10968 7296
rect 11020 7284 11026 7336
rect 11882 7284 11888 7336
rect 11940 7324 11946 7336
rect 12161 7327 12219 7333
rect 12161 7324 12173 7327
rect 11940 7296 12173 7324
rect 11940 7284 11946 7296
rect 12161 7293 12173 7296
rect 12207 7293 12219 7327
rect 12161 7287 12219 7293
rect 14642 7284 14648 7336
rect 14700 7324 14706 7336
rect 16945 7327 17003 7333
rect 16945 7324 16957 7327
rect 14700 7296 16957 7324
rect 14700 7284 14706 7296
rect 16945 7293 16957 7296
rect 16991 7293 17003 7327
rect 16945 7287 17003 7293
rect 1578 7216 1584 7268
rect 1636 7256 1642 7268
rect 2317 7259 2375 7265
rect 2317 7256 2329 7259
rect 1636 7228 2329 7256
rect 1636 7216 1642 7228
rect 2317 7225 2329 7228
rect 2363 7225 2375 7259
rect 3418 7256 3424 7268
rect 3379 7228 3424 7256
rect 2317 7219 2375 7225
rect 3418 7216 3424 7228
rect 3476 7216 3482 7268
rect 3970 7216 3976 7268
rect 4028 7256 4034 7268
rect 6273 7259 6331 7265
rect 4028 7228 5948 7256
rect 4028 7216 4034 7228
rect 2409 7191 2467 7197
rect 2409 7157 2421 7191
rect 2455 7188 2467 7191
rect 3053 7191 3111 7197
rect 3053 7188 3065 7191
rect 2455 7160 3065 7188
rect 2455 7157 2467 7160
rect 2409 7151 2467 7157
rect 3053 7157 3065 7160
rect 3099 7157 3111 7191
rect 3510 7188 3516 7200
rect 3471 7160 3516 7188
rect 3053 7151 3111 7157
rect 3510 7148 3516 7160
rect 3568 7148 3574 7200
rect 4706 7148 4712 7200
rect 4764 7188 4770 7200
rect 5813 7191 5871 7197
rect 5813 7188 5825 7191
rect 4764 7160 5825 7188
rect 4764 7148 4770 7160
rect 5813 7157 5825 7160
rect 5859 7157 5871 7191
rect 5920 7188 5948 7228
rect 6273 7225 6285 7259
rect 6319 7256 6331 7259
rect 7098 7256 7104 7268
rect 6319 7228 7104 7256
rect 6319 7225 6331 7228
rect 6273 7219 6331 7225
rect 7098 7216 7104 7228
rect 7156 7216 7162 7268
rect 7190 7216 7196 7268
rect 7248 7256 7254 7268
rect 9214 7256 9220 7268
rect 7248 7228 7293 7256
rect 7392 7228 9220 7256
rect 7248 7216 7254 7228
rect 7392 7188 7420 7228
rect 9214 7216 9220 7228
rect 9272 7216 9278 7268
rect 10042 7216 10048 7268
rect 10100 7256 10106 7268
rect 10226 7256 10232 7268
rect 10100 7228 10232 7256
rect 10100 7216 10106 7228
rect 10226 7216 10232 7228
rect 10284 7216 10290 7268
rect 10594 7265 10600 7268
rect 10588 7256 10600 7265
rect 10555 7228 10600 7256
rect 10588 7219 10600 7228
rect 10594 7216 10600 7219
rect 10652 7216 10658 7268
rect 14090 7216 14096 7268
rect 14148 7256 14154 7268
rect 14737 7259 14795 7265
rect 14737 7256 14749 7259
rect 14148 7228 14749 7256
rect 14148 7216 14154 7228
rect 14737 7225 14749 7228
rect 14783 7225 14795 7259
rect 14737 7219 14795 7225
rect 17221 7259 17279 7265
rect 17221 7225 17233 7259
rect 17267 7256 17279 7259
rect 17770 7256 17776 7268
rect 17267 7228 17776 7256
rect 17267 7225 17279 7228
rect 17221 7219 17279 7225
rect 17770 7216 17776 7228
rect 17828 7216 17834 7268
rect 5920 7160 7420 7188
rect 8573 7191 8631 7197
rect 5813 7151 5871 7157
rect 8573 7157 8585 7191
rect 8619 7188 8631 7191
rect 10502 7188 10508 7200
rect 8619 7160 10508 7188
rect 8619 7157 8631 7160
rect 8573 7151 8631 7157
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 11698 7188 11704 7200
rect 11659 7160 11704 7188
rect 11698 7148 11704 7160
rect 11756 7148 11762 7200
rect 11882 7148 11888 7200
rect 11940 7188 11946 7200
rect 11977 7191 12035 7197
rect 11977 7188 11989 7191
rect 11940 7160 11989 7188
rect 11940 7148 11946 7160
rect 11977 7157 11989 7160
rect 12023 7157 12035 7191
rect 11977 7151 12035 7157
rect 12434 7148 12440 7200
rect 12492 7188 12498 7200
rect 13633 7191 13691 7197
rect 12492 7160 12537 7188
rect 12492 7148 12498 7160
rect 13633 7157 13645 7191
rect 13679 7188 13691 7191
rect 14182 7188 14188 7200
rect 13679 7160 14188 7188
rect 13679 7157 13691 7160
rect 13633 7151 13691 7157
rect 14182 7148 14188 7160
rect 14240 7148 14246 7200
rect 14366 7148 14372 7200
rect 14424 7188 14430 7200
rect 14645 7191 14703 7197
rect 14645 7188 14657 7191
rect 14424 7160 14657 7188
rect 14424 7148 14430 7160
rect 14645 7157 14657 7160
rect 14691 7157 14703 7191
rect 15562 7188 15568 7200
rect 15523 7160 15568 7188
rect 14645 7151 14703 7157
rect 15562 7148 15568 7160
rect 15620 7148 15626 7200
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 1302 6944 1308 6996
rect 1360 6984 1366 6996
rect 1360 6956 2820 6984
rect 1360 6944 1366 6956
rect 2682 6916 2688 6928
rect 1964 6888 2688 6916
rect 1854 6740 1860 6792
rect 1912 6780 1918 6792
rect 1964 6789 1992 6888
rect 2682 6876 2688 6888
rect 2740 6876 2746 6928
rect 2792 6916 2820 6956
rect 3418 6944 3424 6996
rect 3476 6984 3482 6996
rect 4065 6987 4123 6993
rect 4065 6984 4077 6987
rect 3476 6956 4077 6984
rect 3476 6944 3482 6956
rect 4065 6953 4077 6956
rect 4111 6953 4123 6987
rect 4065 6947 4123 6953
rect 6178 6944 6184 6996
rect 6236 6984 6242 6996
rect 8478 6984 8484 6996
rect 6236 6956 8484 6984
rect 6236 6944 6242 6956
rect 8478 6944 8484 6956
rect 8536 6944 8542 6996
rect 9674 6944 9680 6996
rect 9732 6984 9738 6996
rect 10505 6987 10563 6993
rect 10505 6984 10517 6987
rect 9732 6956 10517 6984
rect 9732 6944 9738 6956
rect 10505 6953 10517 6956
rect 10551 6984 10563 6987
rect 10870 6984 10876 6996
rect 10551 6956 10876 6984
rect 10551 6953 10563 6956
rect 10505 6947 10563 6953
rect 10870 6944 10876 6956
rect 10928 6944 10934 6996
rect 12437 6987 12495 6993
rect 12437 6984 12449 6987
rect 10980 6956 12449 6984
rect 3234 6916 3240 6928
rect 2792 6888 3240 6916
rect 3234 6876 3240 6888
rect 3292 6916 3298 6928
rect 4433 6919 4491 6925
rect 4433 6916 4445 6919
rect 3292 6888 4445 6916
rect 3292 6876 3298 6888
rect 4433 6885 4445 6888
rect 4479 6885 4491 6919
rect 4433 6879 4491 6885
rect 5350 6876 5356 6928
rect 5408 6916 5414 6928
rect 10413 6919 10471 6925
rect 10413 6916 10425 6919
rect 5408 6888 10425 6916
rect 5408 6876 5414 6888
rect 10413 6885 10425 6888
rect 10459 6885 10471 6919
rect 10980 6916 11008 6956
rect 12437 6953 12449 6956
rect 12483 6953 12495 6987
rect 12437 6947 12495 6953
rect 10413 6879 10471 6885
rect 10520 6888 11008 6916
rect 11324 6919 11382 6925
rect 2216 6851 2274 6857
rect 2216 6817 2228 6851
rect 2262 6848 2274 6851
rect 2498 6848 2504 6860
rect 2262 6820 2504 6848
rect 2262 6817 2274 6820
rect 2216 6811 2274 6817
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 2958 6808 2964 6860
rect 3016 6848 3022 6860
rect 3326 6848 3332 6860
rect 3016 6820 3332 6848
rect 3016 6808 3022 6820
rect 3326 6808 3332 6820
rect 3384 6848 3390 6860
rect 4525 6851 4583 6857
rect 4525 6848 4537 6851
rect 3384 6820 4537 6848
rect 3384 6808 3390 6820
rect 4525 6817 4537 6820
rect 4571 6817 4583 6851
rect 4525 6811 4583 6817
rect 5166 6808 5172 6860
rect 5224 6848 5230 6860
rect 5626 6857 5632 6860
rect 5261 6851 5319 6857
rect 5261 6848 5273 6851
rect 5224 6820 5273 6848
rect 5224 6808 5230 6820
rect 5261 6817 5273 6820
rect 5307 6817 5319 6851
rect 5620 6848 5632 6857
rect 5587 6820 5632 6848
rect 5261 6811 5319 6817
rect 5620 6811 5632 6820
rect 5626 6808 5632 6811
rect 5684 6808 5690 6860
rect 7282 6857 7288 6860
rect 7265 6851 7288 6857
rect 7265 6848 7277 6851
rect 6748 6820 7277 6848
rect 1949 6783 2007 6789
rect 1949 6780 1961 6783
rect 1912 6752 1961 6780
rect 1912 6740 1918 6752
rect 1949 6749 1961 6752
rect 1995 6749 2007 6783
rect 4706 6780 4712 6792
rect 4667 6752 4712 6780
rect 1949 6743 2007 6749
rect 4706 6740 4712 6752
rect 4764 6740 4770 6792
rect 5360 6783 5418 6789
rect 5360 6780 5372 6783
rect 5092 6752 5372 6780
rect 3329 6715 3387 6721
rect 3329 6681 3341 6715
rect 3375 6712 3387 6715
rect 4798 6712 4804 6724
rect 3375 6684 4804 6712
rect 3375 6681 3387 6684
rect 3329 6675 3387 6681
rect 4798 6672 4804 6684
rect 4856 6672 4862 6724
rect 5092 6656 5120 6752
rect 5360 6749 5372 6752
rect 5406 6749 5418 6783
rect 5360 6743 5418 6749
rect 6748 6721 6776 6820
rect 7265 6817 7277 6820
rect 7340 6848 7346 6860
rect 7340 6820 7413 6848
rect 7265 6811 7288 6817
rect 7282 6808 7288 6811
rect 7340 6808 7346 6820
rect 10226 6808 10232 6860
rect 10284 6848 10290 6860
rect 10520 6848 10548 6888
rect 11324 6885 11336 6919
rect 11370 6916 11382 6919
rect 11698 6916 11704 6928
rect 11370 6888 11704 6916
rect 11370 6885 11382 6888
rect 11324 6879 11382 6885
rect 11698 6876 11704 6888
rect 11756 6876 11762 6928
rect 12710 6876 12716 6928
rect 12768 6916 12774 6928
rect 12768 6888 13124 6916
rect 12768 6876 12774 6888
rect 10284 6820 10548 6848
rect 10284 6808 10290 6820
rect 10594 6808 10600 6860
rect 10652 6848 10658 6860
rect 13096 6857 13124 6888
rect 13081 6851 13139 6857
rect 10652 6820 13032 6848
rect 10652 6808 10658 6820
rect 10704 6789 10732 6820
rect 7009 6783 7067 6789
rect 7009 6749 7021 6783
rect 7055 6749 7067 6783
rect 7009 6743 7067 6749
rect 10689 6783 10747 6789
rect 10689 6749 10701 6783
rect 10735 6749 10747 6783
rect 10689 6743 10747 6749
rect 6733 6715 6791 6721
rect 6733 6681 6745 6715
rect 6779 6681 6791 6715
rect 6733 6675 6791 6681
rect 5074 6644 5080 6656
rect 5035 6616 5080 6644
rect 5074 6604 5080 6616
rect 5132 6604 5138 6656
rect 7024 6644 7052 6743
rect 10962 6740 10968 6792
rect 11020 6780 11026 6792
rect 11057 6783 11115 6789
rect 11057 6780 11069 6783
rect 11020 6752 11069 6780
rect 11020 6740 11026 6752
rect 11057 6749 11069 6752
rect 11103 6749 11115 6783
rect 11057 6743 11115 6749
rect 8294 6644 8300 6656
rect 7024 6616 8300 6644
rect 8294 6604 8300 6616
rect 8352 6604 8358 6656
rect 8389 6647 8447 6653
rect 8389 6613 8401 6647
rect 8435 6644 8447 6647
rect 8478 6644 8484 6656
rect 8435 6616 8484 6644
rect 8435 6613 8447 6616
rect 8389 6607 8447 6613
rect 8478 6604 8484 6616
rect 8536 6604 8542 6656
rect 10045 6647 10103 6653
rect 10045 6613 10057 6647
rect 10091 6644 10103 6647
rect 11790 6644 11796 6656
rect 10091 6616 11796 6644
rect 10091 6613 10103 6616
rect 10045 6607 10103 6613
rect 11790 6604 11796 6616
rect 11848 6604 11854 6656
rect 13004 6644 13032 6820
rect 13081 6817 13093 6851
rect 13127 6817 13139 6851
rect 13081 6811 13139 6817
rect 13348 6851 13406 6857
rect 13348 6817 13360 6851
rect 13394 6848 13406 6851
rect 13906 6848 13912 6860
rect 13394 6820 13912 6848
rect 13394 6817 13406 6820
rect 13348 6811 13406 6817
rect 13906 6808 13912 6820
rect 13964 6808 13970 6860
rect 15194 6808 15200 6860
rect 15252 6848 15258 6860
rect 15556 6851 15614 6857
rect 15556 6848 15568 6851
rect 15252 6820 15568 6848
rect 15252 6808 15258 6820
rect 15556 6817 15568 6820
rect 15602 6848 15614 6851
rect 16022 6848 16028 6860
rect 15602 6820 16028 6848
rect 15602 6817 15614 6820
rect 15556 6811 15614 6817
rect 16022 6808 16028 6820
rect 16080 6808 16086 6860
rect 16942 6848 16948 6860
rect 16903 6820 16948 6848
rect 16942 6808 16948 6820
rect 17000 6808 17006 6860
rect 15010 6740 15016 6792
rect 15068 6780 15074 6792
rect 15289 6783 15347 6789
rect 15289 6780 15301 6783
rect 15068 6752 15301 6780
rect 15068 6740 15074 6752
rect 15289 6749 15301 6752
rect 15335 6749 15347 6783
rect 15289 6743 15347 6749
rect 17221 6783 17279 6789
rect 17221 6749 17233 6783
rect 17267 6780 17279 6783
rect 17678 6780 17684 6792
rect 17267 6752 17684 6780
rect 17267 6749 17279 6752
rect 17221 6743 17279 6749
rect 17678 6740 17684 6752
rect 17736 6740 17742 6792
rect 14461 6647 14519 6653
rect 14461 6644 14473 6647
rect 13004 6616 14473 6644
rect 14461 6613 14473 6616
rect 14507 6613 14519 6647
rect 14461 6607 14519 6613
rect 15930 6604 15936 6656
rect 15988 6644 15994 6656
rect 16669 6647 16727 6653
rect 16669 6644 16681 6647
rect 15988 6616 16681 6644
rect 15988 6604 15994 6616
rect 16669 6613 16681 6616
rect 16715 6613 16727 6647
rect 16669 6607 16727 6613
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 2498 6400 2504 6452
rect 2556 6440 2562 6452
rect 2777 6443 2835 6449
rect 2777 6440 2789 6443
rect 2556 6412 2789 6440
rect 2556 6400 2562 6412
rect 2777 6409 2789 6412
rect 2823 6409 2835 6443
rect 2777 6403 2835 6409
rect 4062 6400 4068 6452
rect 4120 6440 4126 6452
rect 4120 6412 9168 6440
rect 4120 6400 4126 6412
rect 5626 6332 5632 6384
rect 5684 6372 5690 6384
rect 9140 6372 9168 6412
rect 9766 6400 9772 6452
rect 9824 6449 9830 6452
rect 9824 6440 9834 6449
rect 13906 6440 13912 6452
rect 9824 6412 9869 6440
rect 13867 6412 13912 6440
rect 9824 6403 9834 6412
rect 9824 6400 9830 6403
rect 13906 6400 13912 6412
rect 13964 6400 13970 6452
rect 15197 6443 15255 6449
rect 15197 6409 15209 6443
rect 15243 6440 15255 6443
rect 16942 6440 16948 6452
rect 15243 6412 16948 6440
rect 15243 6409 15255 6412
rect 15197 6403 15255 6409
rect 16942 6400 16948 6412
rect 17000 6400 17006 6452
rect 9677 6375 9735 6381
rect 9677 6372 9689 6375
rect 5684 6344 7512 6372
rect 9140 6344 9689 6372
rect 5684 6332 5690 6344
rect 4890 6264 4896 6316
rect 4948 6304 4954 6316
rect 5810 6304 5816 6316
rect 4948 6276 5816 6304
rect 4948 6264 4954 6276
rect 5810 6264 5816 6276
rect 5868 6264 5874 6316
rect 6288 6313 6316 6344
rect 6273 6307 6331 6313
rect 6273 6273 6285 6307
rect 6319 6273 6331 6307
rect 6273 6267 6331 6273
rect 7282 6264 7288 6316
rect 7340 6304 7346 6316
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 7340 6276 7389 6304
rect 7340 6264 7346 6276
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 7377 6267 7435 6273
rect 1394 6236 1400 6248
rect 1355 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6236 1458 6248
rect 3697 6239 3755 6245
rect 3697 6236 3709 6239
rect 1452 6208 3709 6236
rect 1452 6196 1458 6208
rect 3697 6205 3709 6208
rect 3743 6205 3755 6239
rect 3697 6199 3755 6205
rect 3964 6239 4022 6245
rect 3964 6205 3976 6239
rect 4010 6236 4022 6239
rect 4706 6236 4712 6248
rect 4010 6208 4712 6236
rect 4010 6205 4022 6208
rect 3964 6199 4022 6205
rect 1664 6171 1722 6177
rect 1664 6137 1676 6171
rect 1710 6168 1722 6171
rect 2774 6168 2780 6180
rect 1710 6140 2780 6168
rect 1710 6137 1722 6140
rect 1664 6131 1722 6137
rect 2774 6128 2780 6140
rect 2832 6168 2838 6180
rect 3712 6168 3740 6199
rect 4706 6196 4712 6208
rect 4764 6196 4770 6248
rect 5074 6196 5080 6248
rect 5132 6196 5138 6248
rect 5718 6196 5724 6248
rect 5776 6236 5782 6248
rect 5997 6239 6055 6245
rect 5997 6236 6009 6239
rect 5776 6208 6009 6236
rect 5776 6196 5782 6208
rect 5997 6205 6009 6208
rect 6043 6205 6055 6239
rect 5997 6199 6055 6205
rect 7098 6196 7104 6248
rect 7156 6236 7162 6248
rect 7193 6239 7251 6245
rect 7193 6236 7205 6239
rect 7156 6208 7205 6236
rect 7156 6196 7162 6208
rect 7193 6205 7205 6208
rect 7239 6205 7251 6239
rect 7193 6199 7251 6205
rect 5092 6168 5120 6196
rect 7285 6171 7343 6177
rect 7285 6168 7297 6171
rect 2832 6140 3648 6168
rect 3712 6140 5120 6168
rect 5644 6140 7297 6168
rect 2832 6128 2838 6140
rect 3620 6112 3648 6140
rect 1946 6060 1952 6112
rect 2004 6100 2010 6112
rect 3053 6103 3111 6109
rect 3053 6100 3065 6103
rect 2004 6072 3065 6100
rect 2004 6060 2010 6072
rect 3053 6069 3065 6072
rect 3099 6069 3111 6103
rect 3053 6063 3111 6069
rect 3602 6060 3608 6112
rect 3660 6100 3666 6112
rect 5644 6109 5672 6140
rect 7285 6137 7297 6140
rect 7331 6137 7343 6171
rect 7484 6168 7512 6344
rect 9677 6341 9689 6344
rect 9723 6341 9735 6375
rect 9858 6372 9864 6384
rect 9819 6344 9864 6372
rect 9677 6335 9735 6341
rect 9858 6332 9864 6344
rect 9916 6332 9922 6384
rect 9214 6264 9220 6316
rect 9272 6304 9278 6316
rect 9766 6304 9772 6316
rect 9272 6276 9772 6304
rect 9272 6264 9278 6276
rect 9766 6264 9772 6276
rect 9824 6264 9830 6316
rect 10413 6307 10471 6313
rect 10413 6304 10425 6307
rect 10051 6276 10425 6304
rect 8205 6239 8263 6245
rect 8205 6205 8217 6239
rect 8251 6236 8263 6239
rect 8294 6236 8300 6248
rect 8251 6208 8300 6236
rect 8251 6205 8263 6208
rect 8205 6199 8263 6205
rect 8294 6196 8300 6208
rect 8352 6196 8358 6248
rect 8478 6245 8484 6248
rect 8472 6236 8484 6245
rect 8391 6208 8484 6236
rect 8472 6199 8484 6208
rect 8536 6236 8542 6248
rect 10051 6236 10079 6276
rect 10413 6273 10425 6276
rect 10459 6273 10471 6307
rect 11698 6304 11704 6316
rect 11659 6276 11704 6304
rect 10413 6267 10471 6273
rect 11698 6264 11704 6276
rect 11756 6264 11762 6316
rect 13538 6264 13544 6316
rect 13596 6304 13602 6316
rect 14737 6307 14795 6313
rect 14737 6304 14749 6307
rect 13596 6276 14749 6304
rect 13596 6264 13602 6276
rect 14737 6273 14749 6276
rect 14783 6273 14795 6307
rect 15746 6304 15752 6316
rect 15707 6276 15752 6304
rect 14737 6267 14795 6273
rect 15746 6264 15752 6276
rect 15804 6264 15810 6316
rect 8536 6208 10079 6236
rect 8478 6196 8484 6199
rect 8536 6196 8542 6208
rect 10134 6196 10140 6248
rect 10192 6236 10198 6248
rect 10229 6239 10287 6245
rect 10229 6236 10241 6239
rect 10192 6208 10241 6236
rect 10192 6196 10198 6208
rect 10229 6205 10241 6208
rect 10275 6205 10287 6239
rect 10229 6199 10287 6205
rect 11517 6239 11575 6245
rect 11517 6205 11529 6239
rect 11563 6236 11575 6239
rect 12342 6236 12348 6248
rect 11563 6208 12348 6236
rect 11563 6205 11575 6208
rect 11517 6199 11575 6205
rect 12342 6196 12348 6208
rect 12400 6196 12406 6248
rect 12529 6239 12587 6245
rect 12529 6205 12541 6239
rect 12575 6205 12587 6239
rect 14550 6236 14556 6248
rect 14511 6208 14556 6236
rect 12529 6199 12587 6205
rect 12544 6168 12572 6199
rect 14550 6196 14556 6208
rect 14608 6196 14614 6248
rect 15562 6236 15568 6248
rect 15523 6208 15568 6236
rect 15562 6196 15568 6208
rect 15620 6196 15626 6248
rect 15654 6196 15660 6248
rect 15712 6236 15718 6248
rect 15712 6208 15757 6236
rect 15712 6196 15718 6208
rect 15930 6196 15936 6248
rect 15988 6236 15994 6248
rect 16301 6239 16359 6245
rect 16301 6236 16313 6239
rect 15988 6208 16313 6236
rect 15988 6196 15994 6208
rect 16301 6205 16313 6208
rect 16347 6205 16359 6239
rect 16301 6199 16359 6205
rect 12618 6168 12624 6180
rect 7484 6140 9904 6168
rect 12544 6140 12624 6168
rect 7285 6131 7343 6137
rect 5077 6103 5135 6109
rect 5077 6100 5089 6103
rect 3660 6072 5089 6100
rect 3660 6060 3666 6072
rect 5077 6069 5089 6072
rect 5123 6069 5135 6103
rect 5077 6063 5135 6069
rect 5629 6103 5687 6109
rect 5629 6069 5641 6103
rect 5675 6069 5687 6103
rect 5629 6063 5687 6069
rect 5718 6060 5724 6112
rect 5776 6100 5782 6112
rect 6089 6103 6147 6109
rect 6089 6100 6101 6103
rect 5776 6072 6101 6100
rect 5776 6060 5782 6072
rect 6089 6069 6101 6072
rect 6135 6069 6147 6103
rect 6822 6100 6828 6112
rect 6783 6072 6828 6100
rect 6089 6063 6147 6069
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 9585 6103 9643 6109
rect 9585 6069 9597 6103
rect 9631 6100 9643 6103
rect 9677 6103 9735 6109
rect 9677 6100 9689 6103
rect 9631 6072 9689 6100
rect 9631 6069 9643 6072
rect 9585 6063 9643 6069
rect 9677 6069 9689 6072
rect 9723 6100 9735 6103
rect 9766 6100 9772 6112
rect 9723 6072 9772 6100
rect 9723 6069 9735 6072
rect 9677 6063 9735 6069
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 9876 6100 9904 6140
rect 12618 6128 12624 6140
rect 12676 6128 12682 6180
rect 12796 6171 12854 6177
rect 12796 6137 12808 6171
rect 12842 6168 12854 6171
rect 13538 6168 13544 6180
rect 12842 6140 13544 6168
rect 12842 6137 12854 6140
rect 12796 6131 12854 6137
rect 13538 6128 13544 6140
rect 13596 6128 13602 6180
rect 14090 6128 14096 6180
rect 14148 6168 14154 6180
rect 14645 6171 14703 6177
rect 14645 6168 14657 6171
rect 14148 6140 14657 6168
rect 14148 6128 14154 6140
rect 14645 6137 14657 6140
rect 14691 6137 14703 6171
rect 14645 6131 14703 6137
rect 16568 6171 16626 6177
rect 16568 6137 16580 6171
rect 16614 6168 16626 6171
rect 17402 6168 17408 6180
rect 16614 6140 17408 6168
rect 16614 6137 16626 6140
rect 16568 6131 16626 6137
rect 17402 6128 17408 6140
rect 17460 6128 17466 6180
rect 10226 6100 10232 6112
rect 9876 6072 10232 6100
rect 10226 6060 10232 6072
rect 10284 6060 10290 6112
rect 10321 6103 10379 6109
rect 10321 6069 10333 6103
rect 10367 6100 10379 6103
rect 10410 6100 10416 6112
rect 10367 6072 10416 6100
rect 10367 6069 10379 6072
rect 10321 6063 10379 6069
rect 10410 6060 10416 6072
rect 10468 6060 10474 6112
rect 11146 6100 11152 6112
rect 11107 6072 11152 6100
rect 11146 6060 11152 6072
rect 11204 6060 11210 6112
rect 11609 6103 11667 6109
rect 11609 6069 11621 6103
rect 11655 6100 11667 6103
rect 11790 6100 11796 6112
rect 11655 6072 11796 6100
rect 11655 6069 11667 6072
rect 11609 6063 11667 6069
rect 11790 6060 11796 6072
rect 11848 6060 11854 6112
rect 14185 6103 14243 6109
rect 14185 6069 14197 6103
rect 14231 6100 14243 6103
rect 14274 6100 14280 6112
rect 14231 6072 14280 6100
rect 14231 6069 14243 6072
rect 14185 6063 14243 6069
rect 14274 6060 14280 6072
rect 14332 6060 14338 6112
rect 16022 6060 16028 6112
rect 16080 6100 16086 6112
rect 17681 6103 17739 6109
rect 17681 6100 17693 6103
rect 16080 6072 17693 6100
rect 16080 6060 16086 6072
rect 17681 6069 17693 6072
rect 17727 6069 17739 6103
rect 17681 6063 17739 6069
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 1578 5896 1584 5908
rect 1539 5868 1584 5896
rect 1578 5856 1584 5868
rect 1636 5856 1642 5908
rect 1946 5896 1952 5908
rect 1907 5868 1952 5896
rect 1946 5856 1952 5868
rect 2004 5856 2010 5908
rect 3510 5856 3516 5908
rect 3568 5896 3574 5908
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 3568 5868 4077 5896
rect 3568 5856 3574 5868
rect 4065 5865 4077 5868
rect 4111 5865 4123 5899
rect 4065 5859 4123 5865
rect 4154 5856 4160 5908
rect 4212 5896 4218 5908
rect 8386 5896 8392 5908
rect 4212 5868 8392 5896
rect 4212 5856 4218 5868
rect 8386 5856 8392 5868
rect 8444 5856 8450 5908
rect 9033 5899 9091 5905
rect 9033 5865 9045 5899
rect 9079 5896 9091 5899
rect 9858 5896 9864 5908
rect 9079 5868 9864 5896
rect 9079 5865 9091 5868
rect 9033 5859 9091 5865
rect 9858 5856 9864 5868
rect 9916 5856 9922 5908
rect 10229 5899 10287 5905
rect 10229 5865 10241 5899
rect 10275 5896 10287 5899
rect 12069 5899 12127 5905
rect 12069 5896 12081 5899
rect 10275 5868 12081 5896
rect 10275 5865 10287 5868
rect 10229 5859 10287 5865
rect 12069 5865 12081 5868
rect 12115 5865 12127 5899
rect 12069 5859 12127 5865
rect 5626 5828 5632 5840
rect 2976 5800 5632 5828
rect 2976 5772 3004 5800
rect 5626 5788 5632 5800
rect 5684 5788 5690 5840
rect 7282 5828 7288 5840
rect 5736 5800 7288 5828
rect 2958 5760 2964 5772
rect 2056 5732 2636 5760
rect 2919 5732 2964 5760
rect 1670 5652 1676 5704
rect 1728 5692 1734 5704
rect 2056 5701 2084 5732
rect 2041 5695 2099 5701
rect 2041 5692 2053 5695
rect 1728 5664 2053 5692
rect 1728 5652 1734 5664
rect 2041 5661 2053 5664
rect 2087 5661 2099 5695
rect 2041 5655 2099 5661
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5661 2283 5695
rect 2608 5692 2636 5732
rect 2958 5720 2964 5732
rect 3016 5720 3022 5772
rect 3602 5720 3608 5772
rect 3660 5760 3666 5772
rect 4433 5763 4491 5769
rect 4433 5760 4445 5763
rect 3660 5732 4445 5760
rect 3660 5720 3666 5732
rect 4433 5729 4445 5732
rect 4479 5760 4491 5763
rect 4890 5760 4896 5772
rect 4479 5732 4896 5760
rect 4479 5729 4491 5732
rect 4433 5723 4491 5729
rect 4890 5720 4896 5732
rect 4948 5720 4954 5772
rect 5074 5720 5080 5772
rect 5132 5760 5138 5772
rect 5537 5763 5595 5769
rect 5537 5760 5549 5763
rect 5132 5732 5549 5760
rect 5132 5720 5138 5732
rect 5537 5729 5549 5732
rect 5583 5760 5595 5763
rect 5736 5760 5764 5800
rect 7282 5788 7288 5800
rect 7340 5788 7346 5840
rect 7392 5800 7696 5828
rect 5810 5769 5816 5772
rect 5583 5732 5764 5760
rect 5583 5729 5595 5732
rect 5537 5723 5595 5729
rect 5804 5723 5816 5769
rect 5868 5760 5874 5772
rect 5868 5732 5904 5760
rect 5810 5720 5816 5723
rect 5868 5720 5874 5732
rect 6546 5720 6552 5772
rect 6604 5760 6610 5772
rect 7392 5760 7420 5800
rect 7558 5760 7564 5772
rect 6604 5732 7420 5760
rect 7519 5732 7564 5760
rect 6604 5720 6610 5732
rect 7558 5720 7564 5732
rect 7616 5720 7622 5772
rect 7668 5760 7696 5800
rect 8294 5788 8300 5840
rect 8352 5828 8358 5840
rect 8754 5828 8760 5840
rect 8352 5800 8760 5828
rect 8352 5788 8358 5800
rect 8754 5788 8760 5800
rect 8812 5828 8818 5840
rect 10244 5828 10272 5859
rect 12158 5856 12164 5908
rect 12216 5896 12222 5908
rect 14090 5896 14096 5908
rect 12216 5868 14096 5896
rect 12216 5856 12222 5868
rect 14090 5856 14096 5868
rect 14148 5856 14154 5908
rect 14274 5896 14280 5908
rect 14235 5868 14280 5896
rect 14274 5856 14280 5868
rect 14332 5856 14338 5908
rect 17402 5896 17408 5908
rect 17363 5868 17408 5896
rect 17402 5856 17408 5868
rect 17460 5856 17466 5908
rect 11882 5828 11888 5840
rect 8812 5800 10272 5828
rect 8812 5788 8818 5800
rect 8846 5760 8852 5772
rect 7668 5732 8852 5760
rect 8846 5720 8852 5732
rect 8904 5720 8910 5772
rect 8941 5763 8999 5769
rect 8941 5729 8953 5763
rect 8987 5760 8999 5763
rect 9677 5763 9735 5769
rect 9677 5760 9689 5763
rect 8987 5732 9689 5760
rect 8987 5729 8999 5732
rect 8941 5723 8999 5729
rect 9677 5729 9689 5732
rect 9723 5729 9735 5763
rect 9677 5723 9735 5729
rect 3050 5692 3056 5704
rect 2608 5664 2912 5692
rect 3011 5664 3056 5692
rect 2225 5655 2283 5661
rect 2240 5624 2268 5655
rect 2774 5624 2780 5636
rect 2240 5596 2780 5624
rect 2774 5584 2780 5596
rect 2832 5584 2838 5636
rect 2884 5624 2912 5664
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5692 3295 5695
rect 3510 5692 3516 5704
rect 3283 5664 3516 5692
rect 3283 5661 3295 5664
rect 3237 5655 3295 5661
rect 3510 5652 3516 5664
rect 3568 5652 3574 5704
rect 3694 5652 3700 5704
rect 3752 5692 3758 5704
rect 4525 5695 4583 5701
rect 4525 5692 4537 5695
rect 3752 5664 4537 5692
rect 3752 5652 3758 5664
rect 4525 5661 4537 5664
rect 4571 5661 4583 5695
rect 4706 5692 4712 5704
rect 4667 5664 4712 5692
rect 4525 5655 4583 5661
rect 4706 5652 4712 5664
rect 4764 5652 4770 5704
rect 7650 5692 7656 5704
rect 7611 5664 7656 5692
rect 7650 5652 7656 5664
rect 7708 5652 7714 5704
rect 7837 5695 7895 5701
rect 7837 5661 7849 5695
rect 7883 5692 7895 5695
rect 8294 5692 8300 5704
rect 7883 5664 8300 5692
rect 7883 5661 7895 5664
rect 7837 5655 7895 5661
rect 8294 5652 8300 5664
rect 8352 5652 8358 5704
rect 9217 5695 9275 5701
rect 9217 5661 9229 5695
rect 9263 5692 9275 5695
rect 9766 5692 9772 5704
rect 9263 5664 9772 5692
rect 9263 5661 9275 5664
rect 9217 5655 9275 5661
rect 9766 5652 9772 5664
rect 9824 5652 9830 5704
rect 10244 5692 10272 5800
rect 10428 5800 11888 5828
rect 10428 5769 10456 5800
rect 11882 5788 11888 5800
rect 11940 5828 11946 5840
rect 14182 5828 14188 5840
rect 11940 5800 13492 5828
rect 14143 5800 14188 5828
rect 11940 5788 11946 5800
rect 10778 5769 10784 5772
rect 10413 5763 10471 5769
rect 10413 5729 10425 5763
rect 10459 5729 10471 5763
rect 10772 5760 10784 5769
rect 10739 5732 10784 5760
rect 10413 5723 10471 5729
rect 10772 5723 10784 5732
rect 10778 5720 10784 5723
rect 10836 5720 10842 5772
rect 12428 5763 12486 5769
rect 12428 5760 12440 5763
rect 11900 5732 12440 5760
rect 10505 5695 10563 5701
rect 10505 5692 10517 5695
rect 10244 5664 10517 5692
rect 10505 5661 10517 5664
rect 10551 5661 10563 5695
rect 10505 5655 10563 5661
rect 3142 5624 3148 5636
rect 2884 5596 3148 5624
rect 3142 5584 3148 5596
rect 3200 5584 3206 5636
rect 6822 5584 6828 5636
rect 6880 5624 6886 5636
rect 11900 5633 11928 5732
rect 12428 5729 12440 5732
rect 12474 5760 12486 5763
rect 12986 5760 12992 5772
rect 12474 5732 12992 5760
rect 12474 5729 12486 5732
rect 12428 5723 12486 5729
rect 12986 5720 12992 5732
rect 13044 5720 13050 5772
rect 13464 5760 13492 5800
rect 14182 5788 14188 5800
rect 14240 5788 14246 5840
rect 16292 5831 16350 5837
rect 16292 5797 16304 5831
rect 16338 5828 16350 5831
rect 16482 5828 16488 5840
rect 16338 5800 16488 5828
rect 16338 5797 16350 5800
rect 16292 5791 16350 5797
rect 16482 5788 16488 5800
rect 16540 5788 16546 5840
rect 15013 5763 15071 5769
rect 15013 5760 15025 5763
rect 13464 5732 15025 5760
rect 15013 5729 15025 5732
rect 15059 5729 15071 5763
rect 15013 5723 15071 5729
rect 15289 5763 15347 5769
rect 15289 5729 15301 5763
rect 15335 5729 15347 5763
rect 17678 5760 17684 5772
rect 17639 5732 17684 5760
rect 15289 5723 15347 5729
rect 12069 5695 12127 5701
rect 12069 5661 12081 5695
rect 12115 5692 12127 5695
rect 12161 5695 12219 5701
rect 12161 5692 12173 5695
rect 12115 5664 12173 5692
rect 12115 5661 12127 5664
rect 12069 5655 12127 5661
rect 12161 5661 12173 5664
rect 12207 5661 12219 5695
rect 12161 5655 12219 5661
rect 13906 5652 13912 5704
rect 13964 5692 13970 5704
rect 14369 5695 14427 5701
rect 14369 5692 14381 5695
rect 13964 5664 14381 5692
rect 13964 5652 13970 5664
rect 14369 5661 14381 5664
rect 14415 5661 14427 5695
rect 14369 5655 14427 5661
rect 11885 5627 11943 5633
rect 6880 5596 10364 5624
rect 6880 5584 6886 5596
rect 2590 5556 2596 5568
rect 2551 5528 2596 5556
rect 2590 5516 2596 5528
rect 2648 5516 2654 5568
rect 4062 5516 4068 5568
rect 4120 5556 4126 5568
rect 6270 5556 6276 5568
rect 4120 5528 6276 5556
rect 4120 5516 4126 5528
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 6917 5559 6975 5565
rect 6917 5525 6929 5559
rect 6963 5556 6975 5559
rect 7098 5556 7104 5568
rect 6963 5528 7104 5556
rect 6963 5525 6975 5528
rect 6917 5519 6975 5525
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 7193 5559 7251 5565
rect 7193 5525 7205 5559
rect 7239 5556 7251 5559
rect 8478 5556 8484 5568
rect 7239 5528 8484 5556
rect 7239 5525 7251 5528
rect 7193 5519 7251 5525
rect 8478 5516 8484 5528
rect 8536 5516 8542 5568
rect 8573 5559 8631 5565
rect 8573 5525 8585 5559
rect 8619 5556 8631 5559
rect 10226 5556 10232 5568
rect 8619 5528 10232 5556
rect 8619 5525 8631 5528
rect 8573 5519 8631 5525
rect 10226 5516 10232 5528
rect 10284 5516 10290 5568
rect 10336 5556 10364 5596
rect 11885 5593 11897 5627
rect 11931 5593 11943 5627
rect 15304 5624 15332 5723
rect 17678 5720 17684 5732
rect 17736 5720 17742 5772
rect 15470 5692 15476 5704
rect 15431 5664 15476 5692
rect 15470 5652 15476 5664
rect 15528 5652 15534 5704
rect 15930 5692 15936 5704
rect 15571 5664 15936 5692
rect 11885 5587 11943 5593
rect 13280 5596 15332 5624
rect 13280 5556 13308 5596
rect 13538 5556 13544 5568
rect 10336 5528 13308 5556
rect 13499 5528 13544 5556
rect 13538 5516 13544 5528
rect 13596 5516 13602 5568
rect 13814 5556 13820 5568
rect 13775 5528 13820 5556
rect 13814 5516 13820 5528
rect 13872 5516 13878 5568
rect 14829 5559 14887 5565
rect 14829 5525 14841 5559
rect 14875 5556 14887 5559
rect 15010 5556 15016 5568
rect 14875 5528 15016 5556
rect 14875 5525 14887 5528
rect 14829 5519 14887 5525
rect 15010 5516 15016 5528
rect 15068 5556 15074 5568
rect 15571 5556 15599 5664
rect 15930 5652 15936 5664
rect 15988 5692 15994 5704
rect 16025 5695 16083 5701
rect 16025 5692 16037 5695
rect 15988 5664 16037 5692
rect 15988 5652 15994 5664
rect 16025 5661 16037 5664
rect 16071 5661 16083 5695
rect 16025 5655 16083 5661
rect 15068 5528 15599 5556
rect 17865 5559 17923 5565
rect 15068 5516 15074 5528
rect 17865 5525 17877 5559
rect 17911 5556 17923 5559
rect 17954 5556 17960 5568
rect 17911 5528 17960 5556
rect 17911 5525 17923 5528
rect 17865 5519 17923 5525
rect 17954 5516 17960 5528
rect 18012 5516 18018 5568
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 2866 5312 2872 5364
rect 2924 5352 2930 5364
rect 5626 5352 5632 5364
rect 2924 5324 5632 5352
rect 2924 5312 2930 5324
rect 5626 5312 5632 5324
rect 5684 5312 5690 5364
rect 5721 5355 5779 5361
rect 5721 5321 5733 5355
rect 5767 5352 5779 5355
rect 7650 5352 7656 5364
rect 5767 5324 7656 5352
rect 5767 5321 5779 5324
rect 5721 5315 5779 5321
rect 7650 5312 7656 5324
rect 7708 5312 7714 5364
rect 8294 5352 8300 5364
rect 8255 5324 8300 5352
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 8662 5312 8668 5364
rect 8720 5352 8726 5364
rect 8720 5324 11836 5352
rect 8720 5312 8726 5324
rect 3050 5244 3056 5296
rect 3108 5284 3114 5296
rect 6546 5284 6552 5296
rect 3108 5256 6552 5284
rect 3108 5244 3114 5256
rect 6546 5244 6552 5256
rect 6604 5244 6610 5296
rect 2409 5219 2467 5225
rect 2409 5185 2421 5219
rect 2455 5216 2467 5219
rect 2682 5216 2688 5228
rect 2455 5188 2688 5216
rect 2455 5185 2467 5188
rect 2409 5179 2467 5185
rect 2682 5176 2688 5188
rect 2740 5176 2746 5228
rect 3329 5219 3387 5225
rect 3329 5185 3341 5219
rect 3375 5216 3387 5219
rect 3510 5216 3516 5228
rect 3375 5188 3516 5216
rect 3375 5185 3387 5188
rect 3329 5179 3387 5185
rect 3510 5176 3516 5188
rect 3568 5176 3574 5228
rect 4706 5216 4712 5228
rect 4667 5188 4712 5216
rect 4706 5176 4712 5188
rect 4764 5176 4770 5228
rect 6365 5219 6423 5225
rect 6365 5185 6377 5219
rect 6411 5185 6423 5219
rect 8312 5216 8340 5312
rect 10137 5287 10195 5293
rect 10137 5253 10149 5287
rect 10183 5253 10195 5287
rect 10137 5247 10195 5253
rect 10413 5287 10471 5293
rect 10413 5253 10425 5287
rect 10459 5284 10471 5287
rect 11808 5284 11836 5324
rect 11882 5312 11888 5364
rect 11940 5352 11946 5364
rect 11940 5324 15792 5352
rect 11940 5312 11946 5324
rect 12161 5287 12219 5293
rect 12161 5284 12173 5287
rect 10459 5256 11744 5284
rect 11808 5256 12173 5284
rect 10459 5253 10471 5256
rect 10413 5247 10471 5253
rect 10152 5216 10180 5247
rect 10778 5216 10784 5228
rect 8312 5188 8892 5216
rect 10152 5188 10784 5216
rect 6365 5179 6423 5185
rect 2774 5108 2780 5160
rect 2832 5148 2838 5160
rect 3145 5151 3203 5157
rect 3145 5148 3157 5151
rect 2832 5120 3157 5148
rect 2832 5108 2838 5120
rect 3145 5117 3157 5120
rect 3191 5117 3203 5151
rect 3145 5111 3203 5117
rect 3418 5108 3424 5160
rect 3476 5148 3482 5160
rect 4525 5151 4583 5157
rect 4525 5148 4537 5151
rect 3476 5120 4537 5148
rect 3476 5108 3482 5120
rect 4525 5117 4537 5120
rect 4571 5117 4583 5151
rect 4525 5111 4583 5117
rect 5626 5108 5632 5160
rect 5684 5148 5690 5160
rect 6181 5151 6239 5157
rect 6181 5148 6193 5151
rect 5684 5120 6193 5148
rect 5684 5108 5690 5120
rect 6181 5117 6193 5120
rect 6227 5117 6239 5151
rect 6181 5111 6239 5117
rect 6380 5080 6408 5179
rect 6917 5151 6975 5157
rect 6917 5117 6929 5151
rect 6963 5148 6975 5151
rect 8754 5148 8760 5160
rect 6963 5120 7328 5148
rect 8715 5120 8760 5148
rect 6963 5117 6975 5120
rect 6917 5111 6975 5117
rect 7300 5092 7328 5120
rect 8754 5108 8760 5120
rect 8812 5108 8818 5160
rect 8864 5148 8892 5188
rect 10778 5176 10784 5188
rect 10836 5216 10842 5228
rect 10965 5219 11023 5225
rect 10965 5216 10977 5219
rect 10836 5188 10977 5216
rect 10836 5176 10842 5188
rect 10965 5185 10977 5188
rect 11011 5185 11023 5219
rect 11716 5216 11744 5256
rect 12161 5253 12173 5256
rect 12207 5253 12219 5287
rect 12161 5247 12219 5253
rect 12986 5216 12992 5228
rect 11716 5188 12388 5216
rect 12947 5188 12992 5216
rect 10965 5179 11023 5185
rect 9013 5151 9071 5157
rect 9013 5148 9025 5151
rect 8864 5120 9025 5148
rect 9013 5117 9025 5120
rect 9059 5117 9071 5151
rect 9013 5111 9071 5117
rect 10226 5108 10232 5160
rect 10284 5148 10290 5160
rect 11609 5151 11667 5157
rect 11609 5148 11621 5151
rect 10284 5120 11621 5148
rect 10284 5108 10290 5120
rect 11609 5117 11621 5120
rect 11655 5117 11667 5151
rect 12360 5148 12388 5188
rect 12986 5176 12992 5188
rect 13044 5176 13050 5228
rect 15764 5225 15792 5324
rect 15749 5219 15807 5225
rect 15749 5185 15761 5219
rect 15795 5185 15807 5219
rect 15749 5179 15807 5185
rect 15933 5219 15991 5225
rect 15933 5185 15945 5219
rect 15979 5216 15991 5219
rect 16482 5216 16488 5228
rect 15979 5188 16488 5216
rect 15979 5185 15991 5188
rect 15933 5179 15991 5185
rect 16482 5176 16488 5188
rect 16540 5176 16546 5228
rect 16945 5219 17003 5225
rect 16945 5185 16957 5219
rect 16991 5216 17003 5219
rect 17402 5216 17408 5228
rect 16991 5188 17408 5216
rect 16991 5185 17003 5188
rect 16945 5179 17003 5185
rect 17402 5176 17408 5188
rect 17460 5176 17466 5228
rect 12897 5151 12955 5157
rect 12897 5148 12909 5151
rect 12360 5120 12909 5148
rect 11609 5111 11667 5117
rect 12897 5117 12909 5120
rect 12943 5117 12955 5151
rect 12897 5111 12955 5117
rect 13633 5151 13691 5157
rect 13633 5117 13645 5151
rect 13679 5148 13691 5151
rect 13814 5148 13820 5160
rect 13679 5120 13820 5148
rect 13679 5117 13691 5120
rect 13633 5111 13691 5117
rect 13814 5108 13820 5120
rect 13872 5108 13878 5160
rect 14366 5148 14372 5160
rect 14327 5120 14372 5148
rect 14366 5108 14372 5120
rect 14424 5108 14430 5160
rect 15657 5151 15715 5157
rect 15657 5117 15669 5151
rect 15703 5148 15715 5151
rect 17313 5151 17371 5157
rect 17313 5148 17325 5151
rect 15703 5120 17325 5148
rect 15703 5117 15715 5120
rect 15657 5111 15715 5117
rect 17313 5117 17325 5120
rect 17359 5117 17371 5151
rect 17313 5111 17371 5117
rect 7190 5089 7196 5092
rect 7184 5080 7196 5089
rect 6380 5052 7196 5080
rect 7184 5043 7196 5052
rect 7190 5040 7196 5043
rect 7248 5040 7254 5092
rect 7282 5040 7288 5092
rect 7340 5040 7346 5092
rect 8386 5040 8392 5092
rect 8444 5080 8450 5092
rect 10781 5083 10839 5089
rect 10781 5080 10793 5083
rect 8444 5052 10793 5080
rect 8444 5040 8450 5052
rect 10781 5049 10793 5052
rect 10827 5049 10839 5083
rect 11882 5080 11888 5092
rect 11843 5052 11888 5080
rect 10781 5043 10839 5049
rect 11882 5040 11888 5052
rect 11940 5040 11946 5092
rect 12161 5083 12219 5089
rect 12161 5049 12173 5083
rect 12207 5080 12219 5083
rect 13262 5080 13268 5092
rect 12207 5052 13268 5080
rect 12207 5049 12219 5052
rect 12161 5043 12219 5049
rect 13262 5040 13268 5052
rect 13320 5040 13326 5092
rect 13906 5080 13912 5092
rect 13867 5052 13912 5080
rect 13906 5040 13912 5052
rect 13964 5040 13970 5092
rect 14550 5040 14556 5092
rect 14608 5080 14614 5092
rect 14645 5083 14703 5089
rect 14645 5080 14657 5083
rect 14608 5052 14657 5080
rect 14608 5040 14614 5052
rect 14645 5049 14657 5052
rect 14691 5049 14703 5083
rect 16669 5083 16727 5089
rect 16669 5080 16681 5083
rect 14645 5043 14703 5049
rect 15304 5052 16681 5080
rect 1762 5012 1768 5024
rect 1723 4984 1768 5012
rect 1762 4972 1768 4984
rect 1820 4972 1826 5024
rect 2130 5012 2136 5024
rect 2091 4984 2136 5012
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 2222 4972 2228 5024
rect 2280 5012 2286 5024
rect 2280 4984 2325 5012
rect 2280 4972 2286 4984
rect 2498 4972 2504 5024
rect 2556 5012 2562 5024
rect 2777 5015 2835 5021
rect 2777 5012 2789 5015
rect 2556 4984 2789 5012
rect 2556 4972 2562 4984
rect 2777 4981 2789 4984
rect 2823 4981 2835 5015
rect 2777 4975 2835 4981
rect 3237 5015 3295 5021
rect 3237 4981 3249 5015
rect 3283 5012 3295 5015
rect 3786 5012 3792 5024
rect 3283 4984 3792 5012
rect 3283 4981 3295 4984
rect 3237 4975 3295 4981
rect 3786 4972 3792 4984
rect 3844 4972 3850 5024
rect 4154 5012 4160 5024
rect 4115 4984 4160 5012
rect 4154 4972 4160 4984
rect 4212 4972 4218 5024
rect 4617 5015 4675 5021
rect 4617 4981 4629 5015
rect 4663 5012 4675 5015
rect 5166 5012 5172 5024
rect 4663 4984 5172 5012
rect 4663 4981 4675 4984
rect 4617 4975 4675 4981
rect 5166 4972 5172 4984
rect 5224 4972 5230 5024
rect 6086 5012 6092 5024
rect 6047 4984 6092 5012
rect 6086 4972 6092 4984
rect 6144 4972 6150 5024
rect 6730 4972 6736 5024
rect 6788 5012 6794 5024
rect 10594 5012 10600 5024
rect 6788 4984 10600 5012
rect 6788 4972 6794 4984
rect 10594 4972 10600 4984
rect 10652 4972 10658 5024
rect 10870 5012 10876 5024
rect 10831 4984 10876 5012
rect 10870 4972 10876 4984
rect 10928 4972 10934 5024
rect 11698 4972 11704 5024
rect 11756 5012 11762 5024
rect 12437 5015 12495 5021
rect 12437 5012 12449 5015
rect 11756 4984 12449 5012
rect 11756 4972 11762 4984
rect 12437 4981 12449 4984
rect 12483 4981 12495 5015
rect 12802 5012 12808 5024
rect 12763 4984 12808 5012
rect 12437 4975 12495 4981
rect 12802 4972 12808 4984
rect 12860 4972 12866 5024
rect 15304 5021 15332 5052
rect 16669 5049 16681 5052
rect 16715 5049 16727 5083
rect 16669 5043 16727 5049
rect 15289 5015 15347 5021
rect 15289 4981 15301 5015
rect 15335 4981 15347 5015
rect 15289 4975 15347 4981
rect 16301 5015 16359 5021
rect 16301 4981 16313 5015
rect 16347 5012 16359 5015
rect 16574 5012 16580 5024
rect 16347 4984 16580 5012
rect 16347 4981 16359 4984
rect 16301 4975 16359 4981
rect 16574 4972 16580 4984
rect 16632 4972 16638 5024
rect 16758 5012 16764 5024
rect 16719 4984 16764 5012
rect 16758 4972 16764 4984
rect 16816 4972 16822 5024
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 2130 4768 2136 4820
rect 2188 4808 2194 4820
rect 3421 4811 3479 4817
rect 3421 4808 3433 4811
rect 2188 4780 3433 4808
rect 2188 4768 2194 4780
rect 3421 4777 3433 4780
rect 3467 4777 3479 4811
rect 3421 4771 3479 4777
rect 4154 4768 4160 4820
rect 4212 4808 4218 4820
rect 4985 4811 5043 4817
rect 4985 4808 4997 4811
rect 4212 4780 4997 4808
rect 4212 4768 4218 4780
rect 4985 4777 4997 4780
rect 5031 4777 5043 4811
rect 4985 4771 5043 4777
rect 5537 4811 5595 4817
rect 5537 4777 5549 4811
rect 5583 4808 5595 4811
rect 5626 4808 5632 4820
rect 5583 4780 5632 4808
rect 5583 4777 5595 4780
rect 5537 4771 5595 4777
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 5718 4768 5724 4820
rect 5776 4808 5782 4820
rect 5905 4811 5963 4817
rect 5905 4808 5917 4811
rect 5776 4780 5917 4808
rect 5776 4768 5782 4780
rect 5905 4777 5917 4780
rect 5951 4777 5963 4811
rect 5905 4771 5963 4777
rect 6549 4811 6607 4817
rect 6549 4777 6561 4811
rect 6595 4808 6607 4811
rect 7558 4808 7564 4820
rect 6595 4780 7564 4808
rect 6595 4777 6607 4780
rect 6549 4771 6607 4777
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 8478 4768 8484 4820
rect 8536 4808 8542 4820
rect 12253 4811 12311 4817
rect 12253 4808 12265 4811
rect 8536 4780 12265 4808
rect 8536 4768 8542 4780
rect 12253 4777 12265 4780
rect 12299 4777 12311 4811
rect 12253 4771 12311 4777
rect 13262 4768 13268 4820
rect 13320 4808 13326 4820
rect 14093 4811 14151 4817
rect 14093 4808 14105 4811
rect 13320 4780 14105 4808
rect 13320 4768 13326 4780
rect 14093 4777 14105 4780
rect 14139 4777 14151 4811
rect 14093 4771 14151 4777
rect 2032 4743 2090 4749
rect 2032 4709 2044 4743
rect 2078 4740 2090 4743
rect 2682 4740 2688 4752
rect 2078 4712 2688 4740
rect 2078 4709 2090 4712
rect 2032 4703 2090 4709
rect 2682 4700 2688 4712
rect 2740 4700 2746 4752
rect 4062 4700 4068 4752
rect 4120 4740 4126 4752
rect 8205 4743 8263 4749
rect 8205 4740 8217 4743
rect 4120 4712 8217 4740
rect 4120 4700 4126 4712
rect 8205 4709 8217 4712
rect 8251 4709 8263 4743
rect 8205 4703 8263 4709
rect 9766 4700 9772 4752
rect 9824 4740 9830 4752
rect 9922 4743 9980 4749
rect 9922 4740 9934 4743
rect 9824 4712 9934 4740
rect 9824 4700 9830 4712
rect 9922 4709 9934 4712
rect 9968 4709 9980 4743
rect 9922 4703 9980 4709
rect 10594 4700 10600 4752
rect 10652 4740 10658 4752
rect 14185 4743 14243 4749
rect 14185 4740 14197 4743
rect 10652 4712 14197 4740
rect 10652 4700 10658 4712
rect 14185 4709 14197 4712
rect 14231 4709 14243 4743
rect 18224 4743 18282 4749
rect 14185 4703 14243 4709
rect 15396 4712 18000 4740
rect 1394 4632 1400 4684
rect 1452 4672 1458 4684
rect 1765 4675 1823 4681
rect 1765 4672 1777 4675
rect 1452 4644 1777 4672
rect 1452 4632 1458 4644
rect 1765 4641 1777 4644
rect 1811 4641 1823 4675
rect 4890 4672 4896 4684
rect 4851 4644 4896 4672
rect 1765 4635 1823 4641
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 5997 4675 6055 4681
rect 5997 4641 6009 4675
rect 6043 4672 6055 4675
rect 6546 4672 6552 4684
rect 6043 4644 6552 4672
rect 6043 4641 6055 4644
rect 5997 4635 6055 4641
rect 6546 4632 6552 4644
rect 6604 4632 6610 4684
rect 6914 4672 6920 4684
rect 6875 4644 6920 4672
rect 6914 4632 6920 4644
rect 6972 4632 6978 4684
rect 7650 4632 7656 4684
rect 7708 4672 7714 4684
rect 11698 4672 11704 4684
rect 7708 4644 10916 4672
rect 11659 4644 11704 4672
rect 7708 4632 7714 4644
rect 5169 4607 5227 4613
rect 5169 4573 5181 4607
rect 5215 4604 5227 4607
rect 5350 4604 5356 4616
rect 5215 4576 5356 4604
rect 5215 4573 5227 4576
rect 5169 4567 5227 4573
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 6181 4607 6239 4613
rect 6181 4573 6193 4607
rect 6227 4573 6239 4607
rect 6181 4567 6239 4573
rect 5810 4496 5816 4548
rect 5868 4536 5874 4548
rect 6196 4536 6224 4567
rect 6270 4564 6276 4616
rect 6328 4604 6334 4616
rect 7009 4607 7067 4613
rect 7009 4604 7021 4607
rect 6328 4576 7021 4604
rect 6328 4564 6334 4576
rect 7009 4573 7021 4576
rect 7055 4573 7067 4607
rect 7190 4604 7196 4616
rect 7151 4576 7196 4604
rect 7009 4567 7067 4573
rect 7190 4564 7196 4576
rect 7248 4564 7254 4616
rect 8297 4607 8355 4613
rect 8297 4604 8309 4607
rect 7392 4576 8309 4604
rect 5868 4508 6224 4536
rect 5868 4496 5874 4508
rect 2406 4428 2412 4480
rect 2464 4468 2470 4480
rect 3145 4471 3203 4477
rect 3145 4468 3157 4471
rect 2464 4440 3157 4468
rect 2464 4428 2470 4440
rect 3145 4437 3157 4440
rect 3191 4468 3203 4471
rect 3234 4468 3240 4480
rect 3191 4440 3240 4468
rect 3191 4437 3203 4440
rect 3145 4431 3203 4437
rect 3234 4428 3240 4440
rect 3292 4428 3298 4480
rect 4525 4471 4583 4477
rect 4525 4437 4537 4471
rect 4571 4468 4583 4471
rect 5074 4468 5080 4480
rect 4571 4440 5080 4468
rect 4571 4437 4583 4440
rect 4525 4431 4583 4437
rect 5074 4428 5080 4440
rect 5132 4428 5138 4480
rect 5166 4428 5172 4480
rect 5224 4468 5230 4480
rect 7392 4468 7420 4576
rect 8297 4573 8309 4576
rect 8343 4604 8355 4607
rect 8386 4604 8392 4616
rect 8343 4576 8392 4604
rect 8343 4573 8355 4576
rect 8297 4567 8355 4573
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 8496 4613 8524 4644
rect 8481 4607 8539 4613
rect 8481 4573 8493 4607
rect 8527 4573 8539 4607
rect 8481 4567 8539 4573
rect 8754 4564 8760 4616
rect 8812 4604 8818 4616
rect 9582 4604 9588 4616
rect 8812 4576 9588 4604
rect 8812 4564 8818 4576
rect 9582 4564 9588 4576
rect 9640 4604 9646 4616
rect 9677 4607 9735 4613
rect 9677 4604 9689 4607
rect 9640 4576 9689 4604
rect 9640 4564 9646 4576
rect 9677 4573 9689 4576
rect 9723 4573 9735 4607
rect 9677 4567 9735 4573
rect 10888 4548 10916 4644
rect 11698 4632 11704 4644
rect 11756 4632 11762 4684
rect 12253 4675 12311 4681
rect 12253 4641 12265 4675
rect 12299 4672 12311 4675
rect 12437 4675 12495 4681
rect 12437 4672 12449 4675
rect 12299 4644 12449 4672
rect 12299 4641 12311 4644
rect 12253 4635 12311 4641
rect 12437 4641 12449 4644
rect 12483 4641 12495 4675
rect 12437 4635 12495 4641
rect 11977 4607 12035 4613
rect 11977 4573 11989 4607
rect 12023 4604 12035 4607
rect 12526 4604 12532 4616
rect 12023 4576 12532 4604
rect 12023 4573 12035 4576
rect 11977 4567 12035 4573
rect 12526 4564 12532 4576
rect 12584 4564 12590 4616
rect 12713 4607 12771 4613
rect 12713 4573 12725 4607
rect 12759 4604 12771 4607
rect 13722 4604 13728 4616
rect 12759 4576 13728 4604
rect 12759 4573 12771 4576
rect 12713 4567 12771 4573
rect 13722 4564 13728 4576
rect 13780 4564 13786 4616
rect 14366 4604 14372 4616
rect 14327 4576 14372 4604
rect 14366 4564 14372 4576
rect 14424 4564 14430 4616
rect 14642 4564 14648 4616
rect 14700 4604 14706 4616
rect 15010 4604 15016 4616
rect 14700 4576 15016 4604
rect 14700 4564 14706 4576
rect 15010 4564 15016 4576
rect 15068 4604 15074 4616
rect 15396 4613 15424 4712
rect 15648 4675 15706 4681
rect 15648 4641 15660 4675
rect 15694 4672 15706 4675
rect 16114 4672 16120 4684
rect 15694 4644 16120 4672
rect 15694 4641 15706 4644
rect 15648 4635 15706 4641
rect 16114 4632 16120 4644
rect 16172 4632 16178 4684
rect 16574 4632 16580 4684
rect 16632 4672 16638 4684
rect 17972 4681 18000 4712
rect 18224 4709 18236 4743
rect 18270 4740 18282 4743
rect 18598 4740 18604 4752
rect 18270 4712 18604 4740
rect 18270 4709 18282 4712
rect 18224 4703 18282 4709
rect 18598 4700 18604 4712
rect 18656 4700 18662 4752
rect 17037 4675 17095 4681
rect 17037 4672 17049 4675
rect 16632 4644 17049 4672
rect 16632 4632 16638 4644
rect 17037 4641 17049 4644
rect 17083 4641 17095 4675
rect 17037 4635 17095 4641
rect 17957 4675 18015 4681
rect 17957 4641 17969 4675
rect 18003 4641 18015 4675
rect 17957 4635 18015 4641
rect 15381 4607 15439 4613
rect 15381 4604 15393 4607
rect 15068 4576 15393 4604
rect 15068 4564 15074 4576
rect 15381 4573 15393 4576
rect 15427 4573 15439 4607
rect 17218 4604 17224 4616
rect 17179 4576 17224 4604
rect 15381 4567 15439 4573
rect 17218 4564 17224 4576
rect 17276 4564 17282 4616
rect 10870 4496 10876 4548
rect 10928 4536 10934 4548
rect 10928 4508 15424 4536
rect 10928 4496 10934 4508
rect 7834 4468 7840 4480
rect 5224 4440 7420 4468
rect 7795 4440 7840 4468
rect 5224 4428 5230 4440
rect 7834 4428 7840 4440
rect 7892 4428 7898 4480
rect 10042 4428 10048 4480
rect 10100 4468 10106 4480
rect 11057 4471 11115 4477
rect 11057 4468 11069 4471
rect 10100 4440 11069 4468
rect 10100 4428 10106 4440
rect 11057 4437 11069 4440
rect 11103 4437 11115 4471
rect 11057 4431 11115 4437
rect 13725 4471 13783 4477
rect 13725 4437 13737 4471
rect 13771 4468 13783 4471
rect 14458 4468 14464 4480
rect 13771 4440 14464 4468
rect 13771 4437 13783 4440
rect 13725 4431 13783 4437
rect 14458 4428 14464 4440
rect 14516 4428 14522 4480
rect 15396 4468 15424 4508
rect 16316 4508 16896 4536
rect 16316 4468 16344 4508
rect 15396 4440 16344 4468
rect 16482 4428 16488 4480
rect 16540 4468 16546 4480
rect 16761 4471 16819 4477
rect 16761 4468 16773 4471
rect 16540 4440 16773 4468
rect 16540 4428 16546 4440
rect 16761 4437 16773 4440
rect 16807 4437 16819 4471
rect 16868 4468 16896 4508
rect 19337 4471 19395 4477
rect 19337 4468 19349 4471
rect 16868 4440 19349 4468
rect 16761 4431 16819 4437
rect 19337 4437 19349 4440
rect 19383 4437 19395 4471
rect 19337 4431 19395 4437
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 2406 4224 2412 4276
rect 2464 4224 2470 4276
rect 4982 4264 4988 4276
rect 4632 4236 4988 4264
rect 2424 4196 2452 4224
rect 4632 4208 4660 4236
rect 4982 4224 4988 4236
rect 5040 4224 5046 4276
rect 5810 4224 5816 4276
rect 5868 4264 5874 4276
rect 6454 4264 6460 4276
rect 5868 4236 6460 4264
rect 5868 4224 5874 4236
rect 6454 4224 6460 4236
rect 6512 4224 6518 4276
rect 8202 4224 8208 4276
rect 8260 4224 8266 4276
rect 11790 4264 11796 4276
rect 9324 4236 11796 4264
rect 2424 4168 2636 4196
rect 1394 4088 1400 4140
rect 1452 4128 1458 4140
rect 2406 4128 2412 4140
rect 1452 4100 2412 4128
rect 1452 4088 1458 4100
rect 2406 4088 2412 4100
rect 2464 4128 2470 4140
rect 2608 4137 2636 4168
rect 4614 4156 4620 4208
rect 4672 4156 4678 4208
rect 8220 4196 8248 4224
rect 8220 4168 8340 4196
rect 2593 4131 2651 4137
rect 2464 4100 2544 4128
rect 2464 4088 2470 4100
rect 1762 4020 1768 4072
rect 1820 4060 1826 4072
rect 2317 4063 2375 4069
rect 2317 4060 2329 4063
rect 1820 4032 2329 4060
rect 1820 4020 1826 4032
rect 2317 4029 2329 4032
rect 2363 4029 2375 4063
rect 2516 4060 2544 4100
rect 2593 4097 2605 4131
rect 2639 4097 2651 4131
rect 4985 4131 5043 4137
rect 4985 4128 4997 4131
rect 2593 4091 2651 4097
rect 3988 4100 4997 4128
rect 3234 4069 3240 4072
rect 2961 4063 3019 4069
rect 2961 4060 2973 4063
rect 2516 4032 2973 4060
rect 2317 4023 2375 4029
rect 2961 4029 2973 4032
rect 3007 4029 3019 4063
rect 3228 4060 3240 4069
rect 3195 4032 3240 4060
rect 2961 4023 3019 4029
rect 3228 4023 3240 4032
rect 3234 4020 3240 4023
rect 3292 4020 3298 4072
rect 3786 4020 3792 4072
rect 3844 4060 3850 4072
rect 3988 4060 4016 4100
rect 4985 4097 4997 4100
rect 5031 4097 5043 4131
rect 6914 4128 6920 4140
rect 6875 4100 6920 4128
rect 4985 4091 5043 4097
rect 6914 4088 6920 4100
rect 6972 4088 6978 4140
rect 7834 4088 7840 4140
rect 7892 4128 7898 4140
rect 8312 4137 8340 4168
rect 8205 4131 8263 4137
rect 8205 4128 8217 4131
rect 7892 4100 8217 4128
rect 7892 4088 7898 4100
rect 8205 4097 8217 4100
rect 8251 4097 8263 4131
rect 8205 4091 8263 4097
rect 8297 4131 8355 4137
rect 8297 4097 8309 4131
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 8386 4088 8392 4140
rect 8444 4128 8450 4140
rect 9324 4128 9352 4236
rect 11790 4224 11796 4236
rect 11848 4224 11854 4276
rect 13262 4224 13268 4276
rect 13320 4264 13326 4276
rect 13320 4236 14320 4264
rect 13320 4224 13326 4236
rect 8444 4100 9352 4128
rect 9401 4131 9459 4137
rect 8444 4088 8450 4100
rect 9401 4097 9413 4131
rect 9447 4128 9459 4131
rect 12437 4131 12495 4137
rect 9447 4100 9904 4128
rect 9447 4097 9459 4100
rect 9401 4091 9459 4097
rect 3844 4032 4016 4060
rect 3844 4020 3850 4032
rect 4522 4020 4528 4072
rect 4580 4060 4586 4072
rect 5077 4063 5135 4069
rect 5077 4060 5089 4063
rect 4580 4032 5089 4060
rect 4580 4020 4586 4032
rect 5077 4029 5089 4032
rect 5123 4029 5135 4063
rect 5077 4023 5135 4029
rect 5184 4032 8524 4060
rect 5184 3992 5212 4032
rect 1964 3964 5212 3992
rect 1964 3933 1992 3964
rect 5258 3952 5264 4004
rect 5316 4001 5322 4004
rect 5316 3995 5380 4001
rect 5316 3961 5334 3995
rect 5368 3961 5380 3995
rect 5316 3955 5380 3961
rect 5316 3952 5322 3955
rect 5626 3952 5632 4004
rect 5684 3992 5690 4004
rect 5994 3992 6000 4004
rect 5684 3964 6000 3992
rect 5684 3952 5690 3964
rect 5994 3952 6000 3964
rect 6052 3952 6058 4004
rect 8386 3992 8392 4004
rect 7760 3964 8392 3992
rect 1949 3927 2007 3933
rect 1949 3893 1961 3927
rect 1995 3893 2007 3927
rect 1949 3887 2007 3893
rect 2038 3884 2044 3936
rect 2096 3924 2102 3936
rect 2409 3927 2467 3933
rect 2409 3924 2421 3927
rect 2096 3896 2421 3924
rect 2096 3884 2102 3896
rect 2409 3893 2421 3896
rect 2455 3893 2467 3927
rect 2409 3887 2467 3893
rect 4154 3884 4160 3936
rect 4212 3924 4218 3936
rect 4341 3927 4399 3933
rect 4341 3924 4353 3927
rect 4212 3896 4353 3924
rect 4212 3884 4218 3896
rect 4341 3893 4353 3896
rect 4387 3924 4399 3927
rect 4706 3924 4712 3936
rect 4387 3896 4712 3924
rect 4387 3893 4399 3896
rect 4341 3887 4399 3893
rect 4706 3884 4712 3896
rect 4764 3884 4770 3936
rect 4985 3927 5043 3933
rect 4985 3893 4997 3927
rect 5031 3924 5043 3927
rect 6822 3924 6828 3936
rect 5031 3896 6828 3924
rect 5031 3893 5043 3896
rect 4985 3887 5043 3893
rect 6822 3884 6828 3896
rect 6880 3884 6886 3936
rect 7760 3933 7788 3964
rect 8386 3952 8392 3964
rect 8444 3952 8450 4004
rect 8496 3992 8524 4032
rect 8662 4020 8668 4072
rect 8720 4060 8726 4072
rect 9217 4063 9275 4069
rect 9217 4060 9229 4063
rect 8720 4032 9229 4060
rect 8720 4020 8726 4032
rect 9217 4029 9229 4032
rect 9263 4029 9275 4063
rect 9217 4023 9275 4029
rect 9582 4020 9588 4072
rect 9640 4060 9646 4072
rect 9769 4063 9827 4069
rect 9769 4060 9781 4063
rect 9640 4032 9781 4060
rect 9640 4020 9646 4032
rect 9769 4029 9781 4032
rect 9815 4029 9827 4063
rect 9876 4060 9904 4100
rect 12437 4097 12449 4131
rect 12483 4128 12495 4131
rect 12802 4128 12808 4140
rect 12483 4100 12808 4128
rect 12483 4097 12495 4100
rect 12437 4091 12495 4097
rect 12802 4088 12808 4100
rect 12860 4088 12866 4140
rect 14292 4128 14320 4236
rect 14366 4224 14372 4276
rect 14424 4264 14430 4276
rect 14645 4267 14703 4273
rect 14645 4264 14657 4267
rect 14424 4236 14657 4264
rect 14424 4224 14430 4236
rect 14645 4233 14657 4236
rect 14691 4264 14703 4267
rect 14734 4264 14740 4276
rect 14691 4236 14740 4264
rect 14691 4233 14703 4236
rect 14645 4227 14703 4233
rect 14734 4224 14740 4236
rect 14792 4224 14798 4276
rect 16114 4224 16120 4276
rect 16172 4264 16178 4276
rect 16301 4267 16359 4273
rect 16301 4264 16313 4267
rect 16172 4236 16313 4264
rect 16172 4224 16178 4236
rect 16301 4233 16313 4236
rect 16347 4233 16359 4267
rect 16301 4227 16359 4233
rect 16577 4267 16635 4273
rect 16577 4233 16589 4267
rect 16623 4264 16635 4267
rect 16758 4264 16764 4276
rect 16623 4236 16764 4264
rect 16623 4233 16635 4236
rect 16577 4227 16635 4233
rect 16758 4224 16764 4236
rect 16816 4224 16822 4276
rect 16482 4156 16488 4208
rect 16540 4196 16546 4208
rect 16540 4168 17172 4196
rect 16540 4156 16546 4168
rect 14642 4128 14648 4140
rect 14292 4100 14648 4128
rect 14642 4088 14648 4100
rect 14700 4128 14706 4140
rect 17144 4137 17172 4168
rect 14921 4131 14979 4137
rect 14921 4128 14933 4131
rect 14700 4100 14933 4128
rect 14700 4088 14706 4100
rect 14921 4097 14933 4100
rect 14967 4097 14979 4131
rect 14921 4091 14979 4097
rect 17129 4131 17187 4137
rect 17129 4097 17141 4131
rect 17175 4097 17187 4131
rect 17129 4091 17187 4097
rect 10042 4069 10048 4072
rect 10036 4060 10048 4069
rect 9876 4032 10048 4060
rect 9769 4023 9827 4029
rect 10036 4023 10048 4032
rect 10042 4020 10048 4023
rect 10100 4020 10106 4072
rect 11425 4063 11483 4069
rect 11425 4029 11437 4063
rect 11471 4029 11483 4063
rect 11425 4023 11483 4029
rect 11440 3992 11468 4023
rect 12342 4020 12348 4072
rect 12400 4060 12406 4072
rect 12710 4060 12716 4072
rect 12400 4032 12716 4060
rect 12400 4020 12406 4032
rect 12710 4020 12716 4032
rect 12768 4060 12774 4072
rect 13262 4060 13268 4072
rect 12768 4032 13268 4060
rect 12768 4020 12774 4032
rect 13262 4020 13268 4032
rect 13320 4020 13326 4072
rect 15010 4020 15016 4072
rect 15068 4060 15074 4072
rect 15177 4063 15235 4069
rect 15177 4060 15189 4063
rect 15068 4032 15189 4060
rect 15068 4020 15074 4032
rect 15177 4029 15189 4032
rect 15223 4029 15235 4063
rect 15177 4023 15235 4029
rect 8496 3964 11468 3992
rect 11701 3995 11759 4001
rect 11701 3961 11713 3995
rect 11747 3992 11759 3995
rect 12618 3992 12624 4004
rect 11747 3964 12624 3992
rect 11747 3961 11759 3964
rect 11701 3955 11759 3961
rect 12618 3952 12624 3964
rect 12676 3952 12682 4004
rect 13532 3995 13590 4001
rect 13532 3961 13544 3995
rect 13578 3992 13590 3995
rect 13814 3992 13820 4004
rect 13578 3964 13820 3992
rect 13578 3961 13590 3964
rect 13532 3955 13590 3961
rect 13814 3952 13820 3964
rect 13872 3952 13878 4004
rect 16206 3992 16212 4004
rect 14200 3964 16212 3992
rect 7745 3927 7803 3933
rect 7745 3893 7757 3927
rect 7791 3893 7803 3927
rect 7745 3887 7803 3893
rect 8113 3927 8171 3933
rect 8113 3893 8125 3927
rect 8159 3924 8171 3927
rect 8294 3924 8300 3936
rect 8159 3896 8300 3924
rect 8159 3893 8171 3896
rect 8113 3887 8171 3893
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 8754 3924 8760 3936
rect 8715 3896 8760 3924
rect 8754 3884 8760 3896
rect 8812 3884 8818 3936
rect 9125 3927 9183 3933
rect 9125 3893 9137 3927
rect 9171 3924 9183 3927
rect 9306 3924 9312 3936
rect 9171 3896 9312 3924
rect 9171 3893 9183 3896
rect 9125 3887 9183 3893
rect 9306 3884 9312 3896
rect 9364 3884 9370 3936
rect 9582 3884 9588 3936
rect 9640 3924 9646 3936
rect 10594 3924 10600 3936
rect 9640 3896 10600 3924
rect 9640 3884 9646 3896
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 11146 3924 11152 3936
rect 11107 3896 11152 3924
rect 11146 3884 11152 3896
rect 11204 3884 11210 3936
rect 11238 3884 11244 3936
rect 11296 3924 11302 3936
rect 14200 3924 14228 3964
rect 16206 3952 16212 3964
rect 16264 3952 16270 4004
rect 11296 3896 14228 3924
rect 11296 3884 11302 3896
rect 14274 3884 14280 3936
rect 14332 3924 14338 3936
rect 16945 3927 17003 3933
rect 16945 3924 16957 3927
rect 14332 3896 16957 3924
rect 14332 3884 14338 3896
rect 16945 3893 16957 3896
rect 16991 3893 17003 3927
rect 16945 3887 17003 3893
rect 17034 3884 17040 3936
rect 17092 3924 17098 3936
rect 21174 3924 21180 3936
rect 17092 3896 21180 3924
rect 17092 3884 17098 3896
rect 21174 3884 21180 3896
rect 21232 3884 21238 3936
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 1026 3680 1032 3732
rect 1084 3720 1090 3732
rect 2958 3720 2964 3732
rect 1084 3692 2964 3720
rect 1084 3680 1090 3692
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 4065 3723 4123 3729
rect 4065 3689 4077 3723
rect 4111 3720 4123 3723
rect 4890 3720 4896 3732
rect 4111 3692 4896 3720
rect 4111 3689 4123 3692
rect 4065 3683 4123 3689
rect 4890 3680 4896 3692
rect 4948 3680 4954 3732
rect 6086 3680 6092 3732
rect 6144 3720 6150 3732
rect 6365 3723 6423 3729
rect 6365 3720 6377 3723
rect 6144 3692 6377 3720
rect 6144 3680 6150 3692
rect 6365 3689 6377 3692
rect 6411 3689 6423 3723
rect 6822 3720 6828 3732
rect 6735 3692 6828 3720
rect 6365 3683 6423 3689
rect 6822 3680 6828 3692
rect 6880 3720 6886 3732
rect 8662 3720 8668 3732
rect 6880 3692 8668 3720
rect 6880 3680 6886 3692
rect 8662 3680 8668 3692
rect 8720 3680 8726 3732
rect 8754 3680 8760 3732
rect 8812 3720 8818 3732
rect 10229 3723 10287 3729
rect 10229 3720 10241 3723
rect 8812 3692 10241 3720
rect 8812 3680 8818 3692
rect 10229 3689 10241 3692
rect 10275 3689 10287 3723
rect 11238 3720 11244 3732
rect 10229 3683 10287 3689
rect 10336 3692 11244 3720
rect 1946 3612 1952 3664
rect 2004 3652 2010 3664
rect 3786 3652 3792 3664
rect 2004 3624 3792 3652
rect 2004 3612 2010 3624
rect 3786 3612 3792 3624
rect 3844 3612 3850 3664
rect 3970 3612 3976 3664
rect 4028 3652 4034 3664
rect 10336 3652 10364 3692
rect 11238 3680 11244 3692
rect 11296 3680 11302 3732
rect 12161 3723 12219 3729
rect 12161 3689 12173 3723
rect 12207 3689 12219 3723
rect 13814 3720 13820 3732
rect 13775 3692 13820 3720
rect 12161 3683 12219 3689
rect 11048 3655 11106 3661
rect 11048 3652 11060 3655
rect 4028 3624 10364 3652
rect 10428 3624 11060 3652
rect 4028 3612 4034 3624
rect 1394 3544 1400 3596
rect 1452 3584 1458 3596
rect 1581 3587 1639 3593
rect 1581 3584 1593 3587
rect 1452 3556 1593 3584
rect 1452 3544 1458 3556
rect 1581 3553 1593 3556
rect 1627 3553 1639 3587
rect 1581 3547 1639 3553
rect 1848 3587 1906 3593
rect 1848 3553 1860 3587
rect 1894 3584 1906 3587
rect 3510 3584 3516 3596
rect 1894 3556 3516 3584
rect 1894 3553 1906 3556
rect 1848 3547 1906 3553
rect 3510 3544 3516 3556
rect 3568 3544 3574 3596
rect 3878 3544 3884 3596
rect 3936 3584 3942 3596
rect 4522 3584 4528 3596
rect 3936 3556 4528 3584
rect 3936 3544 3942 3556
rect 4522 3544 4528 3556
rect 4580 3544 4586 3596
rect 4792 3587 4850 3593
rect 4792 3553 4804 3587
rect 4838 3584 4850 3587
rect 5350 3584 5356 3596
rect 4838 3556 5356 3584
rect 4838 3553 4850 3556
rect 4792 3547 4850 3553
rect 5350 3544 5356 3556
rect 5408 3544 5414 3596
rect 6730 3584 6736 3596
rect 6691 3556 6736 3584
rect 6730 3544 6736 3556
rect 6788 3544 6794 3596
rect 7650 3544 7656 3596
rect 7708 3584 7714 3596
rect 8001 3587 8059 3593
rect 8001 3584 8013 3587
rect 7708 3556 8013 3584
rect 7708 3544 7714 3556
rect 8001 3553 8013 3556
rect 8047 3553 8059 3587
rect 8001 3547 8059 3553
rect 10137 3587 10195 3593
rect 10137 3553 10149 3587
rect 10183 3553 10195 3587
rect 10137 3547 10195 3553
rect 6454 3476 6460 3528
rect 6512 3516 6518 3528
rect 6917 3519 6975 3525
rect 6917 3516 6929 3519
rect 6512 3488 6929 3516
rect 6512 3476 6518 3488
rect 6917 3485 6929 3488
rect 6963 3485 6975 3519
rect 6917 3479 6975 3485
rect 7282 3476 7288 3528
rect 7340 3516 7346 3528
rect 7745 3519 7803 3525
rect 7745 3516 7757 3519
rect 7340 3488 7757 3516
rect 7340 3476 7346 3488
rect 7745 3485 7757 3488
rect 7791 3485 7803 3519
rect 7745 3479 7803 3485
rect 3970 3448 3976 3460
rect 2608 3420 3976 3448
rect 566 3340 572 3392
rect 624 3380 630 3392
rect 2608 3380 2636 3420
rect 3970 3408 3976 3420
rect 4028 3408 4034 3460
rect 10152 3448 10180 3547
rect 10428 3525 10456 3624
rect 11048 3621 11060 3624
rect 11094 3652 11106 3655
rect 11146 3652 11152 3664
rect 11094 3624 11152 3652
rect 11094 3621 11106 3624
rect 11048 3615 11106 3621
rect 11146 3612 11152 3624
rect 11204 3612 11210 3664
rect 11974 3612 11980 3664
rect 12032 3652 12038 3664
rect 12176 3652 12204 3683
rect 13814 3680 13820 3692
rect 13872 3680 13878 3732
rect 14458 3680 14464 3732
rect 14516 3720 14522 3732
rect 15841 3723 15899 3729
rect 15841 3720 15853 3723
rect 14516 3692 15853 3720
rect 14516 3680 14522 3692
rect 15841 3689 15853 3692
rect 15887 3689 15899 3723
rect 15841 3683 15899 3689
rect 12682 3655 12740 3661
rect 12682 3652 12694 3655
rect 12032 3624 12694 3652
rect 12032 3612 12038 3624
rect 12682 3621 12694 3624
rect 12728 3621 12740 3655
rect 13832 3652 13860 3680
rect 16114 3652 16120 3664
rect 13832 3624 14688 3652
rect 12682 3615 12740 3621
rect 12066 3584 12072 3596
rect 10520 3556 12072 3584
rect 10413 3519 10471 3525
rect 10413 3485 10425 3519
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 10520 3448 10548 3556
rect 12066 3544 12072 3556
rect 12124 3544 12130 3596
rect 14274 3584 14280 3596
rect 12176 3556 14280 3584
rect 10594 3476 10600 3528
rect 10652 3516 10658 3528
rect 10781 3519 10839 3525
rect 10781 3516 10793 3519
rect 10652 3488 10793 3516
rect 10652 3476 10658 3488
rect 10781 3485 10793 3488
rect 10827 3485 10839 3519
rect 10781 3479 10839 3485
rect 11790 3476 11796 3528
rect 11848 3516 11854 3528
rect 12176 3516 12204 3556
rect 14274 3544 14280 3556
rect 14332 3544 14338 3596
rect 14458 3584 14464 3596
rect 14419 3556 14464 3584
rect 14458 3544 14464 3556
rect 14516 3544 14522 3596
rect 11848 3488 12204 3516
rect 11848 3476 11854 3488
rect 12342 3476 12348 3528
rect 12400 3516 12406 3528
rect 12437 3519 12495 3525
rect 12437 3516 12449 3519
rect 12400 3488 12449 3516
rect 12400 3476 12406 3488
rect 12437 3485 12449 3488
rect 12483 3485 12495 3519
rect 12437 3479 12495 3485
rect 13446 3476 13452 3528
rect 13504 3516 13510 3528
rect 14660 3525 14688 3624
rect 15948 3624 16120 3652
rect 15746 3584 15752 3596
rect 15707 3556 15752 3584
rect 15746 3544 15752 3556
rect 15804 3544 15810 3596
rect 15948 3525 15976 3624
rect 16114 3612 16120 3624
rect 16172 3612 16178 3664
rect 16206 3612 16212 3664
rect 16264 3652 16270 3664
rect 16264 3624 20024 3652
rect 16264 3612 16270 3624
rect 16393 3587 16451 3593
rect 16393 3584 16405 3587
rect 16040 3556 16405 3584
rect 14553 3519 14611 3525
rect 14553 3516 14565 3519
rect 13504 3488 14565 3516
rect 13504 3476 13510 3488
rect 14553 3485 14565 3488
rect 14599 3485 14611 3519
rect 14553 3479 14611 3485
rect 14645 3519 14703 3525
rect 14645 3485 14657 3519
rect 14691 3485 14703 3519
rect 14645 3479 14703 3485
rect 15933 3519 15991 3525
rect 15933 3485 15945 3519
rect 15979 3485 15991 3519
rect 15933 3479 15991 3485
rect 10152 3420 10548 3448
rect 15381 3451 15439 3457
rect 15381 3417 15393 3451
rect 15427 3448 15439 3451
rect 16040 3448 16068 3556
rect 16393 3553 16405 3556
rect 16439 3553 16451 3587
rect 17218 3584 17224 3596
rect 17179 3556 17224 3584
rect 16393 3547 16451 3553
rect 17218 3544 17224 3556
rect 17276 3544 17282 3596
rect 17770 3584 17776 3596
rect 17731 3556 17776 3584
rect 17770 3544 17776 3556
rect 17828 3544 17834 3596
rect 19996 3593 20024 3624
rect 19981 3587 20039 3593
rect 19981 3553 19993 3587
rect 20027 3553 20039 3587
rect 19981 3547 20039 3553
rect 16666 3516 16672 3528
rect 16627 3488 16672 3516
rect 16666 3476 16672 3488
rect 16724 3476 16730 3528
rect 15427 3420 16068 3448
rect 15427 3417 15439 3420
rect 15381 3411 15439 3417
rect 624 3352 2636 3380
rect 624 3340 630 3352
rect 2682 3340 2688 3392
rect 2740 3380 2746 3392
rect 2961 3383 3019 3389
rect 2961 3380 2973 3383
rect 2740 3352 2973 3380
rect 2740 3340 2746 3352
rect 2961 3349 2973 3352
rect 3007 3349 3019 3383
rect 2961 3343 3019 3349
rect 3234 3340 3240 3392
rect 3292 3380 3298 3392
rect 5166 3380 5172 3392
rect 3292 3352 5172 3380
rect 3292 3340 3298 3352
rect 5166 3340 5172 3352
rect 5224 3340 5230 3392
rect 5258 3340 5264 3392
rect 5316 3380 5322 3392
rect 5905 3383 5963 3389
rect 5905 3380 5917 3383
rect 5316 3352 5917 3380
rect 5316 3340 5322 3352
rect 5905 3349 5917 3352
rect 5951 3349 5963 3383
rect 5905 3343 5963 3349
rect 5994 3340 6000 3392
rect 6052 3380 6058 3392
rect 6914 3380 6920 3392
rect 6052 3352 6920 3380
rect 6052 3340 6058 3352
rect 6914 3340 6920 3352
rect 6972 3340 6978 3392
rect 8110 3340 8116 3392
rect 8168 3380 8174 3392
rect 9125 3383 9183 3389
rect 9125 3380 9137 3383
rect 8168 3352 9137 3380
rect 8168 3340 8174 3352
rect 9125 3349 9137 3352
rect 9171 3380 9183 3383
rect 9490 3380 9496 3392
rect 9171 3352 9496 3380
rect 9171 3349 9183 3352
rect 9125 3343 9183 3349
rect 9490 3340 9496 3352
rect 9548 3340 9554 3392
rect 9769 3383 9827 3389
rect 9769 3349 9781 3383
rect 9815 3380 9827 3383
rect 13630 3380 13636 3392
rect 9815 3352 13636 3380
rect 9815 3349 9827 3352
rect 9769 3343 9827 3349
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 14093 3383 14151 3389
rect 14093 3349 14105 3383
rect 14139 3380 14151 3383
rect 15654 3380 15660 3392
rect 14139 3352 15660 3380
rect 14139 3349 14151 3352
rect 14093 3343 14151 3349
rect 15654 3340 15660 3352
rect 15712 3340 15718 3392
rect 17405 3383 17463 3389
rect 17405 3349 17417 3383
rect 17451 3380 17463 3383
rect 17678 3380 17684 3392
rect 17451 3352 17684 3380
rect 17451 3349 17463 3352
rect 17405 3343 17463 3349
rect 17678 3340 17684 3352
rect 17736 3340 17742 3392
rect 17957 3383 18015 3389
rect 17957 3349 17969 3383
rect 18003 3380 18015 3383
rect 18598 3380 18604 3392
rect 18003 3352 18604 3380
rect 18003 3349 18015 3352
rect 17957 3343 18015 3349
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 20165 3383 20223 3389
rect 20165 3349 20177 3383
rect 20211 3380 20223 3383
rect 20806 3380 20812 3392
rect 20211 3352 20812 3380
rect 20211 3349 20223 3352
rect 20165 3343 20223 3349
rect 20806 3340 20812 3352
rect 20864 3340 20870 3392
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 2406 3136 2412 3188
rect 2464 3176 2470 3188
rect 3878 3176 3884 3188
rect 2464 3148 3884 3176
rect 2464 3136 2470 3148
rect 3878 3136 3884 3148
rect 3936 3136 3942 3188
rect 11333 3179 11391 3185
rect 11333 3145 11345 3179
rect 11379 3176 11391 3179
rect 13446 3176 13452 3188
rect 11379 3148 13452 3176
rect 11379 3145 11391 3148
rect 11333 3139 11391 3145
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 15746 3136 15752 3188
rect 15804 3176 15810 3188
rect 17405 3179 17463 3185
rect 17405 3176 17417 3179
rect 15804 3148 17417 3176
rect 15804 3136 15810 3148
rect 17405 3145 17417 3148
rect 17451 3145 17463 3179
rect 17405 3139 17463 3145
rect 3510 3108 3516 3120
rect 3471 3080 3516 3108
rect 3510 3068 3516 3080
rect 3568 3068 3574 3120
rect 4890 3068 4896 3120
rect 4948 3108 4954 3120
rect 5166 3108 5172 3120
rect 4948 3080 5172 3108
rect 4948 3068 4954 3080
rect 5166 3068 5172 3080
rect 5224 3068 5230 3120
rect 5261 3111 5319 3117
rect 5261 3077 5273 3111
rect 5307 3108 5319 3111
rect 5350 3108 5356 3120
rect 5307 3080 5356 3108
rect 5307 3077 5319 3080
rect 5261 3071 5319 3077
rect 5350 3068 5356 3080
rect 5408 3068 5414 3120
rect 5994 3108 6000 3120
rect 5460 3080 6000 3108
rect 1854 3000 1860 3052
rect 1912 3040 1918 3052
rect 2133 3043 2191 3049
rect 2133 3040 2145 3043
rect 1912 3012 2145 3040
rect 1912 3000 1918 3012
rect 2133 3009 2145 3012
rect 2179 3009 2191 3043
rect 3878 3040 3884 3052
rect 3839 3012 3884 3040
rect 2133 3003 2191 3009
rect 3878 3000 3884 3012
rect 3936 3000 3942 3052
rect 4982 3000 4988 3052
rect 5040 3040 5046 3052
rect 5460 3040 5488 3080
rect 5994 3068 6000 3080
rect 6052 3068 6058 3120
rect 9766 3108 9772 3120
rect 9727 3080 9772 3108
rect 9766 3068 9772 3080
rect 9824 3068 9830 3120
rect 10318 3068 10324 3120
rect 10376 3108 10382 3120
rect 10376 3080 11008 3108
rect 10376 3068 10382 3080
rect 6273 3043 6331 3049
rect 6273 3040 6285 3043
rect 5040 3012 5488 3040
rect 5552 3012 6285 3040
rect 5040 3000 5046 3012
rect 2400 2975 2458 2981
rect 2400 2941 2412 2975
rect 2446 2972 2458 2975
rect 3786 2972 3792 2984
rect 2446 2944 3792 2972
rect 2446 2941 2458 2944
rect 2400 2935 2458 2941
rect 3786 2932 3792 2944
rect 3844 2932 3850 2984
rect 4154 2981 4160 2984
rect 4148 2972 4160 2981
rect 4067 2944 4160 2972
rect 4148 2935 4160 2944
rect 4212 2972 4218 2984
rect 5552 2972 5580 3012
rect 6273 3009 6285 3012
rect 6319 3009 6331 3043
rect 9490 3040 9496 3052
rect 9451 3012 9496 3040
rect 6273 3003 6331 3009
rect 9490 3000 9496 3012
rect 9548 3000 9554 3052
rect 9674 3000 9680 3052
rect 9732 3040 9738 3052
rect 10410 3040 10416 3052
rect 9732 3012 10416 3040
rect 9732 3000 9738 3012
rect 10410 3000 10416 3012
rect 10468 3000 10474 3052
rect 10594 3040 10600 3052
rect 10507 3012 10600 3040
rect 10594 3000 10600 3012
rect 10652 3040 10658 3052
rect 10870 3040 10876 3052
rect 10652 3012 10876 3040
rect 10652 3000 10658 3012
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 10980 3040 11008 3080
rect 12526 3068 12532 3120
rect 12584 3108 12590 3120
rect 14093 3111 14151 3117
rect 14093 3108 14105 3111
rect 12584 3080 14105 3108
rect 12584 3068 12590 3080
rect 14093 3077 14105 3080
rect 14139 3077 14151 3111
rect 14093 3071 14151 3077
rect 15930 3068 15936 3120
rect 15988 3108 15994 3120
rect 16577 3111 16635 3117
rect 16577 3108 16589 3111
rect 15988 3080 16589 3108
rect 15988 3068 15994 3080
rect 16577 3077 16589 3080
rect 16623 3077 16635 3111
rect 16577 3071 16635 3077
rect 10980 3012 11928 3040
rect 7282 2972 7288 2984
rect 4212 2944 5580 2972
rect 7243 2944 7288 2972
rect 4154 2932 4160 2935
rect 4212 2932 4218 2944
rect 7282 2932 7288 2944
rect 7340 2932 7346 2984
rect 7552 2975 7610 2981
rect 7552 2941 7564 2975
rect 7598 2972 7610 2975
rect 8110 2972 8116 2984
rect 7598 2944 8116 2972
rect 7598 2941 7610 2944
rect 7552 2935 7610 2941
rect 8110 2932 8116 2944
rect 8168 2932 8174 2984
rect 8754 2932 8760 2984
rect 8812 2972 8818 2984
rect 10321 2975 10379 2981
rect 10321 2972 10333 2975
rect 8812 2944 10333 2972
rect 8812 2932 8818 2944
rect 10321 2941 10333 2944
rect 10367 2972 10379 2975
rect 11793 2975 11851 2981
rect 11793 2972 11805 2975
rect 10367 2944 11805 2972
rect 10367 2941 10379 2944
rect 10321 2935 10379 2941
rect 11793 2941 11805 2944
rect 11839 2941 11851 2975
rect 11900 2972 11928 3012
rect 11974 3000 11980 3052
rect 12032 3040 12038 3052
rect 12032 3012 12077 3040
rect 12032 3000 12038 3012
rect 13630 3000 13636 3052
rect 13688 3040 13694 3052
rect 18417 3043 18475 3049
rect 18417 3040 18429 3043
rect 13688 3012 14964 3040
rect 13688 3000 13694 3012
rect 11900 2944 12112 2972
rect 11793 2935 11851 2941
rect 198 2864 204 2916
rect 256 2904 262 2916
rect 3050 2904 3056 2916
rect 256 2876 3056 2904
rect 256 2864 262 2876
rect 3050 2864 3056 2876
rect 3108 2864 3114 2916
rect 7374 2904 7380 2916
rect 5736 2876 7380 2904
rect 1486 2796 1492 2848
rect 1544 2836 1550 2848
rect 3418 2836 3424 2848
rect 1544 2808 3424 2836
rect 1544 2796 1550 2808
rect 3418 2796 3424 2808
rect 3476 2796 3482 2848
rect 3602 2796 3608 2848
rect 3660 2836 3666 2848
rect 3970 2836 3976 2848
rect 3660 2808 3976 2836
rect 3660 2796 3666 2808
rect 3970 2796 3976 2808
rect 4028 2796 4034 2848
rect 4062 2796 4068 2848
rect 4120 2836 4126 2848
rect 5626 2836 5632 2848
rect 4120 2808 5632 2836
rect 4120 2796 4126 2808
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 5736 2845 5764 2876
rect 7374 2864 7380 2876
rect 7432 2864 7438 2916
rect 9309 2907 9367 2913
rect 9309 2873 9321 2907
rect 9355 2904 9367 2907
rect 9355 2876 9996 2904
rect 9355 2873 9367 2876
rect 9309 2867 9367 2873
rect 5721 2839 5779 2845
rect 5721 2805 5733 2839
rect 5767 2805 5779 2839
rect 6086 2836 6092 2848
rect 6047 2808 6092 2836
rect 5721 2799 5779 2805
rect 6086 2796 6092 2808
rect 6144 2796 6150 2848
rect 6181 2839 6239 2845
rect 6181 2805 6193 2839
rect 6227 2836 6239 2839
rect 7006 2836 7012 2848
rect 6227 2808 7012 2836
rect 6227 2805 6239 2808
rect 6181 2799 6239 2805
rect 7006 2796 7012 2808
rect 7064 2796 7070 2848
rect 7282 2796 7288 2848
rect 7340 2836 7346 2848
rect 8662 2836 8668 2848
rect 7340 2808 8668 2836
rect 7340 2796 7346 2808
rect 8662 2796 8668 2808
rect 8720 2796 8726 2848
rect 8938 2836 8944 2848
rect 8899 2808 8944 2836
rect 8938 2796 8944 2808
rect 8996 2796 9002 2848
rect 9968 2845 9996 2876
rect 10502 2864 10508 2916
rect 10560 2904 10566 2916
rect 11974 2904 11980 2916
rect 10560 2876 11980 2904
rect 10560 2864 10566 2876
rect 11974 2864 11980 2876
rect 12032 2864 12038 2916
rect 12084 2904 12112 2944
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 12713 2975 12771 2981
rect 12492 2944 12537 2972
rect 12492 2932 12498 2944
rect 12713 2941 12725 2975
rect 12759 2972 12771 2975
rect 13173 2975 13231 2981
rect 13173 2972 13185 2975
rect 12759 2944 13185 2972
rect 12759 2941 12771 2944
rect 12713 2935 12771 2941
rect 13173 2941 13185 2944
rect 13219 2941 13231 2975
rect 13722 2972 13728 2984
rect 13683 2944 13728 2972
rect 13173 2935 13231 2941
rect 13722 2932 13728 2944
rect 13780 2932 13786 2984
rect 14936 2981 14964 3012
rect 15120 3012 18429 3040
rect 14093 2975 14151 2981
rect 14093 2941 14105 2975
rect 14139 2972 14151 2975
rect 14277 2975 14335 2981
rect 14277 2972 14289 2975
rect 14139 2944 14289 2972
rect 14139 2941 14151 2944
rect 14093 2935 14151 2941
rect 14277 2941 14289 2944
rect 14323 2941 14335 2975
rect 14277 2935 14335 2941
rect 14921 2975 14979 2981
rect 14921 2941 14933 2975
rect 14967 2941 14979 2975
rect 14921 2935 14979 2941
rect 15120 2904 15148 3012
rect 18417 3009 18429 3012
rect 18463 3009 18475 3043
rect 18417 3003 18475 3009
rect 15654 2972 15660 2984
rect 15615 2944 15660 2972
rect 15654 2932 15660 2944
rect 15712 2932 15718 2984
rect 16390 2972 16396 2984
rect 16351 2944 16396 2972
rect 16390 2932 16396 2944
rect 16448 2932 16454 2984
rect 16945 2975 17003 2981
rect 16945 2941 16957 2975
rect 16991 2941 17003 2975
rect 16945 2935 17003 2941
rect 17405 2975 17463 2981
rect 17405 2941 17417 2975
rect 17451 2972 17463 2975
rect 17497 2975 17555 2981
rect 17497 2972 17509 2975
rect 17451 2944 17509 2972
rect 17451 2941 17463 2944
rect 17405 2935 17463 2941
rect 17497 2941 17509 2944
rect 17543 2941 17555 2975
rect 17497 2935 17555 2941
rect 18233 2975 18291 2981
rect 18233 2941 18245 2975
rect 18279 2941 18291 2975
rect 18233 2935 18291 2941
rect 20533 2975 20591 2981
rect 20533 2941 20545 2975
rect 20579 2972 20591 2975
rect 21634 2972 21640 2984
rect 20579 2944 21640 2972
rect 20579 2941 20591 2944
rect 20533 2935 20591 2941
rect 12084 2876 15148 2904
rect 15197 2907 15255 2913
rect 15197 2873 15209 2907
rect 15243 2873 15255 2907
rect 15197 2867 15255 2873
rect 15933 2907 15991 2913
rect 15933 2873 15945 2907
rect 15979 2904 15991 2907
rect 16960 2904 16988 2935
rect 15979 2876 16988 2904
rect 18248 2904 18276 2935
rect 21634 2932 21640 2944
rect 21692 2932 21698 2984
rect 22554 2904 22560 2916
rect 18248 2876 22560 2904
rect 15979 2873 15991 2876
rect 15933 2867 15991 2873
rect 9401 2839 9459 2845
rect 9401 2805 9413 2839
rect 9447 2836 9459 2839
rect 9769 2839 9827 2845
rect 9769 2836 9781 2839
rect 9447 2808 9781 2836
rect 9447 2805 9459 2808
rect 9401 2799 9459 2805
rect 9769 2805 9781 2808
rect 9815 2805 9827 2839
rect 9769 2799 9827 2805
rect 9953 2839 10011 2845
rect 9953 2805 9965 2839
rect 9999 2805 10011 2839
rect 9953 2799 10011 2805
rect 11701 2839 11759 2845
rect 11701 2805 11713 2839
rect 11747 2836 11759 2839
rect 12250 2836 12256 2848
rect 11747 2808 12256 2836
rect 11747 2805 11759 2808
rect 11701 2799 11759 2805
rect 12250 2796 12256 2808
rect 12308 2796 12314 2848
rect 13354 2836 13360 2848
rect 13315 2808 13360 2836
rect 13354 2796 13360 2808
rect 13412 2796 13418 2848
rect 13722 2796 13728 2848
rect 13780 2836 13786 2848
rect 13909 2839 13967 2845
rect 13909 2836 13921 2839
rect 13780 2808 13921 2836
rect 13780 2796 13786 2808
rect 13909 2805 13921 2808
rect 13955 2805 13967 2839
rect 13909 2799 13967 2805
rect 14182 2796 14188 2848
rect 14240 2836 14246 2848
rect 14461 2839 14519 2845
rect 14461 2836 14473 2839
rect 14240 2808 14473 2836
rect 14240 2796 14246 2808
rect 14461 2805 14473 2808
rect 14507 2805 14519 2839
rect 15212 2836 15240 2867
rect 22554 2864 22560 2876
rect 22612 2864 22618 2916
rect 16022 2836 16028 2848
rect 15212 2808 16028 2836
rect 14461 2799 14519 2805
rect 16022 2796 16028 2808
rect 16080 2796 16086 2848
rect 16850 2796 16856 2848
rect 16908 2836 16914 2848
rect 17129 2839 17187 2845
rect 17129 2836 17141 2839
rect 16908 2808 17141 2836
rect 16908 2796 16914 2808
rect 17129 2805 17141 2808
rect 17175 2805 17187 2839
rect 17129 2799 17187 2805
rect 20717 2839 20775 2845
rect 20717 2805 20729 2839
rect 20763 2836 20775 2839
rect 22094 2836 22100 2848
rect 20763 2808 22100 2836
rect 20763 2805 20775 2808
rect 20717 2799 20775 2805
rect 22094 2796 22100 2808
rect 22152 2796 22158 2848
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 1949 2635 2007 2641
rect 1949 2601 1961 2635
rect 1995 2632 2007 2635
rect 2038 2632 2044 2644
rect 1995 2604 2044 2632
rect 1995 2601 2007 2604
rect 1949 2595 2007 2601
rect 2038 2592 2044 2604
rect 2096 2592 2102 2644
rect 2409 2635 2467 2641
rect 2409 2601 2421 2635
rect 2455 2632 2467 2635
rect 2590 2632 2596 2644
rect 2455 2604 2596 2632
rect 2455 2601 2467 2604
rect 2409 2595 2467 2601
rect 2590 2592 2596 2604
rect 2648 2592 2654 2644
rect 2961 2635 3019 2641
rect 2961 2601 2973 2635
rect 3007 2601 3019 2635
rect 3418 2632 3424 2644
rect 3379 2604 3424 2632
rect 2961 2595 3019 2601
rect 2317 2567 2375 2573
rect 2317 2533 2329 2567
rect 2363 2564 2375 2567
rect 2498 2564 2504 2576
rect 2363 2536 2504 2564
rect 2363 2533 2375 2536
rect 2317 2527 2375 2533
rect 2498 2524 2504 2536
rect 2556 2524 2562 2576
rect 2976 2564 3004 2595
rect 3418 2592 3424 2604
rect 3476 2632 3482 2644
rect 4890 2632 4896 2644
rect 3476 2604 4896 2632
rect 3476 2592 3482 2604
rect 4890 2592 4896 2604
rect 4948 2592 4954 2644
rect 5074 2592 5080 2644
rect 5132 2632 5138 2644
rect 5353 2635 5411 2641
rect 5353 2632 5365 2635
rect 5132 2604 5365 2632
rect 5132 2592 5138 2604
rect 5353 2601 5365 2604
rect 5399 2601 5411 2635
rect 5353 2595 5411 2601
rect 5445 2635 5503 2641
rect 5445 2601 5457 2635
rect 5491 2632 5503 2635
rect 6917 2635 6975 2641
rect 6917 2632 6929 2635
rect 5491 2604 6929 2632
rect 5491 2601 5503 2604
rect 5445 2595 5503 2601
rect 6917 2601 6929 2604
rect 6963 2601 6975 2635
rect 7374 2632 7380 2644
rect 7335 2604 7380 2632
rect 6917 2595 6975 2601
rect 7374 2592 7380 2604
rect 7432 2592 7438 2644
rect 8386 2632 8392 2644
rect 8347 2604 8392 2632
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 8481 2635 8539 2641
rect 8481 2601 8493 2635
rect 8527 2632 8539 2635
rect 8938 2632 8944 2644
rect 8527 2604 8944 2632
rect 8527 2601 8539 2604
rect 8481 2595 8539 2601
rect 8938 2592 8944 2604
rect 8996 2592 9002 2644
rect 9766 2632 9772 2644
rect 9727 2604 9772 2632
rect 9766 2592 9772 2604
rect 9824 2592 9830 2644
rect 10134 2592 10140 2644
rect 10192 2632 10198 2644
rect 10229 2635 10287 2641
rect 10229 2632 10241 2635
rect 10192 2604 10241 2632
rect 10192 2592 10198 2604
rect 10229 2601 10241 2604
rect 10275 2632 10287 2635
rect 10778 2632 10784 2644
rect 10275 2604 10784 2632
rect 10275 2601 10287 2604
rect 10229 2595 10287 2601
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 12066 2632 12072 2644
rect 12027 2604 12072 2632
rect 12066 2592 12072 2604
rect 12124 2592 12130 2644
rect 13725 2635 13783 2641
rect 13725 2601 13737 2635
rect 13771 2632 13783 2635
rect 14458 2632 14464 2644
rect 13771 2604 14464 2632
rect 13771 2601 13783 2604
rect 13725 2595 13783 2601
rect 14458 2592 14464 2604
rect 14516 2592 14522 2644
rect 7285 2567 7343 2573
rect 7285 2564 7297 2567
rect 2976 2536 7297 2564
rect 7285 2533 7297 2536
rect 7331 2533 7343 2567
rect 7285 2527 7343 2533
rect 8294 2524 8300 2576
rect 8352 2564 8358 2576
rect 9033 2567 9091 2573
rect 9033 2564 9045 2567
rect 8352 2536 9045 2564
rect 8352 2524 8358 2536
rect 9033 2533 9045 2536
rect 9079 2533 9091 2567
rect 12434 2564 12440 2576
rect 9033 2527 9091 2533
rect 9140 2536 12440 2564
rect 3329 2499 3387 2505
rect 3329 2496 3341 2499
rect 2332 2468 3341 2496
rect 2332 2440 2360 2468
rect 3329 2465 3341 2468
rect 3375 2496 3387 2499
rect 3418 2496 3424 2508
rect 3375 2468 3424 2496
rect 3375 2465 3387 2468
rect 3329 2459 3387 2465
rect 3418 2456 3424 2468
rect 3476 2456 3482 2508
rect 3878 2456 3884 2508
rect 3936 2496 3942 2508
rect 5166 2496 5172 2508
rect 3936 2468 5172 2496
rect 3936 2456 3942 2468
rect 5166 2456 5172 2468
rect 5224 2456 5230 2508
rect 5350 2456 5356 2508
rect 5408 2496 5414 2508
rect 9140 2496 9168 2536
rect 12434 2524 12440 2536
rect 12492 2524 12498 2576
rect 5408 2468 7512 2496
rect 5408 2456 5414 2468
rect 2314 2388 2320 2440
rect 2372 2388 2378 2440
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2428 2651 2431
rect 2682 2428 2688 2440
rect 2639 2400 2688 2428
rect 2639 2397 2651 2400
rect 2593 2391 2651 2397
rect 2682 2388 2688 2400
rect 2740 2388 2746 2440
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2428 3663 2431
rect 4154 2428 4160 2440
rect 3651 2400 4160 2428
rect 3651 2397 3663 2400
rect 3605 2391 3663 2397
rect 4154 2388 4160 2400
rect 4212 2388 4218 2440
rect 5258 2388 5264 2440
rect 5316 2428 5322 2440
rect 7484 2437 7512 2468
rect 7944 2468 9168 2496
rect 5537 2431 5595 2437
rect 5537 2428 5549 2431
rect 5316 2400 5549 2428
rect 5316 2388 5322 2400
rect 5537 2397 5549 2400
rect 5583 2397 5595 2431
rect 5537 2391 5595 2397
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2397 7527 2431
rect 7469 2391 7527 2397
rect 4985 2363 5043 2369
rect 4985 2329 4997 2363
rect 5031 2360 5043 2363
rect 7944 2360 7972 2468
rect 9674 2456 9680 2508
rect 9732 2496 9738 2508
rect 10137 2499 10195 2505
rect 10137 2496 10149 2499
rect 9732 2468 10149 2496
rect 9732 2456 9738 2468
rect 10137 2465 10149 2468
rect 10183 2465 10195 2499
rect 10137 2459 10195 2465
rect 10781 2499 10839 2505
rect 10781 2465 10793 2499
rect 10827 2465 10839 2499
rect 10781 2459 10839 2465
rect 11057 2499 11115 2505
rect 11057 2465 11069 2499
rect 11103 2496 11115 2499
rect 11517 2499 11575 2505
rect 11517 2496 11529 2499
rect 11103 2468 11529 2496
rect 11103 2465 11115 2468
rect 11057 2459 11115 2465
rect 11517 2465 11529 2468
rect 11563 2465 11575 2499
rect 12618 2496 12624 2508
rect 12579 2468 12624 2496
rect 11517 2459 11575 2465
rect 8662 2428 8668 2440
rect 8623 2400 8668 2428
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2428 10471 2431
rect 10594 2428 10600 2440
rect 10459 2400 10600 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 10594 2388 10600 2400
rect 10652 2388 10658 2440
rect 5031 2332 7972 2360
rect 8021 2363 8079 2369
rect 5031 2329 5043 2332
rect 4985 2323 5043 2329
rect 8021 2329 8033 2363
rect 8067 2360 8079 2363
rect 10796 2360 10824 2459
rect 12618 2456 12624 2468
rect 12676 2456 12682 2508
rect 13906 2456 13912 2508
rect 13964 2496 13970 2508
rect 14185 2499 14243 2505
rect 14185 2496 14197 2499
rect 13964 2468 14197 2496
rect 13964 2456 13970 2468
rect 14185 2465 14197 2468
rect 14231 2465 14243 2499
rect 14185 2459 14243 2465
rect 14550 2456 14556 2508
rect 14608 2496 14614 2508
rect 14737 2499 14795 2505
rect 14737 2496 14749 2499
rect 14608 2468 14749 2496
rect 14608 2456 14614 2468
rect 14737 2465 14749 2468
rect 14783 2465 14795 2499
rect 15470 2496 15476 2508
rect 15431 2468 15476 2496
rect 14737 2459 14795 2465
rect 15470 2456 15476 2468
rect 15528 2456 15534 2508
rect 16022 2496 16028 2508
rect 15983 2468 16028 2496
rect 16022 2456 16028 2468
rect 16080 2456 16086 2508
rect 16666 2496 16672 2508
rect 16627 2468 16672 2496
rect 16666 2456 16672 2468
rect 16724 2456 16730 2508
rect 8067 2332 10824 2360
rect 8067 2329 8079 2332
rect 8021 2323 8079 2329
rect 7006 2252 7012 2304
rect 7064 2292 7070 2304
rect 10134 2292 10140 2304
rect 7064 2264 10140 2292
rect 7064 2252 7070 2264
rect 10134 2252 10140 2264
rect 10192 2252 10198 2304
rect 11701 2295 11759 2301
rect 11701 2261 11713 2295
rect 11747 2292 11759 2295
rect 12434 2292 12440 2304
rect 11747 2264 12440 2292
rect 11747 2261 11759 2264
rect 11701 2255 11759 2261
rect 12434 2252 12440 2264
rect 12492 2252 12498 2304
rect 12805 2295 12863 2301
rect 12805 2261 12817 2295
rect 12851 2292 12863 2295
rect 12894 2292 12900 2304
rect 12851 2264 12900 2292
rect 12851 2261 12863 2264
rect 12805 2255 12863 2261
rect 12894 2252 12900 2264
rect 12952 2252 12958 2304
rect 14369 2295 14427 2301
rect 14369 2261 14381 2295
rect 14415 2292 14427 2295
rect 14642 2292 14648 2304
rect 14415 2264 14648 2292
rect 14415 2261 14427 2264
rect 14369 2255 14427 2261
rect 14642 2252 14648 2264
rect 14700 2252 14706 2304
rect 14921 2295 14979 2301
rect 14921 2261 14933 2295
rect 14967 2292 14979 2295
rect 15102 2292 15108 2304
rect 14967 2264 15108 2292
rect 14967 2261 14979 2264
rect 14921 2255 14979 2261
rect 15102 2252 15108 2264
rect 15160 2252 15166 2304
rect 15470 2252 15476 2304
rect 15528 2292 15534 2304
rect 15657 2295 15715 2301
rect 15657 2292 15669 2295
rect 15528 2264 15669 2292
rect 15528 2252 15534 2264
rect 15657 2261 15669 2264
rect 15703 2261 15715 2295
rect 15657 2255 15715 2261
rect 16209 2295 16267 2301
rect 16209 2261 16221 2295
rect 16255 2292 16267 2295
rect 16390 2292 16396 2304
rect 16255 2264 16396 2292
rect 16255 2261 16267 2264
rect 16209 2255 16267 2261
rect 16390 2252 16396 2264
rect 16448 2252 16454 2304
rect 16853 2295 16911 2301
rect 16853 2261 16865 2295
rect 16899 2292 16911 2295
rect 17310 2292 17316 2304
rect 16899 2264 17316 2292
rect 16899 2261 16911 2264
rect 16853 2255 16911 2261
rect 17310 2252 17316 2264
rect 17368 2252 17374 2304
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 2866 1844 2872 1896
rect 2924 1884 2930 1896
rect 4706 1884 4712 1896
rect 2924 1856 4712 1884
rect 2924 1844 2930 1856
rect 4706 1844 4712 1856
rect 4764 1844 4770 1896
rect 3326 892 3332 944
rect 3384 932 3390 944
rect 6178 932 6184 944
rect 3384 904 6184 932
rect 3384 892 3390 904
rect 6178 892 6184 904
rect 6236 892 6242 944
<< via1 >>
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 1952 20043 2004 20052
rect 1952 20009 1961 20043
rect 1961 20009 1995 20043
rect 1995 20009 2004 20043
rect 1952 20000 2004 20009
rect 2228 19864 2280 19916
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 3700 19456 3752 19508
rect 2044 19252 2096 19304
rect 2320 19295 2372 19304
rect 2320 19261 2329 19295
rect 2329 19261 2363 19295
rect 2363 19261 2372 19295
rect 2320 19252 2372 19261
rect 6828 19295 6880 19304
rect 6828 19261 6837 19295
rect 6837 19261 6871 19295
rect 6871 19261 6880 19295
rect 6828 19252 6880 19261
rect 2872 19184 2924 19236
rect 2780 19116 2832 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 4068 18912 4120 18964
rect 2320 18844 2372 18896
rect 6828 18844 6880 18896
rect 2228 18708 2280 18760
rect 7656 18776 7708 18828
rect 8208 18776 8260 18828
rect 8576 18708 8628 18760
rect 7196 18640 7248 18692
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 2780 18368 2832 18420
rect 3056 18411 3108 18420
rect 3056 18377 3065 18411
rect 3065 18377 3099 18411
rect 3099 18377 3108 18411
rect 3056 18368 3108 18377
rect 3608 18411 3660 18420
rect 3608 18377 3617 18411
rect 3617 18377 3651 18411
rect 3651 18377 3660 18411
rect 3608 18368 3660 18377
rect 2320 18207 2372 18216
rect 2320 18173 2329 18207
rect 2329 18173 2363 18207
rect 2363 18173 2372 18207
rect 2320 18164 2372 18173
rect 2412 18096 2464 18148
rect 8668 18164 8720 18216
rect 10416 18096 10468 18148
rect 1952 18071 2004 18080
rect 1952 18037 1961 18071
rect 1961 18037 1995 18071
rect 1995 18037 2004 18071
rect 1952 18028 2004 18037
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 1860 17867 1912 17876
rect 1860 17833 1869 17867
rect 1869 17833 1903 17867
rect 1903 17833 1912 17867
rect 1860 17824 1912 17833
rect 2320 17756 2372 17808
rect 8208 17799 8260 17808
rect 8208 17765 8217 17799
rect 8217 17765 8251 17799
rect 8251 17765 8260 17799
rect 8208 17756 8260 17765
rect 10416 17799 10468 17808
rect 10416 17765 10425 17799
rect 10425 17765 10459 17799
rect 10459 17765 10468 17799
rect 10416 17756 10468 17765
rect 7012 17688 7064 17740
rect 3056 17620 3108 17672
rect 10784 17688 10836 17740
rect 10416 17620 10468 17672
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 3792 17323 3844 17332
rect 3792 17289 3801 17323
rect 3801 17289 3835 17323
rect 3835 17289 3844 17323
rect 3792 17280 3844 17289
rect 10784 17323 10836 17332
rect 10784 17289 10793 17323
rect 10793 17289 10827 17323
rect 10827 17289 10836 17323
rect 10784 17280 10836 17289
rect 3056 17187 3108 17196
rect 1952 17076 2004 17128
rect 3056 17153 3065 17187
rect 3065 17153 3099 17187
rect 3099 17153 3108 17187
rect 3056 17144 3108 17153
rect 6184 17187 6236 17196
rect 6184 17153 6193 17187
rect 6193 17153 6227 17187
rect 6227 17153 6236 17187
rect 6184 17144 6236 17153
rect 8668 17187 8720 17196
rect 8668 17153 8677 17187
rect 8677 17153 8711 17187
rect 8711 17153 8720 17187
rect 8668 17144 8720 17153
rect 9864 17187 9916 17196
rect 9864 17153 9873 17187
rect 9873 17153 9907 17187
rect 9907 17153 9916 17187
rect 9864 17144 9916 17153
rect 11428 17187 11480 17196
rect 11428 17153 11437 17187
rect 11437 17153 11471 17187
rect 11471 17153 11480 17187
rect 11428 17144 11480 17153
rect 2412 17119 2464 17128
rect 2412 17085 2421 17119
rect 2421 17085 2455 17119
rect 2455 17085 2464 17119
rect 2412 17076 2464 17085
rect 2688 17008 2740 17060
rect 1768 16983 1820 16992
rect 1768 16949 1777 16983
rect 1777 16949 1811 16983
rect 1811 16949 1820 16983
rect 1768 16940 1820 16949
rect 5724 17008 5776 17060
rect 4160 16983 4212 16992
rect 4160 16949 4169 16983
rect 4169 16949 4203 16983
rect 4203 16949 4212 16983
rect 4160 16940 4212 16949
rect 5908 16983 5960 16992
rect 5908 16949 5917 16983
rect 5917 16949 5951 16983
rect 5951 16949 5960 16983
rect 5908 16940 5960 16949
rect 6000 16983 6052 16992
rect 6000 16949 6009 16983
rect 6009 16949 6043 16983
rect 6043 16949 6052 16983
rect 6000 16940 6052 16949
rect 9588 16983 9640 16992
rect 9588 16949 9597 16983
rect 9597 16949 9631 16983
rect 9631 16949 9640 16983
rect 9588 16940 9640 16949
rect 9680 16983 9732 16992
rect 9680 16949 9689 16983
rect 9689 16949 9723 16983
rect 9723 16949 9732 16983
rect 9680 16940 9732 16949
rect 11060 16940 11112 16992
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 2044 16668 2096 16720
rect 4068 16668 4120 16720
rect 2688 16643 2740 16652
rect 2688 16609 2697 16643
rect 2697 16609 2731 16643
rect 2731 16609 2740 16643
rect 2688 16600 2740 16609
rect 3148 16643 3200 16652
rect 3148 16609 3157 16643
rect 3157 16609 3191 16643
rect 3191 16609 3200 16643
rect 3148 16600 3200 16609
rect 3608 16600 3660 16652
rect 4988 16600 5040 16652
rect 6184 16736 6236 16788
rect 9588 16736 9640 16788
rect 9864 16736 9916 16788
rect 10508 16736 10560 16788
rect 11428 16736 11480 16788
rect 17960 16736 18012 16788
rect 6276 16668 6328 16720
rect 7288 16600 7340 16652
rect 10232 16600 10284 16652
rect 10324 16600 10376 16652
rect 11612 16643 11664 16652
rect 11612 16609 11646 16643
rect 11646 16609 11664 16643
rect 11612 16600 11664 16609
rect 6092 16575 6144 16584
rect 6092 16541 6101 16575
rect 6101 16541 6135 16575
rect 6135 16541 6144 16575
rect 6092 16532 6144 16541
rect 8116 16575 8168 16584
rect 8116 16541 8125 16575
rect 8125 16541 8159 16575
rect 8159 16541 8168 16575
rect 8116 16532 8168 16541
rect 3332 16507 3384 16516
rect 3332 16473 3341 16507
rect 3341 16473 3375 16507
rect 3375 16473 3384 16507
rect 3332 16464 3384 16473
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 4988 16235 5040 16244
rect 4988 16201 4997 16235
rect 4997 16201 5031 16235
rect 5031 16201 5040 16235
rect 4988 16192 5040 16201
rect 6000 16192 6052 16244
rect 7288 16235 7340 16244
rect 7288 16201 7297 16235
rect 7297 16201 7331 16235
rect 7331 16201 7340 16235
rect 7288 16192 7340 16201
rect 11612 16235 11664 16244
rect 11612 16201 11621 16235
rect 11621 16201 11655 16235
rect 11655 16201 11664 16235
rect 11612 16192 11664 16201
rect 2872 16124 2924 16176
rect 3148 16056 3200 16108
rect 3608 16099 3660 16108
rect 3608 16065 3617 16099
rect 3617 16065 3651 16099
rect 3651 16065 3660 16099
rect 3608 16056 3660 16065
rect 5908 16056 5960 16108
rect 6276 16099 6328 16108
rect 6276 16065 6285 16099
rect 6285 16065 6319 16099
rect 6319 16065 6328 16099
rect 6276 16056 6328 16065
rect 1492 16031 1544 16040
rect 1492 15997 1501 16031
rect 1501 15997 1535 16031
rect 1535 15997 1544 16031
rect 1492 15988 1544 15997
rect 2780 16031 2832 16040
rect 2780 15997 2789 16031
rect 2789 15997 2823 16031
rect 2823 15997 2832 16031
rect 2780 15988 2832 15997
rect 8116 15988 8168 16040
rect 8208 15988 8260 16040
rect 1676 15895 1728 15904
rect 1676 15861 1685 15895
rect 1685 15861 1719 15895
rect 1719 15861 1728 15895
rect 1676 15852 1728 15861
rect 2964 15895 3016 15904
rect 2964 15861 2973 15895
rect 2973 15861 3007 15895
rect 3007 15861 3016 15895
rect 2964 15852 3016 15861
rect 4252 15920 4304 15972
rect 6828 15920 6880 15972
rect 10324 15988 10376 16040
rect 10508 16031 10560 16040
rect 10508 15997 10542 16031
rect 10542 15997 10560 16031
rect 10508 15988 10560 15997
rect 9128 15920 9180 15972
rect 4804 15852 4856 15904
rect 6276 15852 6328 15904
rect 7748 15895 7800 15904
rect 7748 15861 7757 15895
rect 7757 15861 7791 15895
rect 7791 15861 7800 15895
rect 7748 15852 7800 15861
rect 10232 15852 10284 15904
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 4068 15691 4120 15700
rect 1952 15580 2004 15632
rect 4068 15657 4077 15691
rect 4077 15657 4111 15691
rect 4111 15657 4120 15691
rect 4068 15648 4120 15657
rect 4160 15648 4212 15700
rect 6276 15648 6328 15700
rect 6552 15648 6604 15700
rect 9128 15691 9180 15700
rect 6184 15623 6236 15632
rect 6184 15589 6218 15623
rect 6218 15589 6236 15623
rect 6184 15580 6236 15589
rect 4712 15512 4764 15564
rect 6000 15512 6052 15564
rect 8208 15580 8260 15632
rect 9128 15657 9137 15691
rect 9137 15657 9171 15691
rect 9171 15657 9180 15691
rect 9128 15648 9180 15657
rect 9680 15691 9732 15700
rect 9680 15657 9689 15691
rect 9689 15657 9723 15691
rect 9723 15657 9732 15691
rect 9680 15648 9732 15657
rect 11060 15691 11112 15700
rect 11060 15657 11069 15691
rect 11069 15657 11103 15691
rect 11103 15657 11112 15691
rect 11060 15648 11112 15657
rect 11704 15580 11756 15632
rect 8852 15512 8904 15564
rect 11060 15512 11112 15564
rect 2504 15444 2556 15496
rect 3332 15487 3384 15496
rect 3332 15453 3341 15487
rect 3341 15453 3375 15487
rect 3375 15453 3384 15487
rect 3332 15444 3384 15453
rect 3516 15487 3568 15496
rect 3516 15453 3525 15487
rect 3525 15453 3559 15487
rect 3559 15453 3568 15487
rect 3516 15444 3568 15453
rect 4988 15444 5040 15496
rect 10232 15487 10284 15496
rect 10232 15453 10241 15487
rect 10241 15453 10275 15487
rect 10275 15453 10284 15487
rect 10232 15444 10284 15453
rect 12072 15512 12124 15564
rect 11612 15487 11664 15496
rect 11612 15453 11621 15487
rect 11621 15453 11655 15487
rect 11655 15453 11664 15487
rect 11612 15444 11664 15453
rect 1768 15351 1820 15360
rect 1768 15317 1777 15351
rect 1777 15317 1811 15351
rect 1811 15317 1820 15351
rect 1768 15308 1820 15317
rect 7564 15308 7616 15360
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 4252 15104 4304 15156
rect 4712 15104 4764 15156
rect 5724 15147 5776 15156
rect 5724 15113 5733 15147
rect 5733 15113 5767 15147
rect 5767 15113 5776 15147
rect 5724 15104 5776 15113
rect 7748 15104 7800 15156
rect 8852 15104 8904 15156
rect 2780 15036 2832 15088
rect 5264 14968 5316 15020
rect 6368 15011 6420 15020
rect 1952 14900 2004 14952
rect 2872 14900 2924 14952
rect 5724 14900 5776 14952
rect 6368 14977 6377 15011
rect 6377 14977 6411 15011
rect 6411 14977 6420 15011
rect 6368 14968 6420 14977
rect 7564 15011 7616 15020
rect 7564 14977 7573 15011
rect 7573 14977 7607 15011
rect 7607 14977 7616 15011
rect 7564 14968 7616 14977
rect 8208 14968 8260 15020
rect 3516 14832 3568 14884
rect 7748 14832 7800 14884
rect 9404 14832 9456 14884
rect 1676 14807 1728 14816
rect 1676 14773 1685 14807
rect 1685 14773 1719 14807
rect 1719 14773 1728 14807
rect 1676 14764 1728 14773
rect 5264 14764 5316 14816
rect 5816 14764 5868 14816
rect 7380 14807 7432 14816
rect 7380 14773 7389 14807
rect 7389 14773 7423 14807
rect 7423 14773 7432 14807
rect 7380 14764 7432 14773
rect 7472 14807 7524 14816
rect 7472 14773 7481 14807
rect 7481 14773 7515 14807
rect 7515 14773 7524 14807
rect 7472 14764 7524 14773
rect 10692 14764 10744 14816
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 3516 14603 3568 14612
rect 3516 14569 3525 14603
rect 3525 14569 3559 14603
rect 3559 14569 3568 14603
rect 3516 14560 3568 14569
rect 4804 14560 4856 14612
rect 5816 14603 5868 14612
rect 5816 14569 5825 14603
rect 5825 14569 5859 14603
rect 5859 14569 5868 14603
rect 5816 14560 5868 14569
rect 6368 14560 6420 14612
rect 7104 14560 7156 14612
rect 8576 14603 8628 14612
rect 8576 14569 8585 14603
rect 8585 14569 8619 14603
rect 8619 14569 8628 14603
rect 8576 14560 8628 14569
rect 1492 14492 1544 14544
rect 4252 14492 4304 14544
rect 7564 14492 7616 14544
rect 3976 14424 4028 14476
rect 5816 14424 5868 14476
rect 6092 14424 6144 14476
rect 6920 14424 6972 14476
rect 7380 14424 7432 14476
rect 11060 14560 11112 14612
rect 9680 14492 9732 14544
rect 9588 14424 9640 14476
rect 4896 14399 4948 14408
rect 4896 14365 4905 14399
rect 4905 14365 4939 14399
rect 4939 14365 4948 14399
rect 4896 14356 4948 14365
rect 5080 14399 5132 14408
rect 5080 14365 5089 14399
rect 5089 14365 5123 14399
rect 5123 14365 5132 14399
rect 5080 14356 5132 14365
rect 9404 14356 9456 14408
rect 10324 14492 10376 14544
rect 9956 14467 10008 14476
rect 9956 14433 9990 14467
rect 9990 14433 10008 14467
rect 9956 14424 10008 14433
rect 2872 14220 2924 14272
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 3332 14016 3384 14068
rect 3976 14016 4028 14068
rect 9956 14059 10008 14068
rect 9956 14025 9965 14059
rect 9965 14025 9999 14059
rect 9999 14025 10008 14059
rect 9956 14016 10008 14025
rect 3424 13880 3476 13932
rect 1768 13812 1820 13864
rect 2504 13855 2556 13864
rect 2504 13821 2513 13855
rect 2513 13821 2547 13855
rect 2547 13821 2556 13855
rect 2504 13812 2556 13821
rect 3332 13812 3384 13864
rect 9588 13880 9640 13932
rect 3700 13812 3752 13864
rect 2872 13744 2924 13796
rect 4068 13744 4120 13796
rect 6920 13812 6972 13864
rect 7104 13855 7156 13864
rect 7104 13821 7138 13855
rect 7138 13821 7156 13855
rect 7104 13812 7156 13821
rect 5080 13744 5132 13796
rect 5816 13787 5868 13796
rect 5816 13753 5825 13787
rect 5825 13753 5859 13787
rect 5859 13753 5868 13787
rect 5816 13744 5868 13753
rect 7564 13812 7616 13864
rect 9036 13744 9088 13796
rect 5356 13676 5408 13728
rect 8208 13719 8260 13728
rect 8208 13685 8217 13719
rect 8217 13685 8251 13719
rect 8251 13685 8260 13719
rect 8208 13676 8260 13685
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 3608 13515 3660 13524
rect 3608 13481 3617 13515
rect 3617 13481 3651 13515
rect 3651 13481 3660 13515
rect 3608 13472 3660 13481
rect 5080 13472 5132 13524
rect 5724 13515 5776 13524
rect 5724 13481 5733 13515
rect 5733 13481 5767 13515
rect 5767 13481 5776 13515
rect 5724 13472 5776 13481
rect 6920 13472 6972 13524
rect 7196 13472 7248 13524
rect 9680 13515 9732 13524
rect 9680 13481 9689 13515
rect 9689 13481 9723 13515
rect 9723 13481 9732 13515
rect 9680 13472 9732 13481
rect 5172 13404 5224 13456
rect 5356 13404 5408 13456
rect 1676 13379 1728 13388
rect 1676 13345 1685 13379
rect 1685 13345 1719 13379
rect 1719 13345 1728 13379
rect 1676 13336 1728 13345
rect 2780 13379 2832 13388
rect 2780 13345 2789 13379
rect 2789 13345 2823 13379
rect 2823 13345 2832 13379
rect 3424 13379 3476 13388
rect 2780 13336 2832 13345
rect 3424 13345 3433 13379
rect 3433 13345 3467 13379
rect 3467 13345 3476 13379
rect 3424 13336 3476 13345
rect 4068 13379 4120 13388
rect 4068 13345 4077 13379
rect 4077 13345 4111 13379
rect 4111 13345 4120 13379
rect 4068 13336 4120 13345
rect 4804 13336 4856 13388
rect 7104 13336 7156 13388
rect 1492 13268 1544 13320
rect 2964 13311 3016 13320
rect 2964 13277 2973 13311
rect 2973 13277 3007 13311
rect 3007 13277 3016 13311
rect 6184 13311 6236 13320
rect 2964 13268 3016 13277
rect 6184 13277 6193 13311
rect 6193 13277 6227 13311
rect 6227 13277 6236 13311
rect 6184 13268 6236 13277
rect 6368 13311 6420 13320
rect 6368 13277 6377 13311
rect 6377 13277 6411 13311
rect 6411 13277 6420 13311
rect 6368 13268 6420 13277
rect 7196 13268 7248 13320
rect 9220 13336 9272 13388
rect 9956 13404 10008 13456
rect 9036 13268 9088 13320
rect 2412 13175 2464 13184
rect 2412 13141 2421 13175
rect 2421 13141 2455 13175
rect 2455 13141 2464 13175
rect 2412 13132 2464 13141
rect 10048 13200 10100 13252
rect 3148 13132 3200 13184
rect 7380 13132 7432 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 5172 12928 5224 12980
rect 9036 12971 9088 12980
rect 9036 12937 9045 12971
rect 9045 12937 9079 12971
rect 9079 12937 9088 12971
rect 9036 12928 9088 12937
rect 10324 12928 10376 12980
rect 4712 12860 4764 12912
rect 1952 12792 2004 12844
rect 4804 12792 4856 12844
rect 7196 12835 7248 12844
rect 7196 12801 7205 12835
rect 7205 12801 7239 12835
rect 7239 12801 7248 12835
rect 7196 12792 7248 12801
rect 7564 12792 7616 12844
rect 1860 12767 1912 12776
rect 1860 12733 1869 12767
rect 1869 12733 1903 12767
rect 1903 12733 1912 12767
rect 1860 12724 1912 12733
rect 2688 12724 2740 12776
rect 2872 12767 2924 12776
rect 2872 12733 2881 12767
rect 2881 12733 2915 12767
rect 2915 12733 2924 12767
rect 2872 12724 2924 12733
rect 4988 12767 5040 12776
rect 4988 12733 4997 12767
rect 4997 12733 5031 12767
rect 5031 12733 5040 12767
rect 4988 12724 5040 12733
rect 6368 12724 6420 12776
rect 10416 12724 10468 12776
rect 3516 12656 3568 12708
rect 4804 12656 4856 12708
rect 5356 12656 5408 12708
rect 8668 12656 8720 12708
rect 4160 12588 4212 12640
rect 4988 12588 5040 12640
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 1584 12384 1636 12436
rect 1860 12384 1912 12436
rect 2412 12427 2464 12436
rect 2412 12393 2421 12427
rect 2421 12393 2455 12427
rect 2455 12393 2464 12427
rect 2412 12384 2464 12393
rect 3240 12427 3292 12436
rect 3240 12393 3249 12427
rect 3249 12393 3283 12427
rect 3283 12393 3292 12427
rect 3240 12384 3292 12393
rect 4160 12384 4212 12436
rect 4896 12384 4948 12436
rect 3424 12316 3476 12368
rect 5080 12316 5132 12368
rect 6368 12384 6420 12436
rect 9220 12384 9272 12436
rect 1492 12291 1544 12300
rect 1492 12257 1501 12291
rect 1501 12257 1535 12291
rect 1535 12257 1544 12291
rect 1492 12248 1544 12257
rect 3608 12248 3660 12300
rect 4896 12291 4948 12300
rect 2504 12223 2556 12232
rect 2504 12189 2513 12223
rect 2513 12189 2547 12223
rect 2547 12189 2556 12223
rect 2504 12180 2556 12189
rect 3516 12180 3568 12232
rect 4896 12257 4905 12291
rect 4905 12257 4939 12291
rect 4939 12257 4948 12291
rect 4896 12248 4948 12257
rect 5172 12223 5224 12232
rect 5172 12189 5181 12223
rect 5181 12189 5215 12223
rect 5215 12189 5224 12223
rect 5172 12180 5224 12189
rect 5632 12248 5684 12300
rect 6368 12248 6420 12300
rect 6828 12248 6880 12300
rect 7380 12248 7432 12300
rect 8392 12248 8444 12300
rect 8484 12248 8536 12300
rect 6920 12180 6972 12232
rect 9956 12180 10008 12232
rect 8668 12155 8720 12164
rect 2872 12044 2924 12096
rect 4896 12044 4948 12096
rect 8668 12121 8677 12155
rect 8677 12121 8711 12155
rect 8711 12121 8720 12155
rect 8668 12112 8720 12121
rect 7104 12044 7156 12096
rect 20352 12044 20404 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 2504 11840 2556 11892
rect 4068 11840 4120 11892
rect 6368 11883 6420 11892
rect 3516 11815 3568 11824
rect 3516 11781 3525 11815
rect 3525 11781 3559 11815
rect 3559 11781 3568 11815
rect 3516 11772 3568 11781
rect 6368 11849 6377 11883
rect 6377 11849 6411 11883
rect 6411 11849 6420 11883
rect 6368 11840 6420 11849
rect 7104 11840 7156 11892
rect 7656 11840 7708 11892
rect 3424 11704 3476 11756
rect 1584 11636 1636 11688
rect 2964 11636 3016 11688
rect 4896 11636 4948 11688
rect 7104 11636 7156 11688
rect 8392 11747 8444 11756
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 8392 11704 8444 11713
rect 2688 11568 2740 11620
rect 2780 11568 2832 11620
rect 3240 11568 3292 11620
rect 2320 11500 2372 11552
rect 5632 11568 5684 11620
rect 3608 11500 3660 11552
rect 5540 11500 5592 11552
rect 5724 11500 5776 11552
rect 6276 11500 6328 11552
rect 8576 11500 8628 11552
rect 10324 11636 10376 11688
rect 19064 11679 19116 11688
rect 19064 11645 19073 11679
rect 19073 11645 19107 11679
rect 19107 11645 19116 11679
rect 19064 11636 19116 11645
rect 9588 11611 9640 11620
rect 9588 11577 9622 11611
rect 9622 11577 9640 11611
rect 9588 11568 9640 11577
rect 9680 11568 9732 11620
rect 11152 11500 11204 11552
rect 19892 11500 19944 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 2320 11339 2372 11348
rect 2320 11305 2329 11339
rect 2329 11305 2363 11339
rect 2363 11305 2372 11339
rect 2320 11296 2372 11305
rect 2872 11296 2924 11348
rect 3240 11296 3292 11348
rect 4252 11296 4304 11348
rect 6184 11296 6236 11348
rect 7012 11296 7064 11348
rect 8576 11339 8628 11348
rect 6092 11228 6144 11280
rect 8576 11305 8585 11339
rect 8585 11305 8619 11339
rect 8619 11305 8628 11339
rect 8576 11296 8628 11305
rect 8668 11296 8720 11348
rect 3240 11160 3292 11212
rect 8484 11160 8536 11212
rect 4988 11135 5040 11144
rect 2688 11024 2740 11076
rect 4988 11101 4997 11135
rect 4997 11101 5031 11135
rect 5031 11101 5040 11135
rect 4988 11092 5040 11101
rect 5632 11092 5684 11144
rect 6368 11092 6420 11144
rect 3240 11024 3292 11076
rect 5264 11024 5316 11076
rect 5908 11024 5960 11076
rect 7748 11092 7800 11144
rect 9588 11228 9640 11280
rect 11152 11296 11204 11348
rect 19064 11296 19116 11348
rect 9680 11203 9732 11212
rect 9680 11169 9689 11203
rect 9689 11169 9723 11203
rect 9723 11169 9732 11203
rect 9680 11160 9732 11169
rect 10784 11160 10836 11212
rect 8576 11024 8628 11076
rect 9404 11024 9456 11076
rect 19432 11024 19484 11076
rect 4068 10956 4120 11008
rect 9680 10956 9732 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 2964 10795 3016 10804
rect 2964 10761 2973 10795
rect 2973 10761 3007 10795
rect 3007 10761 3016 10795
rect 2964 10752 3016 10761
rect 3332 10752 3384 10804
rect 5632 10752 5684 10804
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 4344 10659 4396 10668
rect 4344 10625 4353 10659
rect 4353 10625 4387 10659
rect 4387 10625 4396 10659
rect 4344 10616 4396 10625
rect 4896 10616 4948 10668
rect 2688 10548 2740 10600
rect 3056 10548 3108 10600
rect 9496 10752 9548 10804
rect 10508 10795 10560 10804
rect 10508 10761 10517 10795
rect 10517 10761 10551 10795
rect 10551 10761 10560 10795
rect 10508 10752 10560 10761
rect 9036 10727 9088 10736
rect 9036 10693 9045 10727
rect 9045 10693 9079 10727
rect 9079 10693 9088 10727
rect 9036 10684 9088 10693
rect 7656 10591 7708 10600
rect 7656 10557 7665 10591
rect 7665 10557 7699 10591
rect 7699 10557 7708 10591
rect 7656 10548 7708 10557
rect 7748 10548 7800 10600
rect 9128 10548 9180 10600
rect 10784 10548 10836 10600
rect 18236 10591 18288 10600
rect 18236 10557 18245 10591
rect 18245 10557 18279 10591
rect 18279 10557 18288 10591
rect 18236 10548 18288 10557
rect 5080 10480 5132 10532
rect 5448 10480 5500 10532
rect 5724 10480 5776 10532
rect 2780 10412 2832 10464
rect 3424 10412 3476 10464
rect 6828 10412 6880 10464
rect 7104 10412 7156 10464
rect 18696 10412 18748 10464
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 3056 10251 3108 10260
rect 3056 10217 3065 10251
rect 3065 10217 3099 10251
rect 3099 10217 3108 10251
rect 3056 10208 3108 10217
rect 4252 10208 4304 10260
rect 5448 10208 5500 10260
rect 7748 10208 7800 10260
rect 8484 10251 8536 10260
rect 8484 10217 8493 10251
rect 8493 10217 8527 10251
rect 8527 10217 8536 10251
rect 8484 10208 8536 10217
rect 9588 10208 9640 10260
rect 11980 10208 12032 10260
rect 2688 10140 2740 10192
rect 2780 10004 2832 10056
rect 3700 10140 3752 10192
rect 4344 10072 4396 10124
rect 4896 10072 4948 10124
rect 3516 10004 3568 10056
rect 5540 10140 5592 10192
rect 6644 10140 6696 10192
rect 6460 10072 6512 10124
rect 6920 10072 6972 10124
rect 8208 10072 8260 10124
rect 8300 10072 8352 10124
rect 10324 10072 10376 10124
rect 6552 10004 6604 10056
rect 8668 10004 8720 10056
rect 8208 9936 8260 9988
rect 9220 9936 9272 9988
rect 18236 9936 18288 9988
rect 4068 9868 4120 9920
rect 10876 9868 10928 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 2688 9664 2740 9716
rect 3792 9664 3844 9716
rect 3884 9664 3936 9716
rect 4896 9707 4948 9716
rect 4896 9673 4905 9707
rect 4905 9673 4939 9707
rect 4939 9673 4948 9707
rect 4896 9664 4948 9673
rect 10784 9664 10836 9716
rect 10876 9664 10928 9716
rect 14372 9664 14424 9716
rect 4988 9596 5040 9648
rect 6828 9639 6880 9648
rect 6828 9605 6837 9639
rect 6837 9605 6871 9639
rect 6871 9605 6880 9639
rect 6828 9596 6880 9605
rect 10416 9639 10468 9648
rect 10416 9605 10425 9639
rect 10425 9605 10459 9639
rect 10459 9605 10468 9639
rect 10416 9596 10468 9605
rect 5448 9528 5500 9580
rect 1584 9503 1636 9512
rect 1584 9469 1593 9503
rect 1593 9469 1627 9503
rect 1627 9469 1636 9503
rect 3516 9503 3568 9512
rect 1584 9460 1636 9469
rect 3516 9469 3525 9503
rect 3525 9469 3559 9503
rect 3559 9469 3568 9503
rect 3516 9460 3568 9469
rect 4712 9460 4764 9512
rect 5540 9460 5592 9512
rect 2320 9392 2372 9444
rect 2780 9392 2832 9444
rect 8300 9528 8352 9580
rect 7656 9460 7708 9512
rect 9036 9503 9088 9512
rect 9036 9469 9070 9503
rect 9070 9469 9088 9503
rect 9036 9460 9088 9469
rect 11796 9460 11848 9512
rect 6920 9392 6972 9444
rect 9680 9392 9732 9444
rect 11152 9392 11204 9444
rect 4436 9324 4488 9376
rect 4804 9324 4856 9376
rect 4988 9324 5040 9376
rect 5724 9324 5776 9376
rect 6184 9367 6236 9376
rect 6184 9333 6193 9367
rect 6193 9333 6227 9367
rect 6227 9333 6236 9367
rect 6184 9324 6236 9333
rect 6828 9324 6880 9376
rect 8944 9324 8996 9376
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 2780 9163 2832 9172
rect 2780 9129 2789 9163
rect 2789 9129 2823 9163
rect 2823 9129 2832 9163
rect 2780 9120 2832 9129
rect 4436 9163 4488 9172
rect 4436 9129 4445 9163
rect 4445 9129 4479 9163
rect 4479 9129 4488 9163
rect 4436 9120 4488 9129
rect 5080 9163 5132 9172
rect 4712 9052 4764 9104
rect 5080 9129 5089 9163
rect 5089 9129 5123 9163
rect 5123 9129 5132 9163
rect 5080 9120 5132 9129
rect 6184 9120 6236 9172
rect 8576 9163 8628 9172
rect 8576 9129 8585 9163
rect 8585 9129 8619 9163
rect 8619 9129 8628 9163
rect 8576 9120 8628 9129
rect 8944 9163 8996 9172
rect 8944 9129 8953 9163
rect 8953 9129 8987 9163
rect 8987 9129 8996 9163
rect 8944 9120 8996 9129
rect 2504 8984 2556 9036
rect 5816 9052 5868 9104
rect 12256 9052 12308 9104
rect 4712 8959 4764 8968
rect 4712 8925 4721 8959
rect 4721 8925 4755 8959
rect 4755 8925 4764 8959
rect 4712 8916 4764 8925
rect 5264 8916 5316 8968
rect 6184 8984 6236 9036
rect 6736 9027 6788 9036
rect 6736 8993 6745 9027
rect 6745 8993 6779 9027
rect 6779 8993 6788 9027
rect 6736 8984 6788 8993
rect 7012 8984 7064 9036
rect 7748 8984 7800 9036
rect 8208 8984 8260 9036
rect 10876 8984 10928 9036
rect 6552 8916 6604 8968
rect 8116 8959 8168 8968
rect 8116 8925 8125 8959
rect 8125 8925 8159 8959
rect 8159 8925 8168 8959
rect 8116 8916 8168 8925
rect 8576 8916 8628 8968
rect 9220 8959 9272 8968
rect 9220 8925 9229 8959
rect 9229 8925 9263 8959
rect 9263 8925 9272 8959
rect 9220 8916 9272 8925
rect 9680 8916 9732 8968
rect 3976 8848 4028 8900
rect 9312 8848 9364 8900
rect 1584 8780 1636 8832
rect 2596 8780 2648 8832
rect 4804 8780 4856 8832
rect 7196 8780 7248 8832
rect 7288 8780 7340 8832
rect 8852 8780 8904 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 1676 8576 1728 8628
rect 4436 8551 4488 8560
rect 4436 8517 4445 8551
rect 4445 8517 4479 8551
rect 4479 8517 4488 8551
rect 4436 8508 4488 8517
rect 4712 8508 4764 8560
rect 2320 8483 2372 8492
rect 2320 8449 2329 8483
rect 2329 8449 2363 8483
rect 2363 8449 2372 8483
rect 2320 8440 2372 8449
rect 4896 8440 4948 8492
rect 6736 8440 6788 8492
rect 7656 8576 7708 8628
rect 8116 8576 8168 8628
rect 10876 8576 10928 8628
rect 11796 8619 11848 8628
rect 11796 8585 11805 8619
rect 11805 8585 11839 8619
rect 11839 8585 11848 8619
rect 11796 8576 11848 8585
rect 9680 8483 9732 8492
rect 2780 8415 2832 8424
rect 2780 8381 2789 8415
rect 2789 8381 2823 8415
rect 2823 8381 2832 8415
rect 2780 8372 2832 8381
rect 3792 8372 3844 8424
rect 4804 8415 4856 8424
rect 4804 8381 4813 8415
rect 4813 8381 4847 8415
rect 4847 8381 4856 8415
rect 4804 8372 4856 8381
rect 2136 8279 2188 8288
rect 2136 8245 2145 8279
rect 2145 8245 2179 8279
rect 2179 8245 2188 8279
rect 2136 8236 2188 8245
rect 2228 8279 2280 8288
rect 2228 8245 2237 8279
rect 2237 8245 2271 8279
rect 2271 8245 2280 8279
rect 2228 8236 2280 8245
rect 2780 8236 2832 8288
rect 4160 8279 4212 8288
rect 4160 8245 4169 8279
rect 4169 8245 4203 8279
rect 4203 8245 4212 8279
rect 4160 8236 4212 8245
rect 5172 8304 5224 8356
rect 4804 8236 4856 8288
rect 6092 8304 6144 8356
rect 7104 8372 7156 8424
rect 9680 8449 9689 8483
rect 9689 8449 9723 8483
rect 9723 8449 9732 8483
rect 9680 8440 9732 8449
rect 6828 8304 6880 8356
rect 7656 8347 7708 8356
rect 7656 8313 7690 8347
rect 7690 8313 7708 8347
rect 7656 8304 7708 8313
rect 11704 8372 11756 8424
rect 11980 8415 12032 8424
rect 11980 8381 11989 8415
rect 11989 8381 12023 8415
rect 12023 8381 12032 8415
rect 11980 8372 12032 8381
rect 10416 8304 10468 8356
rect 11336 8279 11388 8288
rect 11336 8245 11345 8279
rect 11345 8245 11379 8279
rect 11379 8245 11388 8279
rect 11336 8236 11388 8245
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 2136 8032 2188 8084
rect 5172 8032 5224 8084
rect 7012 8075 7064 8084
rect 7012 8041 7021 8075
rect 7021 8041 7055 8075
rect 7055 8041 7064 8075
rect 7012 8032 7064 8041
rect 5264 7964 5316 8016
rect 6552 7964 6604 8016
rect 2504 7828 2556 7880
rect 2780 7871 2832 7880
rect 2780 7837 2789 7871
rect 2789 7837 2823 7871
rect 2823 7837 2832 7871
rect 2780 7828 2832 7837
rect 4160 7828 4212 7880
rect 4896 7896 4948 7948
rect 6368 7896 6420 7948
rect 7748 8032 7800 8084
rect 11336 7964 11388 8016
rect 11704 7964 11756 8016
rect 15752 7964 15804 8016
rect 4804 7828 4856 7880
rect 2688 7760 2740 7812
rect 3700 7803 3752 7812
rect 3700 7769 3709 7803
rect 3709 7769 3743 7803
rect 3743 7769 3752 7803
rect 7104 7828 7156 7880
rect 11152 7896 11204 7948
rect 7656 7871 7708 7880
rect 7656 7837 7665 7871
rect 7665 7837 7699 7871
rect 7699 7837 7708 7871
rect 7656 7828 7708 7837
rect 8484 7828 8536 7880
rect 8852 7871 8904 7880
rect 8852 7837 8861 7871
rect 8861 7837 8895 7871
rect 8895 7837 8904 7871
rect 8852 7828 8904 7837
rect 10876 7871 10928 7880
rect 10876 7837 10885 7871
rect 10885 7837 10919 7871
rect 10919 7837 10928 7871
rect 10876 7828 10928 7837
rect 10968 7828 11020 7880
rect 15016 7828 15068 7880
rect 3700 7760 3752 7769
rect 4988 7692 5040 7744
rect 14648 7760 14700 7812
rect 6552 7735 6604 7744
rect 6552 7701 6561 7735
rect 6561 7701 6595 7735
rect 6595 7701 6604 7735
rect 6552 7692 6604 7701
rect 7012 7692 7064 7744
rect 7564 7692 7616 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 1768 7488 1820 7540
rect 4068 7488 4120 7540
rect 5724 7488 5776 7540
rect 6460 7488 6512 7540
rect 8208 7488 8260 7540
rect 5448 7420 5500 7472
rect 7104 7420 7156 7472
rect 8668 7420 8720 7472
rect 15660 7420 15712 7472
rect 2504 7395 2556 7404
rect 2504 7361 2513 7395
rect 2513 7361 2547 7395
rect 2547 7361 2556 7395
rect 2504 7352 2556 7361
rect 3608 7395 3660 7404
rect 3608 7361 3617 7395
rect 3617 7361 3651 7395
rect 3651 7361 3660 7395
rect 3608 7352 3660 7361
rect 3700 7352 3752 7404
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 6552 7284 6604 7336
rect 8852 7352 8904 7404
rect 9680 7352 9732 7404
rect 8944 7284 8996 7336
rect 15200 7352 15252 7404
rect 10968 7284 11020 7336
rect 11888 7284 11940 7336
rect 14648 7284 14700 7336
rect 1584 7216 1636 7268
rect 3424 7259 3476 7268
rect 3424 7225 3433 7259
rect 3433 7225 3467 7259
rect 3467 7225 3476 7259
rect 3424 7216 3476 7225
rect 3976 7216 4028 7268
rect 3516 7191 3568 7200
rect 3516 7157 3525 7191
rect 3525 7157 3559 7191
rect 3559 7157 3568 7191
rect 3516 7148 3568 7157
rect 4712 7148 4764 7200
rect 7104 7216 7156 7268
rect 7196 7259 7248 7268
rect 7196 7225 7205 7259
rect 7205 7225 7239 7259
rect 7239 7225 7248 7259
rect 7196 7216 7248 7225
rect 9220 7216 9272 7268
rect 10048 7216 10100 7268
rect 10232 7216 10284 7268
rect 10600 7259 10652 7268
rect 10600 7225 10634 7259
rect 10634 7225 10652 7259
rect 10600 7216 10652 7225
rect 14096 7216 14148 7268
rect 17776 7216 17828 7268
rect 10508 7148 10560 7200
rect 11704 7191 11756 7200
rect 11704 7157 11713 7191
rect 11713 7157 11747 7191
rect 11747 7157 11756 7191
rect 11704 7148 11756 7157
rect 11888 7148 11940 7200
rect 12440 7191 12492 7200
rect 12440 7157 12449 7191
rect 12449 7157 12483 7191
rect 12483 7157 12492 7191
rect 12440 7148 12492 7157
rect 14188 7148 14240 7200
rect 14372 7148 14424 7200
rect 15568 7191 15620 7200
rect 15568 7157 15577 7191
rect 15577 7157 15611 7191
rect 15611 7157 15620 7191
rect 15568 7148 15620 7157
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 1308 6944 1360 6996
rect 1860 6740 1912 6792
rect 2688 6876 2740 6928
rect 3424 6944 3476 6996
rect 6184 6944 6236 6996
rect 8484 6944 8536 6996
rect 9680 6944 9732 6996
rect 10876 6944 10928 6996
rect 3240 6876 3292 6928
rect 5356 6876 5408 6928
rect 2504 6808 2556 6860
rect 2964 6808 3016 6860
rect 3332 6808 3384 6860
rect 5172 6808 5224 6860
rect 5632 6851 5684 6860
rect 5632 6817 5666 6851
rect 5666 6817 5684 6851
rect 5632 6808 5684 6817
rect 7288 6851 7340 6860
rect 4712 6783 4764 6792
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 4712 6740 4764 6749
rect 4804 6672 4856 6724
rect 7288 6817 7311 6851
rect 7311 6817 7340 6851
rect 7288 6808 7340 6817
rect 10232 6808 10284 6860
rect 11704 6876 11756 6928
rect 12716 6876 12768 6928
rect 10600 6808 10652 6860
rect 5080 6647 5132 6656
rect 5080 6613 5089 6647
rect 5089 6613 5123 6647
rect 5123 6613 5132 6647
rect 5080 6604 5132 6613
rect 10968 6740 11020 6792
rect 8300 6604 8352 6656
rect 8484 6604 8536 6656
rect 11796 6604 11848 6656
rect 13912 6808 13964 6860
rect 15200 6808 15252 6860
rect 16028 6808 16080 6860
rect 16948 6851 17000 6860
rect 16948 6817 16957 6851
rect 16957 6817 16991 6851
rect 16991 6817 17000 6851
rect 16948 6808 17000 6817
rect 15016 6740 15068 6792
rect 17684 6740 17736 6792
rect 15936 6604 15988 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 2504 6400 2556 6452
rect 4068 6400 4120 6452
rect 5632 6332 5684 6384
rect 9772 6443 9824 6452
rect 9772 6409 9788 6443
rect 9788 6409 9822 6443
rect 9822 6409 9824 6443
rect 13912 6443 13964 6452
rect 9772 6400 9824 6409
rect 13912 6409 13921 6443
rect 13921 6409 13955 6443
rect 13955 6409 13964 6443
rect 13912 6400 13964 6409
rect 16948 6400 17000 6452
rect 4896 6264 4948 6316
rect 5816 6264 5868 6316
rect 7288 6264 7340 6316
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 2780 6128 2832 6180
rect 4712 6196 4764 6248
rect 5080 6196 5132 6248
rect 5724 6196 5776 6248
rect 7104 6196 7156 6248
rect 1952 6060 2004 6112
rect 3608 6060 3660 6112
rect 9864 6375 9916 6384
rect 9864 6341 9873 6375
rect 9873 6341 9907 6375
rect 9907 6341 9916 6375
rect 9864 6332 9916 6341
rect 9220 6264 9272 6316
rect 9772 6264 9824 6316
rect 8300 6196 8352 6248
rect 8484 6239 8536 6248
rect 8484 6205 8518 6239
rect 8518 6205 8536 6239
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 13544 6264 13596 6316
rect 15752 6307 15804 6316
rect 15752 6273 15761 6307
rect 15761 6273 15795 6307
rect 15795 6273 15804 6307
rect 15752 6264 15804 6273
rect 8484 6196 8536 6205
rect 10140 6196 10192 6248
rect 12348 6196 12400 6248
rect 14556 6239 14608 6248
rect 14556 6205 14565 6239
rect 14565 6205 14599 6239
rect 14599 6205 14608 6239
rect 14556 6196 14608 6205
rect 15568 6239 15620 6248
rect 15568 6205 15577 6239
rect 15577 6205 15611 6239
rect 15611 6205 15620 6239
rect 15568 6196 15620 6205
rect 15660 6239 15712 6248
rect 15660 6205 15669 6239
rect 15669 6205 15703 6239
rect 15703 6205 15712 6239
rect 15660 6196 15712 6205
rect 15936 6196 15988 6248
rect 5724 6060 5776 6112
rect 6828 6103 6880 6112
rect 6828 6069 6837 6103
rect 6837 6069 6871 6103
rect 6871 6069 6880 6103
rect 6828 6060 6880 6069
rect 9772 6103 9824 6112
rect 9772 6069 9781 6103
rect 9781 6069 9815 6103
rect 9815 6069 9824 6103
rect 9772 6060 9824 6069
rect 12624 6128 12676 6180
rect 13544 6128 13596 6180
rect 14096 6128 14148 6180
rect 17408 6128 17460 6180
rect 10232 6060 10284 6112
rect 10416 6060 10468 6112
rect 11152 6103 11204 6112
rect 11152 6069 11161 6103
rect 11161 6069 11195 6103
rect 11195 6069 11204 6103
rect 11152 6060 11204 6069
rect 11796 6060 11848 6112
rect 14280 6060 14332 6112
rect 16028 6060 16080 6112
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 1584 5899 1636 5908
rect 1584 5865 1593 5899
rect 1593 5865 1627 5899
rect 1627 5865 1636 5899
rect 1584 5856 1636 5865
rect 1952 5899 2004 5908
rect 1952 5865 1961 5899
rect 1961 5865 1995 5899
rect 1995 5865 2004 5899
rect 1952 5856 2004 5865
rect 3516 5856 3568 5908
rect 4160 5856 4212 5908
rect 8392 5856 8444 5908
rect 9864 5856 9916 5908
rect 5632 5788 5684 5840
rect 2964 5763 3016 5772
rect 1676 5652 1728 5704
rect 2964 5729 2973 5763
rect 2973 5729 3007 5763
rect 3007 5729 3016 5763
rect 2964 5720 3016 5729
rect 3608 5720 3660 5772
rect 4896 5720 4948 5772
rect 5080 5720 5132 5772
rect 7288 5788 7340 5840
rect 5816 5763 5868 5772
rect 5816 5729 5850 5763
rect 5850 5729 5868 5763
rect 5816 5720 5868 5729
rect 6552 5720 6604 5772
rect 7564 5763 7616 5772
rect 7564 5729 7573 5763
rect 7573 5729 7607 5763
rect 7607 5729 7616 5763
rect 7564 5720 7616 5729
rect 8300 5788 8352 5840
rect 8760 5788 8812 5840
rect 12164 5856 12216 5908
rect 14096 5856 14148 5908
rect 14280 5899 14332 5908
rect 14280 5865 14289 5899
rect 14289 5865 14323 5899
rect 14323 5865 14332 5899
rect 14280 5856 14332 5865
rect 17408 5899 17460 5908
rect 17408 5865 17417 5899
rect 17417 5865 17451 5899
rect 17451 5865 17460 5899
rect 17408 5856 17460 5865
rect 8852 5720 8904 5772
rect 3056 5695 3108 5704
rect 2780 5584 2832 5636
rect 3056 5661 3065 5695
rect 3065 5661 3099 5695
rect 3099 5661 3108 5695
rect 3056 5652 3108 5661
rect 3516 5652 3568 5704
rect 3700 5652 3752 5704
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 7656 5695 7708 5704
rect 7656 5661 7665 5695
rect 7665 5661 7699 5695
rect 7699 5661 7708 5695
rect 7656 5652 7708 5661
rect 8300 5652 8352 5704
rect 9772 5652 9824 5704
rect 11888 5788 11940 5840
rect 14188 5831 14240 5840
rect 10784 5763 10836 5772
rect 10784 5729 10818 5763
rect 10818 5729 10836 5763
rect 10784 5720 10836 5729
rect 3148 5584 3200 5636
rect 6828 5584 6880 5636
rect 12992 5720 13044 5772
rect 14188 5797 14197 5831
rect 14197 5797 14231 5831
rect 14231 5797 14240 5831
rect 14188 5788 14240 5797
rect 16488 5788 16540 5840
rect 17684 5763 17736 5772
rect 13912 5652 13964 5704
rect 2596 5559 2648 5568
rect 2596 5525 2605 5559
rect 2605 5525 2639 5559
rect 2639 5525 2648 5559
rect 2596 5516 2648 5525
rect 4068 5516 4120 5568
rect 6276 5516 6328 5568
rect 7104 5516 7156 5568
rect 8484 5516 8536 5568
rect 10232 5516 10284 5568
rect 17684 5729 17693 5763
rect 17693 5729 17727 5763
rect 17727 5729 17736 5763
rect 17684 5720 17736 5729
rect 15476 5695 15528 5704
rect 15476 5661 15485 5695
rect 15485 5661 15519 5695
rect 15519 5661 15528 5695
rect 15476 5652 15528 5661
rect 13544 5559 13596 5568
rect 13544 5525 13553 5559
rect 13553 5525 13587 5559
rect 13587 5525 13596 5559
rect 13544 5516 13596 5525
rect 13820 5559 13872 5568
rect 13820 5525 13829 5559
rect 13829 5525 13863 5559
rect 13863 5525 13872 5559
rect 13820 5516 13872 5525
rect 15016 5516 15068 5568
rect 15936 5652 15988 5704
rect 17960 5516 18012 5568
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 2872 5312 2924 5364
rect 5632 5312 5684 5364
rect 7656 5312 7708 5364
rect 8300 5355 8352 5364
rect 8300 5321 8309 5355
rect 8309 5321 8343 5355
rect 8343 5321 8352 5355
rect 8300 5312 8352 5321
rect 8668 5312 8720 5364
rect 3056 5244 3108 5296
rect 6552 5244 6604 5296
rect 2688 5176 2740 5228
rect 3516 5176 3568 5228
rect 4712 5219 4764 5228
rect 4712 5185 4721 5219
rect 4721 5185 4755 5219
rect 4755 5185 4764 5219
rect 4712 5176 4764 5185
rect 11888 5312 11940 5364
rect 2780 5108 2832 5160
rect 3424 5108 3476 5160
rect 5632 5108 5684 5160
rect 8760 5151 8812 5160
rect 8760 5117 8769 5151
rect 8769 5117 8803 5151
rect 8803 5117 8812 5151
rect 8760 5108 8812 5117
rect 10784 5176 10836 5228
rect 12992 5219 13044 5228
rect 10232 5108 10284 5160
rect 12992 5185 13001 5219
rect 13001 5185 13035 5219
rect 13035 5185 13044 5219
rect 12992 5176 13044 5185
rect 16488 5176 16540 5228
rect 17408 5176 17460 5228
rect 13820 5108 13872 5160
rect 14372 5151 14424 5160
rect 14372 5117 14381 5151
rect 14381 5117 14415 5151
rect 14415 5117 14424 5151
rect 14372 5108 14424 5117
rect 7196 5083 7248 5092
rect 7196 5049 7230 5083
rect 7230 5049 7248 5083
rect 7196 5040 7248 5049
rect 7288 5040 7340 5092
rect 8392 5040 8444 5092
rect 11888 5083 11940 5092
rect 11888 5049 11897 5083
rect 11897 5049 11931 5083
rect 11931 5049 11940 5083
rect 11888 5040 11940 5049
rect 13268 5040 13320 5092
rect 13912 5083 13964 5092
rect 13912 5049 13921 5083
rect 13921 5049 13955 5083
rect 13955 5049 13964 5083
rect 13912 5040 13964 5049
rect 14556 5040 14608 5092
rect 1768 5015 1820 5024
rect 1768 4981 1777 5015
rect 1777 4981 1811 5015
rect 1811 4981 1820 5015
rect 1768 4972 1820 4981
rect 2136 5015 2188 5024
rect 2136 4981 2145 5015
rect 2145 4981 2179 5015
rect 2179 4981 2188 5015
rect 2136 4972 2188 4981
rect 2228 5015 2280 5024
rect 2228 4981 2237 5015
rect 2237 4981 2271 5015
rect 2271 4981 2280 5015
rect 2228 4972 2280 4981
rect 2504 4972 2556 5024
rect 3792 4972 3844 5024
rect 4160 5015 4212 5024
rect 4160 4981 4169 5015
rect 4169 4981 4203 5015
rect 4203 4981 4212 5015
rect 4160 4972 4212 4981
rect 5172 4972 5224 5024
rect 6092 5015 6144 5024
rect 6092 4981 6101 5015
rect 6101 4981 6135 5015
rect 6135 4981 6144 5015
rect 6092 4972 6144 4981
rect 6736 4972 6788 5024
rect 10600 4972 10652 5024
rect 10876 5015 10928 5024
rect 10876 4981 10885 5015
rect 10885 4981 10919 5015
rect 10919 4981 10928 5015
rect 10876 4972 10928 4981
rect 11704 4972 11756 5024
rect 12808 5015 12860 5024
rect 12808 4981 12817 5015
rect 12817 4981 12851 5015
rect 12851 4981 12860 5015
rect 12808 4972 12860 4981
rect 16580 4972 16632 5024
rect 16764 5015 16816 5024
rect 16764 4981 16773 5015
rect 16773 4981 16807 5015
rect 16807 4981 16816 5015
rect 16764 4972 16816 4981
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 2136 4768 2188 4820
rect 4160 4768 4212 4820
rect 5632 4768 5684 4820
rect 5724 4768 5776 4820
rect 7564 4768 7616 4820
rect 8484 4768 8536 4820
rect 13268 4768 13320 4820
rect 2688 4700 2740 4752
rect 4068 4700 4120 4752
rect 9772 4700 9824 4752
rect 10600 4700 10652 4752
rect 1400 4632 1452 4684
rect 4896 4675 4948 4684
rect 4896 4641 4905 4675
rect 4905 4641 4939 4675
rect 4939 4641 4948 4675
rect 4896 4632 4948 4641
rect 6552 4632 6604 4684
rect 6920 4675 6972 4684
rect 6920 4641 6929 4675
rect 6929 4641 6963 4675
rect 6963 4641 6972 4675
rect 6920 4632 6972 4641
rect 7656 4632 7708 4684
rect 11704 4675 11756 4684
rect 5356 4564 5408 4616
rect 5816 4496 5868 4548
rect 6276 4564 6328 4616
rect 7196 4607 7248 4616
rect 7196 4573 7205 4607
rect 7205 4573 7239 4607
rect 7239 4573 7248 4607
rect 7196 4564 7248 4573
rect 2412 4428 2464 4480
rect 3240 4428 3292 4480
rect 5080 4428 5132 4480
rect 5172 4428 5224 4480
rect 8392 4564 8444 4616
rect 8760 4564 8812 4616
rect 9588 4564 9640 4616
rect 11704 4641 11713 4675
rect 11713 4641 11747 4675
rect 11747 4641 11756 4675
rect 11704 4632 11756 4641
rect 12532 4564 12584 4616
rect 13728 4564 13780 4616
rect 14372 4607 14424 4616
rect 14372 4573 14381 4607
rect 14381 4573 14415 4607
rect 14415 4573 14424 4607
rect 14372 4564 14424 4573
rect 14648 4564 14700 4616
rect 15016 4564 15068 4616
rect 16120 4632 16172 4684
rect 16580 4632 16632 4684
rect 18604 4700 18656 4752
rect 17224 4607 17276 4616
rect 17224 4573 17233 4607
rect 17233 4573 17267 4607
rect 17267 4573 17276 4607
rect 17224 4564 17276 4573
rect 10876 4496 10928 4548
rect 7840 4471 7892 4480
rect 7840 4437 7849 4471
rect 7849 4437 7883 4471
rect 7883 4437 7892 4471
rect 7840 4428 7892 4437
rect 10048 4428 10100 4480
rect 14464 4428 14516 4480
rect 16488 4428 16540 4480
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 2412 4224 2464 4276
rect 4988 4224 5040 4276
rect 5816 4224 5868 4276
rect 6460 4267 6512 4276
rect 6460 4233 6469 4267
rect 6469 4233 6503 4267
rect 6503 4233 6512 4267
rect 6460 4224 6512 4233
rect 8208 4224 8260 4276
rect 1400 4088 1452 4140
rect 2412 4088 2464 4140
rect 4620 4156 4672 4208
rect 1768 4020 1820 4072
rect 3240 4063 3292 4072
rect 3240 4029 3274 4063
rect 3274 4029 3292 4063
rect 3240 4020 3292 4029
rect 3792 4020 3844 4072
rect 6920 4131 6972 4140
rect 6920 4097 6929 4131
rect 6929 4097 6963 4131
rect 6963 4097 6972 4131
rect 6920 4088 6972 4097
rect 7840 4088 7892 4140
rect 8392 4088 8444 4140
rect 11796 4224 11848 4276
rect 13268 4224 13320 4276
rect 4528 4020 4580 4072
rect 5264 3952 5316 4004
rect 5632 3952 5684 4004
rect 6000 3952 6052 4004
rect 2044 3884 2096 3936
rect 4160 3884 4212 3936
rect 4712 3884 4764 3936
rect 6828 3884 6880 3936
rect 8392 3952 8444 4004
rect 8668 4020 8720 4072
rect 9588 4020 9640 4072
rect 12808 4088 12860 4140
rect 14372 4224 14424 4276
rect 14740 4224 14792 4276
rect 16120 4224 16172 4276
rect 16764 4224 16816 4276
rect 16488 4156 16540 4208
rect 14648 4088 14700 4140
rect 10048 4063 10100 4072
rect 10048 4029 10082 4063
rect 10082 4029 10100 4063
rect 10048 4020 10100 4029
rect 12348 4020 12400 4072
rect 12716 4020 12768 4072
rect 13268 4063 13320 4072
rect 13268 4029 13277 4063
rect 13277 4029 13311 4063
rect 13311 4029 13320 4063
rect 13268 4020 13320 4029
rect 15016 4020 15068 4072
rect 12624 3952 12676 4004
rect 13820 3952 13872 4004
rect 8300 3884 8352 3936
rect 8760 3927 8812 3936
rect 8760 3893 8769 3927
rect 8769 3893 8803 3927
rect 8803 3893 8812 3927
rect 8760 3884 8812 3893
rect 9312 3884 9364 3936
rect 9588 3884 9640 3936
rect 10600 3884 10652 3936
rect 11152 3927 11204 3936
rect 11152 3893 11161 3927
rect 11161 3893 11195 3927
rect 11195 3893 11204 3927
rect 11152 3884 11204 3893
rect 11244 3884 11296 3936
rect 16212 3952 16264 4004
rect 14280 3884 14332 3936
rect 17040 3927 17092 3936
rect 17040 3893 17049 3927
rect 17049 3893 17083 3927
rect 17083 3893 17092 3927
rect 17040 3884 17092 3893
rect 21180 3884 21232 3936
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 1032 3680 1084 3732
rect 2964 3680 3016 3732
rect 4896 3680 4948 3732
rect 6092 3680 6144 3732
rect 6828 3723 6880 3732
rect 6828 3689 6837 3723
rect 6837 3689 6871 3723
rect 6871 3689 6880 3723
rect 6828 3680 6880 3689
rect 8668 3680 8720 3732
rect 8760 3680 8812 3732
rect 1952 3612 2004 3664
rect 3792 3612 3844 3664
rect 3976 3612 4028 3664
rect 11244 3680 11296 3732
rect 13820 3723 13872 3732
rect 1400 3544 1452 3596
rect 3516 3544 3568 3596
rect 3884 3544 3936 3596
rect 4528 3587 4580 3596
rect 4528 3553 4537 3587
rect 4537 3553 4571 3587
rect 4571 3553 4580 3587
rect 4528 3544 4580 3553
rect 5356 3544 5408 3596
rect 6736 3587 6788 3596
rect 6736 3553 6745 3587
rect 6745 3553 6779 3587
rect 6779 3553 6788 3587
rect 6736 3544 6788 3553
rect 7656 3544 7708 3596
rect 6460 3476 6512 3528
rect 7288 3476 7340 3528
rect 572 3340 624 3392
rect 3976 3408 4028 3460
rect 11152 3612 11204 3664
rect 11980 3612 12032 3664
rect 13820 3689 13829 3723
rect 13829 3689 13863 3723
rect 13863 3689 13872 3723
rect 13820 3680 13872 3689
rect 14464 3680 14516 3732
rect 12072 3544 12124 3596
rect 10600 3476 10652 3528
rect 11796 3476 11848 3528
rect 14280 3544 14332 3596
rect 14464 3587 14516 3596
rect 14464 3553 14473 3587
rect 14473 3553 14507 3587
rect 14507 3553 14516 3587
rect 14464 3544 14516 3553
rect 12348 3476 12400 3528
rect 13452 3476 13504 3528
rect 15752 3587 15804 3596
rect 15752 3553 15761 3587
rect 15761 3553 15795 3587
rect 15795 3553 15804 3587
rect 15752 3544 15804 3553
rect 16120 3612 16172 3664
rect 16212 3612 16264 3664
rect 17224 3587 17276 3596
rect 17224 3553 17233 3587
rect 17233 3553 17267 3587
rect 17267 3553 17276 3587
rect 17224 3544 17276 3553
rect 17776 3587 17828 3596
rect 17776 3553 17785 3587
rect 17785 3553 17819 3587
rect 17819 3553 17828 3587
rect 17776 3544 17828 3553
rect 16672 3519 16724 3528
rect 16672 3485 16681 3519
rect 16681 3485 16715 3519
rect 16715 3485 16724 3519
rect 16672 3476 16724 3485
rect 2688 3340 2740 3392
rect 3240 3340 3292 3392
rect 5172 3340 5224 3392
rect 5264 3340 5316 3392
rect 6000 3340 6052 3392
rect 6920 3340 6972 3392
rect 8116 3340 8168 3392
rect 9496 3340 9548 3392
rect 13636 3340 13688 3392
rect 15660 3340 15712 3392
rect 17684 3340 17736 3392
rect 18604 3340 18656 3392
rect 20812 3340 20864 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 2412 3136 2464 3188
rect 3884 3136 3936 3188
rect 13452 3136 13504 3188
rect 15752 3136 15804 3188
rect 3516 3111 3568 3120
rect 3516 3077 3525 3111
rect 3525 3077 3559 3111
rect 3559 3077 3568 3111
rect 3516 3068 3568 3077
rect 4896 3068 4948 3120
rect 5172 3068 5224 3120
rect 5356 3068 5408 3120
rect 1860 3000 1912 3052
rect 3884 3043 3936 3052
rect 3884 3009 3893 3043
rect 3893 3009 3927 3043
rect 3927 3009 3936 3043
rect 3884 3000 3936 3009
rect 4988 3000 5040 3052
rect 6000 3068 6052 3120
rect 9772 3111 9824 3120
rect 9772 3077 9781 3111
rect 9781 3077 9815 3111
rect 9815 3077 9824 3111
rect 9772 3068 9824 3077
rect 10324 3068 10376 3120
rect 3792 2932 3844 2984
rect 4160 2975 4212 2984
rect 4160 2941 4194 2975
rect 4194 2941 4212 2975
rect 9496 3043 9548 3052
rect 9496 3009 9505 3043
rect 9505 3009 9539 3043
rect 9539 3009 9548 3043
rect 9496 3000 9548 3009
rect 9680 3000 9732 3052
rect 10416 3043 10468 3052
rect 10416 3009 10425 3043
rect 10425 3009 10459 3043
rect 10459 3009 10468 3043
rect 10416 3000 10468 3009
rect 10600 3043 10652 3052
rect 10600 3009 10609 3043
rect 10609 3009 10643 3043
rect 10643 3009 10652 3043
rect 10600 3000 10652 3009
rect 10876 3000 10928 3052
rect 12532 3068 12584 3120
rect 15936 3068 15988 3120
rect 7288 2975 7340 2984
rect 4160 2932 4212 2941
rect 7288 2941 7297 2975
rect 7297 2941 7331 2975
rect 7331 2941 7340 2975
rect 7288 2932 7340 2941
rect 8116 2932 8168 2984
rect 8760 2932 8812 2984
rect 11980 3043 12032 3052
rect 11980 3009 11989 3043
rect 11989 3009 12023 3043
rect 12023 3009 12032 3043
rect 11980 3000 12032 3009
rect 13636 3000 13688 3052
rect 204 2864 256 2916
rect 3056 2864 3108 2916
rect 1492 2796 1544 2848
rect 3424 2796 3476 2848
rect 3608 2796 3660 2848
rect 3976 2796 4028 2848
rect 4068 2796 4120 2848
rect 5632 2796 5684 2848
rect 7380 2864 7432 2916
rect 6092 2839 6144 2848
rect 6092 2805 6101 2839
rect 6101 2805 6135 2839
rect 6135 2805 6144 2839
rect 6092 2796 6144 2805
rect 7012 2796 7064 2848
rect 7288 2796 7340 2848
rect 8668 2839 8720 2848
rect 8668 2805 8677 2839
rect 8677 2805 8711 2839
rect 8711 2805 8720 2839
rect 8668 2796 8720 2805
rect 8944 2839 8996 2848
rect 8944 2805 8953 2839
rect 8953 2805 8987 2839
rect 8987 2805 8996 2839
rect 8944 2796 8996 2805
rect 10508 2864 10560 2916
rect 11980 2864 12032 2916
rect 12440 2975 12492 2984
rect 12440 2941 12449 2975
rect 12449 2941 12483 2975
rect 12483 2941 12492 2975
rect 12440 2932 12492 2941
rect 13728 2975 13780 2984
rect 13728 2941 13737 2975
rect 13737 2941 13771 2975
rect 13771 2941 13780 2975
rect 13728 2932 13780 2941
rect 15660 2975 15712 2984
rect 15660 2941 15669 2975
rect 15669 2941 15703 2975
rect 15703 2941 15712 2975
rect 15660 2932 15712 2941
rect 16396 2975 16448 2984
rect 16396 2941 16405 2975
rect 16405 2941 16439 2975
rect 16439 2941 16448 2975
rect 16396 2932 16448 2941
rect 21640 2932 21692 2984
rect 12256 2796 12308 2848
rect 13360 2839 13412 2848
rect 13360 2805 13369 2839
rect 13369 2805 13403 2839
rect 13403 2805 13412 2839
rect 13360 2796 13412 2805
rect 13728 2796 13780 2848
rect 14188 2796 14240 2848
rect 22560 2864 22612 2916
rect 16028 2796 16080 2848
rect 16856 2796 16908 2848
rect 22100 2796 22152 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 2044 2592 2096 2644
rect 2596 2592 2648 2644
rect 3424 2635 3476 2644
rect 2504 2524 2556 2576
rect 3424 2601 3433 2635
rect 3433 2601 3467 2635
rect 3467 2601 3476 2635
rect 3424 2592 3476 2601
rect 4896 2592 4948 2644
rect 5080 2592 5132 2644
rect 7380 2635 7432 2644
rect 7380 2601 7389 2635
rect 7389 2601 7423 2635
rect 7423 2601 7432 2635
rect 7380 2592 7432 2601
rect 8392 2635 8444 2644
rect 8392 2601 8401 2635
rect 8401 2601 8435 2635
rect 8435 2601 8444 2635
rect 8392 2592 8444 2601
rect 8944 2592 8996 2644
rect 9772 2635 9824 2644
rect 9772 2601 9781 2635
rect 9781 2601 9815 2635
rect 9815 2601 9824 2635
rect 9772 2592 9824 2601
rect 10140 2592 10192 2644
rect 10784 2592 10836 2644
rect 12072 2635 12124 2644
rect 12072 2601 12081 2635
rect 12081 2601 12115 2635
rect 12115 2601 12124 2635
rect 12072 2592 12124 2601
rect 14464 2592 14516 2644
rect 8300 2524 8352 2576
rect 3424 2456 3476 2508
rect 3884 2456 3936 2508
rect 5172 2456 5224 2508
rect 5356 2456 5408 2508
rect 12440 2524 12492 2576
rect 2320 2388 2372 2440
rect 2688 2388 2740 2440
rect 4160 2388 4212 2440
rect 5264 2388 5316 2440
rect 9680 2456 9732 2508
rect 12624 2499 12676 2508
rect 8668 2431 8720 2440
rect 8668 2397 8677 2431
rect 8677 2397 8711 2431
rect 8711 2397 8720 2431
rect 8668 2388 8720 2397
rect 10600 2388 10652 2440
rect 12624 2465 12633 2499
rect 12633 2465 12667 2499
rect 12667 2465 12676 2499
rect 12624 2456 12676 2465
rect 13912 2456 13964 2508
rect 14556 2456 14608 2508
rect 15476 2499 15528 2508
rect 15476 2465 15485 2499
rect 15485 2465 15519 2499
rect 15519 2465 15528 2499
rect 15476 2456 15528 2465
rect 16028 2499 16080 2508
rect 16028 2465 16037 2499
rect 16037 2465 16071 2499
rect 16071 2465 16080 2499
rect 16028 2456 16080 2465
rect 16672 2499 16724 2508
rect 16672 2465 16681 2499
rect 16681 2465 16715 2499
rect 16715 2465 16724 2499
rect 16672 2456 16724 2465
rect 7012 2252 7064 2304
rect 10140 2252 10192 2304
rect 12440 2252 12492 2304
rect 12900 2252 12952 2304
rect 14648 2252 14700 2304
rect 15108 2252 15160 2304
rect 15476 2252 15528 2304
rect 16396 2252 16448 2304
rect 17316 2252 17368 2304
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 2872 1844 2924 1896
rect 4712 1844 4764 1896
rect 3332 892 3384 944
rect 6184 892 6236 944
<< metal2 >>
rect 3974 22536 4030 22545
rect 3974 22471 4030 22480
rect 3054 22128 3110 22137
rect 3054 22063 3110 22072
rect 2870 21176 2926 21185
rect 2870 21111 2926 21120
rect 2778 20632 2834 20641
rect 2778 20567 2834 20576
rect 1950 20224 2006 20233
rect 1950 20159 2006 20168
rect 1964 20058 1992 20159
rect 1952 20052 2004 20058
rect 1952 19994 2004 20000
rect 2228 19916 2280 19922
rect 2228 19858 2280 19864
rect 2044 19304 2096 19310
rect 2044 19246 2096 19252
rect 1858 18320 1914 18329
rect 1858 18255 1914 18264
rect 1872 17882 1900 18255
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 1964 17921 1992 18022
rect 1950 17912 2006 17921
rect 1860 17876 1912 17882
rect 1950 17847 2006 17856
rect 1860 17818 1912 17824
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 1768 16992 1820 16998
rect 1766 16960 1768 16969
rect 1820 16960 1822 16969
rect 1766 16895 1822 16904
rect 1492 16040 1544 16046
rect 1492 15982 1544 15988
rect 1504 14550 1532 15982
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1688 15609 1716 15846
rect 1964 15638 1992 17070
rect 2056 16726 2084 19246
rect 2240 18766 2268 19858
rect 2320 19304 2372 19310
rect 2320 19246 2372 19252
rect 2332 18902 2360 19246
rect 2792 19174 2820 20567
rect 2884 19242 2912 21111
rect 2872 19236 2924 19242
rect 2872 19178 2924 19184
rect 2780 19168 2832 19174
rect 2780 19110 2832 19116
rect 2320 18896 2372 18902
rect 2320 18838 2372 18844
rect 2778 18864 2834 18873
rect 2778 18799 2834 18808
rect 2228 18760 2280 18766
rect 2228 18702 2280 18708
rect 2792 18426 2820 18799
rect 3068 18426 3096 22063
rect 3606 21584 3662 21593
rect 3606 21519 3662 21528
rect 3620 18426 3648 21519
rect 3698 19816 3754 19825
rect 3698 19751 3754 19760
rect 3712 19514 3740 19751
rect 3700 19508 3752 19514
rect 3700 19450 3752 19456
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 2332 17814 2360 18158
rect 2412 18148 2464 18154
rect 2412 18090 2464 18096
rect 2320 17808 2372 17814
rect 2320 17750 2372 17756
rect 2424 17134 2452 18090
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 3068 17202 3096 17614
rect 3790 17368 3846 17377
rect 3790 17303 3792 17312
rect 3844 17303 3846 17312
rect 3792 17274 3844 17280
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 2412 17128 2464 17134
rect 2412 17070 2464 17076
rect 2688 17060 2740 17066
rect 2688 17002 2740 17008
rect 2044 16720 2096 16726
rect 2044 16662 2096 16668
rect 2700 16658 2728 17002
rect 2688 16652 2740 16658
rect 2688 16594 2740 16600
rect 3148 16652 3200 16658
rect 3148 16594 3200 16600
rect 3608 16652 3660 16658
rect 3608 16594 3660 16600
rect 2872 16176 2924 16182
rect 2872 16118 2924 16124
rect 2780 16040 2832 16046
rect 2780 15982 2832 15988
rect 1952 15632 2004 15638
rect 1674 15600 1730 15609
rect 1952 15574 2004 15580
rect 1674 15535 1730 15544
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 1768 15360 1820 15366
rect 1768 15302 1820 15308
rect 1780 15065 1808 15302
rect 1766 15056 1822 15065
rect 1766 14991 1822 15000
rect 1952 14952 2004 14958
rect 1952 14894 2004 14900
rect 1676 14816 1728 14822
rect 1676 14758 1728 14764
rect 1688 14657 1716 14758
rect 1674 14648 1730 14657
rect 1674 14583 1730 14592
rect 1492 14544 1544 14550
rect 1492 14486 1544 14492
rect 1582 14104 1638 14113
rect 1582 14039 1638 14048
rect 1492 13320 1544 13326
rect 1492 13262 1544 13268
rect 1504 12306 1532 13262
rect 1596 12442 1624 14039
rect 1768 13864 1820 13870
rect 1768 13806 1820 13812
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1492 12300 1544 12306
rect 1492 12242 1544 12248
rect 1584 11688 1636 11694
rect 1584 11630 1636 11636
rect 1596 10674 1624 11630
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1584 9512 1636 9518
rect 1584 9454 1636 9460
rect 1596 8838 1624 9454
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1688 8634 1716 13330
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1780 7546 1808 13806
rect 1964 12850 1992 14894
rect 2516 13870 2544 15438
rect 2792 15094 2820 15982
rect 2780 15088 2832 15094
rect 2780 15030 2832 15036
rect 2884 14958 2912 16118
rect 3160 16114 3188 16594
rect 3330 16552 3386 16561
rect 3330 16487 3332 16496
rect 3384 16487 3386 16496
rect 3332 16458 3384 16464
rect 3620 16114 3648 16594
rect 3148 16108 3200 16114
rect 3148 16050 3200 16056
rect 3608 16108 3660 16114
rect 3608 16050 3660 16056
rect 2962 16008 3018 16017
rect 2962 15943 3018 15952
rect 2976 15910 3004 15943
rect 2964 15904 3016 15910
rect 2964 15846 3016 15852
rect 3332 15496 3384 15502
rect 3332 15438 3384 15444
rect 3516 15496 3568 15502
rect 3516 15438 3568 15444
rect 2872 14952 2924 14958
rect 2872 14894 2924 14900
rect 2884 14278 2912 14894
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 2504 13864 2556 13870
rect 2504 13806 2556 13812
rect 2884 13802 2912 14214
rect 3344 14074 3372 15438
rect 3528 14890 3556 15438
rect 3516 14884 3568 14890
rect 3516 14826 3568 14832
rect 3528 14618 3556 14826
rect 3516 14612 3568 14618
rect 3988 14600 4016 22471
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 6828 19304 6880 19310
rect 4066 19272 4122 19281
rect 6828 19246 6880 19252
rect 4066 19207 4122 19216
rect 4080 18970 4108 19207
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 6840 18902 6868 19246
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 6828 18896 6880 18902
rect 6828 18838 6880 18844
rect 7656 18828 7708 18834
rect 7656 18770 7708 18776
rect 8208 18828 8260 18834
rect 8208 18770 8260 18776
rect 7196 18692 7248 18698
rect 7196 18634 7248 18640
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 7012 17740 7064 17746
rect 7012 17682 7064 17688
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 6184 17196 6236 17202
rect 6184 17138 6236 17144
rect 5724 17060 5776 17066
rect 5724 17002 5776 17008
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 4068 16720 4120 16726
rect 4068 16662 4120 16668
rect 4080 15706 4108 16662
rect 4172 15706 4200 16934
rect 4988 16652 5040 16658
rect 4988 16594 5040 16600
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 5000 16250 5028 16594
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 4252 15972 4304 15978
rect 4252 15914 4304 15920
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4264 15162 4292 15914
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4712 15564 4764 15570
rect 4712 15506 4764 15512
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4724 15162 4752 15506
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 4712 15156 4764 15162
rect 4712 15098 4764 15104
rect 4816 14618 4844 15846
rect 5000 15502 5028 16186
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 5736 15162 5764 17002
rect 5908 16992 5960 16998
rect 5908 16934 5960 16940
rect 6000 16992 6052 16998
rect 6000 16934 6052 16940
rect 5920 16114 5948 16934
rect 6012 16250 6040 16934
rect 6196 16794 6224 17138
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 6092 16584 6144 16590
rect 6092 16526 6144 16532
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 5908 16108 5960 16114
rect 5908 16050 5960 16056
rect 6104 15586 6132 16526
rect 6196 15638 6224 16730
rect 6276 16720 6328 16726
rect 6276 16662 6328 16668
rect 6288 16114 6316 16662
rect 6276 16108 6328 16114
rect 6276 16050 6328 16056
rect 6828 15972 6880 15978
rect 6828 15914 6880 15920
rect 6276 15904 6328 15910
rect 6276 15846 6328 15852
rect 6288 15706 6316 15846
rect 6276 15700 6328 15706
rect 6276 15642 6328 15648
rect 6552 15700 6604 15706
rect 6552 15642 6604 15648
rect 6012 15570 6132 15586
rect 6184 15632 6236 15638
rect 6184 15574 6236 15580
rect 6000 15564 6132 15570
rect 6052 15558 6132 15564
rect 6000 15506 6052 15512
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 5276 14822 5304 14962
rect 5724 14952 5776 14958
rect 5724 14894 5776 14900
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 3516 14554 3568 14560
rect 3896 14572 4016 14600
rect 4804 14612 4856 14618
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 3424 13932 3476 13938
rect 3424 13874 3476 13880
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 2872 13796 2924 13802
rect 2872 13738 2924 13744
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2412 13184 2464 13190
rect 2412 13126 2464 13132
rect 1952 12844 2004 12850
rect 1952 12786 2004 12792
rect 1860 12776 1912 12782
rect 1860 12718 1912 12724
rect 1872 12442 1900 12718
rect 2424 12442 2452 13126
rect 2688 12776 2740 12782
rect 2688 12718 2740 12724
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 2412 12436 2464 12442
rect 2412 12378 2464 12384
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2516 11898 2544 12174
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2700 11626 2728 12718
rect 2792 11626 2820 13330
rect 2884 12782 2912 13738
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 3238 13288 3294 13297
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2688 11620 2740 11626
rect 2688 11562 2740 11568
rect 2780 11620 2832 11626
rect 2780 11562 2832 11568
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2332 11354 2360 11494
rect 2884 11354 2912 12038
rect 2976 11694 3004 13262
rect 3238 13223 3294 13232
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 2964 11688 3016 11694
rect 2964 11630 3016 11636
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 2688 11076 2740 11082
rect 2688 11018 2740 11024
rect 2700 10606 2728 11018
rect 2884 10690 2912 11290
rect 2976 10810 3004 11630
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 2884 10662 3004 10690
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2700 10198 2728 10542
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2688 10192 2740 10198
rect 2688 10134 2740 10140
rect 2700 9722 2728 10134
rect 2792 10062 2820 10406
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2870 10024 2926 10033
rect 2870 9959 2926 9968
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2320 9444 2372 9450
rect 2320 9386 2372 9392
rect 2780 9444 2832 9450
rect 2780 9386 2832 9392
rect 2332 8498 2360 9386
rect 2792 9178 2820 9386
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2504 9036 2556 9042
rect 2504 8978 2556 8984
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2136 8288 2188 8294
rect 2228 8288 2280 8294
rect 2136 8230 2188 8236
rect 2226 8256 2228 8265
rect 2280 8256 2282 8265
rect 2148 8090 2176 8230
rect 2226 8191 2282 8200
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 2516 7886 2544 8978
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 2608 8412 2636 8774
rect 2780 8424 2832 8430
rect 2608 8384 2780 8412
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2700 7818 2728 8384
rect 2780 8366 2832 8372
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 2792 7886 2820 8230
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2688 7812 2740 7818
rect 2688 7754 2740 7760
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 1584 7268 1636 7274
rect 1584 7210 1636 7216
rect 1308 6996 1360 7002
rect 1308 6938 1360 6944
rect 1032 3732 1084 3738
rect 1032 3674 1084 3680
rect 572 3392 624 3398
rect 572 3334 624 3340
rect 204 2916 256 2922
rect 204 2858 256 2864
rect 216 480 244 2858
rect 584 480 612 3334
rect 1044 480 1072 3674
rect 1320 2009 1348 6938
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1412 4690 1440 6190
rect 1596 5914 1624 7210
rect 2516 6866 2544 7346
rect 2700 6934 2728 7754
rect 2688 6928 2740 6934
rect 2688 6870 2740 6876
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 1860 6792 1912 6798
rect 1860 6734 1912 6740
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1676 5704 1728 5710
rect 1676 5646 1728 5652
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1412 4146 1440 4626
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1412 3602 1440 4082
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 1688 2961 1716 5646
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1780 4078 1808 4966
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1872 3058 1900 6734
rect 2516 6458 2544 6802
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2780 6180 2832 6186
rect 2780 6122 2832 6128
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 1964 5914 1992 6054
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 2792 5642 2820 6122
rect 2780 5636 2832 5642
rect 2780 5578 2832 5584
rect 2596 5568 2648 5574
rect 2596 5510 2648 5516
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 2148 4826 2176 4966
rect 2240 4865 2268 4966
rect 2226 4856 2282 4865
rect 2136 4820 2188 4826
rect 2226 4791 2282 4800
rect 2136 4762 2188 4768
rect 2412 4480 2464 4486
rect 2412 4422 2464 4428
rect 2424 4282 2452 4422
rect 2412 4276 2464 4282
rect 2412 4218 2464 4224
rect 2412 4140 2464 4146
rect 2412 4082 2464 4088
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 1952 3664 2004 3670
rect 1952 3606 2004 3612
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 1674 2952 1730 2961
rect 1674 2887 1730 2896
rect 1492 2848 1544 2854
rect 1492 2790 1544 2796
rect 1306 2000 1362 2009
rect 1306 1935 1362 1944
rect 1504 480 1532 2790
rect 1964 480 1992 3606
rect 2056 2650 2084 3878
rect 2424 3194 2452 4082
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 2044 2644 2096 2650
rect 2044 2586 2096 2592
rect 2516 2582 2544 4966
rect 2608 2650 2636 5510
rect 2884 5370 2912 9959
rect 2976 6866 3004 10662
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 3068 10266 3096 10542
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 2964 6860 3016 6866
rect 2964 6802 3016 6808
rect 2964 5772 3016 5778
rect 2964 5714 3016 5720
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2688 5228 2740 5234
rect 2688 5170 2740 5176
rect 2700 4758 2728 5170
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2688 4752 2740 4758
rect 2688 4694 2740 4700
rect 2700 3398 2728 4694
rect 2792 3641 2820 5102
rect 2976 3738 3004 5714
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 3068 5302 3096 5646
rect 3160 5642 3188 13126
rect 3252 12442 3280 13223
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 3240 11620 3292 11626
rect 3240 11562 3292 11568
rect 3252 11354 3280 11562
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3240 11212 3292 11218
rect 3240 11154 3292 11160
rect 3252 11082 3280 11154
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 3252 6934 3280 11018
rect 3344 10810 3372 13806
rect 3436 13394 3464 13874
rect 3700 13864 3752 13870
rect 3700 13806 3752 13812
rect 3606 13696 3662 13705
rect 3606 13631 3662 13640
rect 3620 13530 3648 13631
rect 3608 13524 3660 13530
rect 3608 13466 3660 13472
rect 3424 13388 3476 13394
rect 3424 13330 3476 13336
rect 3422 12744 3478 12753
rect 3422 12679 3478 12688
rect 3516 12708 3568 12714
rect 3436 12374 3464 12679
rect 3516 12650 3568 12656
rect 3424 12368 3476 12374
rect 3424 12310 3476 12316
rect 3528 12238 3556 12650
rect 3608 12300 3660 12306
rect 3608 12242 3660 12248
rect 3516 12232 3568 12238
rect 3516 12174 3568 12180
rect 3528 11830 3556 12174
rect 3516 11824 3568 11830
rect 3516 11766 3568 11772
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3436 10470 3464 11698
rect 3620 11558 3648 12242
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3712 10198 3740 13806
rect 3700 10192 3752 10198
rect 3700 10134 3752 10140
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3528 9518 3556 9998
rect 3896 9738 3924 14572
rect 4804 14554 4856 14560
rect 4252 14544 4304 14550
rect 4252 14486 4304 14492
rect 3976 14476 4028 14482
rect 3976 14418 4028 14424
rect 3988 14074 4016 14418
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 4068 13796 4120 13802
rect 4068 13738 4120 13744
rect 4080 13394 4108 13738
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 4080 13274 4108 13330
rect 4080 13246 4200 13274
rect 4172 12646 4200 13246
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4172 12442 4200 12582
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4066 12336 4122 12345
rect 4066 12271 4122 12280
rect 4080 11898 4108 12271
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4264 11354 4292 14486
rect 4896 14408 4948 14414
rect 4896 14350 4948 14356
rect 5080 14408 5132 14414
rect 5080 14350 5132 14356
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4712 12912 4764 12918
rect 4712 12854 4764 12860
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 4080 10849 4108 10950
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4066 10840 4122 10849
rect 4388 10832 4684 10852
rect 4066 10775 4122 10784
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4066 10432 4122 10441
rect 4066 10367 4122 10376
rect 4080 9926 4108 10367
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 3887 9722 3924 9738
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3804 8430 3832 9658
rect 3882 9480 3938 9489
rect 3882 9415 3938 9424
rect 3792 8424 3844 8430
rect 3792 8366 3844 8372
rect 3700 7812 3752 7818
rect 3700 7754 3752 7760
rect 3712 7410 3740 7754
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3700 7404 3752 7410
rect 3700 7346 3752 7352
rect 3424 7268 3476 7274
rect 3424 7210 3476 7216
rect 3436 7002 3464 7210
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 3240 6928 3292 6934
rect 3240 6870 3292 6876
rect 3332 6860 3384 6866
rect 3332 6802 3384 6808
rect 3148 5636 3200 5642
rect 3148 5578 3200 5584
rect 3056 5296 3108 5302
rect 3056 5238 3108 5244
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2778 3632 2834 3641
rect 2778 3567 2834 3576
rect 2688 3392 2740 3398
rect 2688 3334 2740 3340
rect 2596 2644 2648 2650
rect 2596 2586 2648 2592
rect 2504 2576 2556 2582
rect 2504 2518 2556 2524
rect 2700 2446 2728 3334
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 2688 2440 2740 2446
rect 2688 2382 2740 2388
rect 2332 480 2360 2382
rect 2792 480 2820 3567
rect 3068 2922 3096 5238
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3252 4078 3280 4422
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 3056 2916 3108 2922
rect 3056 2858 3108 2864
rect 2872 1896 2924 1902
rect 2872 1838 2924 1844
rect 2884 1601 2912 1838
rect 2870 1592 2926 1601
rect 2870 1527 2926 1536
rect 3252 480 3280 3334
rect 3344 1057 3372 6802
rect 3528 5914 3556 7142
rect 3620 6118 3648 7346
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3422 5264 3478 5273
rect 3528 5234 3556 5646
rect 3422 5199 3478 5208
rect 3516 5228 3568 5234
rect 3436 5166 3464 5199
rect 3516 5170 3568 5176
rect 3424 5160 3476 5166
rect 3424 5102 3476 5108
rect 3528 3602 3556 5170
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 3528 3126 3556 3538
rect 3516 3120 3568 3126
rect 3516 3062 3568 3068
rect 3620 2854 3648 5714
rect 3700 5704 3752 5710
rect 3896 5681 3924 9415
rect 3976 8900 4028 8906
rect 3976 8842 4028 8848
rect 3988 8537 4016 8842
rect 3974 8528 4030 8537
rect 3974 8463 4030 8472
rect 4158 8392 4214 8401
rect 4158 8327 4214 8336
rect 4172 8294 4200 8327
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 3974 8120 4030 8129
rect 3974 8055 4030 8064
rect 3988 7274 4016 8055
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4066 7576 4122 7585
rect 4066 7511 4068 7520
rect 4120 7511 4122 7520
rect 4068 7482 4120 7488
rect 3976 7268 4028 7274
rect 3976 7210 4028 7216
rect 4066 6760 4122 6769
rect 4066 6695 4122 6704
rect 4080 6458 4108 6695
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4172 6338 4200 7822
rect 3988 6310 4200 6338
rect 3700 5646 3752 5652
rect 3882 5672 3938 5681
rect 3424 2848 3476 2854
rect 3424 2790 3476 2796
rect 3608 2848 3660 2854
rect 3608 2790 3660 2796
rect 3436 2650 3464 2790
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 3436 2417 3464 2450
rect 3422 2408 3478 2417
rect 3422 2343 3478 2352
rect 3330 1048 3386 1057
rect 3330 983 3386 992
rect 3332 944 3384 950
rect 3332 886 3384 892
rect 3344 649 3372 886
rect 3330 640 3386 649
rect 3330 575 3386 584
rect 3712 480 3740 5646
rect 3882 5607 3938 5616
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3804 4078 3832 4966
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3988 4026 4016 6310
rect 4066 6216 4122 6225
rect 4066 6151 4122 6160
rect 4080 5930 4108 6151
rect 4080 5914 4200 5930
rect 4080 5908 4212 5914
rect 4080 5902 4160 5908
rect 4160 5850 4212 5856
rect 4066 5808 4122 5817
rect 4066 5743 4122 5752
rect 4080 5574 4108 5743
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4172 4826 4200 4966
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4068 4752 4120 4758
rect 4068 4694 4120 4700
rect 4080 4321 4108 4694
rect 4066 4312 4122 4321
rect 4066 4247 4122 4256
rect 3804 3670 3832 4014
rect 3988 3998 4108 4026
rect 3974 3904 4030 3913
rect 3974 3839 4030 3848
rect 3988 3670 4016 3839
rect 3792 3664 3844 3670
rect 3792 3606 3844 3612
rect 3976 3664 4028 3670
rect 3976 3606 4028 3612
rect 3884 3596 3936 3602
rect 3884 3538 3936 3544
rect 3896 3194 3924 3538
rect 4080 3505 4108 3998
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 4066 3496 4122 3505
rect 3976 3460 4028 3466
rect 4066 3431 4122 3440
rect 3976 3402 4028 3408
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3896 3058 3924 3130
rect 3988 3097 4016 3402
rect 3974 3088 4030 3097
rect 3884 3052 3936 3058
rect 3974 3023 4030 3032
rect 3884 2994 3936 3000
rect 4172 2990 4200 3878
rect 3792 2984 3844 2990
rect 3792 2926 3844 2932
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 3804 2825 3832 2926
rect 3976 2848 4028 2854
rect 3790 2816 3846 2825
rect 3976 2790 4028 2796
rect 4068 2848 4120 2854
rect 4068 2790 4120 2796
rect 3790 2751 3846 2760
rect 3882 2544 3938 2553
rect 3882 2479 3884 2488
rect 3936 2479 3938 2488
rect 3884 2450 3936 2456
rect 202 0 258 480
rect 570 0 626 480
rect 1030 0 1086 480
rect 1490 0 1546 480
rect 1950 0 2006 480
rect 2318 0 2374 480
rect 2778 0 2834 480
rect 3238 0 3294 480
rect 3698 0 3754 480
rect 3988 241 4016 2790
rect 4080 480 4108 2790
rect 4172 2446 4200 2926
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 4264 1986 4292 10202
rect 4356 10130 4384 10610
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4724 9518 4752 12854
rect 4816 12850 4844 13330
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 4804 12708 4856 12714
rect 4804 12650 4856 12656
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4448 9178 4476 9318
rect 4436 9172 4488 9178
rect 4436 9114 4488 9120
rect 4724 9110 4752 9454
rect 4816 9382 4844 12650
rect 4908 12442 4936 14350
rect 5092 13802 5120 14350
rect 5080 13796 5132 13802
rect 5080 13738 5132 13744
rect 5092 13530 5120 13738
rect 5080 13524 5132 13530
rect 5080 13466 5132 13472
rect 5172 13456 5224 13462
rect 5172 13398 5224 13404
rect 5184 12986 5212 13398
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 4988 12776 5040 12782
rect 4988 12718 5040 12724
rect 5000 12646 5028 12718
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 4896 12436 4948 12442
rect 4896 12378 4948 12384
rect 4894 12336 4950 12345
rect 4894 12271 4896 12280
rect 4948 12271 4950 12280
rect 5000 12322 5028 12582
rect 5080 12368 5132 12374
rect 5000 12316 5080 12322
rect 5000 12310 5132 12316
rect 5000 12294 5120 12310
rect 4896 12242 4948 12248
rect 4908 12102 4936 12242
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 5000 11778 5028 12294
rect 5184 12238 5212 12922
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 4908 11750 5028 11778
rect 4908 11694 4936 11750
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4908 10674 4936 11630
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 4896 10124 4948 10130
rect 4896 10066 4948 10072
rect 4908 9722 4936 10066
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 5000 9654 5028 11086
rect 5276 11082 5304 14758
rect 5356 13728 5408 13734
rect 5356 13670 5408 13676
rect 5368 13462 5396 13670
rect 5736 13530 5764 14894
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5828 14618 5856 14758
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 6104 14482 6132 15558
rect 6368 15020 6420 15026
rect 6368 14962 6420 14968
rect 6380 14618 6408 14962
rect 6368 14612 6420 14618
rect 6368 14554 6420 14560
rect 5816 14476 5868 14482
rect 5816 14418 5868 14424
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 5828 13802 5856 14418
rect 5816 13796 5868 13802
rect 5816 13738 5868 13744
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5356 13456 5408 13462
rect 5356 13398 5408 13404
rect 5368 12714 5396 13398
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 5356 12708 5408 12714
rect 5356 12650 5408 12656
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 5644 11778 5672 12242
rect 5644 11750 5764 11778
rect 5632 11620 5684 11626
rect 5632 11562 5684 11568
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5264 11076 5316 11082
rect 5264 11018 5316 11024
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 5448 10532 5500 10538
rect 5448 10474 5500 10480
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4724 8566 4752 8910
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4436 8560 4488 8566
rect 4436 8502 4488 8508
rect 4712 8560 4764 8566
rect 4712 8502 4764 8508
rect 4448 8265 4476 8502
rect 4434 8256 4490 8265
rect 4724 8242 4752 8502
rect 4816 8430 4844 8774
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4804 8424 4856 8430
rect 4908 8401 4936 8434
rect 4804 8366 4856 8372
rect 4894 8392 4950 8401
rect 4894 8327 4950 8336
rect 4804 8288 4856 8294
rect 4724 8236 4804 8242
rect 4724 8230 4856 8236
rect 4724 8214 4844 8230
rect 4434 8191 4490 8200
rect 4816 7886 4844 8214
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4724 6798 4752 7142
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4724 6254 4752 6734
rect 4816 6730 4844 7822
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4908 6610 4936 7890
rect 5000 7750 5028 9318
rect 5092 9178 5120 10474
rect 5460 10266 5488 10474
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5460 9586 5488 10202
rect 5552 10198 5580 11494
rect 5644 11150 5672 11562
rect 5736 11558 5764 11750
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 6196 11354 6224 13262
rect 6380 12782 6408 13262
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6380 12442 6408 12718
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6380 11898 6408 12242
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 6092 11280 6144 11286
rect 6092 11222 6144 11228
rect 5632 11144 5684 11150
rect 5632 11086 5684 11092
rect 5644 10810 5672 11086
rect 5908 11076 5960 11082
rect 5908 11018 5960 11024
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5724 10532 5776 10538
rect 5724 10474 5776 10480
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 5184 8090 5212 8298
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 4988 7744 5040 7750
rect 4988 7686 5040 7692
rect 4816 6582 4936 6610
rect 4712 6248 4764 6254
rect 4712 6190 4764 6196
rect 4724 5710 4752 6190
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4620 4208 4672 4214
rect 4620 4150 4672 4156
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4540 3602 4568 4014
rect 4632 3754 4660 4150
rect 4724 3942 4752 5170
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4632 3726 4752 3754
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4264 1958 4568 1986
rect 4540 480 4568 1958
rect 4724 1902 4752 3726
rect 4816 3108 4844 6582
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 4908 5778 4936 6258
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4908 3738 4936 4626
rect 5000 4282 5028 7686
rect 5184 6866 5212 8026
rect 5276 8022 5304 8910
rect 5264 8016 5316 8022
rect 5264 7958 5316 7964
rect 5276 7562 5304 7958
rect 5276 7534 5488 7562
rect 5460 7478 5488 7534
rect 5448 7472 5500 7478
rect 5448 7414 5500 7420
rect 5354 7168 5410 7177
rect 5354 7103 5410 7112
rect 5368 6934 5396 7103
rect 5356 6928 5408 6934
rect 5356 6870 5408 6876
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 5092 6254 5120 6598
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 5092 5778 5120 6190
rect 5080 5772 5132 5778
rect 5080 5714 5132 5720
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5184 4486 5212 4966
rect 5552 4706 5580 9454
rect 5736 9382 5764 10474
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5736 7698 5764 9318
rect 5816 9104 5868 9110
rect 5814 9072 5816 9081
rect 5868 9072 5870 9081
rect 5814 9007 5870 9016
rect 5736 7670 5856 7698
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5644 6390 5672 6802
rect 5632 6384 5684 6390
rect 5632 6326 5684 6332
rect 5736 6254 5764 7482
rect 5828 6322 5856 7670
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 5724 6112 5776 6118
rect 5644 6060 5724 6066
rect 5644 6054 5776 6060
rect 5644 6038 5764 6054
rect 5644 5846 5672 6038
rect 5632 5840 5684 5846
rect 5632 5782 5684 5788
rect 5644 5522 5672 5782
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5644 5494 5764 5522
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5644 5273 5672 5306
rect 5630 5264 5686 5273
rect 5630 5199 5686 5208
rect 5632 5160 5684 5166
rect 5632 5102 5684 5108
rect 5644 4826 5672 5102
rect 5736 4826 5764 5494
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5460 4678 5580 4706
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 4988 4276 5040 4282
rect 4988 4218 5040 4224
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 4896 3120 4948 3126
rect 4816 3080 4896 3108
rect 4896 3062 4948 3068
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 4894 2952 4950 2961
rect 4894 2887 4950 2896
rect 4908 2650 4936 2887
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 4712 1896 4764 1902
rect 4712 1838 4764 1844
rect 5000 480 5028 2994
rect 5092 2650 5120 4422
rect 5184 3398 5212 4422
rect 5264 4004 5316 4010
rect 5264 3946 5316 3952
rect 5276 3398 5304 3946
rect 5368 3602 5396 4558
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5172 3120 5224 3126
rect 5172 3062 5224 3068
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 5184 2514 5212 3062
rect 5172 2508 5224 2514
rect 5172 2450 5224 2456
rect 5276 2446 5304 3334
rect 5368 3126 5396 3538
rect 5356 3120 5408 3126
rect 5356 3062 5408 3068
rect 5368 2514 5396 3062
rect 5356 2508 5408 2514
rect 5356 2450 5408 2456
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 5460 480 5488 4678
rect 5828 4554 5856 5714
rect 5816 4548 5868 4554
rect 5816 4490 5868 4496
rect 5828 4282 5856 4490
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5644 2854 5672 3946
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5920 480 5948 11018
rect 6104 9024 6132 11222
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6196 9178 6224 9318
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 6184 9036 6236 9042
rect 6104 8996 6184 9024
rect 6184 8978 6236 8984
rect 6092 8356 6144 8362
rect 6092 8298 6144 8304
rect 6104 5114 6132 8298
rect 6196 7002 6224 8978
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 6012 5086 6132 5114
rect 6012 4010 6040 5086
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6000 4004 6052 4010
rect 6000 3946 6052 3952
rect 6104 3738 6132 4966
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 6012 3126 6040 3334
rect 6000 3120 6052 3126
rect 6000 3062 6052 3068
rect 6090 3088 6146 3097
rect 6090 3023 6146 3032
rect 6104 2854 6132 3023
rect 6092 2848 6144 2854
rect 6092 2790 6144 2796
rect 6196 950 6224 6938
rect 6288 5658 6316 11494
rect 6380 11150 6408 11834
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6564 10282 6592 15642
rect 6840 12306 6868 15914
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 6932 13870 6960 14418
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6932 13530 6960 13806
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 6932 12238 6960 13466
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6642 11384 6698 11393
rect 6642 11319 6698 11328
rect 6380 10254 6592 10282
rect 6380 7954 6408 10254
rect 6656 10198 6684 11319
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6644 10192 6696 10198
rect 6644 10134 6696 10140
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6472 7546 6500 10066
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6564 9058 6592 9998
rect 6840 9654 6868 10406
rect 6932 10130 6960 12174
rect 7024 11354 7052 17682
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7116 13870 7144 14554
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 7208 13530 7236 18634
rect 7288 16652 7340 16658
rect 7288 16594 7340 16600
rect 7300 16250 7328 16594
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7576 15026 7604 15302
rect 7564 15020 7616 15026
rect 7564 14962 7616 14968
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7392 14482 7420 14758
rect 7380 14476 7432 14482
rect 7380 14418 7432 14424
rect 7196 13524 7248 13530
rect 7196 13466 7248 13472
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7116 12102 7144 13330
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 7208 12850 7236 13262
rect 7392 13190 7420 14418
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7116 11898 7144 12038
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 7116 10470 7144 11630
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6564 9030 6684 9058
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6564 8022 6592 8910
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6564 7342 6592 7686
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6288 5630 6408 5658
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6288 4622 6316 5510
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6380 4468 6408 5630
rect 6564 5302 6592 5714
rect 6552 5296 6604 5302
rect 6552 5238 6604 5244
rect 6564 4690 6592 5238
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6288 4440 6408 4468
rect 6184 944 6236 950
rect 6184 886 6236 892
rect 6288 480 6316 4440
rect 6460 4276 6512 4282
rect 6460 4218 6512 4224
rect 6472 3534 6500 4218
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 6656 3482 6684 9030
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6748 8498 6776 8978
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6840 8362 6868 9318
rect 6828 8356 6880 8362
rect 6828 8298 6880 8304
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6840 5642 6868 6054
rect 6828 5636 6880 5642
rect 6828 5578 6880 5584
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6748 3641 6776 4966
rect 6932 4842 6960 9386
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 7024 8090 7052 8978
rect 7116 8430 7144 10406
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6840 4814 6960 4842
rect 6840 4026 6868 4814
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6932 4146 6960 4626
rect 7024 4468 7052 7686
rect 7116 7478 7144 7822
rect 7104 7472 7156 7478
rect 7104 7414 7156 7420
rect 7208 7274 7236 8774
rect 7300 7410 7328 8774
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 7196 7268 7248 7274
rect 7196 7210 7248 7216
rect 7116 6254 7144 7210
rect 7288 6860 7340 6866
rect 7288 6802 7340 6808
rect 7300 6322 7328 6802
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7288 5840 7340 5846
rect 7288 5782 7340 5788
rect 7104 5568 7156 5574
rect 7156 5528 7236 5556
rect 7104 5510 7156 5516
rect 7208 5098 7236 5528
rect 7300 5098 7328 5782
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 7288 5092 7340 5098
rect 7288 5034 7340 5040
rect 7208 4622 7236 5034
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 7024 4440 7236 4468
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6840 3998 6960 4026
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6840 3738 6868 3878
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6734 3632 6790 3641
rect 6734 3567 6736 3576
rect 6788 3567 6790 3576
rect 6736 3538 6788 3544
rect 6656 3454 6776 3482
rect 6748 480 6776 3454
rect 6932 3398 6960 3998
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 7024 2310 7052 2790
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 7208 480 7236 4440
rect 7300 3534 7328 5034
rect 7392 4468 7420 12242
rect 7484 7562 7512 14758
rect 7576 14550 7604 14962
rect 7564 14544 7616 14550
rect 7564 14486 7616 14492
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7576 12850 7604 13806
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7668 11898 7696 18770
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 8220 17814 8248 18770
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8208 17808 8260 17814
rect 8208 17750 8260 17756
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 8128 16046 8156 16526
rect 8116 16040 8168 16046
rect 8116 15982 8168 15988
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 7760 15162 7788 15846
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 8220 15638 8248 15982
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 8220 15026 8248 15574
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 7748 14884 7800 14890
rect 7748 14826 7800 14832
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7760 11234 7788 14826
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 8588 14618 8616 18702
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 8668 18216 8720 18222
rect 8668 18158 8720 18164
rect 8680 17202 8708 18158
rect 10416 18148 10468 18154
rect 10416 18090 10468 18096
rect 10428 17814 10456 18090
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 10416 17808 10468 17814
rect 10416 17750 10468 17756
rect 10784 17740 10836 17746
rect 10784 17682 10836 17688
rect 10416 17672 10468 17678
rect 10416 17614 10468 17620
rect 8668 17196 8720 17202
rect 8668 17138 8720 17144
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9600 16794 9628 16934
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9128 15972 9180 15978
rect 9128 15914 9180 15920
rect 9140 15706 9168 15914
rect 9692 15706 9720 16934
rect 9876 16794 9904 17138
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 10232 16652 10284 16658
rect 10232 16594 10284 16600
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 10244 15910 10272 16594
rect 10336 16046 10364 16594
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 10232 15904 10284 15910
rect 10232 15846 10284 15852
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 8852 15564 8904 15570
rect 8852 15506 8904 15512
rect 8864 15162 8892 15506
rect 10244 15502 10272 15846
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 8852 15156 8904 15162
rect 8852 15098 8904 15104
rect 9404 14884 9456 14890
rect 9404 14826 9456 14832
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 9416 14414 9444 14826
rect 10336 14550 10364 15982
rect 10428 15042 10456 17614
rect 10796 17338 10824 17682
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 17958 17232 18014 17241
rect 11428 17196 11480 17202
rect 17958 17167 18014 17176
rect 11428 17138 11480 17144
rect 11060 16992 11112 16998
rect 11060 16934 11112 16940
rect 10508 16788 10560 16794
rect 10508 16730 10560 16736
rect 10520 16046 10548 16730
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 11072 15706 11100 16934
rect 11440 16794 11468 17138
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 17972 16794 18000 17167
rect 11428 16788 11480 16794
rect 11428 16730 11480 16736
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11624 16250 11652 16594
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 10428 15014 10548 15042
rect 9680 14544 9732 14550
rect 9680 14486 9732 14492
rect 10324 14544 10376 14550
rect 10324 14486 10376 14492
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9404 14408 9456 14414
rect 9404 14350 9456 14356
rect 9600 13938 9628 14418
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9036 13796 9088 13802
rect 9036 13738 9088 13744
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 7576 11206 7788 11234
rect 7576 7750 7604 11206
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 7760 10606 7788 11086
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7668 9518 7696 10542
rect 7760 10266 7788 10542
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 8220 10130 8248 13670
rect 9048 13326 9076 13738
rect 9692 13530 9720 14486
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9968 14074 9996 14418
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9968 13462 9996 14010
rect 9956 13456 10008 13462
rect 9956 13398 10008 13404
rect 9220 13388 9272 13394
rect 9220 13330 9272 13336
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 9048 12986 9076 13262
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 8668 12708 8720 12714
rect 8668 12650 8720 12656
rect 8482 12336 8538 12345
rect 8392 12300 8444 12306
rect 8482 12271 8484 12280
rect 8392 12242 8444 12248
rect 8536 12271 8538 12280
rect 8484 12242 8536 12248
rect 8404 11762 8432 12242
rect 8680 12170 8708 12650
rect 9232 12442 9260 13330
rect 10048 13252 10100 13258
rect 10048 13194 10100 13200
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 8668 12164 8720 12170
rect 8668 12106 8720 12112
rect 8666 11792 8722 11801
rect 8392 11756 8444 11762
rect 8666 11727 8722 11736
rect 8392 11698 8444 11704
rect 8576 11552 8628 11558
rect 8576 11494 8628 11500
rect 8588 11354 8616 11494
rect 8680 11354 8708 11727
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 9600 11286 9628 11562
rect 9588 11280 9640 11286
rect 9588 11222 9640 11228
rect 9692 11218 9720 11562
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 8496 10266 8524 11154
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8220 9994 8248 10066
rect 8208 9988 8260 9994
rect 8208 9930 8260 9936
rect 8312 9586 8340 10066
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7668 8634 7696 9454
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 8588 9178 8616 11018
rect 9036 10736 9088 10742
rect 9036 10678 9088 10684
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 7656 8356 7708 8362
rect 7656 8298 7708 8304
rect 7668 7886 7696 8298
rect 7760 8090 7788 8978
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 8128 8634 8156 8910
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7484 7534 7788 7562
rect 8220 7546 8248 8978
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7576 4826 7604 5714
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 7668 5370 7696 5646
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7656 4684 7708 4690
rect 7656 4626 7708 4632
rect 7392 4440 7604 4468
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7576 3482 7604 4440
rect 7668 3602 7696 4626
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7300 2990 7328 3470
rect 7576 3454 7696 3482
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 7380 2916 7432 2922
rect 7380 2858 7432 2864
rect 7288 2848 7340 2854
rect 7286 2816 7288 2825
rect 7340 2816 7342 2825
rect 7286 2751 7342 2760
rect 7392 2650 7420 2858
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7668 480 7696 3454
rect 7760 2530 7788 7534
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 8496 7002 8524 7822
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8312 6254 8340 6598
rect 8496 6254 8524 6598
rect 8300 6248 8352 6254
rect 8300 6190 8352 6196
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 8312 5846 8340 6190
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8300 5840 8352 5846
rect 8300 5782 8352 5788
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8312 5370 8340 5646
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8404 5098 8432 5850
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8392 5092 8444 5098
rect 8392 5034 8444 5040
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 8496 4826 8524 5510
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7852 4146 7880 4422
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 8116 3392 8168 3398
rect 8220 3380 8248 4218
rect 8404 4146 8432 4558
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8392 4004 8444 4010
rect 8392 3946 8444 3952
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8168 3352 8248 3380
rect 8116 3334 8168 3340
rect 8128 2990 8156 3334
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 8312 2582 8340 3878
rect 8404 2650 8432 3946
rect 8588 2666 8616 8910
rect 8680 7478 8708 9998
rect 9048 9518 9076 10678
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 8956 9178 8984 9318
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8864 7886 8892 8774
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 8864 7410 8892 7822
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 8956 7342 8984 9114
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8760 5840 8812 5846
rect 8760 5782 8812 5788
rect 8850 5808 8906 5817
rect 8666 5672 8722 5681
rect 8666 5607 8722 5616
rect 8680 5370 8708 5607
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8772 5166 8800 5782
rect 8850 5743 8852 5752
rect 8904 5743 8906 5752
rect 8852 5714 8904 5720
rect 8760 5160 8812 5166
rect 8760 5102 8812 5108
rect 8772 4622 8800 5102
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8680 3738 8708 4014
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8772 3738 8800 3878
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 8668 2848 8720 2854
rect 8668 2790 8720 2796
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8496 2638 8616 2666
rect 8300 2576 8352 2582
rect 7760 2502 8064 2530
rect 8300 2518 8352 2524
rect 8036 480 8064 2502
rect 8496 480 8524 2638
rect 8680 2446 8708 2790
rect 8668 2440 8720 2446
rect 8772 2417 8800 2926
rect 8944 2848 8996 2854
rect 8944 2790 8996 2796
rect 8956 2650 8984 2790
rect 8944 2644 8996 2650
rect 8944 2586 8996 2592
rect 9140 2530 9168 10542
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 9232 8974 9260 9930
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9312 8900 9364 8906
rect 9312 8842 9364 8848
rect 9220 7268 9272 7274
rect 9220 7210 9272 7216
rect 9232 6322 9260 7210
rect 9220 6316 9272 6322
rect 9220 6258 9272 6264
rect 9324 3942 9352 8842
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 8956 2502 9168 2530
rect 8668 2382 8720 2388
rect 8758 2408 8814 2417
rect 8758 2343 8814 2352
rect 8956 480 8984 2502
rect 9416 480 9444 11018
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 9508 10248 9536 10746
rect 9588 10260 9640 10266
rect 9508 10220 9588 10248
rect 9588 10202 9640 10208
rect 9692 9450 9720 10950
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9692 8498 9720 8910
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9692 7410 9720 8434
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9692 6202 9720 6938
rect 9770 6488 9826 6497
rect 9770 6423 9772 6432
rect 9824 6423 9826 6432
rect 9772 6394 9824 6400
rect 9864 6384 9916 6390
rect 9770 6352 9826 6361
rect 9864 6326 9916 6332
rect 9770 6287 9772 6296
rect 9824 6287 9826 6296
rect 9772 6258 9824 6264
rect 9600 6174 9720 6202
rect 9600 5930 9628 6174
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9600 5902 9720 5930
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9600 4078 9628 4558
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9600 3942 9628 4014
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9496 3392 9548 3398
rect 9496 3334 9548 3340
rect 9508 3058 9536 3334
rect 9692 3176 9720 5902
rect 9784 5710 9812 6054
rect 9876 5914 9904 6326
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9784 4758 9812 5646
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9600 3148 9720 3176
rect 9600 3097 9628 3148
rect 9772 3120 9824 3126
rect 9586 3088 9642 3097
rect 9496 3052 9548 3058
rect 9772 3062 9824 3068
rect 9586 3023 9642 3032
rect 9680 3052 9732 3058
rect 9496 2994 9548 3000
rect 9600 2802 9628 3023
rect 9680 2994 9732 3000
rect 9692 2961 9720 2994
rect 9678 2952 9734 2961
rect 9678 2887 9734 2896
rect 9600 2774 9720 2802
rect 9692 2514 9720 2774
rect 9784 2650 9812 3062
rect 9772 2644 9824 2650
rect 9772 2586 9824 2592
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 9968 2122 9996 12174
rect 10060 9704 10088 13194
rect 10336 12986 10364 14486
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10336 11694 10364 12922
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10060 9676 10272 9704
rect 10244 7274 10272 9676
rect 10048 7268 10100 7274
rect 10048 7210 10100 7216
rect 10232 7268 10284 7274
rect 10232 7210 10284 7216
rect 10060 6474 10088 7210
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 10051 6446 10088 6474
rect 10051 6338 10079 6446
rect 10138 6352 10194 6361
rect 10051 6310 10088 6338
rect 10060 5148 10088 6310
rect 10138 6287 10194 6296
rect 10152 6254 10180 6287
rect 10140 6248 10192 6254
rect 10140 6190 10192 6196
rect 10244 6118 10272 6802
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10244 5166 10272 5510
rect 10051 5120 10088 5148
rect 10232 5160 10284 5166
rect 10051 5080 10079 5120
rect 10232 5102 10284 5108
rect 10051 5052 10088 5080
rect 10060 4842 10088 5052
rect 10060 4814 10272 4842
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 10060 4078 10088 4422
rect 10048 4072 10100 4078
rect 10048 4014 10100 4020
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 10152 2310 10180 2586
rect 10140 2304 10192 2310
rect 10140 2246 10192 2252
rect 9784 2094 9996 2122
rect 9784 480 9812 2094
rect 10244 480 10272 4814
rect 10336 3126 10364 10066
rect 10428 9654 10456 12718
rect 10520 10810 10548 15014
rect 10692 14816 10744 14822
rect 10692 14758 10744 14764
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10416 9648 10468 9654
rect 10416 9590 10468 9596
rect 10428 8362 10456 9590
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10416 6112 10468 6118
rect 10416 6054 10468 6060
rect 10324 3120 10376 3126
rect 10324 3062 10376 3068
rect 10428 3058 10456 6054
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10520 2922 10548 7142
rect 10612 6866 10640 7210
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 10600 5024 10652 5030
rect 10600 4966 10652 4972
rect 10612 4758 10640 4966
rect 10600 4752 10652 4758
rect 10600 4694 10652 4700
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10612 3534 10640 3878
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10508 2916 10560 2922
rect 10508 2858 10560 2864
rect 10612 2446 10640 2994
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10704 480 10732 14758
rect 11072 14618 11100 15506
rect 11624 15502 11652 16186
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 11704 15632 11756 15638
rect 11704 15574 11756 15580
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11716 15314 11744 15574
rect 12072 15564 12124 15570
rect 12072 15506 12124 15512
rect 11624 15286 11744 15314
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11164 11354 11192 11494
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 10784 11212 10836 11218
rect 10784 11154 10836 11160
rect 10796 10606 10824 11154
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10796 9722 10824 10542
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10888 9722 10916 9862
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 11152 9444 11204 9450
rect 11152 9386 11204 9392
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10888 8634 10916 8978
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10888 7886 10916 8570
rect 11164 7954 11192 9386
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11348 8022 11376 8230
rect 11336 8016 11388 8022
rect 11336 7958 11388 7964
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10980 7426 11008 7822
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 10888 7398 11008 7426
rect 10888 7002 10916 7398
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 10980 6798 11008 7278
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 10796 5234 10824 5714
rect 11164 5681 11192 6054
rect 11150 5672 11206 5681
rect 11150 5607 11206 5616
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 10888 4729 10916 4966
rect 10874 4720 10930 4729
rect 10796 4678 10874 4706
rect 10796 2650 10824 4678
rect 10874 4655 10930 4664
rect 10876 4548 10928 4554
rect 10876 4490 10928 4496
rect 10888 3058 10916 4490
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11164 3670 11192 3878
rect 11256 3738 11284 3878
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11152 3664 11204 3670
rect 11152 3606 11204 3612
rect 11624 3380 11652 15286
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11796 9512 11848 9518
rect 11796 9454 11848 9460
rect 11808 8634 11836 9454
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11808 8514 11836 8570
rect 11808 8486 11928 8514
rect 11704 8424 11756 8430
rect 11704 8366 11756 8372
rect 11716 8022 11744 8366
rect 11704 8016 11756 8022
rect 11704 7958 11756 7964
rect 11900 7342 11928 8486
rect 11992 8430 12020 10202
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11716 6934 11744 7142
rect 11704 6928 11756 6934
rect 11704 6870 11756 6876
rect 11716 6322 11744 6870
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11808 6118 11836 6598
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11900 5846 11928 7142
rect 11888 5840 11940 5846
rect 11888 5782 11940 5788
rect 12084 5522 12112 15506
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 19076 11354 19104 11630
rect 19892 11552 19944 11558
rect 19892 11494 19944 11500
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 19432 11076 19484 11082
rect 19432 11018 19484 11024
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 18236 10600 18288 10606
rect 18236 10542 18288 10548
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 18248 9994 18276 10542
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18236 9988 18288 9994
rect 18236 9930 18288 9936
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 12256 9104 12308 9110
rect 12256 9046 12308 9052
rect 12164 5908 12216 5914
rect 12164 5850 12216 5856
rect 12176 5817 12204 5850
rect 12162 5808 12218 5817
rect 12162 5743 12218 5752
rect 11808 5494 12112 5522
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11716 4690 11744 4966
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11808 4434 11836 5494
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11900 5273 11928 5306
rect 11886 5264 11942 5273
rect 11886 5199 11942 5208
rect 11888 5092 11940 5098
rect 11888 5034 11940 5040
rect 11164 3352 11652 3380
rect 11716 4406 11836 4434
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 11164 480 11192 3352
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11716 3210 11744 4406
rect 11796 4276 11848 4282
rect 11796 4218 11848 4224
rect 11808 3534 11836 4218
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11624 3182 11744 3210
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11624 480 11652 3182
rect 11900 3097 11928 5034
rect 11980 3664 12032 3670
rect 11980 3606 12032 3612
rect 11886 3088 11942 3097
rect 11992 3058 12020 3606
rect 12072 3596 12124 3602
rect 12072 3538 12124 3544
rect 11886 3023 11942 3032
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 11980 2916 12032 2922
rect 11980 2858 12032 2864
rect 11992 480 12020 2858
rect 12084 2650 12112 3538
rect 12268 2854 12296 9046
rect 14096 7268 14148 7274
rect 14096 7210 14148 7216
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12348 6248 12400 6254
rect 12452 6202 12480 7142
rect 12716 6928 12768 6934
rect 12716 6870 12768 6876
rect 12400 6196 12480 6202
rect 12348 6190 12480 6196
rect 12360 6174 12480 6190
rect 12624 6180 12676 6186
rect 12728 6168 12756 6870
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 13924 6458 13952 6802
rect 13912 6452 13964 6458
rect 13912 6394 13964 6400
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13556 6186 13584 6258
rect 12676 6140 12756 6168
rect 12624 6122 12676 6128
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12348 4072 12400 4078
rect 12348 4014 12400 4020
rect 12360 3534 12388 4014
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12544 3126 12572 4558
rect 12728 4078 12756 6140
rect 13544 6180 13596 6186
rect 13544 6122 13596 6128
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 13004 5234 13032 5714
rect 13556 5574 13584 6122
rect 13924 5710 13952 6394
rect 14108 6186 14136 7210
rect 14384 7206 14412 9658
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 15752 8016 15804 8022
rect 15752 7958 15804 7964
rect 15016 7880 15068 7886
rect 15016 7822 15068 7828
rect 14648 7812 14700 7818
rect 14648 7754 14700 7760
rect 14660 7342 14688 7754
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14096 6180 14148 6186
rect 14096 6122 14148 6128
rect 14108 5914 14136 6122
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 14200 5846 14228 7142
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 15028 6798 15056 7822
rect 15660 7472 15712 7478
rect 15660 7414 15712 7420
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15212 6866 15240 7346
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 15016 6792 15068 6798
rect 15016 6734 15068 6740
rect 14554 6352 14610 6361
rect 14554 6287 14610 6296
rect 14568 6254 14596 6287
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14292 5914 14320 6054
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 14188 5840 14240 5846
rect 14188 5782 14240 5788
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 14370 5672 14426 5681
rect 14370 5607 14426 5616
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 13832 5166 13860 5510
rect 14384 5166 14412 5607
rect 15028 5574 15056 6734
rect 15580 6254 15608 7142
rect 15672 6254 15700 7414
rect 15764 6610 15792 7958
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 17776 7268 17828 7274
rect 17776 7210 17828 7216
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 15936 6656 15988 6662
rect 15764 6604 15936 6610
rect 15764 6598 15988 6604
rect 15764 6582 15976 6598
rect 15764 6322 15792 6582
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15660 6248 15712 6254
rect 15660 6190 15712 6196
rect 15936 6248 15988 6254
rect 15936 6190 15988 6196
rect 15948 5710 15976 6190
rect 16040 6118 16068 6802
rect 16960 6458 16988 6802
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 17408 6180 17460 6186
rect 17408 6122 17460 6128
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 17420 5914 17448 6122
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 16488 5840 16540 5846
rect 16488 5782 16540 5788
rect 15476 5704 15528 5710
rect 15476 5646 15528 5652
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 15016 5568 15068 5574
rect 15016 5510 15068 5516
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 13268 5092 13320 5098
rect 13268 5034 13320 5040
rect 13912 5092 13964 5098
rect 13912 5034 13964 5040
rect 14556 5092 14608 5098
rect 14556 5034 14608 5040
rect 12808 5024 12860 5030
rect 12808 4966 12860 4972
rect 12820 4146 12848 4966
rect 13280 4826 13308 5034
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 13280 4078 13308 4218
rect 12716 4072 12768 4078
rect 12716 4014 12768 4020
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 12624 4004 12676 4010
rect 12624 3946 12676 3952
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12256 2848 12308 2854
rect 12256 2790 12308 2796
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 12452 2582 12480 2926
rect 12440 2576 12492 2582
rect 12440 2518 12492 2524
rect 12636 2514 12664 3946
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13464 3194 13492 3470
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13648 3058 13676 3334
rect 13636 3052 13688 3058
rect 13636 2994 13688 3000
rect 13740 2990 13768 4558
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13832 3738 13860 3946
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 13360 2848 13412 2854
rect 13360 2790 13412 2796
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 12452 480 12480 2246
rect 12912 480 12940 2246
rect 13372 480 13400 2790
rect 13740 480 13768 2790
rect 13924 2514 13952 5034
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 14384 4282 14412 4558
rect 14464 4480 14516 4486
rect 14464 4422 14516 4428
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 14292 3602 14320 3878
rect 14476 3738 14504 4422
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 13912 2508 13964 2514
rect 13912 2450 13964 2456
rect 14200 480 14228 2790
rect 14476 2650 14504 3538
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 14568 2514 14596 5034
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 15028 4622 15056 5510
rect 14648 4616 14700 4622
rect 14648 4558 14700 4564
rect 15016 4616 15068 4622
rect 15016 4558 15068 4564
rect 14660 4146 14688 4558
rect 14740 4276 14792 4282
rect 14740 4218 14792 4224
rect 14648 4140 14700 4146
rect 14648 4082 14700 4088
rect 14752 4060 14780 4218
rect 15016 4072 15068 4078
rect 14752 4032 15016 4060
rect 15016 4014 15068 4020
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 15488 2514 15516 5646
rect 16500 5234 16528 5782
rect 17420 5234 17448 5850
rect 17696 5778 17724 6734
rect 17684 5772 17736 5778
rect 17684 5714 17736 5720
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 16132 4282 16160 4626
rect 16500 4486 16528 5170
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 16592 4690 16620 4966
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 16488 4480 16540 4486
rect 16488 4422 16540 4428
rect 16120 4276 16172 4282
rect 16120 4218 16172 4224
rect 16132 3670 16160 4218
rect 16500 4214 16528 4422
rect 16776 4282 16804 4966
rect 17038 4720 17094 4729
rect 17038 4655 17094 4664
rect 16764 4276 16816 4282
rect 16764 4218 16816 4224
rect 16488 4208 16540 4214
rect 16488 4150 16540 4156
rect 16212 4004 16264 4010
rect 16212 3946 16264 3952
rect 16224 3670 16252 3946
rect 17052 3942 17080 4655
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 16212 3664 16264 3670
rect 16212 3606 16264 3612
rect 17236 3602 17264 4558
rect 17788 3602 17816 7210
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 18602 5808 18658 5817
rect 18602 5743 18658 5752
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 15752 3596 15804 3602
rect 15752 3538 15804 3544
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 15660 3392 15712 3398
rect 15660 3334 15712 3340
rect 15672 2990 15700 3334
rect 15764 3194 15792 3538
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 15752 3188 15804 3194
rect 15752 3130 15804 3136
rect 15936 3120 15988 3126
rect 15936 3062 15988 3068
rect 16394 3088 16450 3097
rect 15660 2984 15712 2990
rect 15660 2926 15712 2932
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 14648 2304 14700 2310
rect 14648 2246 14700 2252
rect 15108 2304 15160 2310
rect 15108 2246 15160 2252
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 14660 480 14688 2246
rect 15120 480 15148 2246
rect 15488 480 15516 2246
rect 15948 480 15976 3062
rect 16394 3023 16450 3032
rect 16408 2990 16436 3023
rect 16396 2984 16448 2990
rect 16396 2926 16448 2932
rect 16028 2848 16080 2854
rect 16028 2790 16080 2796
rect 16040 2514 16068 2790
rect 16684 2514 16712 3470
rect 17684 3392 17736 3398
rect 17684 3334 17736 3340
rect 16856 2848 16908 2854
rect 16856 2790 16908 2796
rect 16028 2508 16080 2514
rect 16028 2450 16080 2456
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 16396 2304 16448 2310
rect 16396 2246 16448 2252
rect 16408 480 16436 2246
rect 16868 480 16896 2790
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 17328 480 17356 2246
rect 17696 480 17724 3334
rect 17972 1986 18000 5510
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 18616 4758 18644 5743
rect 18604 4752 18656 4758
rect 18604 4694 18656 4700
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 17972 1958 18184 1986
rect 18156 480 18184 1958
rect 18616 480 18644 3334
rect 18708 626 18736 10406
rect 18708 598 19104 626
rect 19076 480 19104 598
rect 19444 480 19472 11018
rect 19904 480 19932 11494
rect 20364 480 20392 12038
rect 21180 3936 21232 3942
rect 21180 3878 21232 3884
rect 20812 3392 20864 3398
rect 20812 3334 20864 3340
rect 20824 480 20852 3334
rect 21192 480 21220 3878
rect 21640 2984 21692 2990
rect 21640 2926 21692 2932
rect 21652 480 21680 2926
rect 22560 2916 22612 2922
rect 22560 2858 22612 2864
rect 22100 2848 22152 2854
rect 22100 2790 22152 2796
rect 22112 480 22140 2790
rect 22572 480 22600 2858
rect 3974 232 4030 241
rect 3974 167 4030 176
rect 4066 0 4122 480
rect 4526 0 4582 480
rect 4986 0 5042 480
rect 5446 0 5502 480
rect 5906 0 5962 480
rect 6274 0 6330 480
rect 6734 0 6790 480
rect 7194 0 7250 480
rect 7654 0 7710 480
rect 8022 0 8078 480
rect 8482 0 8538 480
rect 8942 0 8998 480
rect 9402 0 9458 480
rect 9770 0 9826 480
rect 10230 0 10286 480
rect 10690 0 10746 480
rect 11150 0 11206 480
rect 11610 0 11666 480
rect 11978 0 12034 480
rect 12438 0 12494 480
rect 12898 0 12954 480
rect 13358 0 13414 480
rect 13726 0 13782 480
rect 14186 0 14242 480
rect 14646 0 14702 480
rect 15106 0 15162 480
rect 15474 0 15530 480
rect 15934 0 15990 480
rect 16394 0 16450 480
rect 16854 0 16910 480
rect 17314 0 17370 480
rect 17682 0 17738 480
rect 18142 0 18198 480
rect 18602 0 18658 480
rect 19062 0 19118 480
rect 19430 0 19486 480
rect 19890 0 19946 480
rect 20350 0 20406 480
rect 20810 0 20866 480
rect 21178 0 21234 480
rect 21638 0 21694 480
rect 22098 0 22154 480
rect 22558 0 22614 480
<< via2 >>
rect 3974 22480 4030 22536
rect 3054 22072 3110 22128
rect 2870 21120 2926 21176
rect 2778 20576 2834 20632
rect 1950 20168 2006 20224
rect 1858 18264 1914 18320
rect 1950 17856 2006 17912
rect 1766 16940 1768 16960
rect 1768 16940 1820 16960
rect 1820 16940 1822 16960
rect 1766 16904 1822 16940
rect 2778 18808 2834 18864
rect 3606 21528 3662 21584
rect 3698 19760 3754 19816
rect 3790 17332 3846 17368
rect 3790 17312 3792 17332
rect 3792 17312 3844 17332
rect 3844 17312 3846 17332
rect 1674 15544 1730 15600
rect 1766 15000 1822 15056
rect 1674 14592 1730 14648
rect 1582 14048 1638 14104
rect 3330 16516 3386 16552
rect 3330 16496 3332 16516
rect 3332 16496 3384 16516
rect 3384 16496 3386 16516
rect 2962 15952 3018 16008
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 4066 19216 4122 19272
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 3238 13232 3294 13288
rect 2870 9968 2926 10024
rect 2226 8236 2228 8256
rect 2228 8236 2280 8256
rect 2280 8236 2282 8256
rect 2226 8200 2282 8236
rect 2226 4800 2282 4856
rect 1674 2896 1730 2952
rect 1306 1944 1362 2000
rect 3606 13640 3662 13696
rect 3422 12688 3478 12744
rect 4066 12280 4122 12336
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4066 10784 4122 10840
rect 4066 10376 4122 10432
rect 3882 9424 3938 9480
rect 2778 3576 2834 3632
rect 2870 1536 2926 1592
rect 3422 5208 3478 5264
rect 3974 8472 4030 8528
rect 4158 8336 4214 8392
rect 3974 8064 4030 8120
rect 4066 7540 4122 7576
rect 4066 7520 4068 7540
rect 4068 7520 4120 7540
rect 4120 7520 4122 7540
rect 4066 6704 4122 6760
rect 3422 2352 3478 2408
rect 3330 992 3386 1048
rect 3330 584 3386 640
rect 3882 5616 3938 5672
rect 4066 6160 4122 6216
rect 4066 5752 4122 5808
rect 4066 4256 4122 4312
rect 3974 3848 4030 3904
rect 4066 3440 4122 3496
rect 3974 3032 4030 3088
rect 3790 2760 3846 2816
rect 3882 2508 3938 2544
rect 3882 2488 3884 2508
rect 3884 2488 3936 2508
rect 3936 2488 3938 2508
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4894 12300 4950 12336
rect 4894 12280 4896 12300
rect 4896 12280 4948 12300
rect 4948 12280 4950 12300
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4434 8200 4490 8256
rect 4894 8336 4950 8392
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 5354 7112 5410 7168
rect 5814 9052 5816 9072
rect 5816 9052 5868 9072
rect 5868 9052 5870 9072
rect 5814 9016 5870 9052
rect 5630 5208 5686 5264
rect 4894 2896 4950 2952
rect 6090 3032 6146 3088
rect 6642 11328 6698 11384
rect 6734 3596 6790 3632
rect 6734 3576 6736 3596
rect 6736 3576 6788 3596
rect 6788 3576 6790 3596
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 17958 17176 18014 17232
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 8482 12300 8538 12336
rect 8482 12280 8484 12300
rect 8484 12280 8536 12300
rect 8536 12280 8538 12300
rect 8666 11736 8722 11792
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7286 2796 7288 2816
rect 7288 2796 7340 2816
rect 7340 2796 7342 2816
rect 7286 2760 7342 2796
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 8666 5616 8722 5672
rect 8850 5772 8906 5808
rect 8850 5752 8852 5772
rect 8852 5752 8904 5772
rect 8904 5752 8906 5772
rect 8758 2352 8814 2408
rect 9770 6452 9826 6488
rect 9770 6432 9772 6452
rect 9772 6432 9824 6452
rect 9824 6432 9826 6452
rect 9770 6316 9826 6352
rect 9770 6296 9772 6316
rect 9772 6296 9824 6316
rect 9824 6296 9826 6316
rect 9586 3032 9642 3088
rect 9678 2896 9734 2952
rect 10138 6296 10194 6352
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 11150 5616 11206 5672
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 10874 4664 10930 4720
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 12162 5752 12218 5808
rect 11886 5208 11942 5264
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 11886 3032 11942 3088
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14554 6296 14610 6352
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 14370 5616 14426 5672
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 17038 4664 17094 4720
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 18602 5752 18658 5808
rect 16394 3032 16450 3088
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 3974 176 4030 232
<< metal3 >>
rect 0 22538 480 22568
rect 3969 22538 4035 22541
rect 0 22536 4035 22538
rect 0 22480 3974 22536
rect 4030 22480 4035 22536
rect 0 22478 4035 22480
rect 0 22448 480 22478
rect 3969 22475 4035 22478
rect 0 22130 480 22160
rect 3049 22130 3115 22133
rect 0 22128 3115 22130
rect 0 22072 3054 22128
rect 3110 22072 3115 22128
rect 0 22070 3115 22072
rect 0 22040 480 22070
rect 3049 22067 3115 22070
rect 0 21586 480 21616
rect 3601 21586 3667 21589
rect 0 21584 3667 21586
rect 0 21528 3606 21584
rect 3662 21528 3667 21584
rect 0 21526 3667 21528
rect 0 21496 480 21526
rect 3601 21523 3667 21526
rect 0 21178 480 21208
rect 2865 21178 2931 21181
rect 0 21176 2931 21178
rect 0 21120 2870 21176
rect 2926 21120 2931 21176
rect 0 21118 2931 21120
rect 0 21088 480 21118
rect 2865 21115 2931 21118
rect 0 20634 480 20664
rect 2773 20634 2839 20637
rect 0 20632 2839 20634
rect 0 20576 2778 20632
rect 2834 20576 2839 20632
rect 0 20574 2839 20576
rect 0 20544 480 20574
rect 2773 20571 2839 20574
rect 0 20226 480 20256
rect 1945 20226 2011 20229
rect 0 20224 2011 20226
rect 0 20168 1950 20224
rect 2006 20168 2011 20224
rect 0 20166 2011 20168
rect 0 20136 480 20166
rect 1945 20163 2011 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 20095 14992 20096
rect 0 19818 480 19848
rect 3693 19818 3759 19821
rect 0 19816 3759 19818
rect 0 19760 3698 19816
rect 3754 19760 3759 19816
rect 0 19758 3759 19760
rect 0 19728 480 19758
rect 3693 19755 3759 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 0 19274 480 19304
rect 4061 19274 4127 19277
rect 0 19272 4127 19274
rect 0 19216 4066 19272
rect 4122 19216 4127 19272
rect 0 19214 4127 19216
rect 0 19184 480 19214
rect 4061 19211 4127 19214
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 0 18866 480 18896
rect 2773 18866 2839 18869
rect 0 18864 2839 18866
rect 0 18808 2778 18864
rect 2834 18808 2839 18864
rect 0 18806 2839 18808
rect 0 18776 480 18806
rect 2773 18803 2839 18806
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 0 18322 480 18352
rect 1853 18322 1919 18325
rect 0 18320 1919 18322
rect 0 18264 1858 18320
rect 1914 18264 1919 18320
rect 0 18262 1919 18264
rect 0 18232 480 18262
rect 1853 18259 1919 18262
rect 7808 17984 8128 17985
rect 0 17914 480 17944
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 1945 17914 2011 17917
rect 0 17912 2011 17914
rect 0 17856 1950 17912
rect 2006 17856 2011 17912
rect 0 17854 2011 17856
rect 0 17824 480 17854
rect 1945 17851 2011 17854
rect 4376 17440 4696 17441
rect 0 17370 480 17400
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 3785 17370 3851 17373
rect 0 17368 3851 17370
rect 0 17312 3790 17368
rect 3846 17312 3851 17368
rect 0 17310 3851 17312
rect 0 17280 480 17310
rect 3785 17307 3851 17310
rect 17953 17234 18019 17237
rect 22320 17234 22800 17264
rect 17953 17232 22800 17234
rect 17953 17176 17958 17232
rect 18014 17176 22800 17232
rect 17953 17174 22800 17176
rect 17953 17171 18019 17174
rect 22320 17144 22800 17174
rect 0 16962 480 16992
rect 1761 16962 1827 16965
rect 0 16960 1827 16962
rect 0 16904 1766 16960
rect 1822 16904 1827 16960
rect 0 16902 1827 16904
rect 0 16872 480 16902
rect 1761 16899 1827 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 16831 14992 16832
rect 0 16554 480 16584
rect 3325 16554 3391 16557
rect 0 16552 3391 16554
rect 0 16496 3330 16552
rect 3386 16496 3391 16552
rect 0 16494 3391 16496
rect 0 16464 480 16494
rect 3325 16491 3391 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 0 16010 480 16040
rect 2957 16010 3023 16013
rect 0 16008 3023 16010
rect 0 15952 2962 16008
rect 3018 15952 3023 16008
rect 0 15950 3023 15952
rect 0 15920 480 15950
rect 2957 15947 3023 15950
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 0 15602 480 15632
rect 1669 15602 1735 15605
rect 0 15600 1735 15602
rect 0 15544 1674 15600
rect 1730 15544 1735 15600
rect 0 15542 1735 15544
rect 0 15512 480 15542
rect 1669 15539 1735 15542
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 0 15058 480 15088
rect 1761 15058 1827 15061
rect 0 15056 1827 15058
rect 0 15000 1766 15056
rect 1822 15000 1827 15056
rect 0 14998 1827 15000
rect 0 14968 480 14998
rect 1761 14995 1827 14998
rect 7808 14720 8128 14721
rect 0 14650 480 14680
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 1669 14650 1735 14653
rect 0 14648 1735 14650
rect 0 14592 1674 14648
rect 1730 14592 1735 14648
rect 0 14590 1735 14592
rect 0 14560 480 14590
rect 1669 14587 1735 14590
rect 4376 14176 4696 14177
rect 0 14106 480 14136
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 1577 14106 1643 14109
rect 0 14104 1643 14106
rect 0 14048 1582 14104
rect 1638 14048 1643 14104
rect 0 14046 1643 14048
rect 0 14016 480 14046
rect 1577 14043 1643 14046
rect 0 13698 480 13728
rect 3601 13698 3667 13701
rect 0 13696 3667 13698
rect 0 13640 3606 13696
rect 3662 13640 3667 13696
rect 0 13638 3667 13640
rect 0 13608 480 13638
rect 3601 13635 3667 13638
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 13567 14992 13568
rect 0 13290 480 13320
rect 3233 13290 3299 13293
rect 0 13288 3299 13290
rect 0 13232 3238 13288
rect 3294 13232 3299 13288
rect 0 13230 3299 13232
rect 0 13200 480 13230
rect 3233 13227 3299 13230
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 0 12746 480 12776
rect 3417 12746 3483 12749
rect 0 12744 3483 12746
rect 0 12688 3422 12744
rect 3478 12688 3483 12744
rect 0 12686 3483 12688
rect 0 12656 480 12686
rect 3417 12683 3483 12686
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 0 12338 480 12368
rect 4061 12338 4127 12341
rect 0 12336 4127 12338
rect 0 12280 4066 12336
rect 4122 12280 4127 12336
rect 0 12278 4127 12280
rect 0 12248 480 12278
rect 4061 12275 4127 12278
rect 4889 12338 4955 12341
rect 8477 12338 8543 12341
rect 4889 12336 8543 12338
rect 4889 12280 4894 12336
rect 4950 12280 8482 12336
rect 8538 12280 8543 12336
rect 4889 12278 8543 12280
rect 4889 12275 4955 12278
rect 8477 12275 8543 12278
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 0 11794 480 11824
rect 8661 11794 8727 11797
rect 0 11792 8727 11794
rect 0 11736 8666 11792
rect 8722 11736 8727 11792
rect 0 11734 8727 11736
rect 0 11704 480 11734
rect 8661 11731 8727 11734
rect 7808 11456 8128 11457
rect 0 11386 480 11416
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 6637 11386 6703 11389
rect 0 11384 6703 11386
rect 0 11328 6642 11384
rect 6698 11328 6703 11384
rect 0 11326 6703 11328
rect 0 11296 480 11326
rect 6637 11323 6703 11326
rect 4376 10912 4696 10913
rect 0 10842 480 10872
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 4061 10842 4127 10845
rect 0 10840 4127 10842
rect 0 10784 4066 10840
rect 4122 10784 4127 10840
rect 0 10782 4127 10784
rect 0 10752 480 10782
rect 4061 10779 4127 10782
rect 0 10434 480 10464
rect 4061 10434 4127 10437
rect 0 10432 4127 10434
rect 0 10376 4066 10432
rect 4122 10376 4127 10432
rect 0 10374 4127 10376
rect 0 10344 480 10374
rect 4061 10371 4127 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 10303 14992 10304
rect 0 10026 480 10056
rect 2865 10026 2931 10029
rect 0 10024 2931 10026
rect 0 9968 2870 10024
rect 2926 9968 2931 10024
rect 0 9966 2931 9968
rect 0 9936 480 9966
rect 2865 9963 2931 9966
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 0 9482 480 9512
rect 3877 9482 3943 9485
rect 0 9480 3943 9482
rect 0 9424 3882 9480
rect 3938 9424 3943 9480
rect 0 9422 3943 9424
rect 0 9392 480 9422
rect 3877 9419 3943 9422
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 0 9074 480 9104
rect 5809 9074 5875 9077
rect 0 9072 5875 9074
rect 0 9016 5814 9072
rect 5870 9016 5875 9072
rect 0 9014 5875 9016
rect 0 8984 480 9014
rect 5809 9011 5875 9014
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 0 8530 480 8560
rect 3969 8530 4035 8533
rect 0 8528 4035 8530
rect 0 8472 3974 8528
rect 4030 8472 4035 8528
rect 0 8470 4035 8472
rect 0 8440 480 8470
rect 3969 8467 4035 8470
rect 4153 8394 4219 8397
rect 4889 8394 4955 8397
rect 4153 8392 4955 8394
rect 4153 8336 4158 8392
rect 4214 8336 4894 8392
rect 4950 8336 4955 8392
rect 4153 8334 4955 8336
rect 4153 8331 4219 8334
rect 4889 8331 4955 8334
rect 2221 8258 2287 8261
rect 4429 8258 4495 8261
rect 2221 8256 4495 8258
rect 2221 8200 2226 8256
rect 2282 8200 4434 8256
rect 4490 8200 4495 8256
rect 2221 8198 4495 8200
rect 2221 8195 2287 8198
rect 4429 8195 4495 8198
rect 7808 8192 8128 8193
rect 0 8122 480 8152
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 3969 8122 4035 8125
rect 0 8120 4035 8122
rect 0 8064 3974 8120
rect 4030 8064 4035 8120
rect 0 8062 4035 8064
rect 0 8032 480 8062
rect 3969 8059 4035 8062
rect 4376 7648 4696 7649
rect 0 7578 480 7608
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 4061 7578 4127 7581
rect 0 7576 4127 7578
rect 0 7520 4066 7576
rect 4122 7520 4127 7576
rect 0 7518 4127 7520
rect 0 7488 480 7518
rect 4061 7515 4127 7518
rect 0 7170 480 7200
rect 5349 7170 5415 7173
rect 0 7168 5415 7170
rect 0 7112 5354 7168
rect 5410 7112 5415 7168
rect 0 7110 5415 7112
rect 0 7080 480 7110
rect 5349 7107 5415 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 7039 14992 7040
rect 0 6762 480 6792
rect 4061 6762 4127 6765
rect 0 6760 4127 6762
rect 0 6704 4066 6760
rect 4122 6704 4127 6760
rect 0 6702 4127 6704
rect 0 6672 480 6702
rect 4061 6699 4127 6702
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 9765 6490 9831 6493
rect 9765 6488 10426 6490
rect 9765 6432 9770 6488
rect 9826 6432 10426 6488
rect 9765 6430 10426 6432
rect 9765 6427 9831 6430
rect 9765 6354 9831 6357
rect 10133 6354 10199 6357
rect 9765 6352 10199 6354
rect 9765 6296 9770 6352
rect 9826 6296 10138 6352
rect 10194 6296 10199 6352
rect 9765 6294 10199 6296
rect 10366 6354 10426 6430
rect 14549 6354 14615 6357
rect 10366 6352 14615 6354
rect 10366 6296 14554 6352
rect 14610 6296 14615 6352
rect 10366 6294 14615 6296
rect 9765 6291 9831 6294
rect 10133 6291 10199 6294
rect 14549 6291 14615 6294
rect 0 6218 480 6248
rect 4061 6218 4127 6221
rect 0 6216 4127 6218
rect 0 6160 4066 6216
rect 4122 6160 4127 6216
rect 0 6158 4127 6160
rect 0 6128 480 6158
rect 4061 6155 4127 6158
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 0 5810 480 5840
rect 4061 5810 4127 5813
rect 0 5808 4127 5810
rect 0 5752 4066 5808
rect 4122 5752 4127 5808
rect 0 5750 4127 5752
rect 0 5720 480 5750
rect 4061 5747 4127 5750
rect 8845 5810 8911 5813
rect 12157 5810 12223 5813
rect 8845 5808 12223 5810
rect 8845 5752 8850 5808
rect 8906 5752 12162 5808
rect 12218 5752 12223 5808
rect 8845 5750 12223 5752
rect 8845 5747 8911 5750
rect 12157 5747 12223 5750
rect 18597 5810 18663 5813
rect 22320 5810 22800 5840
rect 18597 5808 22800 5810
rect 18597 5752 18602 5808
rect 18658 5752 22800 5808
rect 18597 5750 22800 5752
rect 18597 5747 18663 5750
rect 22320 5720 22800 5750
rect 3877 5674 3943 5677
rect 8661 5674 8727 5677
rect 3877 5672 8727 5674
rect 3877 5616 3882 5672
rect 3938 5616 8666 5672
rect 8722 5616 8727 5672
rect 3877 5614 8727 5616
rect 3877 5611 3943 5614
rect 8661 5611 8727 5614
rect 11145 5674 11211 5677
rect 14365 5674 14431 5677
rect 11145 5672 14431 5674
rect 11145 5616 11150 5672
rect 11206 5616 14370 5672
rect 14426 5616 14431 5672
rect 11145 5614 14431 5616
rect 11145 5611 11211 5614
rect 14365 5611 14431 5614
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 0 5266 480 5296
rect 3417 5266 3483 5269
rect 0 5264 3483 5266
rect 0 5208 3422 5264
rect 3478 5208 3483 5264
rect 0 5206 3483 5208
rect 0 5176 480 5206
rect 3417 5203 3483 5206
rect 5625 5266 5691 5269
rect 11881 5266 11947 5269
rect 5625 5264 11947 5266
rect 5625 5208 5630 5264
rect 5686 5208 11886 5264
rect 11942 5208 11947 5264
rect 5625 5206 11947 5208
rect 5625 5203 5691 5206
rect 11881 5203 11947 5206
rect 7808 4928 8128 4929
rect 0 4858 480 4888
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 2221 4858 2287 4861
rect 0 4856 2287 4858
rect 0 4800 2226 4856
rect 2282 4800 2287 4856
rect 0 4798 2287 4800
rect 0 4768 480 4798
rect 2221 4795 2287 4798
rect 10869 4722 10935 4725
rect 17033 4722 17099 4725
rect 10869 4720 17099 4722
rect 10869 4664 10874 4720
rect 10930 4664 17038 4720
rect 17094 4664 17099 4720
rect 10869 4662 17099 4664
rect 10869 4659 10935 4662
rect 17033 4659 17099 4662
rect 4376 4384 4696 4385
rect 0 4314 480 4344
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 4061 4314 4127 4317
rect 0 4312 4127 4314
rect 0 4256 4066 4312
rect 4122 4256 4127 4312
rect 0 4254 4127 4256
rect 0 4224 480 4254
rect 4061 4251 4127 4254
rect 0 3906 480 3936
rect 3969 3906 4035 3909
rect 0 3904 4035 3906
rect 0 3848 3974 3904
rect 4030 3848 4035 3904
rect 0 3846 4035 3848
rect 0 3816 480 3846
rect 3969 3843 4035 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 3775 14992 3776
rect 2773 3634 2839 3637
rect 6729 3634 6795 3637
rect 2773 3632 6795 3634
rect 2773 3576 2778 3632
rect 2834 3576 6734 3632
rect 6790 3576 6795 3632
rect 2773 3574 6795 3576
rect 2773 3571 2839 3574
rect 6729 3571 6795 3574
rect 0 3498 480 3528
rect 4061 3498 4127 3501
rect 0 3496 4127 3498
rect 0 3440 4066 3496
rect 4122 3440 4127 3496
rect 0 3438 4127 3440
rect 0 3408 480 3438
rect 4061 3435 4127 3438
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 3969 3090 4035 3093
rect 6085 3090 6151 3093
rect 9581 3090 9647 3093
rect 3969 3088 9647 3090
rect 3969 3032 3974 3088
rect 4030 3032 6090 3088
rect 6146 3032 9586 3088
rect 9642 3032 9647 3088
rect 3969 3030 9647 3032
rect 3969 3027 4035 3030
rect 6085 3027 6151 3030
rect 9581 3027 9647 3030
rect 11881 3090 11947 3093
rect 16389 3090 16455 3093
rect 11881 3088 16455 3090
rect 11881 3032 11886 3088
rect 11942 3032 16394 3088
rect 16450 3032 16455 3088
rect 11881 3030 16455 3032
rect 11881 3027 11947 3030
rect 16389 3027 16455 3030
rect 0 2954 480 2984
rect 1669 2954 1735 2957
rect 0 2952 1735 2954
rect 0 2896 1674 2952
rect 1730 2896 1735 2952
rect 0 2894 1735 2896
rect 0 2864 480 2894
rect 1669 2891 1735 2894
rect 4889 2954 4955 2957
rect 9673 2954 9739 2957
rect 4889 2952 9739 2954
rect 4889 2896 4894 2952
rect 4950 2896 9678 2952
rect 9734 2896 9739 2952
rect 4889 2894 9739 2896
rect 4889 2891 4955 2894
rect 9673 2891 9739 2894
rect 3785 2818 3851 2821
rect 7281 2818 7347 2821
rect 3785 2816 7347 2818
rect 3785 2760 3790 2816
rect 3846 2760 7286 2816
rect 7342 2760 7347 2816
rect 3785 2758 7347 2760
rect 3785 2755 3851 2758
rect 7281 2755 7347 2758
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 0 2546 480 2576
rect 3877 2546 3943 2549
rect 0 2544 3943 2546
rect 0 2488 3882 2544
rect 3938 2488 3943 2544
rect 0 2486 3943 2488
rect 0 2456 480 2486
rect 3877 2483 3943 2486
rect 3417 2410 3483 2413
rect 8753 2410 8819 2413
rect 3417 2408 8819 2410
rect 3417 2352 3422 2408
rect 3478 2352 8758 2408
rect 8814 2352 8819 2408
rect 3417 2350 8819 2352
rect 3417 2347 3483 2350
rect 8753 2347 8819 2350
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 0 2002 480 2032
rect 1301 2002 1367 2005
rect 0 2000 1367 2002
rect 0 1944 1306 2000
rect 1362 1944 1367 2000
rect 0 1942 1367 1944
rect 0 1912 480 1942
rect 1301 1939 1367 1942
rect 0 1594 480 1624
rect 2865 1594 2931 1597
rect 0 1592 2931 1594
rect 0 1536 2870 1592
rect 2926 1536 2931 1592
rect 0 1534 2931 1536
rect 0 1504 480 1534
rect 2865 1531 2931 1534
rect 0 1050 480 1080
rect 3325 1050 3391 1053
rect 0 1048 3391 1050
rect 0 992 3330 1048
rect 3386 992 3391 1048
rect 0 990 3391 992
rect 0 960 480 990
rect 3325 987 3391 990
rect 0 642 480 672
rect 3325 642 3391 645
rect 0 640 3391 642
rect 0 584 3330 640
rect 3386 584 3391 640
rect 0 582 3391 584
rect 0 552 480 582
rect 3325 579 3391 582
rect 0 234 480 264
rect 3969 234 4035 237
rect 0 232 4035 234
rect 0 176 3974 232
rect 4030 176 4035 232
rect 0 174 4035 176
rect 0 144 480 174
rect 3969 171 4035 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2116 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1932 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1606821651
transform 1 0 2944 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606821651
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2760 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 3864 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1606821651
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32
timestamp 1606821651
transform 1 0 4048 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40
timestamp 1606821651
transform 1 0 4784 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_27
timestamp 1606821651
transform 1 0 3588 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5704 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4968 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606821651
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606821651
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51
timestamp 1606821651
transform 1 0 5796 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59
timestamp 1606821651
transform 1 0 6532 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_46 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 5336 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1606821651
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1606821651
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7268 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1606821651
transform 1 0 8004 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72
timestamp 1606821651
transform 1 0 7728 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 7176 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_83
timestamp 1606821651
transform 1 0 8740 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _058_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 9016 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1606821651
transform 1 0 9936 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8924 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606821651
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_84
timestamp 1606821651
transform 1 0 8832 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89
timestamp 1606821651
transform 1 0 9292 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1606821651
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_94
timestamp 1606821651
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1606821651
transform 1 0 10764 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_111
timestamp 1606821651
transform 1 0 11316 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11316 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 10764 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _110_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 11500 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1606821651
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1606821651
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117
timestamp 1606821651
transform 1 0 11868 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606821651
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 12420 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1606821651
transform 1 0 12052 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606821651
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1606821651
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_129
timestamp 1606821651
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_129
timestamp 1606821651
transform 1 0 12972 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1606821651
transform 1 0 13156 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_141
timestamp 1606821651
transform 1 0 14076 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_135
timestamp 1606821651
transform 1 0 13524 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_140
timestamp 1606821651
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1606821651
transform 1 0 13708 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1606821651
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1606821651
transform 1 0 13708 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1606821651
transform 1 0 14260 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_147
timestamp 1606821651
transform 1 0 14628 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_152
timestamp 1606821651
transform 1 0 15088 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_146
timestamp 1606821651
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 14904 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1606821651
transform 1 0 14720 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_156
timestamp 1606821651
transform 1 0 15456 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606821651
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 15640 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1606821651
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_164
timestamp 1606821651
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_166
timestamp 1606821651
transform 1 0 16376 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_160
timestamp 1606821651
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1606821651
transform 1 0 16376 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1606821651
transform 1 0 16008 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_176
timestamp 1606821651
transform 1 0 17296 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_170
timestamp 1606821651
transform 1 0 16744 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1606821651
transform 1 0 16928 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1606821651
transform 1 0 16652 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1606821651
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1606821651
transform 1 0 18124 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606821651
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606821651
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1606821651
transform 1 0 17480 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_173
timestamp 1606821651
transform 1 0 17020 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1606821651
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1606821651
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_208
timestamp 1606821651
transform 1 0 20240 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1606821651
transform 1 0 20516 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606821651
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606821651
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606821651
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1606821651
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1606821651
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1606821651
transform 1 0 20884 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_219
timestamp 1606821651
transform 1 0 21252 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 1564 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606821651
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1606821651
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1606821651
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 4508 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606821651
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_21
timestamp 1606821651
transform 1 0 3036 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1606821651
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_35
timestamp 1606821651
transform 1 0 4324 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1606821651
transform 1 0 6348 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_53
timestamp 1606821651
transform 1 0 5980 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7728 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_2_66
timestamp 1606821651
transform 1 0 7176 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9752 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606821651
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_88
timestamp 1606821651
transform 1 0 9200 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_93
timestamp 1606821651
transform 1 0 9660 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_103
timestamp 1606821651
transform 1 0 10580 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10764 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 12420 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_121
timestamp 1606821651
transform 1 0 12236 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1606821651
transform 1 0 14076 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_139
timestamp 1606821651
transform 1 0 13892 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1606821651
transform 1 0 15364 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 16376 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606821651
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_150
timestamp 1606821651
transform 1 0 14904 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_154
timestamp 1606821651
transform 1 0 15272 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_164
timestamp 1606821651
transform 1 0 16192 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1606821651
transform 1 0 17756 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1606821651
transform 1 0 17204 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_172
timestamp 1606821651
transform 1 0 16928 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_179
timestamp 1606821651
transform 1 0 17572 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_185
timestamp 1606821651
transform 1 0 18124 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1606821651
transform 1 0 19964 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_197
timestamp 1606821651
transform 1 0 19228 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606821651
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606821651
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1606821651
transform 1 0 20332 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1606821651
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1606821651
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1606821651
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2944 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1606821651
transform 1 0 1932 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606821651
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1606821651
transform 1 0 1380 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_18
timestamp 1606821651
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_36
timestamp 1606821651
transform 1 0 4416 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5060 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606821651
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_42
timestamp 1606821651
transform 1 0 4968 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1606821651
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_62
timestamp 1606821651
transform 1 0 6808 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1606821651
transform 1 0 6900 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1606821651
transform 1 0 7728 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8740 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_3_66
timestamp 1606821651
transform 1 0 7176 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_81
timestamp 1606821651
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9752 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_92
timestamp 1606821651
transform 1 0 9568 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1606821651
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 11408 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606821651
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1606821651
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_118
timestamp 1606821651
transform 1 0 11960 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13248 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_3_126
timestamp 1606821651
transform 1 0 12696 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 14904 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_148
timestamp 1606821651
transform 1 0 14720 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1606821651
transform 1 0 16376 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16560 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606821651
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_177
timestamp 1606821651
transform 1 0 17388 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1606821651
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1606821651
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1606821651
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606821651
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 1748 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606821651
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1606821651
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _069_
timestamp 1606821651
transform 1 0 3404 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1606821651
transform 1 0 4508 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606821651
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_23
timestamp 1606821651
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_28
timestamp 1606821651
transform 1 0 3680 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1606821651
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_36
timestamp 1606821651
transform 1 0 4416 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5520 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1606821651
transform 1 0 6532 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_46
timestamp 1606821651
transform 1 0 5336 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_57
timestamp 1606821651
transform 1 0 6348 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1606821651
transform 1 0 7820 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_68
timestamp 1606821651
transform 1 0 7360 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_72
timestamp 1606821651
transform 1 0 7728 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_82
timestamp 1606821651
transform 1 0 8648 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9660 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606821651
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1606821651
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 12420 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 11684 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_109
timestamp 1606821651
transform 1 0 11132 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_121
timestamp 1606821651
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13708 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_4_129
timestamp 1606821651
transform 1 0 12972 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15364 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606821651
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_146
timestamp 1606821651
transform 1 0 14536 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 1606821651
transform 1 0 15088 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_154
timestamp 1606821651
transform 1 0 15272 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 17940 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 17020 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_171
timestamp 1606821651
transform 1 0 16836 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_179
timestamp 1606821651
transform 1 0 17572 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_199
timestamp 1606821651
transform 1 0 19412 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606821651
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606821651
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_211
timestamp 1606821651
transform 1 0 20516 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1606821651
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1606821651
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1606821651
transform 1 0 2760 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1606821651
transform 1 0 1748 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606821651
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1606821651
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_16
timestamp 1606821651
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1606821651
transform 1 0 4140 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_5_27
timestamp 1606821651
transform 1 0 3588 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5704 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606821651
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_42
timestamp 1606821651
transform 1 0 4968 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1606821651
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_62
timestamp 1606821651
transform 1 0 6808 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 6900 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 8740 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_79
timestamp 1606821651
transform 1 0 8372 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10396 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_5_99
timestamp 1606821651
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 11592 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606821651
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_110
timestamp 1606821651
transform 1 0 11224 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1606821651
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 13616 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 14352 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_132
timestamp 1606821651
transform 1 0 13248 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_142
timestamp 1606821651
transform 1 0 14168 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1606821651
transform 1 0 15272 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16284 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_150
timestamp 1606821651
transform 1 0 14904 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_163
timestamp 1606821651
transform 1 0 16100 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _066_
timestamp 1606821651
transform 1 0 17296 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606821651
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_174
timestamp 1606821651
transform 1 0 17112 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_179
timestamp 1606821651
transform 1 0 17572 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1606821651
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1606821651
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1606821651
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606821651
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 1380 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1606821651
transform 1 0 2576 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1606821651
transform 1 0 1564 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606821651
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606821651
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1606821651
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_14
timestamp 1606821651
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_19
timestamp 1606821651
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1606821651
transform 1 0 3036 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 3680 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606821651
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_25
timestamp 1606821651
transform 1 0 3404 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_41
timestamp 1606821651
transform 1 0 4876 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_24
timestamp 1606821651
transform 1 0 3312 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 5520 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5612 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606821651
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_47
timestamp 1606821651
transform 1 0 5428 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_44
timestamp 1606821651
transform 1 0 5152 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_48
timestamp 1606821651
transform 1 0 5520 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_58
timestamp 1606821651
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8188 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8556 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1606821651
transform 1 0 7176 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_64
timestamp 1606821651
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_75
timestamp 1606821651
transform 1 0 8004 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_71
timestamp 1606821651
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1606821651
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10488 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9844 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606821651
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 10212 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1606821651
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_96
timestamp 1606821651
transform 1 0 9936 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_93
timestamp 1606821651
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_104
timestamp 1606821651
transform 1 0 10672 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 12144 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 12512 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1606821651
transform 1 0 11132 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606821651
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_118
timestamp 1606821651
transform 1 0 11960 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_108
timestamp 1606821651
transform 1 0 11040 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_118
timestamp 1606821651
transform 1 0 11960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_123
timestamp 1606821651
transform 1 0 12420 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1606821651
transform 1 0 14168 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13800 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_136
timestamp 1606821651
transform 1 0 13616 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_140
timestamp 1606821651
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_151
timestamp 1606821651
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_152
timestamp 1606821651
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_147
timestamp 1606821651
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 14812 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606821651
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1606821651
transform 1 0 15180 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 15272 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_7_162
timestamp 1606821651
transform 1 0 16008 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_160
timestamp 1606821651
transform 1 0 15824 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 16284 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 16008 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1606821651
transform 1 0 17664 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606821651
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_178
timestamp 1606821651
transform 1 0 17480 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_184
timestamp 1606821651
transform 1 0 18032 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1606821651
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1606821651
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_196
timestamp 1606821651
transform 1 0 19136 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_208
timestamp 1606821651
transform 1 0 20240 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1606821651
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1606821651
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606821651
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606821651
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606821651
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1606821651
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1606821651
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 1932 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606821651
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1606821651
transform 1 0 1380 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1606821651
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606821651
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_25
timestamp 1606821651
transform 1 0 3404 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_41
timestamp 1606821651
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 5336 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 5060 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_62
timestamp 1606821651
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6992 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1606821651
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10028 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606821651
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_93
timestamp 1606821651
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 11040 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_106
timestamp 1606821651
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_124
timestamp 1606821651
transform 1 0 12512 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13064 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15272 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606821651
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_146
timestamp 1606821651
transform 1 0 14536 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1606821651
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 16928 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_170
timestamp 1606821651
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1606821651
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1606821651
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1606821651
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606821651
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606821651
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1606821651
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1606821651
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1606821651
transform 1 0 1932 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606821651
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1606821651
transform 1 0 1380 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_9_18
timestamp 1606821651
transform 1 0 2760 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4416 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1606821651
transform 1 0 3036 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_9_30
timestamp 1606821651
transform 1 0 3864 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1606821651
transform 1 0 6256 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606821651
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1606821651
transform 1 0 5888 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1606821651
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8096 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_71
timestamp 1606821651
transform 1 0 7636 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_75
timestamp 1606821651
transform 1 0 8004 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10304 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_9_85
timestamp 1606821651
transform 1 0 8924 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_97
timestamp 1606821651
transform 1 0 10028 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1606821651
transform 1 0 12420 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606821651
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 11960 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_116
timestamp 1606821651
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1606821651
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1606821651
transform 1 0 13616 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1606821651
transform 1 0 14260 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_126
timestamp 1606821651
transform 1 0 12696 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_134
timestamp 1606821651
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_139
timestamp 1606821651
transform 1 0 13892 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _067_
timestamp 1606821651
transform 1 0 15548 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_152
timestamp 1606821651
transform 1 0 15088 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_156
timestamp 1606821651
transform 1 0 15456 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_160
timestamp 1606821651
transform 1 0 15824 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 16928 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606821651
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_178
timestamp 1606821651
transform 1 0 17480 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1606821651
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1606821651
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1606821651
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1606821651
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606821651
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1606821651
transform 1 0 2208 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606821651
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1606821651
transform 1 0 1380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_11
timestamp 1606821651
transform 1 0 2116 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1606821651
transform 1 0 3220 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1606821651
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606821651
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 3680 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_21
timestamp 1606821651
transform 1 0 3036 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1606821651
transform 1 0 3496 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_41
timestamp 1606821651
transform 1 0 4876 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 5152 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_60
timestamp 1606821651
transform 1 0 6624 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1606821651
transform 1 0 8188 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1606821651
transform 1 0 6992 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_10_73
timestamp 1606821651
transform 1 0 7820 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10212 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606821651
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_86
timestamp 1606821651
transform 1 0 9016 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_93
timestamp 1606821651
transform 1 0 9660 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11224 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_108
timestamp 1606821651
transform 1 0 11040 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_119
timestamp 1606821651
transform 1 0 12052 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_131
timestamp 1606821651
transform 1 0 13156 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_143
timestamp 1606821651
transform 1 0 14260 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15272 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606821651
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1606821651
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_170
timestamp 1606821651
transform 1 0 16744 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_182
timestamp 1606821651
transform 1 0 17848 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_194
timestamp 1606821651
transform 1 0 18952 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_206
timestamp 1606821651
transform 1 0 20056 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606821651
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606821651
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1606821651
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1606821651
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 2760 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1606821651
transform 1 0 1748 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606821651
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1606821651
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_16
timestamp 1606821651
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4416 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_34
timestamp 1606821651
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1606821651
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5428 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606821651
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 6440 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_45
timestamp 1606821651
transform 1 0 5244 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_56
timestamp 1606821651
transform 1 0 6256 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7360 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_11_65
timestamp 1606821651
transform 1 0 7084 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9660 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 9200 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_84
timestamp 1606821651
transform 1 0 8832 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_91
timestamp 1606821651
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _068_
timestamp 1606821651
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606821651
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 11776 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_109
timestamp 1606821651
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_114
timestamp 1606821651
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_119
timestamp 1606821651
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1606821651
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1606821651
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1606821651
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1606821651
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606821651
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1606821651
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1606821651
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1606821651
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1606821651
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606821651
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 1380 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606821651
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_19
timestamp 1606821651
transform 1 0 2852 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1606821651
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606821651
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1606821651
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1606821651
transform 1 0 6348 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1606821651
transform 1 0 5060 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_52
timestamp 1606821651
transform 1 0 5888 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_56
timestamp 1606821651
transform 1 0 6256 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 7544 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8556 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_66
timestamp 1606821651
transform 1 0 7176 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_79
timestamp 1606821651
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10028 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606821651
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1606821651
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1606821651
transform 1 0 9660 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_113
timestamp 1606821651
transform 1 0 11500 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_125
timestamp 1606821651
transform 1 0 12604 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_137
timestamp 1606821651
transform 1 0 13708 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606821651
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1606821651
transform 1 0 14812 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1606821651
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1606821651
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1606821651
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1606821651
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1606821651
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606821651
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606821651
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1606821651
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1606821651
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 1564 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1606821651
transform 1 0 2668 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606821651
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606821651
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1606821651
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1606821651
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_15
timestamp 1606821651
transform 1 0 2484 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4232 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 3496 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606821651
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_21
timestamp 1606821651
transform 1 0 3036 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_25
timestamp 1606821651
transform 1 0 3404 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_26
timestamp 1606821651
transform 1 0 3496 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_30
timestamp 1606821651
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 1606821651
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_50
timestamp 1606821651
transform 1 0 5704 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_42
timestamp 1606821651
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 5888 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_58
timestamp 1606821651
transform 1 0 6440 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_58
timestamp 1606821651
transform 1 0 6440 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_53
timestamp 1606821651
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606821651
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1606821651
transform 1 0 6164 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6808 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1606821651
transform 1 0 7820 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8740 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1606821651
transform 1 0 8464 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_71
timestamp 1606821651
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_76
timestamp 1606821651
transform 1 0 8096 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_82
timestamp 1606821651
transform 1 0 8648 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_78
timestamp 1606821651
transform 1 0 8280 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606821651
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 9844 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 10396 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_99
timestamp 1606821651
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_104
timestamp 1606821651
transform 1 0 10672 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_89
timestamp 1606821651
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1606821651
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606821651
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_116
timestamp 1606821651
transform 1 0 11776 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1606821651
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_115
timestamp 1606821651
transform 1 0 11684 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1606821651
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_127
timestamp 1606821651
transform 1 0 12788 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_139
timestamp 1606821651
transform 1 0 13892 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606821651
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_147
timestamp 1606821651
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_159
timestamp 1606821651
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1606821651
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1606821651
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1606821651
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606821651
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_171
timestamp 1606821651
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1606821651
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1606821651
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1606821651
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1606821651
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_190
timestamp 1606821651
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_202
timestamp 1606821651
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606821651
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606821651
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606821651
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1606821651
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1606821651
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 1564 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606821651
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1606821651
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1606821651
transform 1 0 3680 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_15_21
timestamp 1606821651
transform 1 0 3036 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_27
timestamp 1606821651
transform 1 0 3588 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_37
timestamp 1606821651
transform 1 0 4508 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_41
timestamp 1606821651
transform 1 0 4876 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4968 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606821651
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_58
timestamp 1606821651
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_62
timestamp 1606821651
transform 1 0 6808 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7636 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 7176 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_69
timestamp 1606821651
transform 1 0 7452 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1606821651
transform 1 0 9384 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9660 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10488 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_87
timestamp 1606821651
transform 1 0 9108 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606821651
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_111
timestamp 1606821651
transform 1 0 11316 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_119
timestamp 1606821651
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1606821651
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1606821651
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_147
timestamp 1606821651
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_159
timestamp 1606821651
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1606821651
transform 1 0 18216 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606821651
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_171
timestamp 1606821651
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_184
timestamp 1606821651
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_190
timestamp 1606821651
transform 1 0 18584 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_202
timestamp 1606821651
transform 1 0 19688 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606821651
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_214
timestamp 1606821651
transform 1 0 20792 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1606821651
transform 1 0 2300 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606821651
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1606821651
transform 1 0 1380 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_11
timestamp 1606821651
transform 1 0 2116 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1606821651
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1606821651
transform 1 0 3312 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4508 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606821651
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_22
timestamp 1606821651
transform 1 0 3128 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1606821651
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_35
timestamp 1606821651
transform 1 0 4324 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5520 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_46
timestamp 1606821651
transform 1 0 5336 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_57
timestamp 1606821651
transform 1 0 6348 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6900 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8556 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_72
timestamp 1606821651
transform 1 0 7728 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_80
timestamp 1606821651
transform 1 0 8464 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9660 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606821651
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1606821651
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1606821651
transform 1 0 11132 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1606821651
transform 1 0 12236 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_133
timestamp 1606821651
transform 1 0 13340 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_145
timestamp 1606821651
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606821651
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1606821651
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1606821651
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1606821651
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1606821651
transform 1 0 18584 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_194
timestamp 1606821651
transform 1 0 18952 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_206
timestamp 1606821651
transform 1 0 20056 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606821651
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606821651
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1606821651
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1606821651
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 2116 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606821651
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1606821651
transform 1 0 1380 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1606821651
transform 1 0 3772 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_27
timestamp 1606821651
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_38
timestamp 1606821651
transform 1 0 4600 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4968 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606821651
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_58
timestamp 1606821651
transform 1 0 6440 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1606821651
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1606821651
transform 1 0 8740 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1606821651
transform 1 0 7728 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 6992 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_67
timestamp 1606821651
transform 1 0 7268 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_71
timestamp 1606821651
transform 1 0 7636 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_81
timestamp 1606821651
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9292 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_17_86
timestamp 1606821651
transform 1 0 9016 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606821651
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_105
timestamp 1606821651
transform 1 0 10764 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_117
timestamp 1606821651
transform 1 0 11868 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1606821651
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1606821651
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1606821651
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_147
timestamp 1606821651
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_159
timestamp 1606821651
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606821651
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_171
timestamp 1606821651
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_184
timestamp 1606821651
transform 1 0 18032 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1606821651
transform 1 0 19044 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_192
timestamp 1606821651
transform 1 0 18768 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_199
timestamp 1606821651
transform 1 0 19412 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606821651
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_211
timestamp 1606821651
transform 1 0 20516 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_219
timestamp 1606821651
transform 1 0 21252 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1606821651
transform 1 0 1472 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1606821651
transform 1 0 2024 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606821651
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1606821651
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_8
timestamp 1606821651
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_19
timestamp 1606821651
transform 1 0 2852 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1606821651
transform 1 0 3036 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4508 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606821651
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 4232 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_25
timestamp 1606821651
transform 1 0 3404 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_32
timestamp 1606821651
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 5520 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_46
timestamp 1606821651
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7268 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_64
timestamp 1606821651
transform 1 0 6992 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_83
timestamp 1606821651
transform 1 0 8740 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606821651
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1606821651
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_102
timestamp 1606821651
transform 1 0 10488 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_114
timestamp 1606821651
transform 1 0 11592 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_126
timestamp 1606821651
transform 1 0 12696 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_138
timestamp 1606821651
transform 1 0 13800 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606821651
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_150
timestamp 1606821651
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1606821651
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1606821651
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1606821651
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1606821651
transform 1 0 19504 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_190
timestamp 1606821651
transform 1 0 18584 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_198
timestamp 1606821651
transform 1 0 19320 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_204
timestamp 1606821651
transform 1 0 19872 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606821651
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606821651
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1606821651
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1606821651
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1606821651
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1606821651
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1606821651
transform 1 0 1748 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1606821651
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606821651
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606821651
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1840 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1656 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_12
timestamp 1606821651
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_18
timestamp 1606821651
transform 1 0 2760 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_14
timestamp 1606821651
transform 1 0 2392 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1606821651
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2852 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1606821651
transform 1 0 4508 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1606821651
transform 1 0 3404 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4048 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606821651
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_35
timestamp 1606821651
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_40
timestamp 1606821651
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1606821651
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1606821651
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4968 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5704 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606821651
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_58
timestamp 1606821651
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_62
timestamp 1606821651
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_48
timestamp 1606821651
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_59
timestamp 1606821651
transform 1 0 6532 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1606821651
transform 1 0 7176 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7636 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1606821651
transform 1 0 7544 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 7084 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_69
timestamp 1606821651
transform 1 0 7452 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_68
timestamp 1606821651
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_79
timestamp 1606821651
transform 1 0 8372 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606821651
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 10028 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_87
timestamp 1606821651
transform 1 0 9108 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_95
timestamp 1606821651
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_100
timestamp 1606821651
transform 1 0 10304 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1606821651
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_102
timestamp 1606821651
transform 1 0 10488 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606821651
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_112
timestamp 1606821651
transform 1 0 11408 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1606821651
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1606821651
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_114
timestamp 1606821651
transform 1 0 11592 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1606821651
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_126
timestamp 1606821651
transform 1 0 12696 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_138
timestamp 1606821651
transform 1 0 13800 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606821651
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1606821651
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_159
timestamp 1606821651
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_150
timestamp 1606821651
transform 1 0 14904 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1606821651
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1606821651
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606821651
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_171
timestamp 1606821651
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1606821651
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1606821651
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1606821651
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1606821651
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_190
timestamp 1606821651
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1606821651
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606821651
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606821651
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606821651
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1606821651
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1606821651
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1656 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2208 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606821651
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1606821651
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_18
timestamp 1606821651
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4140 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1606821651
transform 1 0 3128 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_31
timestamp 1606821651
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1606821651
transform 1 0 5796 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6808 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606821651
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_49
timestamp 1606821651
transform 1 0 5612 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_54
timestamp 1606821651
transform 1 0 6072 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp 1606821651
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 8556 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_21_78
timestamp 1606821651
transform 1 0 8280 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1606821651
transform 1 0 10212 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_97
timestamp 1606821651
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_102
timestamp 1606821651
transform 1 0 10488 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606821651
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_114
timestamp 1606821651
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1606821651
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1606821651
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1606821651
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_159
timestamp 1606821651
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606821651
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_171
timestamp 1606821651
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1606821651
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1606821651
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1606821651
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606821651
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 2116 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1380 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606821651
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_9
timestamp 1606821651
transform 1 0 1932 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4416 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606821651
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1606821651
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_32
timestamp 1606821651
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1606821651
transform 1 0 5796 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6256 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_22_45
timestamp 1606821651
transform 1 0 5244 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_54
timestamp 1606821651
transform 1 0 6072 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8556 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_72
timestamp 1606821651
transform 1 0 7728 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_80
timestamp 1606821651
transform 1 0 8464 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9660 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606821651
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 1606821651
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1606821651
transform 1 0 11132 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1606821651
transform 1 0 12236 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_133
timestamp 1606821651
transform 1 0 13340 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_145
timestamp 1606821651
transform 1 0 14444 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606821651
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1606821651
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1606821651
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1606821651
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1606821651
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1606821651
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606821651
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606821651
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1606821651
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1606821651
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1606821651
transform 1 0 1472 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2760 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2024 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606821651
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_3
timestamp 1606821651
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_8
timestamp 1606821651
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_16
timestamp 1606821651
transform 1 0 2576 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4600 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1606821651
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_34
timestamp 1606821651
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5704 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606821651
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_47
timestamp 1606821651
transform 1 0 5428 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1606821651
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_62
timestamp 1606821651
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1606821651
transform 1 0 6992 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8188 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1606821651
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_75
timestamp 1606821651
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9200 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1606821651
transform 1 0 9016 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_104
timestamp 1606821651
transform 1 0 10672 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606821651
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_116
timestamp 1606821651
transform 1 0 11776 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1606821651
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1606821651
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1606821651
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1606821651
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606821651
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1606821651
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1606821651
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1606821651
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1606821651
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606821651
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1606821651
transform 1 0 1564 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1606821651
transform 1 0 2852 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2116 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606821651
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1606821651
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_9
timestamp 1606821651
transform 1 0 1932 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_17
timestamp 1606821651
transform 1 0 2668 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606821651
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_28
timestamp 1606821651
transform 1 0 3680 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_41
timestamp 1606821651
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1606821651
transform 1 0 5060 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5888 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_24_46
timestamp 1606821651
transform 1 0 5336 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7728 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_68
timestamp 1606821651
transform 1 0 7360 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606821651
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1606821651
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_88
timestamp 1606821651
transform 1 0 9200 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_104
timestamp 1606821651
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11040 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1606821651
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1606821651
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1606821651
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1606821651
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606821651
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1606821651
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1606821651
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1606821651
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1606821651
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1606821651
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606821651
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606821651
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1606821651
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1606821651
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1606821651
transform 1 0 2760 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1606821651
transform 1 0 1472 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2024 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606821651
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1606821651
transform 1 0 1380 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_8
timestamp 1606821651
transform 1 0 1840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_16
timestamp 1606821651
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 3588 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_22
timestamp 1606821651
transform 1 0 3128 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_26
timestamp 1606821651
transform 1 0 3496 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1606821651
transform 1 0 5244 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5704 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606821651
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_43
timestamp 1606821651
transform 1 0 5060 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_48
timestamp 1606821651
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1606821651
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_62
timestamp 1606821651
transform 1 0 6808 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 8280 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1606821651
transform 1 0 7268 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_25_66
timestamp 1606821651
transform 1 0 7176 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_76
timestamp 1606821651
transform 1 0 8096 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10212 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_94
timestamp 1606821651
transform 1 0 9752 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_98
timestamp 1606821651
transform 1 0 10120 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606821651
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_115
timestamp 1606821651
transform 1 0 11684 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1606821651
transform 1 0 12236 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1606821651
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1606821651
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1606821651
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_159
timestamp 1606821651
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606821651
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_171
timestamp 1606821651
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1606821651
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1606821651
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1606821651
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606821651
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1606821651
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1606821651
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606821651
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606821651
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1656 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1606821651
transform 1 0 1564 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_9
timestamp 1606821651
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_12
timestamp 1606821651
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2116 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_17
timestamp 1606821651
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_20
timestamp 1606821651
transform 1 0 2944 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2852 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2392 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_31
timestamp 1606821651
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_25
timestamp 1606821651
transform 1 0 3404 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_30
timestamp 1606821651
transform 1 0 3864 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_26
timestamp 1606821651
transform 1 0 3496 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606821651
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1606821651
transform 1 0 3128 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1606821651
transform 1 0 3588 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_32
timestamp 1606821651
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1606821651
transform 1 0 4140 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_36
timestamp 1606821651
transform 1 0 4416 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4416 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6072 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5520 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606821651
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_52
timestamp 1606821651
transform 1 0 5888 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1606821651
transform 1 0 6348 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1606821651
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1606821651
transform 1 0 8096 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 8464 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_70
timestamp 1606821651
transform 1 0 7544 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_79
timestamp 1606821651
transform 1 0 8372 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_74
timestamp 1606821651
transform 1 0 7912 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1606821651
transform 1 0 9108 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9660 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1606821651
transform 1 0 9200 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606821651
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1606821651
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_86
timestamp 1606821651
transform 1 0 9016 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_97
timestamp 1606821651
transform 1 0 10028 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1606821651
transform 1 0 11776 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 11316 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10764 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606821651
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_109
timestamp 1606821651
transform 1 0 11132 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_114
timestamp 1606821651
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_119
timestamp 1606821651
transform 1 0 12052 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1606821651
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_127
timestamp 1606821651
transform 1 0 12788 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_139
timestamp 1606821651
transform 1 0 13892 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1606821651
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606821651
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_151
timestamp 1606821651
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1606821651
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1606821651
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1606821651
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1606821651
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606821651
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1606821651
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1606821651
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1606821651
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1606821651
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1606821651
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1606821651
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1606821651
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606821651
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606821651
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606821651
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1606821651
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1606821651
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1606821651
transform 1 0 1656 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2208 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606821651
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_3
timestamp 1606821651
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_10
timestamp 1606821651
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_18
timestamp 1606821651
transform 1 0 2760 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606821651
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_30
timestamp 1606821651
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1606821651
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1606821651
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1606821651
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 7912 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_68
timestamp 1606821651
transform 1 0 7360 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1606821651
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 10120 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606821651
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_93
timestamp 1606821651
transform 1 0 9660 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_97
timestamp 1606821651
transform 1 0 10028 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_104
timestamp 1606821651
transform 1 0 10672 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_116
timestamp 1606821651
transform 1 0 11776 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_128
timestamp 1606821651
transform 1 0 12880 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_140
timestamp 1606821651
transform 1 0 13984 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606821651
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_152
timestamp 1606821651
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1606821651
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1606821651
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1606821651
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1606821651
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1606821651
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606821651
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606821651
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1606821651
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1606821651
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1606821651
transform 1 0 2852 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1606821651
transform 1 0 2300 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1606821651
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606821651
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1606821651
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_11
timestamp 1606821651
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_17
timestamp 1606821651
transform 1 0 2668 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1606821651
transform 1 0 3404 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_23
timestamp 1606821651
transform 1 0 3220 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_29
timestamp 1606821651
transform 1 0 3772 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_41
timestamp 1606821651
transform 1 0 4876 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606821651
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_53
timestamp 1606821651
transform 1 0 5980 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1606821651
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1606821651
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1606821651
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1606821651
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606821651
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_110
timestamp 1606821651
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1606821651
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1606821651
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1606821651
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1606821651
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606821651
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1606821651
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1606821651
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1606821651
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1606821651
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606821651
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2116 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2852 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606821651
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1606821651
transform 1 0 1380 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_17
timestamp 1606821651
transform 1 0 2668 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606821651
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_25
timestamp 1606821651
transform 1 0 3404 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1606821651
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1606821651
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_56
timestamp 1606821651
transform 1 0 6256 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1606821651
transform 1 0 7820 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 7084 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_64
timestamp 1606821651
transform 1 0 6992 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_71
timestamp 1606821651
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_77
timestamp 1606821651
transform 1 0 8188 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606821651
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_89
timestamp 1606821651
transform 1 0 9292 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1606821651
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1606821651
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1606821651
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1606821651
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1606821651
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606821651
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1606821651
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1606821651
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_178
timestamp 1606821651
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_190
timestamp 1606821651
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1606821651
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606821651
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606821651
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1606821651
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1606821651
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1606821651
transform 1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1606821651
transform 1 0 2300 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606821651
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1606821651
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1606821651
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_17
timestamp 1606821651
transform 1 0 2668 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_29
timestamp 1606821651
transform 1 0 3772 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_41
timestamp 1606821651
transform 1 0 4876 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1606821651
transform 1 0 6808 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606821651
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_53
timestamp 1606821651
transform 1 0 5980 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_66
timestamp 1606821651
transform 1 0 7176 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_78
timestamp 1606821651
transform 1 0 8280 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_90
timestamp 1606821651
transform 1 0 9384 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_102
timestamp 1606821651
transform 1 0 10488 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606821651
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_114
timestamp 1606821651
transform 1 0 11592 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1606821651
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1606821651
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1606821651
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1606821651
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606821651
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1606821651
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1606821651
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1606821651
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1606821651
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606821651
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1606821651
transform 1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606821651
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1606821651
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_11
timestamp 1606821651
transform 1 0 2116 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606821651
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_23
timestamp 1606821651
transform 1 0 3220 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1606821651
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606821651
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1606821651
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1606821651
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1606821651
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_75
timestamp 1606821651
transform 1 0 8004 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606821651
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_87
timestamp 1606821651
transform 1 0 9108 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1606821651
transform 1 0 9752 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606821651
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_106
timestamp 1606821651
transform 1 0 10856 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_118
timestamp 1606821651
transform 1 0 11960 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_125
timestamp 1606821651
transform 1 0 12604 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_137
timestamp 1606821651
transform 1 0 13708 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606821651
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_149
timestamp 1606821651
transform 1 0 14812 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1606821651
transform 1 0 15456 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606821651
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1606821651
transform 1 0 16560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_180
timestamp 1606821651
transform 1 0 17664 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_187
timestamp 1606821651
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_199
timestamp 1606821651
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606821651
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606821651
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_211
timestamp 1606821651
transform 1 0 20516 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1606821651
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 21638 0 21694 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 22098 0 22154 480 6 SC_OUT_BOT
port 1 nsew default tristate
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_42_
port 2 nsew default input
rlabel metal2 s 570 0 626 480 6 bottom_left_grid_pin_43_
port 3 nsew default input
rlabel metal2 s 1030 0 1086 480 6 bottom_left_grid_pin_44_
port 4 nsew default input
rlabel metal2 s 1490 0 1546 480 6 bottom_left_grid_pin_45_
port 5 nsew default input
rlabel metal2 s 1950 0 2006 480 6 bottom_left_grid_pin_46_
port 6 nsew default input
rlabel metal2 s 2318 0 2374 480 6 bottom_left_grid_pin_47_
port 7 nsew default input
rlabel metal2 s 2778 0 2834 480 6 bottom_left_grid_pin_48_
port 8 nsew default input
rlabel metal2 s 3238 0 3294 480 6 bottom_left_grid_pin_49_
port 9 nsew default input
rlabel metal2 s 21178 0 21234 480 6 bottom_right_grid_pin_1_
port 10 nsew default input
rlabel metal3 s 22320 5720 22800 5840 6 ccff_head
port 11 nsew default input
rlabel metal3 s 22320 17144 22800 17264 6 ccff_tail
port 12 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_in[0]
port 13 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[10]
port 14 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[11]
port 15 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[12]
port 16 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[13]
port 17 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[14]
port 18 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[15]
port 19 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[16]
port 20 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[17]
port 21 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[18]
port 22 nsew default input
rlabel metal3 s 0 12656 480 12776 6 chanx_left_in[19]
port 23 nsew default input
rlabel metal3 s 0 4224 480 4344 6 chanx_left_in[1]
port 24 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[2]
port 25 nsew default input
rlabel metal3 s 0 5176 480 5296 6 chanx_left_in[3]
port 26 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[4]
port 27 nsew default input
rlabel metal3 s 0 6128 480 6248 6 chanx_left_in[5]
port 28 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[6]
port 29 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[7]
port 30 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[8]
port 31 nsew default input
rlabel metal3 s 0 8032 480 8152 6 chanx_left_in[9]
port 32 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chanx_left_out[0]
port 33 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[10]
port 34 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chanx_left_out[11]
port 35 nsew default tristate
rlabel metal3 s 0 18776 480 18896 6 chanx_left_out[12]
port 36 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chanx_left_out[13]
port 37 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_left_out[14]
port 38 nsew default tristate
rlabel metal3 s 0 20136 480 20256 6 chanx_left_out[15]
port 39 nsew default tristate
rlabel metal3 s 0 20544 480 20664 6 chanx_left_out[16]
port 40 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[17]
port 41 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[18]
port 42 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[19]
port 43 nsew default tristate
rlabel metal3 s 0 13608 480 13728 6 chanx_left_out[1]
port 44 nsew default tristate
rlabel metal3 s 0 14016 480 14136 6 chanx_left_out[2]
port 45 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[3]
port 46 nsew default tristate
rlabel metal3 s 0 14968 480 15088 6 chanx_left_out[4]
port 47 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[5]
port 48 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[6]
port 49 nsew default tristate
rlabel metal3 s 0 16464 480 16584 6 chanx_left_out[7]
port 50 nsew default tristate
rlabel metal3 s 0 16872 480 16992 6 chanx_left_out[8]
port 51 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[9]
port 52 nsew default tristate
rlabel metal2 s 3698 0 3754 480 6 chany_bottom_in[0]
port 53 nsew default input
rlabel metal2 s 8022 0 8078 480 6 chany_bottom_in[10]
port 54 nsew default input
rlabel metal2 s 8482 0 8538 480 6 chany_bottom_in[11]
port 55 nsew default input
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_in[12]
port 56 nsew default input
rlabel metal2 s 9402 0 9458 480 6 chany_bottom_in[13]
port 57 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[14]
port 58 nsew default input
rlabel metal2 s 10230 0 10286 480 6 chany_bottom_in[15]
port 59 nsew default input
rlabel metal2 s 10690 0 10746 480 6 chany_bottom_in[16]
port 60 nsew default input
rlabel metal2 s 11150 0 11206 480 6 chany_bottom_in[17]
port 61 nsew default input
rlabel metal2 s 11610 0 11666 480 6 chany_bottom_in[18]
port 62 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chany_bottom_in[19]
port 63 nsew default input
rlabel metal2 s 4066 0 4122 480 6 chany_bottom_in[1]
port 64 nsew default input
rlabel metal2 s 4526 0 4582 480 6 chany_bottom_in[2]
port 65 nsew default input
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_in[3]
port 66 nsew default input
rlabel metal2 s 5446 0 5502 480 6 chany_bottom_in[4]
port 67 nsew default input
rlabel metal2 s 5906 0 5962 480 6 chany_bottom_in[5]
port 68 nsew default input
rlabel metal2 s 6274 0 6330 480 6 chany_bottom_in[6]
port 69 nsew default input
rlabel metal2 s 6734 0 6790 480 6 chany_bottom_in[7]
port 70 nsew default input
rlabel metal2 s 7194 0 7250 480 6 chany_bottom_in[8]
port 71 nsew default input
rlabel metal2 s 7654 0 7710 480 6 chany_bottom_in[9]
port 72 nsew default input
rlabel metal2 s 12438 0 12494 480 6 chany_bottom_out[0]
port 73 nsew default tristate
rlabel metal2 s 16854 0 16910 480 6 chany_bottom_out[10]
port 74 nsew default tristate
rlabel metal2 s 17314 0 17370 480 6 chany_bottom_out[11]
port 75 nsew default tristate
rlabel metal2 s 17682 0 17738 480 6 chany_bottom_out[12]
port 76 nsew default tristate
rlabel metal2 s 18142 0 18198 480 6 chany_bottom_out[13]
port 77 nsew default tristate
rlabel metal2 s 18602 0 18658 480 6 chany_bottom_out[14]
port 78 nsew default tristate
rlabel metal2 s 19062 0 19118 480 6 chany_bottom_out[15]
port 79 nsew default tristate
rlabel metal2 s 19430 0 19486 480 6 chany_bottom_out[16]
port 80 nsew default tristate
rlabel metal2 s 19890 0 19946 480 6 chany_bottom_out[17]
port 81 nsew default tristate
rlabel metal2 s 20350 0 20406 480 6 chany_bottom_out[18]
port 82 nsew default tristate
rlabel metal2 s 20810 0 20866 480 6 chany_bottom_out[19]
port 83 nsew default tristate
rlabel metal2 s 12898 0 12954 480 6 chany_bottom_out[1]
port 84 nsew default tristate
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_out[2]
port 85 nsew default tristate
rlabel metal2 s 13726 0 13782 480 6 chany_bottom_out[3]
port 86 nsew default tristate
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_out[4]
port 87 nsew default tristate
rlabel metal2 s 14646 0 14702 480 6 chany_bottom_out[5]
port 88 nsew default tristate
rlabel metal2 s 15106 0 15162 480 6 chany_bottom_out[6]
port 89 nsew default tristate
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_out[7]
port 90 nsew default tristate
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_out[8]
port 91 nsew default tristate
rlabel metal2 s 16394 0 16450 480 6 chany_bottom_out[9]
port 92 nsew default tristate
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_34_
port 93 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_35_
port 94 nsew default input
rlabel metal3 s 0 960 480 1080 6 left_bottom_grid_pin_36_
port 95 nsew default input
rlabel metal3 s 0 1504 480 1624 6 left_bottom_grid_pin_37_
port 96 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_38_
port 97 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_39_
port 98 nsew default input
rlabel metal3 s 0 2864 480 2984 6 left_bottom_grid_pin_40_
port 99 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_bottom_grid_pin_41_
port 100 nsew default input
rlabel metal3 s 0 22448 480 22568 6 left_top_grid_pin_1_
port 101 nsew default input
rlabel metal2 s 22558 0 22614 480 6 prog_clk_0_S_in
port 102 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 103 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 104 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22568
<< end >>
