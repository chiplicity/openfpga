magic
tech EFS8A
magscale 1 2
timestamp 1602076530
<< locali >>
rect 20223 20553 20361 20587
rect 15243 18785 15370 18819
rect 12811 18071 12845 18139
rect 18423 18071 18457 18139
rect 12811 18037 12817 18071
rect 18423 18037 18429 18071
rect 6779 17765 6824 17799
rect 17083 17697 17118 17731
rect 12719 16745 12725 16779
rect 12719 16677 12753 16745
rect 6377 16609 6538 16643
rect 6377 16575 6411 16609
rect 6653 16031 6687 16133
rect 12081 15895 12115 16065
rect 19211 15589 19257 15623
rect 10051 14569 10057 14603
rect 10051 14501 10085 14569
rect 13369 13787 13403 13957
rect 6831 13481 6837 13515
rect 11615 13481 11621 13515
rect 6831 13413 6865 13481
rect 11615 13413 11649 13481
rect 10183 13345 10310 13379
rect 13645 12835 13679 12937
rect 19291 12257 19418 12291
rect 19067 11305 19073 11339
rect 19067 11237 19101 11305
rect 5727 9129 5733 9163
rect 18331 9129 18337 9163
rect 5727 9061 5761 9129
rect 18331 9061 18365 9129
rect 4387 8993 4422 9027
rect 8671 8279 8705 8347
rect 8671 8245 8677 8279
rect 9999 7905 10034 7939
rect 14139 7905 14266 7939
rect 6503 6817 6538 6851
rect 3151 6103 3185 6171
rect 4899 6103 4933 6171
rect 3151 6069 3157 6103
rect 4899 6069 4905 6103
rect 4905 5627 4939 5729
rect 18607 4777 18613 4811
rect 18607 4709 18641 4777
rect 2915 4641 3042 4675
rect 5583 4029 5710 4063
rect 10517 3383 10551 3553
rect 2145 2499 2179 2601
rect 3709 2295 3743 2533
rect 9723 2465 9850 2499
<< viali >>
rect 8217 20893 8251 20927
rect 18337 20893 18371 20927
rect 1593 20553 1627 20587
rect 5503 20553 5537 20587
rect 8309 20553 8343 20587
rect 11161 20553 11195 20587
rect 19165 20553 19199 20587
rect 20361 20553 20395 20587
rect 7619 20485 7653 20519
rect 2053 20417 2087 20451
rect 8585 20417 8619 20451
rect 1409 20349 1443 20383
rect 5432 20349 5466 20383
rect 5825 20349 5859 20383
rect 7532 20349 7566 20383
rect 10977 20349 11011 20383
rect 11529 20349 11563 20383
rect 12516 20349 12550 20383
rect 18981 20349 19015 20383
rect 20120 20349 20154 20383
rect 20545 20349 20579 20383
rect 8033 20281 8067 20315
rect 8677 20281 8711 20315
rect 9229 20281 9263 20315
rect 19533 20281 19567 20315
rect 7389 20213 7423 20247
rect 12587 20213 12621 20247
rect 13001 20213 13035 20247
rect 8769 20009 8803 20043
rect 5273 19941 5307 19975
rect 8211 19941 8245 19975
rect 10793 19941 10827 19975
rect 18429 19941 18463 19975
rect 18521 19941 18555 19975
rect 4077 19805 4111 19839
rect 5181 19805 5215 19839
rect 5549 19805 5583 19839
rect 7849 19805 7883 19839
rect 10701 19805 10735 19839
rect 11345 19805 11379 19839
rect 19073 19805 19107 19839
rect 9965 19669 9999 19703
rect 18061 19669 18095 19703
rect 5273 19465 5307 19499
rect 10885 19465 10919 19499
rect 11161 19465 11195 19499
rect 17509 19465 17543 19499
rect 18981 19465 19015 19499
rect 21051 19465 21085 19499
rect 4997 19397 5031 19431
rect 5641 19397 5675 19431
rect 7573 19329 7607 19363
rect 9965 19329 9999 19363
rect 4077 19261 4111 19295
rect 7665 19261 7699 19295
rect 8217 19261 8251 19295
rect 16681 19261 16715 19295
rect 16865 19261 16899 19295
rect 18061 19261 18095 19295
rect 20980 19261 21014 19295
rect 21373 19261 21407 19295
rect 4398 19193 4432 19227
rect 7205 19193 7239 19227
rect 10286 19193 10320 19227
rect 17141 19193 17175 19227
rect 18382 19193 18416 19227
rect 3617 19125 3651 19159
rect 3985 19125 4019 19159
rect 7941 19125 7975 19159
rect 8677 19125 8711 19159
rect 9781 19125 9815 19159
rect 11529 19125 11563 19159
rect 16221 19125 16255 19159
rect 17785 19125 17819 19159
rect 1593 18921 1627 18955
rect 6469 18921 6503 18955
rect 9965 18921 9999 18955
rect 18429 18921 18463 18955
rect 4997 18853 5031 18887
rect 11529 18853 11563 18887
rect 17325 18853 17359 18887
rect 18797 18853 18831 18887
rect 1409 18785 1443 18819
rect 6653 18785 6687 18819
rect 6837 18785 6871 18819
rect 8309 18785 8343 18819
rect 8585 18785 8619 18819
rect 9965 18785 9999 18819
rect 10149 18785 10183 18819
rect 15209 18785 15243 18819
rect 16865 18785 16899 18819
rect 17049 18785 17083 18819
rect 4905 18717 4939 18751
rect 5549 18717 5583 18751
rect 8769 18717 8803 18751
rect 11437 18717 11471 18751
rect 11713 18717 11747 18751
rect 18705 18717 18739 18751
rect 19257 18649 19291 18683
rect 3433 18581 3467 18615
rect 7665 18581 7699 18615
rect 10793 18581 10827 18615
rect 12541 18581 12575 18615
rect 15439 18581 15473 18615
rect 16497 18581 16531 18615
rect 1593 18377 1627 18411
rect 4721 18377 4755 18411
rect 6101 18377 6135 18411
rect 17417 18377 17451 18411
rect 18981 18377 19015 18411
rect 19257 18377 19291 18411
rect 5549 18309 5583 18343
rect 9781 18309 9815 18343
rect 11713 18309 11747 18343
rect 13369 18309 13403 18343
rect 16589 18309 16623 18343
rect 6377 18241 6411 18275
rect 7205 18241 7239 18275
rect 8861 18241 8895 18275
rect 11345 18241 11379 18275
rect 15945 18241 15979 18275
rect 18061 18241 18095 18275
rect 3525 18173 3559 18207
rect 3801 18173 3835 18207
rect 10057 18173 10091 18207
rect 12449 18173 12483 18207
rect 19625 18173 19659 18207
rect 19809 18173 19843 18207
rect 20269 18173 20303 18207
rect 4997 18105 5031 18139
rect 5089 18105 5123 18139
rect 6929 18105 6963 18139
rect 7021 18105 7055 18139
rect 9182 18105 9216 18139
rect 10701 18105 10735 18139
rect 10793 18105 10827 18139
rect 15025 18105 15059 18139
rect 15117 18105 15151 18139
rect 15669 18105 15703 18139
rect 3157 18037 3191 18071
rect 3617 18037 3651 18071
rect 4445 18037 4479 18071
rect 8125 18037 8159 18071
rect 8677 18037 8711 18071
rect 10425 18037 10459 18071
rect 12265 18037 12299 18071
rect 12817 18037 12851 18071
rect 14841 18037 14875 18071
rect 16957 18037 16991 18071
rect 17785 18037 17819 18071
rect 18429 18037 18463 18071
rect 19901 18037 19935 18071
rect 4997 17833 5031 17867
rect 6377 17833 6411 17867
rect 8355 17833 8389 17867
rect 8861 17833 8895 17867
rect 11437 17833 11471 17867
rect 15025 17833 15059 17867
rect 16221 17833 16255 17867
rect 19349 17833 19383 17867
rect 21097 17833 21131 17867
rect 4398 17765 4432 17799
rect 6745 17765 6779 17799
rect 10057 17765 10091 17799
rect 12541 17765 12575 17799
rect 15622 17765 15656 17799
rect 18474 17765 18508 17799
rect 2605 17697 2639 17731
rect 2881 17697 2915 17731
rect 5641 17697 5675 17731
rect 6469 17697 6503 17731
rect 8284 17697 8318 17731
rect 11897 17697 11931 17731
rect 12265 17697 12299 17731
rect 13921 17697 13955 17731
rect 14197 17697 14231 17731
rect 17049 17697 17083 17731
rect 18153 17697 18187 17731
rect 20913 17697 20947 17731
rect 3157 17629 3191 17663
rect 4077 17629 4111 17663
rect 9965 17629 9999 17663
rect 14381 17629 14415 17663
rect 15301 17629 15335 17663
rect 10517 17561 10551 17595
rect 13277 17561 13311 17595
rect 19809 17561 19843 17595
rect 5365 17493 5399 17527
rect 7389 17493 7423 17527
rect 7665 17493 7699 17527
rect 8125 17493 8159 17527
rect 10885 17493 10919 17527
rect 12817 17493 12851 17527
rect 17187 17493 17221 17527
rect 19073 17493 19107 17527
rect 3157 17289 3191 17323
rect 4997 17289 5031 17323
rect 6193 17289 6227 17323
rect 8217 17289 8251 17323
rect 8907 17289 8941 17323
rect 9689 17289 9723 17323
rect 11161 17289 11195 17323
rect 11483 17289 11517 17323
rect 14427 17289 14461 17323
rect 16497 17289 16531 17323
rect 17877 17289 17911 17323
rect 21097 17289 21131 17323
rect 13369 17221 13403 17255
rect 17141 17221 17175 17255
rect 7113 17153 7147 17187
rect 8585 17153 8619 17187
rect 15577 17153 15611 17187
rect 18245 17153 18279 17187
rect 18889 17153 18923 17187
rect 19257 17153 19291 17187
rect 4077 17085 4111 17119
rect 8836 17085 8870 17119
rect 11380 17085 11414 17119
rect 11805 17085 11839 17119
rect 14356 17085 14390 17119
rect 14749 17085 14783 17119
rect 20913 17085 20947 17119
rect 21465 17085 21499 17119
rect 2513 17017 2547 17051
rect 4398 17017 4432 17051
rect 7205 17017 7239 17051
rect 7757 17017 7791 17051
rect 9873 17017 9907 17051
rect 9965 17017 9999 17051
rect 10517 17017 10551 17051
rect 12817 17017 12851 17051
rect 12909 17017 12943 17051
rect 13829 17017 13863 17051
rect 15669 17017 15703 17051
rect 16221 17017 16255 17051
rect 18981 17017 19015 17051
rect 2789 16949 2823 16983
rect 3617 16949 3651 16983
rect 3893 16949 3927 16983
rect 5273 16949 5307 16983
rect 6469 16949 6503 16983
rect 9321 16949 9355 16983
rect 10793 16949 10827 16983
rect 12265 16949 12299 16983
rect 14105 16949 14139 16983
rect 15301 16949 15335 16983
rect 18705 16949 18739 16983
rect 20729 16949 20763 16983
rect 7113 16745 7147 16779
rect 12725 16745 12759 16779
rect 13277 16745 13311 16779
rect 15117 16745 15151 16779
rect 4813 16677 4847 16711
rect 7619 16677 7653 16711
rect 10149 16677 10183 16711
rect 10701 16677 10735 16711
rect 15853 16677 15887 16711
rect 18337 16677 18371 16711
rect 4261 16609 4295 16643
rect 4629 16609 4663 16643
rect 7532 16609 7566 16643
rect 8620 16609 8654 16643
rect 14140 16609 14174 16643
rect 6377 16541 6411 16575
rect 8723 16541 8757 16575
rect 10057 16541 10091 16575
rect 12357 16541 12391 16575
rect 15761 16541 15795 16575
rect 18245 16541 18279 16575
rect 16313 16473 16347 16507
rect 18797 16473 18831 16507
rect 19165 16473 19199 16507
rect 5089 16405 5123 16439
rect 6607 16405 6641 16439
rect 9045 16405 9079 16439
rect 9505 16405 9539 16439
rect 10977 16405 11011 16439
rect 11805 16405 11839 16439
rect 14243 16405 14277 16439
rect 15577 16405 15611 16439
rect 6193 16201 6227 16235
rect 6561 16201 6595 16235
rect 9505 16201 9539 16235
rect 10057 16201 10091 16235
rect 14105 16201 14139 16235
rect 16497 16201 16531 16235
rect 19441 16201 19475 16235
rect 4261 16133 4295 16167
rect 6653 16133 6687 16167
rect 10977 16133 11011 16167
rect 18705 16133 18739 16167
rect 3479 16065 3513 16099
rect 4445 16065 4479 16099
rect 4721 16065 4755 16099
rect 6929 16065 6963 16099
rect 7205 16065 7239 16099
rect 8585 16065 8619 16099
rect 11805 16065 11839 16099
rect 12081 16065 12115 16099
rect 14657 16065 14691 16099
rect 17095 16065 17129 16099
rect 18153 16065 18187 16099
rect 19073 16065 19107 16099
rect 3392 15997 3426 16031
rect 6653 15997 6687 16031
rect 3249 15929 3283 15963
rect 4537 15929 4571 15963
rect 7021 15929 7055 15963
rect 8906 15929 8940 15963
rect 10425 15929 10459 15963
rect 10517 15929 10551 15963
rect 11529 15929 11563 15963
rect 12449 15997 12483 16031
rect 13001 15997 13035 16031
rect 14841 15997 14875 16031
rect 17008 15997 17042 16031
rect 15162 15929 15196 15963
rect 17877 15929 17911 15963
rect 18245 15929 18279 15963
rect 3801 15861 3835 15895
rect 5365 15861 5399 15895
rect 7941 15861 7975 15895
rect 8401 15861 8435 15895
rect 12081 15861 12115 15895
rect 12173 15861 12207 15895
rect 12541 15861 12575 15895
rect 15761 15861 15795 15895
rect 16037 15861 16071 15895
rect 17509 15861 17543 15895
rect 19993 15861 20027 15895
rect 4997 15657 5031 15691
rect 6745 15657 6779 15691
rect 7021 15657 7055 15691
rect 8953 15657 8987 15691
rect 10057 15657 10091 15691
rect 12449 15657 12483 15691
rect 18245 15657 18279 15691
rect 18521 15657 18555 15691
rect 4398 15589 4432 15623
rect 6146 15589 6180 15623
rect 8677 15589 8711 15623
rect 10333 15589 10367 15623
rect 14381 15589 14415 15623
rect 14841 15589 14875 15623
rect 15485 15589 15519 15623
rect 16037 15589 16071 15623
rect 17646 15589 17680 15623
rect 18889 15589 18923 15623
rect 19257 15589 19291 15623
rect 2697 15521 2731 15555
rect 2881 15521 2915 15555
rect 7941 15521 7975 15555
rect 8401 15521 8435 15555
rect 13829 15521 13863 15555
rect 14105 15521 14139 15555
rect 19108 15521 19142 15555
rect 3157 15453 3191 15487
rect 4077 15453 4111 15487
rect 5825 15453 5859 15487
rect 10241 15453 10275 15487
rect 10609 15453 10643 15487
rect 15393 15453 15427 15487
rect 17325 15453 17359 15487
rect 13001 15385 13035 15419
rect 7389 15317 7423 15351
rect 11161 15317 11195 15351
rect 16405 15317 16439 15351
rect 2789 15113 2823 15147
rect 3157 15113 3191 15147
rect 5825 15113 5859 15147
rect 6653 15113 6687 15147
rect 8999 15113 9033 15147
rect 9781 15113 9815 15147
rect 10011 15113 10045 15147
rect 10701 15113 10735 15147
rect 15393 15113 15427 15147
rect 18705 15113 18739 15147
rect 20453 15113 20487 15147
rect 2513 15045 2547 15079
rect 4997 15045 5031 15079
rect 7481 15045 7515 15079
rect 11023 15045 11057 15079
rect 11437 15045 11471 15079
rect 15669 15045 15703 15079
rect 3479 14977 3513 15011
rect 4445 14977 4479 15011
rect 5365 14977 5399 15011
rect 6929 14977 6963 15011
rect 14565 14977 14599 15011
rect 16221 14977 16255 15011
rect 17141 14977 17175 15011
rect 17785 14977 17819 15011
rect 20729 14977 20763 15011
rect 21373 14977 21407 15011
rect 3376 14909 3410 14943
rect 3801 14909 3835 14943
rect 8896 14909 8930 14943
rect 9321 14909 9355 14943
rect 9940 14909 9974 14943
rect 10425 14909 10459 14943
rect 10952 14909 10986 14943
rect 16405 14909 16439 14943
rect 16865 14909 16899 14943
rect 18889 14909 18923 14943
rect 4537 14841 4571 14875
rect 7021 14841 7055 14875
rect 11897 14841 11931 14875
rect 12541 14841 12575 14875
rect 12633 14841 12667 14875
rect 13185 14841 13219 14875
rect 13737 14841 13771 14875
rect 14289 14841 14323 14875
rect 14381 14841 14415 14875
rect 19210 14841 19244 14875
rect 20821 14841 20855 14875
rect 4169 14773 4203 14807
rect 6193 14773 6227 14807
rect 8033 14773 8067 14807
rect 8309 14773 8343 14807
rect 12173 14773 12207 14807
rect 14013 14773 14047 14807
rect 17417 14773 17451 14807
rect 18337 14773 18371 14807
rect 19809 14773 19843 14807
rect 1593 14569 1627 14603
rect 4537 14569 4571 14603
rect 6975 14569 7009 14603
rect 10057 14569 10091 14603
rect 10609 14569 10643 14603
rect 10885 14569 10919 14603
rect 20637 14569 20671 14603
rect 21097 14569 21131 14603
rect 6009 14501 6043 14535
rect 11758 14501 11792 14535
rect 17877 14501 17911 14535
rect 1409 14433 1443 14467
rect 4144 14433 4178 14467
rect 5273 14433 5307 14467
rect 5733 14433 5767 14467
rect 6904 14433 6938 14467
rect 7884 14433 7918 14467
rect 13369 14433 13403 14467
rect 13645 14433 13679 14467
rect 15577 14433 15611 14467
rect 16037 14433 16071 14467
rect 17141 14433 17175 14467
rect 17601 14433 17635 14467
rect 18981 14433 19015 14467
rect 19165 14433 19199 14467
rect 20913 14433 20947 14467
rect 9689 14365 9723 14399
rect 11437 14365 11471 14399
rect 13737 14365 13771 14399
rect 16129 14365 16163 14399
rect 19257 14365 19291 14399
rect 4215 14229 4249 14263
rect 7481 14229 7515 14263
rect 7987 14229 8021 14263
rect 12357 14229 12391 14263
rect 14289 14229 14323 14263
rect 14565 14229 14599 14263
rect 20177 14229 20211 14263
rect 1593 14025 1627 14059
rect 4077 14025 4111 14059
rect 8401 14025 8435 14059
rect 12771 14025 12805 14059
rect 19073 14025 19107 14059
rect 4813 13957 4847 13991
rect 8033 13957 8067 13991
rect 13369 13957 13403 13991
rect 13461 13957 13495 13991
rect 14565 13957 14599 13991
rect 19441 13957 19475 13991
rect 3341 13889 3375 13923
rect 4261 13889 4295 13923
rect 7481 13889 7515 13923
rect 8861 13889 8895 13923
rect 1409 13821 1443 13855
rect 5733 13821 5767 13855
rect 9229 13821 9263 13855
rect 9505 13821 9539 13855
rect 10057 13821 10091 13855
rect 10517 13821 10551 13855
rect 10793 13821 10827 13855
rect 11069 13821 11103 13855
rect 11621 13821 11655 13855
rect 12668 13821 12702 13855
rect 13093 13821 13127 13855
rect 13645 13889 13679 13923
rect 15761 13889 15795 13923
rect 21097 13889 21131 13923
rect 17024 13821 17058 13855
rect 17417 13821 17451 13855
rect 18061 13821 18095 13855
rect 18613 13821 18647 13855
rect 20821 13821 20855 13855
rect 3709 13753 3743 13787
rect 4353 13753 4387 13787
rect 5365 13753 5399 13787
rect 7573 13753 7607 13787
rect 9689 13753 9723 13787
rect 13369 13753 13403 13787
rect 13966 13753 14000 13787
rect 15485 13753 15519 13787
rect 15577 13753 15611 13787
rect 17785 13753 17819 13787
rect 18797 13753 18831 13787
rect 20177 13753 20211 13787
rect 20269 13753 20303 13787
rect 2053 13685 2087 13719
rect 7021 13685 7055 13719
rect 10885 13685 10919 13719
rect 11989 13685 12023 13719
rect 14933 13685 14967 13719
rect 15301 13685 15335 13719
rect 16405 13685 16439 13719
rect 16773 13685 16807 13719
rect 17095 13685 17129 13719
rect 19993 13685 20027 13719
rect 6837 13481 6871 13515
rect 7665 13481 7699 13515
rect 9045 13481 9079 13515
rect 9873 13481 9907 13515
rect 11069 13481 11103 13515
rect 11621 13481 11655 13515
rect 12173 13481 12207 13515
rect 14381 13481 14415 13515
rect 15577 13481 15611 13515
rect 15945 13481 15979 13515
rect 17325 13481 17359 13515
rect 18153 13481 18187 13515
rect 19993 13481 20027 13515
rect 4439 13413 4473 13447
rect 13185 13413 13219 13447
rect 16450 13413 16484 13447
rect 19394 13413 19428 13447
rect 21097 13413 21131 13447
rect 2697 13345 2731 13379
rect 2881 13345 2915 13379
rect 7389 13345 7423 13379
rect 8284 13345 8318 13379
rect 10149 13345 10183 13379
rect 11253 13345 11287 13379
rect 16129 13345 16163 13379
rect 3157 13277 3191 13311
rect 4077 13277 4111 13311
rect 6469 13277 6503 13311
rect 13093 13277 13127 13311
rect 13369 13277 13403 13311
rect 19073 13277 19107 13311
rect 21005 13277 21039 13311
rect 21281 13277 21315 13311
rect 5273 13209 5307 13243
rect 10379 13209 10413 13243
rect 1685 13141 1719 13175
rect 4997 13141 5031 13175
rect 8125 13141 8159 13175
rect 8355 13141 8389 13175
rect 10793 13141 10827 13175
rect 12449 13141 12483 13175
rect 14013 13141 14047 13175
rect 17049 13141 17083 13175
rect 2789 12937 2823 12971
rect 3249 12937 3283 12971
rect 5457 12937 5491 12971
rect 7297 12937 7331 12971
rect 13461 12937 13495 12971
rect 13645 12937 13679 12971
rect 15853 12937 15887 12971
rect 18889 12937 18923 12971
rect 19993 12937 20027 12971
rect 20821 12937 20855 12971
rect 21097 12937 21131 12971
rect 13093 12869 13127 12903
rect 14657 12869 14691 12903
rect 20269 12869 20303 12903
rect 3571 12801 3605 12835
rect 4537 12801 4571 12835
rect 7481 12801 7515 12835
rect 9321 12801 9355 12835
rect 13645 12801 13679 12835
rect 14105 12801 14139 12835
rect 15025 12801 15059 12835
rect 16497 12801 16531 12835
rect 17417 12801 17451 12835
rect 19073 12801 19107 12835
rect 3484 12733 3518 12767
rect 10977 12733 11011 12767
rect 11253 12733 11287 12767
rect 11437 12733 11471 12767
rect 16129 12733 16163 12767
rect 18096 12733 18130 12767
rect 18521 12733 18555 12767
rect 20913 12733 20947 12767
rect 21465 12733 21499 12767
rect 4629 12665 4663 12699
rect 5181 12665 5215 12699
rect 7573 12665 7607 12699
rect 8125 12665 8159 12699
rect 9045 12665 9079 12699
rect 9137 12665 9171 12699
rect 12541 12665 12575 12699
rect 12633 12665 12667 12699
rect 14197 12665 14231 12699
rect 16589 12665 16623 12699
rect 17141 12665 17175 12699
rect 19394 12665 19428 12699
rect 2513 12597 2547 12631
rect 3985 12597 4019 12631
rect 4353 12597 4387 12631
rect 6193 12597 6227 12631
rect 6561 12597 6595 12631
rect 8493 12597 8527 12631
rect 8769 12597 8803 12631
rect 10333 12597 10367 12631
rect 11713 12597 11747 12631
rect 12265 12597 12299 12631
rect 13921 12597 13955 12631
rect 18199 12597 18233 12631
rect 6193 12393 6227 12427
rect 9045 12393 9079 12427
rect 9827 12393 9861 12427
rect 11069 12393 11103 12427
rect 15439 12393 15473 12427
rect 19809 12393 19843 12427
rect 21097 12393 21131 12427
rect 4537 12325 4571 12359
rect 8217 12325 8251 12359
rect 11805 12325 11839 12359
rect 12357 12325 12391 12359
rect 13001 12325 13035 12359
rect 13829 12325 13863 12359
rect 16405 12325 16439 12359
rect 17233 12325 17267 12359
rect 17785 12325 17819 12359
rect 2513 12257 2547 12291
rect 2881 12257 2915 12291
rect 5917 12257 5951 12291
rect 6469 12257 6503 12291
rect 9756 12257 9790 12291
rect 15336 12257 15370 12291
rect 19073 12257 19107 12291
rect 19257 12257 19291 12291
rect 3157 12189 3191 12223
rect 4445 12189 4479 12223
rect 4721 12189 4755 12223
rect 8125 12189 8159 12223
rect 8401 12189 8435 12223
rect 11713 12189 11747 12223
rect 13737 12189 13771 12223
rect 14381 12189 14415 12223
rect 17141 12189 17175 12223
rect 5457 12121 5491 12155
rect 7757 12053 7791 12087
rect 10701 12053 10735 12087
rect 11345 12053 11379 12087
rect 13461 12053 13495 12087
rect 16773 12053 16807 12087
rect 19487 12053 19521 12087
rect 4077 11849 4111 11883
rect 4445 11849 4479 11883
rect 6285 11849 6319 11883
rect 8585 11849 8619 11883
rect 8861 11849 8895 11883
rect 10333 11849 10367 11883
rect 11529 11849 11563 11883
rect 11805 11849 11839 11883
rect 17417 11849 17451 11883
rect 17877 11849 17911 11883
rect 21649 11849 21683 11883
rect 17049 11781 17083 11815
rect 21281 11781 21315 11815
rect 3157 11713 3191 11747
rect 5273 11713 5307 11747
rect 12587 11713 12621 11747
rect 15531 11713 15565 11747
rect 16497 11713 16531 11747
rect 20269 11713 20303 11747
rect 2145 11645 2179 11679
rect 7665 11645 7699 11679
rect 9480 11645 9514 11679
rect 10609 11645 10643 11679
rect 12500 11645 12534 11679
rect 12909 11645 12943 11679
rect 13461 11645 13495 11679
rect 15428 11645 15462 11679
rect 15853 11645 15887 11679
rect 18128 11645 18162 11679
rect 21097 11645 21131 11679
rect 3478 11577 3512 11611
rect 4997 11577 5031 11611
rect 5089 11577 5123 11611
rect 6009 11577 6043 11611
rect 8027 11577 8061 11611
rect 10930 11577 10964 11611
rect 13277 11577 13311 11611
rect 13782 11577 13816 11611
rect 16313 11577 16347 11611
rect 16589 11577 16623 11611
rect 19073 11577 19107 11611
rect 19625 11577 19659 11611
rect 19717 11577 19751 11611
rect 2513 11509 2547 11543
rect 2973 11509 3007 11543
rect 4813 11509 4847 11543
rect 7481 11509 7515 11543
rect 9551 11509 9585 11543
rect 9965 11509 9999 11543
rect 12173 11509 12207 11543
rect 14381 11509 14415 11543
rect 15209 11509 15243 11543
rect 18199 11509 18233 11543
rect 18613 11509 18647 11543
rect 19349 11509 19383 11543
rect 3157 11305 3191 11339
rect 3893 11305 3927 11339
rect 4997 11305 5031 11339
rect 5365 11305 5399 11339
rect 8125 11305 8159 11339
rect 13829 11305 13863 11339
rect 17049 11305 17083 11339
rect 18061 11305 18095 11339
rect 19073 11305 19107 11339
rect 19901 11305 19935 11339
rect 21051 11305 21085 11339
rect 4439 11237 4473 11271
rect 7757 11237 7791 11271
rect 11161 11237 11195 11271
rect 12633 11237 12667 11271
rect 13461 11237 13495 11271
rect 14105 11237 14139 11271
rect 16450 11237 16484 11271
rect 1476 11169 1510 11203
rect 5892 11169 5926 11203
rect 7113 11169 7147 11203
rect 7573 11169 7607 11203
rect 8652 11169 8686 11203
rect 10701 11169 10735 11203
rect 10977 11169 11011 11203
rect 13001 11169 13035 11203
rect 13185 11169 13219 11203
rect 19625 11169 19659 11203
rect 20948 11169 20982 11203
rect 2421 11101 2455 11135
rect 4077 11101 4111 11135
rect 16129 11101 16163 11135
rect 18705 11101 18739 11135
rect 10241 11033 10275 11067
rect 1547 10965 1581 10999
rect 1961 10965 1995 10999
rect 5963 10965 5997 10999
rect 6929 10965 6963 10999
rect 8723 10965 8757 10999
rect 9873 10965 9907 10999
rect 6285 10761 6319 10795
rect 6653 10761 6687 10795
rect 8953 10761 8987 10795
rect 9321 10761 9355 10795
rect 11069 10761 11103 10795
rect 11391 10761 11425 10795
rect 14381 10761 14415 10795
rect 16589 10761 16623 10795
rect 17785 10761 17819 10795
rect 19073 10761 19107 10795
rect 19533 10761 19567 10795
rect 2513 10693 2547 10727
rect 7941 10693 7975 10727
rect 10701 10693 10735 10727
rect 13093 10693 13127 10727
rect 14013 10693 14047 10727
rect 1777 10625 1811 10659
rect 1961 10625 1995 10659
rect 3525 10625 3559 10659
rect 4261 10625 4295 10659
rect 6929 10625 6963 10659
rect 8217 10625 8251 10659
rect 16313 10625 16347 10659
rect 16957 10625 16991 10659
rect 18153 10625 18187 10659
rect 18613 10625 18647 10659
rect 19717 10625 19751 10659
rect 20177 10625 20211 10659
rect 3709 10557 3743 10591
rect 4169 10557 4203 10591
rect 5457 10557 5491 10591
rect 5733 10557 5767 10591
rect 8468 10557 8502 10591
rect 11320 10557 11354 10591
rect 12909 10557 12943 10591
rect 13001 10557 13035 10591
rect 13277 10557 13311 10591
rect 14600 10557 14634 10591
rect 15025 10557 15059 10591
rect 15577 10557 15611 10591
rect 16037 10557 16071 10591
rect 2053 10489 2087 10523
rect 4997 10489 5031 10523
rect 7021 10489 7055 10523
rect 7573 10489 7607 10523
rect 9689 10489 9723 10523
rect 9781 10489 9815 10523
rect 10333 10489 10367 10523
rect 12265 10489 12299 10523
rect 18245 10489 18279 10523
rect 19809 10489 19843 10523
rect 4721 10421 4755 10455
rect 5273 10421 5307 10455
rect 8539 10421 8573 10455
rect 11713 10421 11747 10455
rect 13461 10421 13495 10455
rect 14703 10421 14737 10455
rect 15393 10421 15427 10455
rect 20913 10421 20947 10455
rect 1685 10217 1719 10251
rect 2789 10217 2823 10251
rect 3709 10217 3743 10251
rect 4261 10217 4295 10251
rect 5917 10217 5951 10251
rect 12449 10217 12483 10251
rect 13553 10217 13587 10251
rect 14105 10217 14139 10251
rect 15945 10217 15979 10251
rect 19717 10217 19751 10251
rect 2231 10149 2265 10183
rect 5359 10149 5393 10183
rect 6929 10149 6963 10183
rect 9873 10149 9907 10183
rect 18429 10149 18463 10183
rect 18705 10149 18739 10183
rect 4997 10081 5031 10115
rect 8636 10081 8670 10115
rect 11989 10081 12023 10115
rect 12265 10081 12299 10115
rect 13645 10081 13679 10115
rect 13921 10081 13955 10115
rect 16405 10081 16439 10115
rect 16589 10081 16623 10115
rect 17969 10081 18003 10115
rect 18153 10081 18187 10115
rect 19324 10081 19358 10115
rect 20913 10081 20947 10115
rect 1869 10013 1903 10047
rect 6837 10013 6871 10047
rect 8723 10013 8757 10047
rect 9781 10013 9815 10047
rect 10425 10013 10459 10047
rect 11897 10013 11931 10047
rect 14657 10013 14691 10047
rect 16865 10013 16899 10047
rect 7389 9945 7423 9979
rect 12081 9945 12115 9979
rect 13737 9945 13771 9979
rect 21097 9945 21131 9979
rect 4629 9877 4663 9911
rect 13093 9877 13127 9911
rect 15577 9877 15611 9911
rect 19073 9877 19107 9911
rect 19395 9877 19429 9911
rect 6285 9673 6319 9707
rect 8401 9673 8435 9707
rect 9413 9673 9447 9707
rect 9781 9673 9815 9707
rect 10057 9673 10091 9707
rect 11391 9673 11425 9707
rect 17693 9673 17727 9707
rect 12081 9605 12115 9639
rect 16681 9605 16715 9639
rect 2881 9537 2915 9571
rect 3525 9537 3559 9571
rect 6653 9537 6687 9571
rect 12541 9537 12575 9571
rect 13645 9537 13679 9571
rect 14105 9537 14139 9571
rect 14749 9537 14783 9571
rect 16129 9537 16163 9571
rect 18797 9537 18831 9571
rect 2145 9469 2179 9503
rect 2697 9469 2731 9503
rect 4629 9469 4663 9503
rect 5181 9469 5215 9503
rect 6929 9469 6963 9503
rect 7481 9469 7515 9503
rect 8493 9469 8527 9503
rect 10308 9469 10342 9503
rect 11161 9469 11195 9503
rect 11288 9469 11322 9503
rect 12449 9469 12483 9503
rect 12725 9469 12759 9503
rect 14013 9469 14047 9503
rect 14289 9469 14323 9503
rect 15025 9469 15059 9503
rect 3157 9401 3191 9435
rect 4537 9401 4571 9435
rect 5365 9401 5399 9435
rect 7665 9401 7699 9435
rect 7941 9401 7975 9435
rect 8814 9401 8848 9435
rect 10793 9401 10827 9435
rect 15393 9401 15427 9435
rect 16221 9401 16255 9435
rect 18889 9401 18923 9435
rect 19441 9401 19475 9435
rect 19809 9401 19843 9435
rect 1961 9333 1995 9367
rect 5733 9333 5767 9367
rect 10379 9333 10413 9367
rect 12909 9333 12943 9367
rect 15853 9333 15887 9367
rect 17049 9333 17083 9367
rect 18245 9333 18279 9367
rect 20913 9333 20947 9367
rect 2237 9129 2271 9163
rect 2421 9129 2455 9163
rect 4997 9129 5031 9163
rect 5733 9129 5767 9163
rect 6285 9129 6319 9163
rect 8585 9129 8619 9163
rect 12909 9129 12943 9163
rect 16313 9129 16347 9163
rect 16589 9129 16623 9163
rect 18337 9129 18371 9163
rect 18889 9129 18923 9163
rect 19257 9129 19291 9163
rect 6653 9061 6687 9095
rect 6929 9061 6963 9095
rect 7205 9061 7239 9095
rect 7297 9061 7331 9095
rect 9873 9061 9907 9095
rect 10425 9061 10459 9095
rect 13461 9061 13495 9095
rect 15755 9061 15789 9095
rect 2329 8993 2363 9027
rect 2881 8993 2915 9027
rect 4353 8993 4387 9027
rect 11897 8993 11931 9027
rect 12173 8993 12207 9027
rect 13553 8993 13587 9027
rect 17969 8993 18003 9027
rect 19752 8993 19786 9027
rect 5365 8925 5399 8959
rect 7481 8925 7515 8959
rect 9781 8925 9815 8959
rect 12357 8925 12391 8959
rect 14473 8925 14507 8959
rect 15393 8925 15427 8959
rect 4491 8857 4525 8891
rect 11989 8857 12023 8891
rect 11805 8789 11839 8823
rect 13277 8789 13311 8823
rect 19625 8789 19659 8823
rect 19855 8789 19889 8823
rect 2237 8585 2271 8619
rect 5917 8585 5951 8619
rect 6653 8585 6687 8619
rect 11529 8585 11563 8619
rect 11897 8585 11931 8619
rect 12173 8585 12207 8619
rect 15853 8585 15887 8619
rect 16221 8585 16255 8619
rect 17785 8585 17819 8619
rect 18245 8585 18279 8619
rect 19717 8585 19751 8619
rect 2973 8517 3007 8551
rect 8217 8517 8251 8551
rect 10701 8517 10735 8551
rect 2421 8449 2455 8483
rect 3341 8449 3375 8483
rect 4261 8449 4295 8483
rect 10149 8449 10183 8483
rect 11069 8449 11103 8483
rect 13185 8449 13219 8483
rect 16405 8449 16439 8483
rect 18797 8449 18831 8483
rect 19073 8449 19107 8483
rect 4353 8381 4387 8415
rect 5641 8381 5675 8415
rect 6904 8381 6938 8415
rect 7849 8381 7883 8415
rect 8309 8381 8343 8415
rect 9229 8381 9263 8415
rect 12541 8381 12575 8415
rect 14933 8381 14967 8415
rect 15301 8381 15335 8415
rect 2513 8313 2547 8347
rect 4715 8313 4749 8347
rect 7389 8313 7423 8347
rect 9781 8313 9815 8347
rect 10241 8313 10275 8347
rect 14657 8313 14691 8347
rect 15485 8313 15519 8347
rect 16497 8313 16531 8347
rect 17049 8313 17083 8347
rect 18889 8313 18923 8347
rect 1869 8245 1903 8279
rect 3801 8245 3835 8279
rect 5273 8245 5307 8279
rect 6975 8245 7009 8279
rect 8677 8245 8711 8279
rect 13553 8245 13587 8279
rect 1961 8041 1995 8075
rect 2973 8041 3007 8075
rect 4353 8041 4387 8075
rect 5089 8041 5123 8075
rect 7113 8041 7147 8075
rect 7849 8041 7883 8075
rect 9505 8041 9539 8075
rect 10425 8041 10459 8075
rect 12357 8041 12391 8075
rect 13185 8041 13219 8075
rect 15485 8041 15519 8075
rect 18797 8041 18831 8075
rect 2415 7973 2449 8007
rect 6009 7973 6043 8007
rect 6561 7973 6595 8007
rect 15853 7973 15887 8007
rect 16405 7973 16439 8007
rect 19165 7973 19199 8007
rect 4077 7905 4111 7939
rect 4537 7905 4571 7939
rect 7757 7905 7791 7939
rect 8125 7905 8159 7939
rect 9965 7905 9999 7939
rect 11136 7905 11170 7939
rect 12541 7905 12575 7939
rect 14105 7905 14139 7939
rect 17693 7905 17727 7939
rect 17877 7905 17911 7939
rect 2053 7837 2087 7871
rect 5917 7837 5951 7871
rect 12909 7837 12943 7871
rect 14335 7837 14369 7871
rect 15761 7837 15795 7871
rect 18153 7837 18187 7871
rect 19073 7837 19107 7871
rect 12706 7769 12740 7803
rect 13921 7769 13955 7803
rect 19625 7769 19659 7803
rect 5457 7701 5491 7735
rect 8585 7701 8619 7735
rect 10103 7701 10137 7735
rect 10885 7701 10919 7735
rect 11207 7701 11241 7735
rect 11989 7701 12023 7735
rect 12817 7701 12851 7735
rect 13553 7701 13587 7735
rect 14841 7701 14875 7735
rect 16773 7701 16807 7735
rect 2881 7497 2915 7531
rect 4537 7497 4571 7531
rect 5917 7497 5951 7531
rect 6285 7497 6319 7531
rect 8033 7497 8067 7531
rect 8401 7497 8435 7531
rect 11713 7497 11747 7531
rect 12725 7497 12759 7531
rect 13093 7497 13127 7531
rect 13553 7497 13587 7531
rect 15577 7497 15611 7531
rect 17785 7497 17819 7531
rect 18981 7497 19015 7531
rect 7389 7429 7423 7463
rect 16681 7429 16715 7463
rect 19717 7429 19751 7463
rect 2053 7361 2087 7395
rect 4813 7361 4847 7395
rect 9965 7361 9999 7395
rect 10793 7361 10827 7395
rect 11069 7361 11103 7395
rect 13424 7361 13458 7395
rect 13645 7361 13679 7395
rect 15163 7361 15197 7395
rect 16129 7361 16163 7395
rect 17049 7361 17083 7395
rect 19165 7361 19199 7395
rect 20085 7361 20119 7395
rect 3776 7293 3810 7327
rect 4169 7293 4203 7327
rect 7532 7293 7566 7327
rect 8493 7293 8527 7327
rect 12265 7293 12299 7327
rect 13277 7293 13311 7327
rect 15076 7293 15110 7327
rect 4905 7225 4939 7259
rect 5457 7225 5491 7259
rect 7619 7225 7653 7259
rect 8814 7225 8848 7259
rect 10517 7225 10551 7259
rect 10885 7225 10919 7259
rect 14013 7225 14047 7259
rect 14933 7225 14967 7259
rect 15853 7225 15887 7259
rect 16221 7225 16255 7259
rect 19257 7225 19291 7259
rect 2605 7157 2639 7191
rect 3617 7157 3651 7191
rect 3847 7157 3881 7191
rect 9413 7157 9447 7191
rect 14289 7157 14323 7191
rect 17509 7157 17543 7191
rect 18613 7157 18647 7191
rect 20821 7157 20855 7191
rect 3111 6953 3145 6987
rect 6929 6953 6963 6987
rect 7665 6953 7699 6987
rect 16221 6953 16255 6987
rect 16497 6953 16531 6987
rect 17187 6953 17221 6987
rect 19257 6953 19291 6987
rect 19533 6953 19567 6987
rect 21051 6953 21085 6987
rect 4721 6885 4755 6919
rect 5089 6885 5123 6919
rect 8493 6885 8527 6919
rect 10333 6885 10367 6919
rect 10425 6885 10459 6919
rect 15622 6885 15656 6919
rect 18658 6885 18692 6919
rect 1476 6817 1510 6851
rect 3040 6817 3074 6851
rect 6469 6817 6503 6851
rect 7757 6817 7791 6851
rect 8217 6817 8251 6851
rect 11872 6817 11906 6851
rect 13921 6817 13955 6851
rect 14197 6817 14231 6851
rect 17116 6817 17150 6851
rect 20980 6817 21014 6851
rect 4997 6749 5031 6783
rect 5641 6749 5675 6783
rect 10609 6749 10643 6783
rect 14381 6749 14415 6783
rect 15301 6749 15335 6783
rect 18337 6749 18371 6783
rect 13277 6681 13311 6715
rect 1547 6613 1581 6647
rect 2881 6613 2915 6647
rect 6607 6613 6641 6647
rect 10149 6613 10183 6647
rect 11943 6613 11977 6647
rect 12633 6613 12667 6647
rect 12909 6613 12943 6647
rect 14749 6613 14783 6647
rect 1685 6409 1719 6443
rect 2697 6409 2731 6443
rect 3709 6409 3743 6443
rect 5733 6409 5767 6443
rect 8401 6409 8435 6443
rect 9689 6409 9723 6443
rect 11529 6409 11563 6443
rect 12817 6409 12851 6443
rect 13737 6409 13771 6443
rect 15393 6409 15427 6443
rect 16589 6409 16623 6443
rect 17141 6409 17175 6443
rect 17877 6409 17911 6443
rect 18245 6409 18279 6443
rect 19349 6409 19383 6443
rect 21465 6409 21499 6443
rect 6469 6341 6503 6375
rect 11897 6341 11931 6375
rect 12706 6341 12740 6375
rect 6929 6273 6963 6307
rect 7205 6273 7239 6307
rect 10333 6273 10367 6307
rect 10977 6273 11011 6307
rect 12909 6273 12943 6307
rect 14565 6273 14599 6307
rect 16129 6273 16163 6307
rect 18429 6273 18463 6307
rect 2789 6205 2823 6239
rect 4077 6205 4111 6239
rect 4537 6205 4571 6239
rect 5457 6205 5491 6239
rect 8493 6205 8527 6239
rect 9413 6205 9447 6239
rect 10057 6205 10091 6239
rect 12541 6205 12575 6239
rect 14105 6205 14139 6239
rect 14289 6205 14323 6239
rect 15853 6205 15887 6239
rect 16037 6205 16071 6239
rect 20545 6205 20579 6239
rect 7021 6137 7055 6171
rect 8814 6137 8848 6171
rect 10425 6137 10459 6171
rect 12173 6137 12207 6171
rect 13277 6137 13311 6171
rect 17509 6137 17543 6171
rect 18750 6137 18784 6171
rect 21189 6137 21223 6171
rect 3157 6069 3191 6103
rect 4445 6069 4479 6103
rect 4905 6069 4939 6103
rect 7941 6069 7975 6103
rect 14933 6069 14967 6103
rect 20361 6069 20395 6103
rect 4353 5865 4387 5899
rect 5089 5865 5123 5899
rect 7573 5865 7607 5899
rect 10885 5865 10919 5899
rect 12081 5865 12115 5899
rect 15669 5865 15703 5899
rect 15945 5865 15979 5899
rect 18889 5865 18923 5899
rect 5917 5797 5951 5831
rect 6009 5797 6043 5831
rect 6837 5797 6871 5831
rect 8493 5797 8527 5831
rect 8769 5797 8803 5831
rect 10057 5797 10091 5831
rect 10609 5797 10643 5831
rect 12725 5797 12759 5831
rect 13277 5797 13311 5831
rect 16450 5797 16484 5831
rect 18061 5797 18095 5831
rect 21005 5797 21039 5831
rect 21097 5797 21131 5831
rect 4353 5729 4387 5763
rect 4629 5729 4663 5763
rect 4905 5729 4939 5763
rect 6561 5729 6595 5763
rect 7757 5729 7791 5763
rect 8309 5729 8343 5763
rect 11621 5729 11655 5763
rect 11897 5729 11931 5763
rect 13369 5729 13403 5763
rect 13645 5729 13679 5763
rect 16129 5729 16163 5763
rect 17049 5729 17083 5763
rect 9965 5661 9999 5695
rect 14013 5661 14047 5695
rect 17969 5661 18003 5695
rect 19441 5661 19475 5695
rect 21465 5661 21499 5695
rect 4905 5593 4939 5627
rect 11713 5593 11747 5627
rect 13461 5593 13495 5627
rect 18521 5593 18555 5627
rect 2881 5525 2915 5559
rect 7205 5525 7239 5559
rect 11529 5525 11563 5559
rect 14381 5525 14415 5559
rect 20545 5525 20579 5559
rect 4169 5321 4203 5355
rect 4537 5321 4571 5355
rect 5641 5321 5675 5355
rect 6285 5321 6319 5355
rect 9781 5321 9815 5355
rect 11345 5321 11379 5355
rect 12541 5321 12575 5355
rect 15485 5321 15519 5355
rect 17509 5321 17543 5355
rect 19073 5321 19107 5355
rect 20453 5321 20487 5355
rect 21557 5321 21591 5355
rect 1547 5253 1581 5287
rect 5871 5253 5905 5287
rect 14381 5253 14415 5287
rect 2973 5185 3007 5219
rect 6929 5185 6963 5219
rect 7389 5185 7423 5219
rect 10977 5185 11011 5219
rect 12265 5185 12299 5219
rect 14473 5185 14507 5219
rect 16773 5185 16807 5219
rect 17877 5185 17911 5219
rect 21281 5185 21315 5219
rect 1476 5117 1510 5151
rect 3341 5117 3375 5151
rect 3525 5117 3559 5151
rect 4772 5117 4806 5151
rect 5181 5117 5215 5151
rect 5800 5117 5834 5151
rect 8401 5117 8435 5151
rect 8861 5117 8895 5151
rect 12725 5117 12759 5151
rect 12909 5117 12943 5151
rect 13185 5117 13219 5151
rect 14565 5117 14599 5151
rect 16037 5117 16071 5151
rect 16129 5117 16163 5151
rect 16313 5117 16347 5151
rect 18061 5117 18095 5151
rect 18521 5117 18555 5151
rect 2605 5049 2639 5083
rect 4859 5049 4893 5083
rect 7021 5049 7055 5083
rect 9137 5049 9171 5083
rect 10333 5049 10367 5083
rect 10425 5049 10459 5083
rect 20637 5049 20671 5083
rect 20729 5049 20763 5083
rect 1961 4981 1995 5015
rect 3157 4981 3191 5015
rect 6653 4981 6687 5015
rect 7941 4981 7975 5015
rect 8309 4981 8343 5015
rect 10149 4981 10183 5015
rect 11621 4981 11655 5015
rect 14013 4981 14047 5015
rect 15853 4981 15887 5015
rect 17141 4981 17175 5015
rect 18153 4981 18187 5015
rect 3111 4777 3145 4811
rect 5917 4777 5951 4811
rect 6745 4777 6779 4811
rect 7941 4777 7975 4811
rect 8401 4777 8435 4811
rect 8723 4777 8757 4811
rect 10885 4777 10919 4811
rect 11253 4777 11287 4811
rect 12909 4777 12943 4811
rect 14565 4777 14599 4811
rect 15761 4777 15795 4811
rect 16681 4777 16715 4811
rect 18061 4777 18095 4811
rect 18613 4777 18647 4811
rect 19165 4777 19199 4811
rect 20545 4777 20579 4811
rect 5089 4709 5123 4743
rect 7113 4709 7147 4743
rect 9413 4709 9447 4743
rect 10010 4709 10044 4743
rect 11621 4709 11655 4743
rect 13001 4709 13035 4743
rect 2881 4641 2915 4675
rect 8620 4641 8654 4675
rect 9689 4641 9723 4675
rect 10609 4641 10643 4675
rect 13553 4641 13587 4675
rect 16221 4641 16255 4675
rect 16497 4641 16531 4675
rect 20948 4641 20982 4675
rect 4997 4573 5031 4607
rect 5641 4573 5675 4607
rect 7021 4573 7055 4607
rect 7297 4573 7331 4607
rect 11529 4573 11563 4607
rect 11805 4573 11839 4607
rect 18245 4573 18279 4607
rect 16313 4505 16347 4539
rect 20177 4505 20211 4539
rect 21051 4505 21085 4539
rect 3617 4437 3651 4471
rect 12449 4437 12483 4471
rect 14013 4437 14047 4471
rect 16129 4437 16163 4471
rect 4537 4233 4571 4267
rect 4905 4233 4939 4267
rect 5365 4233 5399 4267
rect 6285 4233 6319 4267
rect 7757 4233 7791 4267
rect 8401 4233 8435 4267
rect 10057 4233 10091 4267
rect 11713 4233 11747 4267
rect 21097 4233 21131 4267
rect 3157 4165 3191 4199
rect 8125 4165 8159 4199
rect 12633 4165 12667 4199
rect 18337 4165 18371 4199
rect 10793 4097 10827 4131
rect 12265 4097 12299 4131
rect 16957 4097 16991 4131
rect 20177 4097 20211 4131
rect 20453 4097 20487 4131
rect 2329 4029 2363 4063
rect 2605 4029 2639 4063
rect 2789 4029 2823 4063
rect 3617 4029 3651 4063
rect 5549 4029 5583 4063
rect 6837 4029 6871 4063
rect 8585 4029 8619 4063
rect 9137 4029 9171 4063
rect 12449 4029 12483 4063
rect 13553 4029 13587 4063
rect 14013 4029 14047 4063
rect 14381 4029 14415 4063
rect 14749 4029 14783 4063
rect 16313 4029 16347 4063
rect 17877 4029 17911 4063
rect 18613 4029 18647 4063
rect 1961 3961 1995 3995
rect 3938 3961 3972 3995
rect 5779 3961 5813 3995
rect 7158 3961 7192 3995
rect 9689 3961 9723 3995
rect 10609 3961 10643 3995
rect 10885 3961 10919 3995
rect 11437 3961 11471 3995
rect 15025 3961 15059 3995
rect 19257 3961 19291 3995
rect 19901 3961 19935 3995
rect 20269 3961 20303 3995
rect 3433 3893 3467 3927
rect 6561 3893 6595 3927
rect 8677 3893 8711 3927
rect 13001 3893 13035 3927
rect 13461 3893 13495 3927
rect 15393 3893 15427 3927
rect 15761 3893 15795 3927
rect 16037 3893 16071 3927
rect 17417 3893 17451 3927
rect 2145 3689 2179 3723
rect 3433 3689 3467 3723
rect 5457 3689 5491 3723
rect 7389 3689 7423 3723
rect 7941 3689 7975 3723
rect 8953 3689 8987 3723
rect 9965 3689 9999 3723
rect 10701 3689 10735 3723
rect 11161 3689 11195 3723
rect 12633 3689 12667 3723
rect 13093 3689 13127 3723
rect 16037 3689 16071 3723
rect 17693 3689 17727 3723
rect 19349 3689 19383 3723
rect 19809 3689 19843 3723
rect 4858 3621 4892 3655
rect 5733 3621 5767 3655
rect 6469 3621 6503 3655
rect 11529 3621 11563 3655
rect 18750 3621 18784 3655
rect 8125 3553 8159 3587
rect 8401 3553 8435 3587
rect 9689 3553 9723 3587
rect 10241 3553 10275 3587
rect 10517 3553 10551 3587
rect 13737 3553 13771 3587
rect 15577 3553 15611 3587
rect 15853 3553 15887 3587
rect 17141 3553 17175 3587
rect 18429 3553 18463 3587
rect 20948 3553 20982 3587
rect 4537 3485 4571 3519
rect 6377 3485 6411 3519
rect 6653 3485 6687 3519
rect 9505 3417 9539 3451
rect 11437 3485 11471 3519
rect 11713 3485 11747 3519
rect 13553 3485 13587 3519
rect 14381 3485 14415 3519
rect 15669 3417 15703 3451
rect 7757 3349 7791 3383
rect 10517 3349 10551 3383
rect 15117 3349 15151 3383
rect 16681 3349 16715 3383
rect 17325 3349 17359 3383
rect 18061 3349 18095 3383
rect 20269 3349 20303 3383
rect 21051 3349 21085 3383
rect 5917 3145 5951 3179
rect 6285 3145 6319 3179
rect 7941 3145 7975 3179
rect 9505 3145 9539 3179
rect 10885 3145 10919 3179
rect 11529 3145 11563 3179
rect 12265 3145 12299 3179
rect 19073 3145 19107 3179
rect 20913 3145 20947 3179
rect 9781 3077 9815 3111
rect 12633 3077 12667 3111
rect 15025 3077 15059 3111
rect 17049 3077 17083 3111
rect 17325 3077 17359 3111
rect 17877 3077 17911 3111
rect 3985 3009 4019 3043
rect 5641 3009 5675 3043
rect 8953 3009 8987 3043
rect 9965 3009 9999 3043
rect 11161 3009 11195 3043
rect 15945 3009 15979 3043
rect 19441 3009 19475 3043
rect 19901 3009 19935 3043
rect 20361 3009 20395 3043
rect 3617 2941 3651 2975
rect 3801 2941 3835 2975
rect 7113 2941 7147 2975
rect 12449 2941 12483 2975
rect 13093 2941 13127 2975
rect 13645 2941 13679 2975
rect 14105 2941 14139 2975
rect 14473 2941 14507 2975
rect 15025 2941 15059 2975
rect 16589 2941 16623 2975
rect 18061 2941 18095 2975
rect 18153 2941 18187 2975
rect 18337 2941 18371 2975
rect 3249 2873 3283 2907
rect 4997 2873 5031 2907
rect 5089 2873 5123 2907
rect 7205 2873 7239 2907
rect 8309 2873 8343 2907
rect 8401 2873 8435 2907
rect 10286 2873 10320 2907
rect 19993 2873 20027 2907
rect 4537 2805 4571 2839
rect 13461 2805 13495 2839
rect 15669 2805 15703 2839
rect 18521 2805 18555 2839
rect 2145 2601 2179 2635
rect 2237 2601 2271 2635
rect 5273 2601 5307 2635
rect 5825 2601 5859 2635
rect 6377 2601 6411 2635
rect 7481 2601 7515 2635
rect 8585 2601 8619 2635
rect 10241 2601 10275 2635
rect 10609 2601 10643 2635
rect 11713 2601 11747 2635
rect 12725 2601 12759 2635
rect 13645 2601 13679 2635
rect 14105 2601 14139 2635
rect 16405 2601 16439 2635
rect 19349 2601 19383 2635
rect 20545 2601 20579 2635
rect 1961 2533 1995 2567
rect 3709 2533 3743 2567
rect 4398 2533 4432 2567
rect 7986 2533 8020 2567
rect 8861 2533 8895 2567
rect 11114 2533 11148 2567
rect 12449 2533 12483 2567
rect 2145 2465 2179 2499
rect 2421 2465 2455 2499
rect 2973 2465 3007 2499
rect 3157 2397 3191 2431
rect 3433 2397 3467 2431
rect 4997 2465 5031 2499
rect 5641 2465 5675 2499
rect 7205 2465 7239 2499
rect 7665 2465 7699 2499
rect 9689 2465 9723 2499
rect 10793 2465 10827 2499
rect 12909 2465 12943 2499
rect 13185 2465 13219 2499
rect 14197 2465 14231 2499
rect 14749 2465 14783 2499
rect 15945 2465 15979 2499
rect 16221 2465 16255 2499
rect 17141 2465 17175 2499
rect 18153 2465 18187 2499
rect 18337 2465 18371 2499
rect 18613 2465 18647 2499
rect 19901 2465 19935 2499
rect 21189 2465 21223 2499
rect 21741 2465 21775 2499
rect 4077 2397 4111 2431
rect 9597 2397 9631 2431
rect 12081 2397 12115 2431
rect 18797 2397 18831 2431
rect 9919 2329 9953 2363
rect 14381 2329 14415 2363
rect 16037 2329 16071 2363
rect 18429 2329 18463 2363
rect 19717 2329 19751 2363
rect 20085 2329 20119 2363
rect 21373 2329 21407 2363
rect 3709 2261 3743 2295
rect 3801 2261 3835 2295
rect 15301 2261 15335 2295
rect 15761 2261 15795 2295
rect 17785 2261 17819 2295
<< metal1 >>
rect 13814 23536 13820 23588
rect 13872 23576 13878 23588
rect 14642 23576 14648 23588
rect 13872 23548 14648 23576
rect 13872 23536 13878 23548
rect 14642 23536 14648 23548
rect 14700 23536 14706 23588
rect 1104 21786 22816 21808
rect 1104 21734 4982 21786
rect 5034 21734 5046 21786
rect 5098 21734 5110 21786
rect 5162 21734 5174 21786
rect 5226 21734 12982 21786
rect 13034 21734 13046 21786
rect 13098 21734 13110 21786
rect 13162 21734 13174 21786
rect 13226 21734 20982 21786
rect 21034 21734 21046 21786
rect 21098 21734 21110 21786
rect 21162 21734 21174 21786
rect 21226 21734 22816 21786
rect 1104 21712 22816 21734
rect 1104 21242 22816 21264
rect 1104 21190 8982 21242
rect 9034 21190 9046 21242
rect 9098 21190 9110 21242
rect 9162 21190 9174 21242
rect 9226 21190 16982 21242
rect 17034 21190 17046 21242
rect 17098 21190 17110 21242
rect 17162 21190 17174 21242
rect 17226 21190 22816 21242
rect 1104 21168 22816 21190
rect 8202 20924 8208 20936
rect 8163 20896 8208 20924
rect 8202 20884 8208 20896
rect 8260 20884 8266 20936
rect 18325 20927 18383 20933
rect 18325 20893 18337 20927
rect 18371 20924 18383 20927
rect 18414 20924 18420 20936
rect 18371 20896 18420 20924
rect 18371 20893 18383 20896
rect 18325 20887 18383 20893
rect 18414 20884 18420 20896
rect 18472 20884 18478 20936
rect 1104 20698 22816 20720
rect 1104 20646 4982 20698
rect 5034 20646 5046 20698
rect 5098 20646 5110 20698
rect 5162 20646 5174 20698
rect 5226 20646 12982 20698
rect 13034 20646 13046 20698
rect 13098 20646 13110 20698
rect 13162 20646 13174 20698
rect 13226 20646 20982 20698
rect 21034 20646 21046 20698
rect 21098 20646 21110 20698
rect 21162 20646 21174 20698
rect 21226 20646 22816 20698
rect 1104 20624 22816 20646
rect 1578 20584 1584 20596
rect 1539 20556 1584 20584
rect 1578 20544 1584 20556
rect 1636 20544 1642 20596
rect 5491 20587 5549 20593
rect 5491 20553 5503 20587
rect 5537 20584 5549 20587
rect 6362 20584 6368 20596
rect 5537 20556 6368 20584
rect 5537 20553 5549 20556
rect 5491 20547 5549 20553
rect 6362 20544 6368 20556
rect 6420 20544 6426 20596
rect 8202 20544 8208 20596
rect 8260 20584 8266 20596
rect 8297 20587 8355 20593
rect 8297 20584 8309 20587
rect 8260 20556 8309 20584
rect 8260 20544 8266 20556
rect 8297 20553 8309 20556
rect 8343 20584 8355 20587
rect 8570 20584 8576 20596
rect 8343 20556 8576 20584
rect 8343 20553 8355 20556
rect 8297 20547 8355 20553
rect 8570 20544 8576 20556
rect 8628 20544 8634 20596
rect 11149 20587 11207 20593
rect 11149 20553 11161 20587
rect 11195 20584 11207 20587
rect 11606 20584 11612 20596
rect 11195 20556 11612 20584
rect 11195 20553 11207 20556
rect 11149 20547 11207 20553
rect 11606 20544 11612 20556
rect 11664 20544 11670 20596
rect 19153 20587 19211 20593
rect 19153 20553 19165 20587
rect 19199 20584 19211 20587
rect 19702 20584 19708 20596
rect 19199 20556 19708 20584
rect 19199 20553 19211 20556
rect 19153 20547 19211 20553
rect 19702 20544 19708 20556
rect 19760 20544 19766 20596
rect 20346 20584 20352 20596
rect 20307 20556 20352 20584
rect 20346 20544 20352 20556
rect 20404 20544 20410 20596
rect 4154 20476 4160 20528
rect 4212 20516 4218 20528
rect 7607 20519 7665 20525
rect 7607 20516 7619 20519
rect 4212 20488 7619 20516
rect 4212 20476 4218 20488
rect 7607 20485 7619 20488
rect 7653 20485 7665 20519
rect 9398 20516 9404 20528
rect 7607 20479 7665 20485
rect 7852 20488 9404 20516
rect 2041 20451 2099 20457
rect 2041 20448 2053 20451
rect 1412 20420 2053 20448
rect 1412 20389 1440 20420
rect 2041 20417 2053 20420
rect 2087 20448 2099 20451
rect 7852 20448 7880 20488
rect 9398 20476 9404 20488
rect 9456 20476 9462 20528
rect 2087 20420 7880 20448
rect 2087 20417 2099 20420
rect 2041 20411 2099 20417
rect 8570 20408 8576 20460
rect 8628 20448 8634 20460
rect 8628 20420 8673 20448
rect 8628 20408 8634 20420
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20349 1455 20383
rect 1397 20343 1455 20349
rect 5420 20383 5478 20389
rect 5420 20349 5432 20383
rect 5466 20380 5478 20383
rect 5534 20380 5540 20392
rect 5466 20352 5540 20380
rect 5466 20349 5478 20352
rect 5420 20343 5478 20349
rect 5534 20340 5540 20352
rect 5592 20380 5598 20392
rect 5813 20383 5871 20389
rect 5813 20380 5825 20383
rect 5592 20352 5825 20380
rect 5592 20340 5598 20352
rect 5813 20349 5825 20352
rect 5859 20349 5871 20383
rect 5813 20343 5871 20349
rect 7520 20383 7578 20389
rect 7520 20349 7532 20383
rect 7566 20349 7578 20383
rect 10962 20380 10968 20392
rect 10923 20352 10968 20380
rect 7520 20343 7578 20349
rect 7377 20247 7435 20253
rect 7377 20213 7389 20247
rect 7423 20244 7435 20247
rect 7535 20244 7563 20343
rect 10962 20340 10968 20352
rect 11020 20380 11026 20392
rect 11517 20383 11575 20389
rect 11517 20380 11529 20383
rect 11020 20352 11529 20380
rect 11020 20340 11026 20352
rect 11517 20349 11529 20352
rect 11563 20349 11575 20383
rect 11517 20343 11575 20349
rect 12504 20383 12562 20389
rect 12504 20349 12516 20383
rect 12550 20380 12562 20383
rect 12550 20352 13032 20380
rect 12550 20349 12562 20352
rect 12504 20343 12562 20349
rect 8021 20315 8079 20321
rect 8021 20281 8033 20315
rect 8067 20312 8079 20315
rect 8665 20315 8723 20321
rect 8665 20312 8677 20315
rect 8067 20284 8677 20312
rect 8067 20281 8079 20284
rect 8021 20275 8079 20281
rect 8665 20281 8677 20284
rect 8711 20312 8723 20315
rect 8754 20312 8760 20324
rect 8711 20284 8760 20312
rect 8711 20281 8723 20284
rect 8665 20275 8723 20281
rect 8754 20272 8760 20284
rect 8812 20272 8818 20324
rect 9217 20315 9275 20321
rect 9217 20281 9229 20315
rect 9263 20312 9275 20315
rect 11330 20312 11336 20324
rect 9263 20284 11336 20312
rect 9263 20281 9275 20284
rect 9217 20275 9275 20281
rect 9232 20244 9260 20275
rect 11330 20272 11336 20284
rect 11388 20272 11394 20324
rect 7423 20216 9260 20244
rect 7423 20213 7435 20216
rect 7377 20207 7435 20213
rect 11606 20204 11612 20256
rect 11664 20244 11670 20256
rect 13004 20253 13032 20352
rect 18874 20340 18880 20392
rect 18932 20380 18938 20392
rect 18969 20383 19027 20389
rect 18969 20380 18981 20383
rect 18932 20352 18981 20380
rect 18932 20340 18938 20352
rect 18969 20349 18981 20352
rect 19015 20349 19027 20383
rect 18969 20343 19027 20349
rect 18984 20312 19012 20343
rect 19242 20340 19248 20392
rect 19300 20380 19306 20392
rect 20108 20383 20166 20389
rect 20108 20380 20120 20383
rect 19300 20352 20120 20380
rect 19300 20340 19306 20352
rect 20108 20349 20120 20352
rect 20154 20380 20166 20383
rect 20533 20383 20591 20389
rect 20533 20380 20545 20383
rect 20154 20352 20545 20380
rect 20154 20349 20166 20352
rect 20108 20343 20166 20349
rect 20533 20349 20545 20352
rect 20579 20349 20591 20383
rect 20533 20343 20591 20349
rect 19521 20315 19579 20321
rect 19521 20312 19533 20315
rect 18984 20284 19533 20312
rect 19521 20281 19533 20284
rect 19567 20281 19579 20315
rect 19521 20275 19579 20281
rect 12575 20247 12633 20253
rect 12575 20244 12587 20247
rect 11664 20216 12587 20244
rect 11664 20204 11670 20216
rect 12575 20213 12587 20216
rect 12621 20213 12633 20247
rect 12575 20207 12633 20213
rect 12989 20247 13047 20253
rect 12989 20213 13001 20247
rect 13035 20244 13047 20247
rect 13354 20244 13360 20256
rect 13035 20216 13360 20244
rect 13035 20213 13047 20216
rect 12989 20207 13047 20213
rect 13354 20204 13360 20216
rect 13412 20204 13418 20256
rect 1104 20154 22816 20176
rect 1104 20102 8982 20154
rect 9034 20102 9046 20154
rect 9098 20102 9110 20154
rect 9162 20102 9174 20154
rect 9226 20102 16982 20154
rect 17034 20102 17046 20154
rect 17098 20102 17110 20154
rect 17162 20102 17174 20154
rect 17226 20102 22816 20154
rect 1104 20080 22816 20102
rect 8754 20040 8760 20052
rect 8715 20012 8760 20040
rect 8754 20000 8760 20012
rect 8812 20000 8818 20052
rect 5261 19975 5319 19981
rect 5261 19941 5273 19975
rect 5307 19972 5319 19975
rect 5350 19972 5356 19984
rect 5307 19944 5356 19972
rect 5307 19941 5319 19944
rect 5261 19935 5319 19941
rect 5350 19932 5356 19944
rect 5408 19932 5414 19984
rect 8199 19975 8257 19981
rect 8199 19941 8211 19975
rect 8245 19972 8257 19975
rect 8662 19972 8668 19984
rect 8245 19944 8668 19972
rect 8245 19941 8257 19944
rect 8199 19935 8257 19941
rect 8662 19932 8668 19944
rect 8720 19932 8726 19984
rect 10778 19972 10784 19984
rect 10739 19944 10784 19972
rect 10778 19932 10784 19944
rect 10836 19932 10842 19984
rect 18414 19972 18420 19984
rect 18375 19944 18420 19972
rect 18414 19932 18420 19944
rect 18472 19932 18478 19984
rect 18506 19932 18512 19984
rect 18564 19972 18570 19984
rect 18564 19944 18609 19972
rect 18564 19932 18570 19944
rect 4065 19839 4123 19845
rect 4065 19805 4077 19839
rect 4111 19836 4123 19839
rect 4798 19836 4804 19848
rect 4111 19808 4804 19836
rect 4111 19805 4123 19808
rect 4065 19799 4123 19805
rect 4798 19796 4804 19808
rect 4856 19836 4862 19848
rect 5169 19839 5227 19845
rect 5169 19836 5181 19839
rect 4856 19808 5181 19836
rect 4856 19796 4862 19808
rect 5169 19805 5181 19808
rect 5215 19805 5227 19839
rect 5534 19836 5540 19848
rect 5495 19808 5540 19836
rect 5169 19799 5227 19805
rect 5534 19796 5540 19808
rect 5592 19796 5598 19848
rect 7834 19836 7840 19848
rect 7795 19808 7840 19836
rect 7834 19796 7840 19808
rect 7892 19796 7898 19848
rect 10689 19839 10747 19845
rect 10689 19805 10701 19839
rect 10735 19805 10747 19839
rect 11330 19836 11336 19848
rect 11243 19808 11336 19836
rect 10689 19799 10747 19805
rect 10594 19728 10600 19780
rect 10652 19768 10658 19780
rect 10704 19768 10732 19799
rect 11330 19796 11336 19808
rect 11388 19836 11394 19848
rect 11698 19836 11704 19848
rect 11388 19808 11704 19836
rect 11388 19796 11394 19808
rect 11698 19796 11704 19808
rect 11756 19796 11762 19848
rect 19061 19839 19119 19845
rect 19061 19805 19073 19839
rect 19107 19836 19119 19839
rect 19242 19836 19248 19848
rect 19107 19808 19248 19836
rect 19107 19805 19119 19808
rect 19061 19799 19119 19805
rect 19242 19796 19248 19808
rect 19300 19796 19306 19848
rect 10652 19740 10732 19768
rect 10652 19728 10658 19740
rect 9950 19700 9956 19712
rect 9911 19672 9956 19700
rect 9950 19660 9956 19672
rect 10008 19660 10014 19712
rect 18046 19700 18052 19712
rect 18007 19672 18052 19700
rect 18046 19660 18052 19672
rect 18104 19660 18110 19712
rect 1104 19610 22816 19632
rect 1104 19558 4982 19610
rect 5034 19558 5046 19610
rect 5098 19558 5110 19610
rect 5162 19558 5174 19610
rect 5226 19558 12982 19610
rect 13034 19558 13046 19610
rect 13098 19558 13110 19610
rect 13162 19558 13174 19610
rect 13226 19558 20982 19610
rect 21034 19558 21046 19610
rect 21098 19558 21110 19610
rect 21162 19558 21174 19610
rect 21226 19558 22816 19610
rect 1104 19536 22816 19558
rect 4798 19456 4804 19508
rect 4856 19496 4862 19508
rect 5261 19499 5319 19505
rect 5261 19496 5273 19499
rect 4856 19468 5273 19496
rect 4856 19456 4862 19468
rect 5261 19465 5273 19468
rect 5307 19465 5319 19499
rect 5261 19459 5319 19465
rect 10778 19456 10784 19508
rect 10836 19496 10842 19508
rect 10873 19499 10931 19505
rect 10873 19496 10885 19499
rect 10836 19468 10885 19496
rect 10836 19456 10842 19468
rect 10873 19465 10885 19468
rect 10919 19496 10931 19499
rect 11149 19499 11207 19505
rect 11149 19496 11161 19499
rect 10919 19468 11161 19496
rect 10919 19465 10931 19468
rect 10873 19459 10931 19465
rect 11149 19465 11161 19468
rect 11195 19465 11207 19499
rect 11149 19459 11207 19465
rect 17497 19499 17555 19505
rect 17497 19465 17509 19499
rect 17543 19496 17555 19499
rect 18506 19496 18512 19508
rect 17543 19468 18512 19496
rect 17543 19465 17555 19468
rect 17497 19459 17555 19465
rect 18506 19456 18512 19468
rect 18564 19496 18570 19508
rect 18969 19499 19027 19505
rect 18969 19496 18981 19499
rect 18564 19468 18981 19496
rect 18564 19456 18570 19468
rect 18969 19465 18981 19468
rect 19015 19465 19027 19499
rect 18969 19459 19027 19465
rect 21039 19499 21097 19505
rect 21039 19465 21051 19499
rect 21085 19496 21097 19499
rect 21266 19496 21272 19508
rect 21085 19468 21272 19496
rect 21085 19465 21097 19468
rect 21039 19459 21097 19465
rect 21266 19456 21272 19468
rect 21324 19456 21330 19508
rect 4985 19431 5043 19437
rect 4985 19397 4997 19431
rect 5031 19428 5043 19431
rect 5350 19428 5356 19440
rect 5031 19400 5356 19428
rect 5031 19397 5043 19400
rect 4985 19391 5043 19397
rect 5350 19388 5356 19400
rect 5408 19428 5414 19440
rect 5629 19431 5687 19437
rect 5629 19428 5641 19431
rect 5408 19400 5641 19428
rect 5408 19388 5414 19400
rect 5629 19397 5641 19400
rect 5675 19397 5687 19431
rect 5629 19391 5687 19397
rect 7561 19363 7619 19369
rect 7561 19329 7573 19363
rect 7607 19360 7619 19363
rect 9950 19360 9956 19372
rect 7607 19332 8248 19360
rect 9911 19332 9956 19360
rect 7607 19329 7619 19332
rect 7561 19323 7619 19329
rect 4065 19295 4123 19301
rect 4065 19292 4077 19295
rect 3620 19264 4077 19292
rect 3620 19168 3648 19264
rect 4065 19261 4077 19264
rect 4111 19261 4123 19295
rect 7650 19292 7656 19304
rect 7611 19264 7656 19292
rect 4065 19255 4123 19261
rect 7650 19252 7656 19264
rect 7708 19252 7714 19304
rect 8220 19301 8248 19332
rect 9950 19320 9956 19332
rect 10008 19320 10014 19372
rect 8205 19295 8263 19301
rect 8205 19261 8217 19295
rect 8251 19292 8263 19295
rect 8570 19292 8576 19304
rect 8251 19264 8576 19292
rect 8251 19261 8263 19264
rect 8205 19255 8263 19261
rect 8570 19252 8576 19264
rect 8628 19252 8634 19304
rect 16666 19292 16672 19304
rect 16627 19264 16672 19292
rect 16666 19252 16672 19264
rect 16724 19252 16730 19304
rect 16853 19295 16911 19301
rect 16853 19261 16865 19295
rect 16899 19261 16911 19295
rect 16853 19255 16911 19261
rect 4386 19227 4444 19233
rect 4386 19224 4398 19227
rect 4172 19196 4398 19224
rect 4172 19168 4200 19196
rect 4386 19193 4398 19196
rect 4432 19193 4444 19227
rect 4386 19187 4444 19193
rect 7193 19227 7251 19233
rect 7193 19193 7205 19227
rect 7239 19224 7251 19227
rect 10274 19227 10332 19233
rect 10274 19224 10286 19227
rect 7239 19196 7880 19224
rect 7239 19193 7251 19196
rect 7193 19187 7251 19193
rect 7852 19168 7880 19196
rect 9784 19196 10286 19224
rect 3602 19156 3608 19168
rect 3563 19128 3608 19156
rect 3602 19116 3608 19128
rect 3660 19116 3666 19168
rect 3973 19159 4031 19165
rect 3973 19125 3985 19159
rect 4019 19156 4031 19159
rect 4154 19156 4160 19168
rect 4019 19128 4160 19156
rect 4019 19125 4031 19128
rect 3973 19119 4031 19125
rect 4154 19116 4160 19128
rect 4212 19116 4218 19168
rect 7834 19116 7840 19168
rect 7892 19156 7898 19168
rect 7929 19159 7987 19165
rect 7929 19156 7941 19159
rect 7892 19128 7941 19156
rect 7892 19116 7898 19128
rect 7929 19125 7941 19128
rect 7975 19125 7987 19159
rect 8662 19156 8668 19168
rect 8623 19128 8668 19156
rect 7929 19119 7987 19125
rect 8662 19116 8668 19128
rect 8720 19156 8726 19168
rect 9784 19165 9812 19196
rect 10274 19193 10286 19196
rect 10320 19193 10332 19227
rect 16868 19224 16896 19255
rect 17310 19252 17316 19304
rect 17368 19292 17374 19304
rect 18046 19292 18052 19304
rect 17368 19264 18052 19292
rect 17368 19252 17374 19264
rect 18046 19252 18052 19264
rect 18104 19252 18110 19304
rect 20968 19295 21026 19301
rect 20968 19261 20980 19295
rect 21014 19292 21026 19295
rect 21361 19295 21419 19301
rect 21361 19292 21373 19295
rect 21014 19264 21373 19292
rect 21014 19261 21026 19264
rect 20968 19255 21026 19261
rect 21361 19261 21373 19264
rect 21407 19292 21419 19295
rect 21450 19292 21456 19304
rect 21407 19264 21456 19292
rect 21407 19261 21419 19264
rect 21361 19255 21419 19261
rect 21450 19252 21456 19264
rect 21508 19252 21514 19304
rect 10274 19187 10332 19193
rect 16224 19196 16896 19224
rect 17129 19227 17187 19233
rect 16224 19168 16252 19196
rect 17129 19193 17141 19227
rect 17175 19224 17187 19227
rect 17402 19224 17408 19236
rect 17175 19196 17408 19224
rect 17175 19193 17187 19196
rect 17129 19187 17187 19193
rect 17402 19184 17408 19196
rect 17460 19184 17466 19236
rect 18370 19227 18428 19233
rect 18370 19193 18382 19227
rect 18416 19193 18428 19227
rect 18370 19187 18428 19193
rect 9769 19159 9827 19165
rect 9769 19156 9781 19159
rect 8720 19128 9781 19156
rect 8720 19116 8726 19128
rect 9769 19125 9781 19128
rect 9815 19125 9827 19159
rect 9769 19119 9827 19125
rect 10594 19116 10600 19168
rect 10652 19156 10658 19168
rect 11517 19159 11575 19165
rect 11517 19156 11529 19159
rect 10652 19128 11529 19156
rect 10652 19116 10658 19128
rect 11517 19125 11529 19128
rect 11563 19125 11575 19159
rect 16206 19156 16212 19168
rect 16167 19128 16212 19156
rect 11517 19119 11575 19125
rect 16206 19116 16212 19128
rect 16264 19116 16270 19168
rect 17770 19156 17776 19168
rect 17731 19128 17776 19156
rect 17770 19116 17776 19128
rect 17828 19156 17834 19168
rect 18385 19156 18413 19187
rect 17828 19128 18413 19156
rect 17828 19116 17834 19128
rect 1104 19066 22816 19088
rect 1104 19014 8982 19066
rect 9034 19014 9046 19066
rect 9098 19014 9110 19066
rect 9162 19014 9174 19066
rect 9226 19014 16982 19066
rect 17034 19014 17046 19066
rect 17098 19014 17110 19066
rect 17162 19014 17174 19066
rect 17226 19014 22816 19066
rect 1104 18992 22816 19014
rect 1578 18952 1584 18964
rect 1539 18924 1584 18952
rect 1578 18912 1584 18924
rect 1636 18912 1642 18964
rect 6454 18952 6460 18964
rect 6415 18924 6460 18952
rect 6454 18912 6460 18924
rect 6512 18912 6518 18964
rect 9950 18952 9956 18964
rect 9911 18924 9956 18952
rect 9950 18912 9956 18924
rect 10008 18912 10014 18964
rect 18414 18952 18420 18964
rect 18375 18924 18420 18952
rect 18414 18912 18420 18924
rect 18472 18912 18478 18964
rect 4706 18844 4712 18896
rect 4764 18884 4770 18896
rect 4985 18887 5043 18893
rect 4985 18884 4997 18887
rect 4764 18856 4997 18884
rect 4764 18844 4770 18856
rect 4985 18853 4997 18856
rect 5031 18853 5043 18887
rect 11514 18884 11520 18896
rect 11475 18856 11520 18884
rect 4985 18847 5043 18853
rect 11514 18844 11520 18856
rect 11572 18844 11578 18896
rect 17310 18884 17316 18896
rect 17271 18856 17316 18884
rect 17310 18844 17316 18856
rect 17368 18844 17374 18896
rect 18782 18884 18788 18896
rect 18743 18856 18788 18884
rect 18782 18844 18788 18856
rect 18840 18844 18846 18896
rect 1394 18816 1400 18828
rect 1355 18788 1400 18816
rect 1394 18776 1400 18788
rect 1452 18776 1458 18828
rect 6641 18819 6699 18825
rect 6641 18785 6653 18819
rect 6687 18785 6699 18819
rect 6641 18779 6699 18785
rect 4893 18751 4951 18757
rect 4893 18717 4905 18751
rect 4939 18717 4951 18751
rect 5534 18748 5540 18760
rect 5495 18720 5540 18748
rect 4893 18711 4951 18717
rect 4908 18680 4936 18711
rect 5534 18708 5540 18720
rect 5592 18708 5598 18760
rect 6086 18708 6092 18760
rect 6144 18748 6150 18760
rect 6656 18748 6684 18779
rect 6730 18776 6736 18828
rect 6788 18816 6794 18828
rect 6825 18819 6883 18825
rect 6825 18816 6837 18819
rect 6788 18788 6837 18816
rect 6788 18776 6794 18788
rect 6825 18785 6837 18788
rect 6871 18785 6883 18819
rect 8294 18816 8300 18828
rect 8255 18788 8300 18816
rect 6825 18779 6883 18785
rect 8294 18776 8300 18788
rect 8352 18776 8358 18828
rect 8570 18816 8576 18828
rect 8531 18788 8576 18816
rect 8570 18776 8576 18788
rect 8628 18776 8634 18828
rect 9953 18819 10011 18825
rect 9953 18785 9965 18819
rect 9999 18785 10011 18819
rect 10134 18816 10140 18828
rect 10095 18788 10140 18816
rect 9953 18779 10011 18785
rect 8312 18748 8340 18776
rect 8754 18748 8760 18760
rect 6144 18720 8340 18748
rect 8715 18720 8760 18748
rect 6144 18708 6150 18720
rect 8754 18708 8760 18720
rect 8812 18708 8818 18760
rect 9968 18748 9996 18779
rect 10134 18776 10140 18788
rect 10192 18776 10198 18828
rect 15194 18816 15200 18828
rect 15155 18788 15200 18816
rect 15194 18776 15200 18788
rect 15252 18776 15258 18828
rect 16850 18816 16856 18828
rect 16811 18788 16856 18816
rect 16850 18776 16856 18788
rect 16908 18776 16914 18828
rect 17034 18816 17040 18828
rect 16995 18788 17040 18816
rect 17034 18776 17040 18788
rect 17092 18776 17098 18828
rect 10410 18748 10416 18760
rect 9968 18720 10416 18748
rect 10410 18708 10416 18720
rect 10468 18708 10474 18760
rect 11422 18748 11428 18760
rect 11383 18720 11428 18748
rect 11422 18708 11428 18720
rect 11480 18708 11486 18760
rect 11698 18748 11704 18760
rect 11659 18720 11704 18748
rect 11698 18708 11704 18720
rect 11756 18708 11762 18760
rect 18690 18748 18696 18760
rect 18651 18720 18696 18748
rect 18690 18708 18696 18720
rect 18748 18708 18754 18760
rect 5442 18680 5448 18692
rect 4908 18652 5448 18680
rect 5442 18640 5448 18652
rect 5500 18640 5506 18692
rect 19242 18680 19248 18692
rect 19203 18652 19248 18680
rect 19242 18640 19248 18652
rect 19300 18640 19306 18692
rect 3421 18615 3479 18621
rect 3421 18581 3433 18615
rect 3467 18612 3479 18615
rect 3510 18612 3516 18624
rect 3467 18584 3516 18612
rect 3467 18581 3479 18584
rect 3421 18575 3479 18581
rect 3510 18572 3516 18584
rect 3568 18612 3574 18624
rect 7650 18612 7656 18624
rect 3568 18584 7656 18612
rect 3568 18572 3574 18584
rect 7650 18572 7656 18584
rect 7708 18572 7714 18624
rect 10778 18612 10784 18624
rect 10739 18584 10784 18612
rect 10778 18572 10784 18584
rect 10836 18572 10842 18624
rect 12526 18612 12532 18624
rect 12487 18584 12532 18612
rect 12526 18572 12532 18584
rect 12584 18572 12590 18624
rect 15427 18615 15485 18621
rect 15427 18581 15439 18615
rect 15473 18612 15485 18615
rect 15562 18612 15568 18624
rect 15473 18584 15568 18612
rect 15473 18581 15485 18584
rect 15427 18575 15485 18581
rect 15562 18572 15568 18584
rect 15620 18572 15626 18624
rect 16485 18615 16543 18621
rect 16485 18581 16497 18615
rect 16531 18612 16543 18615
rect 16666 18612 16672 18624
rect 16531 18584 16672 18612
rect 16531 18581 16543 18584
rect 16485 18575 16543 18581
rect 16666 18572 16672 18584
rect 16724 18572 16730 18624
rect 1104 18522 22816 18544
rect 1104 18470 4982 18522
rect 5034 18470 5046 18522
rect 5098 18470 5110 18522
rect 5162 18470 5174 18522
rect 5226 18470 12982 18522
rect 13034 18470 13046 18522
rect 13098 18470 13110 18522
rect 13162 18470 13174 18522
rect 13226 18470 20982 18522
rect 21034 18470 21046 18522
rect 21098 18470 21110 18522
rect 21162 18470 21174 18522
rect 21226 18470 22816 18522
rect 1104 18448 22816 18470
rect 1394 18368 1400 18420
rect 1452 18408 1458 18420
rect 1581 18411 1639 18417
rect 1581 18408 1593 18411
rect 1452 18380 1593 18408
rect 1452 18368 1458 18380
rect 1581 18377 1593 18380
rect 1627 18377 1639 18411
rect 4706 18408 4712 18420
rect 4667 18380 4712 18408
rect 1581 18371 1639 18377
rect 1596 18340 1624 18371
rect 4706 18368 4712 18380
rect 4764 18368 4770 18420
rect 6086 18408 6092 18420
rect 5368 18380 5994 18408
rect 6047 18380 6092 18408
rect 5368 18340 5396 18380
rect 5534 18340 5540 18352
rect 1596 18312 5396 18340
rect 5495 18312 5540 18340
rect 5534 18300 5540 18312
rect 5592 18300 5598 18352
rect 5966 18340 5994 18380
rect 6086 18368 6092 18380
rect 6144 18368 6150 18420
rect 17402 18408 17408 18420
rect 17363 18380 17408 18408
rect 17402 18368 17408 18380
rect 17460 18368 17466 18420
rect 18782 18368 18788 18420
rect 18840 18408 18846 18420
rect 18969 18411 19027 18417
rect 18969 18408 18981 18411
rect 18840 18380 18981 18408
rect 18840 18368 18846 18380
rect 18969 18377 18981 18380
rect 19015 18408 19027 18411
rect 19245 18411 19303 18417
rect 19245 18408 19257 18411
rect 19015 18380 19257 18408
rect 19015 18377 19027 18380
rect 18969 18371 19027 18377
rect 19245 18377 19257 18380
rect 19291 18377 19303 18411
rect 19245 18371 19303 18377
rect 8202 18340 8208 18352
rect 5966 18312 8208 18340
rect 8202 18300 8208 18312
rect 8260 18300 8266 18352
rect 9769 18343 9827 18349
rect 9769 18309 9781 18343
rect 9815 18340 9827 18343
rect 10042 18340 10048 18352
rect 9815 18312 10048 18340
rect 9815 18309 9827 18312
rect 9769 18303 9827 18309
rect 10042 18300 10048 18312
rect 10100 18340 10106 18352
rect 10778 18340 10784 18352
rect 10100 18312 10784 18340
rect 10100 18300 10106 18312
rect 10778 18300 10784 18312
rect 10836 18300 10842 18352
rect 11514 18300 11520 18352
rect 11572 18340 11578 18352
rect 11701 18343 11759 18349
rect 11701 18340 11713 18343
rect 11572 18312 11713 18340
rect 11572 18300 11578 18312
rect 11701 18309 11713 18312
rect 11747 18340 11759 18343
rect 13357 18343 13415 18349
rect 13357 18340 13369 18343
rect 11747 18312 13369 18340
rect 11747 18309 11759 18312
rect 11701 18303 11759 18309
rect 13357 18309 13369 18312
rect 13403 18309 13415 18343
rect 13357 18303 13415 18309
rect 14182 18300 14188 18352
rect 14240 18340 14246 18352
rect 16206 18340 16212 18352
rect 14240 18312 16212 18340
rect 14240 18300 14246 18312
rect 16206 18300 16212 18312
rect 16264 18340 16270 18352
rect 16577 18343 16635 18349
rect 16577 18340 16589 18343
rect 16264 18312 16589 18340
rect 16264 18300 16270 18312
rect 16577 18309 16589 18312
rect 16623 18340 16635 18343
rect 17034 18340 17040 18352
rect 16623 18312 17040 18340
rect 16623 18309 16635 18312
rect 16577 18303 16635 18309
rect 17034 18300 17040 18312
rect 17092 18300 17098 18352
rect 6365 18275 6423 18281
rect 6365 18272 6377 18275
rect 4126 18244 6377 18272
rect 3510 18204 3516 18216
rect 3471 18176 3516 18204
rect 3510 18164 3516 18176
rect 3568 18164 3574 18216
rect 3789 18207 3847 18213
rect 3789 18173 3801 18207
rect 3835 18204 3847 18207
rect 4126 18204 4154 18244
rect 6365 18241 6377 18244
rect 6411 18272 6423 18275
rect 6730 18272 6736 18284
rect 6411 18244 6736 18272
rect 6411 18241 6423 18244
rect 6365 18235 6423 18241
rect 6730 18232 6736 18244
rect 6788 18232 6794 18284
rect 7006 18232 7012 18284
rect 7064 18272 7070 18284
rect 7193 18275 7251 18281
rect 7193 18272 7205 18275
rect 7064 18244 7205 18272
rect 7064 18232 7070 18244
rect 7193 18241 7205 18244
rect 7239 18241 7251 18275
rect 7193 18235 7251 18241
rect 8754 18232 8760 18284
rect 8812 18272 8818 18284
rect 8849 18275 8907 18281
rect 8849 18272 8861 18275
rect 8812 18244 8861 18272
rect 8812 18232 8818 18244
rect 8849 18241 8861 18244
rect 8895 18241 8907 18275
rect 8849 18235 8907 18241
rect 11333 18275 11391 18281
rect 11333 18241 11345 18275
rect 11379 18272 11391 18275
rect 11422 18272 11428 18284
rect 11379 18244 11428 18272
rect 11379 18241 11391 18244
rect 11333 18235 11391 18241
rect 11422 18232 11428 18244
rect 11480 18232 11486 18284
rect 11790 18232 11796 18284
rect 11848 18272 11854 18284
rect 15194 18272 15200 18284
rect 11848 18244 15200 18272
rect 11848 18232 11854 18244
rect 15194 18232 15200 18244
rect 15252 18272 15258 18284
rect 15933 18275 15991 18281
rect 15933 18272 15945 18275
rect 15252 18244 15945 18272
rect 15252 18232 15258 18244
rect 15933 18241 15945 18244
rect 15979 18241 15991 18275
rect 15933 18235 15991 18241
rect 8570 18204 8576 18216
rect 3835 18176 4154 18204
rect 8128 18176 8576 18204
rect 3835 18173 3847 18176
rect 3789 18167 3847 18173
rect 3804 18136 3832 18167
rect 4982 18136 4988 18148
rect 3160 18108 3832 18136
rect 4943 18108 4988 18136
rect 2866 18028 2872 18080
rect 2924 18068 2930 18080
rect 3160 18077 3188 18108
rect 4982 18096 4988 18108
rect 5040 18096 5046 18148
rect 5077 18139 5135 18145
rect 5077 18105 5089 18139
rect 5123 18105 5135 18139
rect 6914 18136 6920 18148
rect 6875 18108 6920 18136
rect 5077 18099 5135 18105
rect 3145 18071 3203 18077
rect 3145 18068 3157 18071
rect 2924 18040 3157 18068
rect 2924 18028 2930 18040
rect 3145 18037 3157 18040
rect 3191 18037 3203 18071
rect 3602 18068 3608 18080
rect 3563 18040 3608 18068
rect 3145 18031 3203 18037
rect 3602 18028 3608 18040
rect 3660 18028 3666 18080
rect 4433 18071 4491 18077
rect 4433 18037 4445 18071
rect 4479 18068 4491 18071
rect 4798 18068 4804 18080
rect 4479 18040 4804 18068
rect 4479 18037 4491 18040
rect 4433 18031 4491 18037
rect 4798 18028 4804 18040
rect 4856 18068 4862 18080
rect 5092 18068 5120 18099
rect 6914 18096 6920 18108
rect 6972 18096 6978 18148
rect 7009 18139 7067 18145
rect 7009 18105 7021 18139
rect 7055 18136 7067 18139
rect 7098 18136 7104 18148
rect 7055 18108 7104 18136
rect 7055 18105 7067 18108
rect 7009 18099 7067 18105
rect 7098 18096 7104 18108
rect 7156 18096 7162 18148
rect 8128 18080 8156 18176
rect 8570 18164 8576 18176
rect 8628 18204 8634 18216
rect 10045 18207 10103 18213
rect 10045 18204 10057 18207
rect 8628 18176 10057 18204
rect 8628 18164 8634 18176
rect 10045 18173 10057 18176
rect 10091 18204 10103 18207
rect 10134 18204 10140 18216
rect 10091 18176 10140 18204
rect 10091 18173 10103 18176
rect 10045 18167 10103 18173
rect 10134 18164 10140 18176
rect 10192 18164 10198 18216
rect 12437 18207 12495 18213
rect 12437 18173 12449 18207
rect 12483 18204 12495 18207
rect 12526 18204 12532 18216
rect 12483 18176 12532 18204
rect 12483 18173 12495 18176
rect 12437 18167 12495 18173
rect 12526 18164 12532 18176
rect 12584 18164 12590 18216
rect 17052 18204 17080 18300
rect 17420 18272 17448 18368
rect 18049 18275 18107 18281
rect 18049 18272 18061 18275
rect 17420 18244 18061 18272
rect 18049 18241 18061 18244
rect 18095 18241 18107 18275
rect 18049 18235 18107 18241
rect 19613 18207 19671 18213
rect 19613 18204 19625 18207
rect 17052 18176 19625 18204
rect 19613 18173 19625 18176
rect 19659 18173 19671 18207
rect 19794 18204 19800 18216
rect 19755 18176 19800 18204
rect 19613 18167 19671 18173
rect 9170 18139 9228 18145
rect 9170 18136 9182 18139
rect 8680 18108 9182 18136
rect 8680 18080 8708 18108
rect 9170 18105 9182 18108
rect 9216 18105 9228 18139
rect 10686 18136 10692 18148
rect 10647 18108 10692 18136
rect 9170 18099 9228 18105
rect 10686 18096 10692 18108
rect 10744 18096 10750 18148
rect 10778 18096 10784 18148
rect 10836 18136 10842 18148
rect 15010 18136 15016 18148
rect 10836 18108 10881 18136
rect 14971 18108 15016 18136
rect 10836 18096 10842 18108
rect 15010 18096 15016 18108
rect 15068 18096 15074 18148
rect 15105 18139 15163 18145
rect 15105 18105 15117 18139
rect 15151 18105 15163 18139
rect 15105 18099 15163 18105
rect 15657 18139 15715 18145
rect 15657 18105 15669 18139
rect 15703 18136 15715 18139
rect 16022 18136 16028 18148
rect 15703 18108 16028 18136
rect 15703 18105 15715 18108
rect 15657 18099 15715 18105
rect 8110 18068 8116 18080
rect 4856 18040 5120 18068
rect 8071 18040 8116 18068
rect 4856 18028 4862 18040
rect 8110 18028 8116 18040
rect 8168 18028 8174 18080
rect 8662 18068 8668 18080
rect 8623 18040 8668 18068
rect 8662 18028 8668 18040
rect 8720 18028 8726 18080
rect 10410 18068 10416 18080
rect 10371 18040 10416 18068
rect 10410 18028 10416 18040
rect 10468 18028 10474 18080
rect 12253 18071 12311 18077
rect 12253 18037 12265 18071
rect 12299 18068 12311 18071
rect 12618 18068 12624 18080
rect 12299 18040 12624 18068
rect 12299 18037 12311 18040
rect 12253 18031 12311 18037
rect 12618 18028 12624 18040
rect 12676 18028 12682 18080
rect 12802 18068 12808 18080
rect 12763 18040 12808 18068
rect 12802 18028 12808 18040
rect 12860 18028 12866 18080
rect 14829 18071 14887 18077
rect 14829 18037 14841 18071
rect 14875 18068 14887 18071
rect 15120 18068 15148 18099
rect 16022 18096 16028 18108
rect 16080 18096 16086 18148
rect 19628 18136 19656 18167
rect 19794 18164 19800 18176
rect 19852 18164 19858 18216
rect 20257 18207 20315 18213
rect 20257 18173 20269 18207
rect 20303 18173 20315 18207
rect 20257 18167 20315 18173
rect 20272 18136 20300 18167
rect 19628 18108 20300 18136
rect 15746 18068 15752 18080
rect 14875 18040 15752 18068
rect 14875 18037 14887 18040
rect 14829 18031 14887 18037
rect 15746 18028 15752 18040
rect 15804 18068 15810 18080
rect 16206 18068 16212 18080
rect 15804 18040 16212 18068
rect 15804 18028 15810 18040
rect 16206 18028 16212 18040
rect 16264 18028 16270 18080
rect 16850 18028 16856 18080
rect 16908 18068 16914 18080
rect 16945 18071 17003 18077
rect 16945 18068 16957 18071
rect 16908 18040 16957 18068
rect 16908 18028 16914 18040
rect 16945 18037 16957 18040
rect 16991 18037 17003 18071
rect 17770 18068 17776 18080
rect 17731 18040 17776 18068
rect 16945 18031 17003 18037
rect 17770 18028 17776 18040
rect 17828 18028 17834 18080
rect 18417 18071 18475 18077
rect 18417 18037 18429 18071
rect 18463 18068 18475 18071
rect 18506 18068 18512 18080
rect 18463 18040 18512 18068
rect 18463 18037 18475 18040
rect 18417 18031 18475 18037
rect 18506 18028 18512 18040
rect 18564 18028 18570 18080
rect 19886 18068 19892 18080
rect 19847 18040 19892 18068
rect 19886 18028 19892 18040
rect 19944 18028 19950 18080
rect 1104 17978 22816 18000
rect 1104 17926 8982 17978
rect 9034 17926 9046 17978
rect 9098 17926 9110 17978
rect 9162 17926 9174 17978
rect 9226 17926 16982 17978
rect 17034 17926 17046 17978
rect 17098 17926 17110 17978
rect 17162 17926 17174 17978
rect 17226 17926 22816 17978
rect 1104 17904 22816 17926
rect 4706 17824 4712 17876
rect 4764 17864 4770 17876
rect 4985 17867 5043 17873
rect 4985 17864 4997 17867
rect 4764 17836 4997 17864
rect 4764 17824 4770 17836
rect 4985 17833 4997 17836
rect 5031 17833 5043 17867
rect 4985 17827 5043 17833
rect 6365 17867 6423 17873
rect 6365 17833 6377 17867
rect 6411 17864 6423 17867
rect 6914 17864 6920 17876
rect 6411 17836 6920 17864
rect 6411 17833 6423 17836
rect 6365 17827 6423 17833
rect 6914 17824 6920 17836
rect 6972 17864 6978 17876
rect 8343 17867 8401 17873
rect 8343 17864 8355 17867
rect 6972 17836 8355 17864
rect 6972 17824 6978 17836
rect 8343 17833 8355 17836
rect 8389 17833 8401 17867
rect 8343 17827 8401 17833
rect 8754 17824 8760 17876
rect 8812 17864 8818 17876
rect 8849 17867 8907 17873
rect 8849 17864 8861 17867
rect 8812 17836 8861 17864
rect 8812 17824 8818 17836
rect 8849 17833 8861 17836
rect 8895 17833 8907 17867
rect 11422 17864 11428 17876
rect 11383 17836 11428 17864
rect 8849 17827 8907 17833
rect 11422 17824 11428 17836
rect 11480 17824 11486 17876
rect 15010 17864 15016 17876
rect 14971 17836 15016 17864
rect 15010 17824 15016 17836
rect 15068 17824 15074 17876
rect 16206 17864 16212 17876
rect 16167 17836 16212 17864
rect 16206 17824 16212 17836
rect 16264 17824 16270 17876
rect 18690 17824 18696 17876
rect 18748 17864 18754 17876
rect 19337 17867 19395 17873
rect 19337 17864 19349 17867
rect 18748 17836 19349 17864
rect 18748 17824 18754 17836
rect 19337 17833 19349 17836
rect 19383 17833 19395 17867
rect 19337 17827 19395 17833
rect 21085 17867 21143 17873
rect 21085 17833 21097 17867
rect 21131 17864 21143 17867
rect 21266 17864 21272 17876
rect 21131 17836 21272 17864
rect 21131 17833 21143 17836
rect 21085 17827 21143 17833
rect 21266 17824 21272 17836
rect 21324 17824 21330 17876
rect 4154 17756 4160 17808
rect 4212 17796 4218 17808
rect 4386 17799 4444 17805
rect 4386 17796 4398 17799
rect 4212 17768 4398 17796
rect 4212 17756 4218 17768
rect 4386 17765 4398 17768
rect 4432 17765 4444 17799
rect 6730 17796 6736 17808
rect 6691 17768 6736 17796
rect 4386 17759 4444 17765
rect 6730 17756 6736 17768
rect 6788 17796 6794 17808
rect 8662 17796 8668 17808
rect 6788 17768 8668 17796
rect 6788 17756 6794 17768
rect 8662 17756 8668 17768
rect 8720 17756 8726 17808
rect 10042 17796 10048 17808
rect 10003 17768 10048 17796
rect 10042 17756 10048 17768
rect 10100 17756 10106 17808
rect 12526 17796 12532 17808
rect 12487 17768 12532 17796
rect 12526 17756 12532 17768
rect 12584 17756 12590 17808
rect 15286 17756 15292 17808
rect 15344 17796 15350 17808
rect 15610 17799 15668 17805
rect 15610 17796 15622 17799
rect 15344 17768 15622 17796
rect 15344 17756 15350 17768
rect 15610 17765 15622 17768
rect 15656 17796 15668 17799
rect 17770 17796 17776 17808
rect 15656 17768 17776 17796
rect 15656 17765 15668 17768
rect 15610 17759 15668 17765
rect 17770 17756 17776 17768
rect 17828 17796 17834 17808
rect 18506 17805 18512 17808
rect 18462 17799 18512 17805
rect 18462 17796 18474 17799
rect 17828 17768 18474 17796
rect 17828 17756 17834 17768
rect 18462 17765 18474 17768
rect 18508 17765 18512 17799
rect 18462 17759 18512 17765
rect 18506 17756 18512 17759
rect 18564 17756 18570 17808
rect 2590 17728 2596 17740
rect 2551 17700 2596 17728
rect 2590 17688 2596 17700
rect 2648 17688 2654 17740
rect 2866 17728 2872 17740
rect 2827 17700 2872 17728
rect 2866 17688 2872 17700
rect 2924 17688 2930 17740
rect 4706 17688 4712 17740
rect 4764 17728 4770 17740
rect 4982 17728 4988 17740
rect 4764 17700 4988 17728
rect 4764 17688 4770 17700
rect 4982 17688 4988 17700
rect 5040 17728 5046 17740
rect 5629 17731 5687 17737
rect 5629 17728 5641 17731
rect 5040 17700 5641 17728
rect 5040 17688 5046 17700
rect 5629 17697 5641 17700
rect 5675 17697 5687 17731
rect 6454 17728 6460 17740
rect 6415 17700 6460 17728
rect 5629 17691 5687 17697
rect 6454 17688 6460 17700
rect 6512 17688 6518 17740
rect 8272 17731 8330 17737
rect 8272 17697 8284 17731
rect 8318 17728 8330 17731
rect 8478 17728 8484 17740
rect 8318 17700 8484 17728
rect 8318 17697 8330 17700
rect 8272 17691 8330 17697
rect 8478 17688 8484 17700
rect 8536 17688 8542 17740
rect 11882 17728 11888 17740
rect 11843 17700 11888 17728
rect 11882 17688 11888 17700
rect 11940 17688 11946 17740
rect 12250 17728 12256 17740
rect 12211 17700 12256 17728
rect 12250 17688 12256 17700
rect 12308 17688 12314 17740
rect 13909 17731 13967 17737
rect 13909 17697 13921 17731
rect 13955 17728 13967 17731
rect 13998 17728 14004 17740
rect 13955 17700 14004 17728
rect 13955 17697 13967 17700
rect 13909 17691 13967 17697
rect 13998 17688 14004 17700
rect 14056 17688 14062 17740
rect 14182 17728 14188 17740
rect 14143 17700 14188 17728
rect 14182 17688 14188 17700
rect 14240 17688 14246 17740
rect 17037 17731 17095 17737
rect 17037 17697 17049 17731
rect 17083 17728 17095 17731
rect 17126 17728 17132 17740
rect 17083 17700 17132 17728
rect 17083 17697 17095 17700
rect 17037 17691 17095 17697
rect 17126 17688 17132 17700
rect 17184 17688 17190 17740
rect 17862 17688 17868 17740
rect 17920 17728 17926 17740
rect 18141 17731 18199 17737
rect 18141 17728 18153 17731
rect 17920 17700 18153 17728
rect 17920 17688 17926 17700
rect 18141 17697 18153 17700
rect 18187 17728 18199 17731
rect 19886 17728 19892 17740
rect 18187 17700 19892 17728
rect 18187 17697 18199 17700
rect 18141 17691 18199 17697
rect 19886 17688 19892 17700
rect 19944 17688 19950 17740
rect 20714 17688 20720 17740
rect 20772 17728 20778 17740
rect 20901 17731 20959 17737
rect 20901 17728 20913 17731
rect 20772 17700 20913 17728
rect 20772 17688 20778 17700
rect 20901 17697 20913 17700
rect 20947 17697 20959 17731
rect 20901 17691 20959 17697
rect 3142 17660 3148 17672
rect 3103 17632 3148 17660
rect 3142 17620 3148 17632
rect 3200 17660 3206 17672
rect 4065 17663 4123 17669
rect 4065 17660 4077 17663
rect 3200 17632 4077 17660
rect 3200 17620 3206 17632
rect 4065 17629 4077 17632
rect 4111 17629 4123 17663
rect 4065 17623 4123 17629
rect 9953 17663 10011 17669
rect 9953 17629 9965 17663
rect 9999 17660 10011 17663
rect 11146 17660 11152 17672
rect 9999 17632 11152 17660
rect 9999 17629 10011 17632
rect 9953 17623 10011 17629
rect 11146 17620 11152 17632
rect 11204 17620 11210 17672
rect 11900 17660 11928 17688
rect 14369 17663 14427 17669
rect 11900 17632 13814 17660
rect 10505 17595 10563 17601
rect 10505 17561 10517 17595
rect 10551 17592 10563 17595
rect 10594 17592 10600 17604
rect 10551 17564 10600 17592
rect 10551 17561 10563 17564
rect 10505 17555 10563 17561
rect 10594 17552 10600 17564
rect 10652 17552 10658 17604
rect 13262 17592 13268 17604
rect 13223 17564 13268 17592
rect 13262 17552 13268 17564
rect 13320 17552 13326 17604
rect 13786 17592 13814 17632
rect 14369 17629 14381 17663
rect 14415 17660 14427 17663
rect 15289 17663 15347 17669
rect 15289 17660 15301 17663
rect 14415 17632 15301 17660
rect 14415 17629 14427 17632
rect 14369 17623 14427 17629
rect 15289 17629 15301 17632
rect 15335 17660 15347 17663
rect 16482 17660 16488 17672
rect 15335 17632 16488 17660
rect 15335 17629 15347 17632
rect 15289 17623 15347 17629
rect 16482 17620 16488 17632
rect 16540 17620 16546 17672
rect 18046 17592 18052 17604
rect 13786 17564 18052 17592
rect 18046 17552 18052 17564
rect 18104 17592 18110 17604
rect 19794 17592 19800 17604
rect 18104 17564 19800 17592
rect 18104 17552 18110 17564
rect 19794 17552 19800 17564
rect 19852 17552 19858 17604
rect 5353 17527 5411 17533
rect 5353 17493 5365 17527
rect 5399 17524 5411 17527
rect 5442 17524 5448 17536
rect 5399 17496 5448 17524
rect 5399 17493 5411 17496
rect 5353 17487 5411 17493
rect 5442 17484 5448 17496
rect 5500 17524 5506 17536
rect 7006 17524 7012 17536
rect 5500 17496 7012 17524
rect 5500 17484 5506 17496
rect 7006 17484 7012 17496
rect 7064 17484 7070 17536
rect 7098 17484 7104 17536
rect 7156 17524 7162 17536
rect 7377 17527 7435 17533
rect 7377 17524 7389 17527
rect 7156 17496 7389 17524
rect 7156 17484 7162 17496
rect 7377 17493 7389 17496
rect 7423 17524 7435 17527
rect 7653 17527 7711 17533
rect 7653 17524 7665 17527
rect 7423 17496 7665 17524
rect 7423 17493 7435 17496
rect 7377 17487 7435 17493
rect 7653 17493 7665 17496
rect 7699 17493 7711 17527
rect 7653 17487 7711 17493
rect 8113 17527 8171 17533
rect 8113 17493 8125 17527
rect 8159 17524 8171 17527
rect 8294 17524 8300 17536
rect 8159 17496 8300 17524
rect 8159 17493 8171 17496
rect 8113 17487 8171 17493
rect 8294 17484 8300 17496
rect 8352 17484 8358 17536
rect 9582 17484 9588 17536
rect 9640 17524 9646 17536
rect 10686 17524 10692 17536
rect 9640 17496 10692 17524
rect 9640 17484 9646 17496
rect 10686 17484 10692 17496
rect 10744 17524 10750 17536
rect 10873 17527 10931 17533
rect 10873 17524 10885 17527
rect 10744 17496 10885 17524
rect 10744 17484 10750 17496
rect 10873 17493 10885 17496
rect 10919 17493 10931 17527
rect 12802 17524 12808 17536
rect 12763 17496 12808 17524
rect 10873 17487 10931 17493
rect 12802 17484 12808 17496
rect 12860 17484 12866 17536
rect 16574 17484 16580 17536
rect 16632 17524 16638 17536
rect 17175 17527 17233 17533
rect 17175 17524 17187 17527
rect 16632 17496 17187 17524
rect 16632 17484 16638 17496
rect 17175 17493 17187 17496
rect 17221 17493 17233 17527
rect 19058 17524 19064 17536
rect 19019 17496 19064 17524
rect 17175 17487 17233 17493
rect 19058 17484 19064 17496
rect 19116 17484 19122 17536
rect 1104 17434 22816 17456
rect 1104 17382 4982 17434
rect 5034 17382 5046 17434
rect 5098 17382 5110 17434
rect 5162 17382 5174 17434
rect 5226 17382 12982 17434
rect 13034 17382 13046 17434
rect 13098 17382 13110 17434
rect 13162 17382 13174 17434
rect 13226 17382 20982 17434
rect 21034 17382 21046 17434
rect 21098 17382 21110 17434
rect 21162 17382 21174 17434
rect 21226 17382 22816 17434
rect 1104 17360 22816 17382
rect 3142 17320 3148 17332
rect 3103 17292 3148 17320
rect 3142 17280 3148 17292
rect 3200 17280 3206 17332
rect 4798 17280 4804 17332
rect 4856 17320 4862 17332
rect 4985 17323 5043 17329
rect 4985 17320 4997 17323
rect 4856 17292 4997 17320
rect 4856 17280 4862 17292
rect 4985 17289 4997 17292
rect 5031 17289 5043 17323
rect 4985 17283 5043 17289
rect 6181 17323 6239 17329
rect 6181 17289 6193 17323
rect 6227 17320 6239 17323
rect 6454 17320 6460 17332
rect 6227 17292 6460 17320
rect 6227 17289 6239 17292
rect 6181 17283 6239 17289
rect 6454 17280 6460 17292
rect 6512 17280 6518 17332
rect 8202 17320 8208 17332
rect 8163 17292 8208 17320
rect 8202 17280 8208 17292
rect 8260 17320 8266 17332
rect 8478 17320 8484 17332
rect 8260 17292 8484 17320
rect 8260 17280 8266 17292
rect 8478 17280 8484 17292
rect 8536 17280 8542 17332
rect 8895 17323 8953 17329
rect 8895 17289 8907 17323
rect 8941 17320 8953 17323
rect 9582 17320 9588 17332
rect 8941 17292 9588 17320
rect 8941 17289 8953 17292
rect 8895 17283 8953 17289
rect 9582 17280 9588 17292
rect 9640 17280 9646 17332
rect 9677 17323 9735 17329
rect 9677 17289 9689 17323
rect 9723 17320 9735 17323
rect 10042 17320 10048 17332
rect 9723 17292 10048 17320
rect 9723 17289 9735 17292
rect 9677 17283 9735 17289
rect 10042 17280 10048 17292
rect 10100 17280 10106 17332
rect 11146 17320 11152 17332
rect 11107 17292 11152 17320
rect 11146 17280 11152 17292
rect 11204 17320 11210 17332
rect 11471 17323 11529 17329
rect 11471 17320 11483 17323
rect 11204 17292 11483 17320
rect 11204 17280 11210 17292
rect 11471 17289 11483 17292
rect 11517 17289 11529 17323
rect 11471 17283 11529 17289
rect 14415 17323 14473 17329
rect 14415 17289 14427 17323
rect 14461 17320 14473 17323
rect 15010 17320 15016 17332
rect 14461 17292 15016 17320
rect 14461 17289 14473 17292
rect 14415 17283 14473 17289
rect 15010 17280 15016 17292
rect 15068 17280 15074 17332
rect 16482 17320 16488 17332
rect 16443 17292 16488 17320
rect 16482 17280 16488 17292
rect 16540 17280 16546 17332
rect 17862 17320 17868 17332
rect 17823 17292 17868 17320
rect 17862 17280 17868 17292
rect 17920 17280 17926 17332
rect 21085 17323 21143 17329
rect 21085 17289 21097 17323
rect 21131 17320 21143 17323
rect 21266 17320 21272 17332
rect 21131 17292 21272 17320
rect 21131 17289 21143 17292
rect 21085 17283 21143 17289
rect 21266 17280 21272 17292
rect 21324 17280 21330 17332
rect 2590 17212 2596 17264
rect 2648 17252 2654 17264
rect 10410 17252 10416 17264
rect 2648 17224 10416 17252
rect 2648 17212 2654 17224
rect 10410 17212 10416 17224
rect 10468 17252 10474 17264
rect 10870 17252 10876 17264
rect 10468 17224 10876 17252
rect 10468 17212 10474 17224
rect 10870 17212 10876 17224
rect 10928 17212 10934 17264
rect 10962 17212 10968 17264
rect 11020 17252 11026 17264
rect 13354 17252 13360 17264
rect 11020 17224 12801 17252
rect 13315 17224 13360 17252
rect 11020 17212 11026 17224
rect 7101 17187 7159 17193
rect 7101 17153 7113 17187
rect 7147 17184 7159 17187
rect 7742 17184 7748 17196
rect 7147 17156 7748 17184
rect 7147 17153 7159 17156
rect 7101 17147 7159 17153
rect 7742 17144 7748 17156
rect 7800 17184 7806 17196
rect 8573 17187 8631 17193
rect 8573 17184 8585 17187
rect 7800 17156 8585 17184
rect 7800 17144 7806 17156
rect 8573 17153 8585 17156
rect 8619 17153 8631 17187
rect 8573 17147 8631 17153
rect 9950 17144 9956 17196
rect 10008 17184 10014 17196
rect 12773 17184 12801 17224
rect 13354 17212 13360 17224
rect 13412 17212 13418 17264
rect 15102 17212 15108 17264
rect 15160 17252 15166 17264
rect 17126 17252 17132 17264
rect 15160 17224 17132 17252
rect 15160 17212 15166 17224
rect 17126 17212 17132 17224
rect 17184 17252 17190 17264
rect 20530 17252 20536 17264
rect 17184 17224 20536 17252
rect 17184 17212 17190 17224
rect 20530 17212 20536 17224
rect 20588 17212 20594 17264
rect 15562 17184 15568 17196
rect 10008 17156 11411 17184
rect 12773 17156 13814 17184
rect 15523 17156 15568 17184
rect 10008 17144 10014 17156
rect 4065 17119 4123 17125
rect 4065 17085 4077 17119
rect 4111 17116 4123 17119
rect 8824 17119 8882 17125
rect 4111 17088 5304 17116
rect 4111 17085 4123 17088
rect 4065 17079 4123 17085
rect 2501 17051 2559 17057
rect 2501 17017 2513 17051
rect 2547 17048 2559 17051
rect 2866 17048 2872 17060
rect 2547 17020 2872 17048
rect 2547 17017 2559 17020
rect 2501 17011 2559 17017
rect 2866 17008 2872 17020
rect 2924 17008 2930 17060
rect 4386 17051 4444 17057
rect 4386 17048 4398 17051
rect 4172 17020 4398 17048
rect 4172 16992 4200 17020
rect 4386 17017 4398 17020
rect 4432 17017 4444 17051
rect 4386 17011 4444 17017
rect 5276 16992 5304 17088
rect 8824 17085 8836 17119
rect 8870 17116 8882 17119
rect 9306 17116 9312 17128
rect 8870 17088 9312 17116
rect 8870 17085 8882 17088
rect 8824 17079 8882 17085
rect 9306 17076 9312 17088
rect 9364 17076 9370 17128
rect 11383 17125 11411 17156
rect 11368 17119 11426 17125
rect 11368 17085 11380 17119
rect 11414 17116 11426 17119
rect 11790 17116 11796 17128
rect 11414 17088 11796 17116
rect 11414 17085 11426 17088
rect 11368 17079 11426 17085
rect 11790 17076 11796 17088
rect 11848 17076 11854 17128
rect 13786 17116 13814 17156
rect 15562 17144 15568 17156
rect 15620 17144 15626 17196
rect 17770 17144 17776 17196
rect 17828 17184 17834 17196
rect 18233 17187 18291 17193
rect 18233 17184 18245 17187
rect 17828 17156 18245 17184
rect 17828 17144 17834 17156
rect 18233 17153 18245 17156
rect 18279 17153 18291 17187
rect 18233 17147 18291 17153
rect 18877 17187 18935 17193
rect 18877 17153 18889 17187
rect 18923 17184 18935 17187
rect 18966 17184 18972 17196
rect 18923 17156 18972 17184
rect 18923 17153 18935 17156
rect 18877 17147 18935 17153
rect 18966 17144 18972 17156
rect 19024 17144 19030 17196
rect 19242 17184 19248 17196
rect 19203 17156 19248 17184
rect 19242 17144 19248 17156
rect 19300 17144 19306 17196
rect 14344 17119 14402 17125
rect 14344 17116 14356 17119
rect 13786 17088 14356 17116
rect 14344 17085 14356 17088
rect 14390 17116 14402 17119
rect 14737 17119 14795 17125
rect 14737 17116 14749 17119
rect 14390 17088 14749 17116
rect 14390 17085 14402 17088
rect 14344 17079 14402 17085
rect 14737 17085 14749 17088
rect 14783 17085 14795 17119
rect 14737 17079 14795 17085
rect 19518 17076 19524 17128
rect 19576 17116 19582 17128
rect 20901 17119 20959 17125
rect 20901 17116 20913 17119
rect 19576 17088 20913 17116
rect 19576 17076 19582 17088
rect 20901 17085 20913 17088
rect 20947 17116 20959 17119
rect 21453 17119 21511 17125
rect 21453 17116 21465 17119
rect 20947 17088 21465 17116
rect 20947 17085 20959 17088
rect 20901 17079 20959 17085
rect 21453 17085 21465 17088
rect 21499 17085 21511 17119
rect 21453 17079 21511 17085
rect 7098 17008 7104 17060
rect 7156 17048 7162 17060
rect 7193 17051 7251 17057
rect 7193 17048 7205 17051
rect 7156 17020 7205 17048
rect 7156 17008 7162 17020
rect 7193 17017 7205 17020
rect 7239 17017 7251 17051
rect 7193 17011 7251 17017
rect 7282 17008 7288 17060
rect 7340 17048 7346 17060
rect 7745 17051 7803 17057
rect 7745 17048 7757 17051
rect 7340 17020 7757 17048
rect 7340 17008 7346 17020
rect 7745 17017 7757 17020
rect 7791 17017 7803 17051
rect 7745 17011 7803 17017
rect 9490 17008 9496 17060
rect 9548 17048 9554 17060
rect 9861 17051 9919 17057
rect 9861 17048 9873 17051
rect 9548 17020 9873 17048
rect 9548 17008 9554 17020
rect 9861 17017 9873 17020
rect 9907 17017 9919 17051
rect 9861 17011 9919 17017
rect 9953 17051 10011 17057
rect 9953 17017 9965 17051
rect 9999 17017 10011 17051
rect 9953 17011 10011 17017
rect 10505 17051 10563 17057
rect 10505 17017 10517 17051
rect 10551 17048 10563 17051
rect 10594 17048 10600 17060
rect 10551 17020 10600 17048
rect 10551 17017 10563 17020
rect 10505 17011 10563 17017
rect 2590 16940 2596 16992
rect 2648 16980 2654 16992
rect 2777 16983 2835 16989
rect 2777 16980 2789 16983
rect 2648 16952 2789 16980
rect 2648 16940 2654 16952
rect 2777 16949 2789 16952
rect 2823 16949 2835 16983
rect 2777 16943 2835 16949
rect 3605 16983 3663 16989
rect 3605 16949 3617 16983
rect 3651 16980 3663 16983
rect 3881 16983 3939 16989
rect 3881 16980 3893 16983
rect 3651 16952 3893 16980
rect 3651 16949 3663 16952
rect 3605 16943 3663 16949
rect 3881 16949 3893 16952
rect 3927 16980 3939 16983
rect 4154 16980 4160 16992
rect 3927 16952 4160 16980
rect 3927 16949 3939 16952
rect 3881 16943 3939 16949
rect 4154 16940 4160 16952
rect 4212 16940 4218 16992
rect 5258 16980 5264 16992
rect 5219 16952 5264 16980
rect 5258 16940 5264 16952
rect 5316 16940 5322 16992
rect 5810 16940 5816 16992
rect 5868 16980 5874 16992
rect 6457 16983 6515 16989
rect 6457 16980 6469 16983
rect 5868 16952 6469 16980
rect 5868 16940 5874 16952
rect 6457 16949 6469 16952
rect 6503 16980 6515 16983
rect 6730 16980 6736 16992
rect 6503 16952 6736 16980
rect 6503 16949 6515 16952
rect 6457 16943 6515 16949
rect 6730 16940 6736 16952
rect 6788 16940 6794 16992
rect 9306 16980 9312 16992
rect 9267 16952 9312 16980
rect 9306 16940 9312 16952
rect 9364 16940 9370 16992
rect 9968 16980 9996 17011
rect 10594 17008 10600 17020
rect 10652 17008 10658 17060
rect 12434 17008 12440 17060
rect 12492 17048 12498 17060
rect 12802 17048 12808 17060
rect 12492 17020 12808 17048
rect 12492 17008 12498 17020
rect 12802 17008 12808 17020
rect 12860 17008 12866 17060
rect 12897 17051 12955 17057
rect 12897 17017 12909 17051
rect 12943 17048 12955 17051
rect 13262 17048 13268 17060
rect 12943 17020 13268 17048
rect 12943 17017 12955 17020
rect 12897 17011 12955 17017
rect 13262 17008 13268 17020
rect 13320 17008 13326 17060
rect 13817 17051 13875 17057
rect 13817 17017 13829 17051
rect 13863 17048 13875 17051
rect 13998 17048 14004 17060
rect 13863 17020 14004 17048
rect 13863 17017 13875 17020
rect 13817 17011 13875 17017
rect 13998 17008 14004 17020
rect 14056 17048 14062 17060
rect 14182 17048 14188 17060
rect 14056 17020 14188 17048
rect 14056 17008 14062 17020
rect 14182 17008 14188 17020
rect 14240 17008 14246 17060
rect 15657 17051 15715 17057
rect 15657 17017 15669 17051
rect 15703 17048 15715 17051
rect 15746 17048 15752 17060
rect 15703 17020 15752 17048
rect 15703 17017 15715 17020
rect 15657 17011 15715 17017
rect 15746 17008 15752 17020
rect 15804 17008 15810 17060
rect 16206 17048 16212 17060
rect 16167 17020 16212 17048
rect 16206 17008 16212 17020
rect 16264 17008 16270 17060
rect 18969 17051 19027 17057
rect 18969 17017 18981 17051
rect 19015 17048 19027 17051
rect 19058 17048 19064 17060
rect 19015 17020 19064 17048
rect 19015 17017 19027 17020
rect 18969 17011 19027 17017
rect 10134 16980 10140 16992
rect 9968 16952 10140 16980
rect 10134 16940 10140 16952
rect 10192 16980 10198 16992
rect 10781 16983 10839 16989
rect 10781 16980 10793 16983
rect 10192 16952 10793 16980
rect 10192 16940 10198 16952
rect 10781 16949 10793 16952
rect 10827 16949 10839 16983
rect 12250 16980 12256 16992
rect 12211 16952 12256 16980
rect 10781 16943 10839 16949
rect 12250 16940 12256 16952
rect 12308 16940 12314 16992
rect 14090 16980 14096 16992
rect 14051 16952 14096 16980
rect 14090 16940 14096 16952
rect 14148 16940 14154 16992
rect 15286 16980 15292 16992
rect 15247 16952 15292 16980
rect 15286 16940 15292 16952
rect 15344 16940 15350 16992
rect 18693 16983 18751 16989
rect 18693 16949 18705 16983
rect 18739 16980 18751 16983
rect 18984 16980 19012 17011
rect 19058 17008 19064 17020
rect 19116 17008 19122 17060
rect 20714 16980 20720 16992
rect 18739 16952 19012 16980
rect 20675 16952 20720 16980
rect 18739 16949 18751 16952
rect 18693 16943 18751 16949
rect 20714 16940 20720 16952
rect 20772 16940 20778 16992
rect 1104 16890 22816 16912
rect 1104 16838 8982 16890
rect 9034 16838 9046 16890
rect 9098 16838 9110 16890
rect 9162 16838 9174 16890
rect 9226 16838 16982 16890
rect 17034 16838 17046 16890
rect 17098 16838 17110 16890
rect 17162 16838 17174 16890
rect 17226 16838 22816 16890
rect 1104 16816 22816 16838
rect 7098 16776 7104 16788
rect 7059 16748 7104 16776
rect 7098 16736 7104 16748
rect 7156 16736 7162 16788
rect 12710 16776 12716 16788
rect 12671 16748 12716 16776
rect 12710 16736 12716 16748
rect 12768 16736 12774 16788
rect 13262 16776 13268 16788
rect 13223 16748 13268 16776
rect 13262 16736 13268 16748
rect 13320 16736 13326 16788
rect 15105 16779 15163 16785
rect 15105 16745 15117 16779
rect 15151 16776 15163 16779
rect 15562 16776 15568 16788
rect 15151 16748 15568 16776
rect 15151 16745 15163 16748
rect 15105 16739 15163 16745
rect 15562 16736 15568 16748
rect 15620 16736 15626 16788
rect 4801 16711 4859 16717
rect 4801 16677 4813 16711
rect 4847 16708 4859 16711
rect 5258 16708 5264 16720
rect 4847 16680 5264 16708
rect 4847 16677 4859 16680
rect 4801 16671 4859 16677
rect 5258 16668 5264 16680
rect 5316 16668 5322 16720
rect 7607 16711 7665 16717
rect 7607 16677 7619 16711
rect 7653 16708 7665 16711
rect 7742 16708 7748 16720
rect 7653 16680 7748 16708
rect 7653 16677 7665 16680
rect 7607 16671 7665 16677
rect 7742 16668 7748 16680
rect 7800 16668 7806 16720
rect 10134 16708 10140 16720
rect 10095 16680 10140 16708
rect 10134 16668 10140 16680
rect 10192 16668 10198 16720
rect 10689 16711 10747 16717
rect 10689 16677 10701 16711
rect 10735 16708 10747 16711
rect 10962 16708 10968 16720
rect 10735 16680 10968 16708
rect 10735 16677 10747 16680
rect 10689 16671 10747 16677
rect 10962 16668 10968 16680
rect 11020 16708 11026 16720
rect 11422 16708 11428 16720
rect 11020 16680 11428 16708
rect 11020 16668 11026 16680
rect 11422 16668 11428 16680
rect 11480 16668 11486 16720
rect 15838 16708 15844 16720
rect 15799 16680 15844 16708
rect 15838 16668 15844 16680
rect 15896 16668 15902 16720
rect 18322 16708 18328 16720
rect 18283 16680 18328 16708
rect 18322 16668 18328 16680
rect 18380 16668 18386 16720
rect 4246 16640 4252 16652
rect 4207 16612 4252 16640
rect 4246 16600 4252 16612
rect 4304 16600 4310 16652
rect 4614 16640 4620 16652
rect 4575 16612 4620 16640
rect 4614 16600 4620 16612
rect 4672 16600 4678 16652
rect 7520 16643 7578 16649
rect 7520 16609 7532 16643
rect 7566 16640 7578 16643
rect 7926 16640 7932 16652
rect 7566 16612 7932 16640
rect 7566 16609 7578 16612
rect 7520 16603 7578 16609
rect 7926 16600 7932 16612
rect 7984 16600 7990 16652
rect 8386 16600 8392 16652
rect 8444 16640 8450 16652
rect 8608 16643 8666 16649
rect 8608 16640 8620 16643
rect 8444 16612 8620 16640
rect 8444 16600 8450 16612
rect 8608 16609 8620 16612
rect 8654 16609 8666 16643
rect 8608 16603 8666 16609
rect 13906 16600 13912 16652
rect 13964 16640 13970 16652
rect 14128 16643 14186 16649
rect 14128 16640 14140 16643
rect 13964 16612 14140 16640
rect 13964 16600 13970 16612
rect 14128 16609 14140 16612
rect 14174 16609 14186 16643
rect 14128 16603 14186 16609
rect 6362 16572 6368 16584
rect 6323 16544 6368 16572
rect 6362 16532 6368 16544
rect 6420 16532 6426 16584
rect 8711 16575 8769 16581
rect 8711 16541 8723 16575
rect 8757 16572 8769 16575
rect 10042 16572 10048 16584
rect 8757 16544 10048 16572
rect 8757 16541 8769 16544
rect 8711 16535 8769 16541
rect 10042 16532 10048 16544
rect 10100 16532 10106 16584
rect 12342 16572 12348 16584
rect 12303 16544 12348 16572
rect 12342 16532 12348 16544
rect 12400 16532 12406 16584
rect 15749 16575 15807 16581
rect 15749 16541 15761 16575
rect 15795 16572 15807 16575
rect 16574 16572 16580 16584
rect 15795 16544 16580 16572
rect 15795 16541 15807 16544
rect 15749 16535 15807 16541
rect 16574 16532 16580 16544
rect 16632 16532 16638 16584
rect 18230 16572 18236 16584
rect 18191 16544 18236 16572
rect 18230 16532 18236 16544
rect 18288 16532 18294 16584
rect 16206 16464 16212 16516
rect 16264 16504 16270 16516
rect 16301 16507 16359 16513
rect 16301 16504 16313 16507
rect 16264 16476 16313 16504
rect 16264 16464 16270 16476
rect 16301 16473 16313 16476
rect 16347 16504 16359 16507
rect 18690 16504 18696 16516
rect 16347 16476 18696 16504
rect 16347 16473 16359 16476
rect 16301 16467 16359 16473
rect 18690 16464 18696 16476
rect 18748 16464 18754 16516
rect 18785 16507 18843 16513
rect 18785 16473 18797 16507
rect 18831 16504 18843 16507
rect 18966 16504 18972 16516
rect 18831 16476 18972 16504
rect 18831 16473 18843 16476
rect 18785 16467 18843 16473
rect 4430 16396 4436 16448
rect 4488 16436 4494 16448
rect 5077 16439 5135 16445
rect 5077 16436 5089 16439
rect 4488 16408 5089 16436
rect 4488 16396 4494 16408
rect 5077 16405 5089 16408
rect 5123 16405 5135 16439
rect 5077 16399 5135 16405
rect 6178 16396 6184 16448
rect 6236 16436 6242 16448
rect 6595 16439 6653 16445
rect 6595 16436 6607 16439
rect 6236 16408 6607 16436
rect 6236 16396 6242 16408
rect 6595 16405 6607 16408
rect 6641 16405 6653 16439
rect 9030 16436 9036 16448
rect 8991 16408 9036 16436
rect 6595 16399 6653 16405
rect 9030 16396 9036 16408
rect 9088 16396 9094 16448
rect 9490 16436 9496 16448
rect 9451 16408 9496 16436
rect 9490 16396 9496 16408
rect 9548 16396 9554 16448
rect 10502 16396 10508 16448
rect 10560 16436 10566 16448
rect 10965 16439 11023 16445
rect 10965 16436 10977 16439
rect 10560 16408 10977 16436
rect 10560 16396 10566 16408
rect 10965 16405 10977 16408
rect 11011 16405 11023 16439
rect 11790 16436 11796 16448
rect 11751 16408 11796 16436
rect 10965 16399 11023 16405
rect 11790 16396 11796 16408
rect 11848 16396 11854 16448
rect 14231 16439 14289 16445
rect 14231 16405 14243 16439
rect 14277 16436 14289 16439
rect 15194 16436 15200 16448
rect 14277 16408 15200 16436
rect 14277 16405 14289 16408
rect 14231 16399 14289 16405
rect 15194 16396 15200 16408
rect 15252 16396 15258 16448
rect 15565 16439 15623 16445
rect 15565 16405 15577 16439
rect 15611 16436 15623 16439
rect 15746 16436 15752 16448
rect 15611 16408 15752 16436
rect 15611 16405 15623 16408
rect 15565 16399 15623 16405
rect 15746 16396 15752 16408
rect 15804 16396 15810 16448
rect 16022 16396 16028 16448
rect 16080 16436 16086 16448
rect 18800 16436 18828 16467
rect 18966 16464 18972 16476
rect 19024 16504 19030 16516
rect 19153 16507 19211 16513
rect 19153 16504 19165 16507
rect 19024 16476 19165 16504
rect 19024 16464 19030 16476
rect 19153 16473 19165 16476
rect 19199 16473 19211 16507
rect 19153 16467 19211 16473
rect 16080 16408 18828 16436
rect 16080 16396 16086 16408
rect 1104 16346 22816 16368
rect 1104 16294 4982 16346
rect 5034 16294 5046 16346
rect 5098 16294 5110 16346
rect 5162 16294 5174 16346
rect 5226 16294 12982 16346
rect 13034 16294 13046 16346
rect 13098 16294 13110 16346
rect 13162 16294 13174 16346
rect 13226 16294 20982 16346
rect 21034 16294 21046 16346
rect 21098 16294 21110 16346
rect 21162 16294 21174 16346
rect 21226 16294 22816 16346
rect 1104 16272 22816 16294
rect 6178 16232 6184 16244
rect 6139 16204 6184 16232
rect 6178 16192 6184 16204
rect 6236 16192 6242 16244
rect 6362 16192 6368 16244
rect 6420 16232 6426 16244
rect 6549 16235 6607 16241
rect 6549 16232 6561 16235
rect 6420 16204 6561 16232
rect 6420 16192 6426 16204
rect 6549 16201 6561 16204
rect 6595 16232 6607 16235
rect 6730 16232 6736 16244
rect 6595 16204 6736 16232
rect 6595 16201 6607 16204
rect 6549 16195 6607 16201
rect 6730 16192 6736 16204
rect 6788 16232 6794 16244
rect 9306 16232 9312 16244
rect 6788 16204 9312 16232
rect 6788 16192 6794 16204
rect 9306 16192 9312 16204
rect 9364 16192 9370 16244
rect 9493 16235 9551 16241
rect 9493 16201 9505 16235
rect 9539 16232 9551 16235
rect 10045 16235 10103 16241
rect 10045 16232 10057 16235
rect 9539 16204 10057 16232
rect 9539 16201 9551 16204
rect 9493 16195 9551 16201
rect 10045 16201 10057 16204
rect 10091 16232 10103 16235
rect 10134 16232 10140 16244
rect 10091 16204 10140 16232
rect 10091 16201 10103 16204
rect 10045 16195 10103 16201
rect 10134 16192 10140 16204
rect 10192 16192 10198 16244
rect 10318 16192 10324 16244
rect 10376 16232 10382 16244
rect 13814 16232 13820 16244
rect 10376 16204 13820 16232
rect 10376 16192 10382 16204
rect 13814 16192 13820 16204
rect 13872 16192 13878 16244
rect 13906 16192 13912 16244
rect 13964 16232 13970 16244
rect 14093 16235 14151 16241
rect 14093 16232 14105 16235
rect 13964 16204 14105 16232
rect 13964 16192 13970 16204
rect 14093 16201 14105 16204
rect 14139 16201 14151 16235
rect 14093 16195 14151 16201
rect 16485 16235 16543 16241
rect 16485 16201 16497 16235
rect 16531 16232 16543 16235
rect 16574 16232 16580 16244
rect 16531 16204 16580 16232
rect 16531 16201 16543 16204
rect 16485 16195 16543 16201
rect 16574 16192 16580 16204
rect 16632 16192 16638 16244
rect 18230 16192 18236 16244
rect 18288 16232 18294 16244
rect 19242 16232 19248 16244
rect 18288 16204 19248 16232
rect 18288 16192 18294 16204
rect 19242 16192 19248 16204
rect 19300 16232 19306 16244
rect 19429 16235 19487 16241
rect 19429 16232 19441 16235
rect 19300 16204 19441 16232
rect 19300 16192 19306 16204
rect 19429 16201 19441 16204
rect 19475 16201 19487 16235
rect 19429 16195 19487 16201
rect 2866 16124 2872 16176
rect 2924 16164 2930 16176
rect 4249 16167 4307 16173
rect 4249 16164 4261 16167
rect 2924 16136 4261 16164
rect 2924 16124 2930 16136
rect 4249 16133 4261 16136
rect 4295 16164 4307 16167
rect 4614 16164 4620 16176
rect 4295 16136 4620 16164
rect 4295 16133 4307 16136
rect 4249 16127 4307 16133
rect 4614 16124 4620 16136
rect 4672 16164 4678 16176
rect 5350 16164 5356 16176
rect 4672 16136 5356 16164
rect 4672 16124 4678 16136
rect 5350 16124 5356 16136
rect 5408 16124 5414 16176
rect 3467 16099 3525 16105
rect 3467 16065 3479 16099
rect 3513 16096 3525 16099
rect 4430 16096 4436 16108
rect 3513 16068 4436 16096
rect 3513 16065 3525 16068
rect 3467 16059 3525 16065
rect 4430 16056 4436 16068
rect 4488 16056 4494 16108
rect 4706 16096 4712 16108
rect 4667 16068 4712 16096
rect 4706 16056 4712 16068
rect 4764 16096 4770 16108
rect 6196 16096 6224 16192
rect 6641 16167 6699 16173
rect 6641 16133 6653 16167
rect 6687 16164 6699 16167
rect 7282 16164 7288 16176
rect 6687 16136 7288 16164
rect 6687 16133 6699 16136
rect 6641 16127 6699 16133
rect 7208 16105 7236 16136
rect 7282 16124 7288 16136
rect 7340 16124 7346 16176
rect 7650 16124 7656 16176
rect 7708 16164 7714 16176
rect 10962 16164 10968 16176
rect 7708 16136 10317 16164
rect 10923 16136 10968 16164
rect 7708 16124 7714 16136
rect 6917 16099 6975 16105
rect 6917 16096 6929 16099
rect 4764 16068 6132 16096
rect 6196 16068 6929 16096
rect 4764 16056 4770 16068
rect 3380 16031 3438 16037
rect 3380 15997 3392 16031
rect 3426 16028 3438 16031
rect 3786 16028 3792 16040
rect 3426 16000 3792 16028
rect 3426 15997 3438 16000
rect 3380 15991 3438 15997
rect 3786 15988 3792 16000
rect 3844 15988 3850 16040
rect 6104 16028 6132 16068
rect 6917 16065 6929 16068
rect 6963 16065 6975 16099
rect 6917 16059 6975 16065
rect 7193 16099 7251 16105
rect 7193 16065 7205 16099
rect 7239 16065 7251 16099
rect 7193 16059 7251 16065
rect 8573 16099 8631 16105
rect 8573 16065 8585 16099
rect 8619 16096 8631 16099
rect 8662 16096 8668 16108
rect 8619 16068 8668 16096
rect 8619 16065 8631 16068
rect 8573 16059 8631 16065
rect 8662 16056 8668 16068
rect 8720 16096 8726 16108
rect 9030 16096 9036 16108
rect 8720 16068 9036 16096
rect 8720 16056 8726 16068
rect 9030 16056 9036 16068
rect 9088 16056 9094 16108
rect 10289 16096 10317 16136
rect 10962 16124 10968 16136
rect 11020 16124 11026 16176
rect 18690 16164 18696 16176
rect 18651 16136 18696 16164
rect 18690 16124 18696 16136
rect 18748 16124 18754 16176
rect 11793 16099 11851 16105
rect 11793 16096 11805 16099
rect 10289 16068 11805 16096
rect 11793 16065 11805 16068
rect 11839 16065 11851 16099
rect 11793 16059 11851 16065
rect 12069 16099 12127 16105
rect 12069 16065 12081 16099
rect 12115 16096 12127 16099
rect 12710 16096 12716 16108
rect 12115 16068 12716 16096
rect 12115 16065 12127 16068
rect 12069 16059 12127 16065
rect 6641 16031 6699 16037
rect 6641 16028 6653 16031
rect 6104 16000 6653 16028
rect 6641 15997 6653 16000
rect 6687 15997 6699 16031
rect 11808 16028 11836 16059
rect 12710 16056 12716 16068
rect 12768 16096 12774 16108
rect 14645 16099 14703 16105
rect 14645 16096 14657 16099
rect 12768 16068 14657 16096
rect 12768 16056 12774 16068
rect 14645 16065 14657 16068
rect 14691 16065 14703 16099
rect 14645 16059 14703 16065
rect 17083 16099 17141 16105
rect 17083 16065 17095 16099
rect 17129 16096 17141 16099
rect 18141 16099 18199 16105
rect 18141 16096 18153 16099
rect 17129 16068 18153 16096
rect 17129 16065 17141 16068
rect 17083 16059 17141 16065
rect 18141 16065 18153 16068
rect 18187 16096 18199 16099
rect 19061 16099 19119 16105
rect 19061 16096 19073 16099
rect 18187 16068 19073 16096
rect 18187 16065 18199 16068
rect 18141 16059 18199 16065
rect 19061 16065 19073 16068
rect 19107 16065 19119 16099
rect 19061 16059 19119 16065
rect 12437 16031 12495 16037
rect 12437 16028 12449 16031
rect 11808 16000 12449 16028
rect 6641 15991 6699 15997
rect 12437 15997 12449 16000
rect 12483 16028 12495 16031
rect 12526 16028 12532 16040
rect 12483 16000 12532 16028
rect 12483 15997 12495 16000
rect 12437 15991 12495 15997
rect 12526 15988 12532 16000
rect 12584 15988 12590 16040
rect 12989 16031 13047 16037
rect 12989 15997 13001 16031
rect 13035 16028 13047 16031
rect 13262 16028 13268 16040
rect 13035 16000 13268 16028
rect 13035 15997 13047 16000
rect 12989 15991 13047 15997
rect 13262 15988 13268 16000
rect 13320 15988 13326 16040
rect 3237 15963 3295 15969
rect 3237 15929 3249 15963
rect 3283 15960 3295 15963
rect 4246 15960 4252 15972
rect 3283 15932 4252 15960
rect 3283 15929 3295 15932
rect 3237 15923 3295 15929
rect 4246 15920 4252 15932
rect 4304 15920 4310 15972
rect 4522 15960 4528 15972
rect 4483 15932 4528 15960
rect 4522 15920 4528 15932
rect 4580 15920 4586 15972
rect 7006 15960 7012 15972
rect 6967 15932 7012 15960
rect 7006 15920 7012 15932
rect 7064 15920 7070 15972
rect 8754 15920 8760 15972
rect 8812 15960 8818 15972
rect 8894 15963 8952 15969
rect 8894 15960 8906 15963
rect 8812 15932 8906 15960
rect 8812 15920 8818 15932
rect 8894 15929 8906 15932
rect 8940 15929 8952 15963
rect 10410 15960 10416 15972
rect 10371 15932 10416 15960
rect 8894 15923 8952 15929
rect 10410 15920 10416 15932
rect 10468 15920 10474 15972
rect 10502 15920 10508 15972
rect 10560 15960 10566 15972
rect 11517 15963 11575 15969
rect 10560 15932 10605 15960
rect 10560 15920 10566 15932
rect 11517 15929 11529 15963
rect 11563 15960 11575 15963
rect 14660 15960 14688 16059
rect 14826 16028 14832 16040
rect 14787 16000 14832 16028
rect 14826 15988 14832 16000
rect 14884 15988 14890 16040
rect 16996 16031 17054 16037
rect 16996 15997 17008 16031
rect 17042 16028 17054 16031
rect 17042 16000 17540 16028
rect 17042 15997 17054 16000
rect 16996 15991 17054 15997
rect 15150 15963 15208 15969
rect 15150 15960 15162 15963
rect 11563 15932 12388 15960
rect 14660 15932 15162 15960
rect 11563 15929 11575 15932
rect 11517 15923 11575 15929
rect 12360 15904 12388 15932
rect 15150 15929 15162 15932
rect 15196 15960 15208 15963
rect 15286 15960 15292 15972
rect 15196 15932 15292 15960
rect 15196 15929 15208 15932
rect 15150 15923 15208 15929
rect 15286 15920 15292 15932
rect 15344 15920 15350 15972
rect 3786 15892 3792 15904
rect 3747 15864 3792 15892
rect 3786 15852 3792 15864
rect 3844 15852 3850 15904
rect 4982 15852 4988 15904
rect 5040 15892 5046 15904
rect 5353 15895 5411 15901
rect 5353 15892 5365 15895
rect 5040 15864 5365 15892
rect 5040 15852 5046 15864
rect 5353 15861 5365 15864
rect 5399 15861 5411 15895
rect 7926 15892 7932 15904
rect 7887 15864 7932 15892
rect 5353 15855 5411 15861
rect 7926 15852 7932 15864
rect 7984 15852 7990 15904
rect 8386 15892 8392 15904
rect 8347 15864 8392 15892
rect 8386 15852 8392 15864
rect 8444 15852 8450 15904
rect 11606 15852 11612 15904
rect 11664 15892 11670 15904
rect 12069 15895 12127 15901
rect 12069 15892 12081 15895
rect 11664 15864 12081 15892
rect 11664 15852 11670 15864
rect 12069 15861 12081 15864
rect 12115 15892 12127 15895
rect 12161 15895 12219 15901
rect 12161 15892 12173 15895
rect 12115 15864 12173 15892
rect 12115 15861 12127 15864
rect 12069 15855 12127 15861
rect 12161 15861 12173 15864
rect 12207 15861 12219 15895
rect 12161 15855 12219 15861
rect 12342 15852 12348 15904
rect 12400 15892 12406 15904
rect 12529 15895 12587 15901
rect 12529 15892 12541 15895
rect 12400 15864 12541 15892
rect 12400 15852 12406 15864
rect 12529 15861 12541 15864
rect 12575 15861 12587 15895
rect 12529 15855 12587 15861
rect 15378 15852 15384 15904
rect 15436 15892 15442 15904
rect 15749 15895 15807 15901
rect 15749 15892 15761 15895
rect 15436 15864 15761 15892
rect 15436 15852 15442 15864
rect 15749 15861 15761 15864
rect 15795 15892 15807 15895
rect 15838 15892 15844 15904
rect 15795 15864 15844 15892
rect 15795 15861 15807 15864
rect 15749 15855 15807 15861
rect 15838 15852 15844 15864
rect 15896 15892 15902 15904
rect 17512 15901 17540 16000
rect 17865 15963 17923 15969
rect 17865 15929 17877 15963
rect 17911 15960 17923 15963
rect 18233 15963 18291 15969
rect 18233 15960 18245 15963
rect 17911 15932 18245 15960
rect 17911 15929 17923 15932
rect 17865 15923 17923 15929
rect 18233 15929 18245 15932
rect 18279 15960 18291 15963
rect 18322 15960 18328 15972
rect 18279 15932 18328 15960
rect 18279 15929 18291 15932
rect 18233 15923 18291 15929
rect 18322 15920 18328 15932
rect 18380 15920 18386 15972
rect 16025 15895 16083 15901
rect 16025 15892 16037 15895
rect 15896 15864 16037 15892
rect 15896 15852 15902 15864
rect 16025 15861 16037 15864
rect 16071 15861 16083 15895
rect 16025 15855 16083 15861
rect 17497 15895 17555 15901
rect 17497 15861 17509 15895
rect 17543 15892 17555 15895
rect 18138 15892 18144 15904
rect 17543 15864 18144 15892
rect 17543 15861 17555 15864
rect 17497 15855 17555 15861
rect 18138 15852 18144 15864
rect 18196 15892 18202 15904
rect 19518 15892 19524 15904
rect 18196 15864 19524 15892
rect 18196 15852 18202 15864
rect 19518 15852 19524 15864
rect 19576 15852 19582 15904
rect 19978 15892 19984 15904
rect 19939 15864 19984 15892
rect 19978 15852 19984 15864
rect 20036 15852 20042 15904
rect 1104 15802 22816 15824
rect 1104 15750 8982 15802
rect 9034 15750 9046 15802
rect 9098 15750 9110 15802
rect 9162 15750 9174 15802
rect 9226 15750 16982 15802
rect 17034 15750 17046 15802
rect 17098 15750 17110 15802
rect 17162 15750 17174 15802
rect 17226 15750 22816 15802
rect 1104 15728 22816 15750
rect 4154 15648 4160 15700
rect 4212 15688 4218 15700
rect 4212 15660 4429 15688
rect 4212 15648 4218 15660
rect 2774 15620 2780 15632
rect 2687 15592 2780 15620
rect 2700 15561 2728 15592
rect 2774 15580 2780 15592
rect 2832 15620 2838 15632
rect 4401 15629 4429 15660
rect 4522 15648 4528 15700
rect 4580 15688 4586 15700
rect 4982 15688 4988 15700
rect 4580 15660 4988 15688
rect 4580 15648 4586 15660
rect 4982 15648 4988 15660
rect 5040 15648 5046 15700
rect 6733 15691 6791 15697
rect 6733 15657 6745 15691
rect 6779 15688 6791 15691
rect 7006 15688 7012 15700
rect 6779 15660 7012 15688
rect 6779 15657 6791 15660
rect 6733 15651 6791 15657
rect 7006 15648 7012 15660
rect 7064 15648 7070 15700
rect 8754 15648 8760 15700
rect 8812 15688 8818 15700
rect 8941 15691 8999 15697
rect 8941 15688 8953 15691
rect 8812 15660 8953 15688
rect 8812 15648 8818 15660
rect 8941 15657 8953 15660
rect 8987 15688 8999 15691
rect 10042 15688 10048 15700
rect 8987 15660 9674 15688
rect 10003 15660 10048 15688
rect 8987 15657 8999 15660
rect 8941 15651 8999 15657
rect 4386 15623 4444 15629
rect 2832 15592 4154 15620
rect 2832 15580 2838 15592
rect 2685 15555 2743 15561
rect 2685 15521 2697 15555
rect 2731 15521 2743 15555
rect 2866 15552 2872 15564
rect 2827 15524 2872 15552
rect 2685 15515 2743 15521
rect 2866 15512 2872 15524
rect 2924 15512 2930 15564
rect 4126 15552 4154 15592
rect 4386 15589 4398 15623
rect 4432 15589 4444 15623
rect 4386 15583 4444 15589
rect 5810 15580 5816 15632
rect 5868 15620 5874 15632
rect 6134 15623 6192 15629
rect 6134 15620 6146 15623
rect 5868 15592 6146 15620
rect 5868 15580 5874 15592
rect 6134 15589 6146 15592
rect 6180 15589 6192 15623
rect 8662 15620 8668 15632
rect 8623 15592 8668 15620
rect 6134 15583 6192 15589
rect 8662 15580 8668 15592
rect 8720 15580 8726 15632
rect 5902 15552 5908 15564
rect 4126 15524 5908 15552
rect 5902 15512 5908 15524
rect 5960 15552 5966 15564
rect 7929 15555 7987 15561
rect 7929 15552 7941 15555
rect 5960 15524 7941 15552
rect 5960 15512 5966 15524
rect 7929 15521 7941 15524
rect 7975 15552 7987 15555
rect 8294 15552 8300 15564
rect 7975 15524 8300 15552
rect 7975 15521 7987 15524
rect 7929 15515 7987 15521
rect 8294 15512 8300 15524
rect 8352 15512 8358 15564
rect 8389 15555 8447 15561
rect 8389 15521 8401 15555
rect 8435 15521 8447 15555
rect 9646 15552 9674 15660
rect 10042 15648 10048 15660
rect 10100 15648 10106 15700
rect 12434 15688 12440 15700
rect 12395 15660 12440 15688
rect 12434 15648 12440 15660
rect 12492 15648 12498 15700
rect 18233 15691 18291 15697
rect 18233 15657 18245 15691
rect 18279 15688 18291 15691
rect 18322 15688 18328 15700
rect 18279 15660 18328 15688
rect 18279 15657 18291 15660
rect 18233 15651 18291 15657
rect 18322 15648 18328 15660
rect 18380 15688 18386 15700
rect 18509 15691 18567 15697
rect 18509 15688 18521 15691
rect 18380 15660 18521 15688
rect 18380 15648 18386 15660
rect 18509 15657 18521 15660
rect 18555 15657 18567 15691
rect 18509 15651 18567 15657
rect 10321 15623 10379 15629
rect 10321 15589 10333 15623
rect 10367 15620 10379 15623
rect 10502 15620 10508 15632
rect 10367 15592 10508 15620
rect 10367 15589 10379 15592
rect 10321 15583 10379 15589
rect 10502 15580 10508 15592
rect 10560 15580 10566 15632
rect 14369 15623 14427 15629
rect 14369 15589 14381 15623
rect 14415 15620 14427 15623
rect 14826 15620 14832 15632
rect 14415 15592 14832 15620
rect 14415 15589 14427 15592
rect 14369 15583 14427 15589
rect 14826 15580 14832 15592
rect 14884 15580 14890 15632
rect 15378 15580 15384 15632
rect 15436 15620 15442 15632
rect 15473 15623 15531 15629
rect 15473 15620 15485 15623
rect 15436 15592 15485 15620
rect 15436 15580 15442 15592
rect 15473 15589 15485 15592
rect 15519 15589 15531 15623
rect 16022 15620 16028 15632
rect 15983 15592 16028 15620
rect 15473 15583 15531 15589
rect 16022 15580 16028 15592
rect 16080 15580 16086 15632
rect 17402 15580 17408 15632
rect 17460 15620 17466 15632
rect 17634 15623 17692 15629
rect 17634 15620 17646 15623
rect 17460 15592 17646 15620
rect 17460 15580 17466 15592
rect 17634 15589 17646 15592
rect 17680 15620 17692 15623
rect 18877 15623 18935 15629
rect 18877 15620 18889 15623
rect 17680 15592 18889 15620
rect 17680 15589 17692 15592
rect 17634 15583 17692 15589
rect 18877 15589 18889 15592
rect 18923 15620 18935 15623
rect 18966 15620 18972 15632
rect 18923 15592 18972 15620
rect 18923 15589 18935 15592
rect 18877 15583 18935 15589
rect 18966 15580 18972 15592
rect 19024 15580 19030 15632
rect 19242 15620 19248 15632
rect 19203 15592 19248 15620
rect 19242 15580 19248 15592
rect 19300 15580 19306 15632
rect 10042 15552 10048 15564
rect 9646 15524 10048 15552
rect 8389 15515 8447 15521
rect 3142 15484 3148 15496
rect 3103 15456 3148 15484
rect 3142 15444 3148 15456
rect 3200 15484 3206 15496
rect 4065 15487 4123 15493
rect 4065 15484 4077 15487
rect 3200 15456 4077 15484
rect 3200 15444 3206 15456
rect 4065 15453 4077 15456
rect 4111 15453 4123 15487
rect 4065 15447 4123 15453
rect 5813 15487 5871 15493
rect 5813 15453 5825 15487
rect 5859 15484 5871 15487
rect 5994 15484 6000 15496
rect 5859 15456 6000 15484
rect 5859 15453 5871 15456
rect 5813 15447 5871 15453
rect 5994 15444 6000 15456
rect 6052 15444 6058 15496
rect 8110 15444 8116 15496
rect 8168 15484 8174 15496
rect 8404 15484 8432 15515
rect 10042 15512 10048 15524
rect 10100 15512 10106 15564
rect 13814 15512 13820 15564
rect 13872 15552 13878 15564
rect 14090 15552 14096 15564
rect 13872 15524 13917 15552
rect 14051 15524 14096 15552
rect 13872 15512 13878 15524
rect 14090 15512 14096 15524
rect 14148 15512 14154 15564
rect 18690 15512 18696 15564
rect 18748 15552 18754 15564
rect 19096 15555 19154 15561
rect 19096 15552 19108 15555
rect 18748 15524 19108 15552
rect 18748 15512 18754 15524
rect 19096 15521 19108 15524
rect 19142 15552 19154 15555
rect 21634 15552 21640 15564
rect 19142 15524 21640 15552
rect 19142 15521 19154 15524
rect 19096 15515 19154 15521
rect 21634 15512 21640 15524
rect 21692 15552 21698 15564
rect 23566 15552 23572 15564
rect 21692 15524 23572 15552
rect 21692 15512 21698 15524
rect 23566 15512 23572 15524
rect 23624 15512 23630 15564
rect 8168 15456 8432 15484
rect 8168 15444 8174 15456
rect 9766 15444 9772 15496
rect 9824 15484 9830 15496
rect 10229 15487 10287 15493
rect 10229 15484 10241 15487
rect 9824 15456 10241 15484
rect 9824 15444 9830 15456
rect 10229 15453 10241 15456
rect 10275 15453 10287 15487
rect 10594 15484 10600 15496
rect 10555 15456 10600 15484
rect 10229 15447 10287 15453
rect 10594 15444 10600 15456
rect 10652 15444 10658 15496
rect 15194 15444 15200 15496
rect 15252 15484 15258 15496
rect 15381 15487 15439 15493
rect 15381 15484 15393 15487
rect 15252 15456 15393 15484
rect 15252 15444 15258 15456
rect 15381 15453 15393 15456
rect 15427 15453 15439 15487
rect 17310 15484 17316 15496
rect 17271 15456 17316 15484
rect 15381 15447 15439 15453
rect 17310 15444 17316 15456
rect 17368 15444 17374 15496
rect 12989 15419 13047 15425
rect 12989 15385 13001 15419
rect 13035 15416 13047 15419
rect 13262 15416 13268 15428
rect 13035 15388 13268 15416
rect 13035 15385 13047 15388
rect 12989 15379 13047 15385
rect 13262 15376 13268 15388
rect 13320 15376 13326 15428
rect 7374 15348 7380 15360
rect 7335 15320 7380 15348
rect 7374 15308 7380 15320
rect 7432 15308 7438 15360
rect 10410 15308 10416 15360
rect 10468 15348 10474 15360
rect 11149 15351 11207 15357
rect 11149 15348 11161 15351
rect 10468 15320 11161 15348
rect 10468 15308 10474 15320
rect 11149 15317 11161 15320
rect 11195 15317 11207 15351
rect 16390 15348 16396 15360
rect 16351 15320 16396 15348
rect 11149 15311 11207 15317
rect 16390 15308 16396 15320
rect 16448 15308 16454 15360
rect 1104 15258 22816 15280
rect 1104 15206 4982 15258
rect 5034 15206 5046 15258
rect 5098 15206 5110 15258
rect 5162 15206 5174 15258
rect 5226 15206 12982 15258
rect 13034 15206 13046 15258
rect 13098 15206 13110 15258
rect 13162 15206 13174 15258
rect 13226 15206 20982 15258
rect 21034 15206 21046 15258
rect 21098 15206 21110 15258
rect 21162 15206 21174 15258
rect 21226 15206 22816 15258
rect 1104 15184 22816 15206
rect 2774 15144 2780 15156
rect 2735 15116 2780 15144
rect 2774 15104 2780 15116
rect 2832 15104 2838 15156
rect 3142 15144 3148 15156
rect 3103 15116 3148 15144
rect 3142 15104 3148 15116
rect 3200 15104 3206 15156
rect 4154 15104 4160 15156
rect 4212 15144 4218 15156
rect 5810 15144 5816 15156
rect 4212 15116 5816 15144
rect 4212 15104 4218 15116
rect 5810 15104 5816 15116
rect 5868 15104 5874 15156
rect 6641 15147 6699 15153
rect 6641 15113 6653 15147
rect 6687 15144 6699 15147
rect 7006 15144 7012 15156
rect 6687 15116 7012 15144
rect 6687 15113 6699 15116
rect 6641 15107 6699 15113
rect 7006 15104 7012 15116
rect 7064 15104 7070 15156
rect 8987 15147 9045 15153
rect 8987 15113 8999 15147
rect 9033 15144 9045 15147
rect 9766 15144 9772 15156
rect 9033 15116 9772 15144
rect 9033 15113 9045 15116
rect 8987 15107 9045 15113
rect 9766 15104 9772 15116
rect 9824 15104 9830 15156
rect 9999 15147 10057 15153
rect 9999 15113 10011 15147
rect 10045 15144 10057 15147
rect 10410 15144 10416 15156
rect 10045 15116 10416 15144
rect 10045 15113 10057 15116
rect 9999 15107 10057 15113
rect 10410 15104 10416 15116
rect 10468 15104 10474 15156
rect 10502 15104 10508 15156
rect 10560 15144 10566 15156
rect 10689 15147 10747 15153
rect 10689 15144 10701 15147
rect 10560 15116 10701 15144
rect 10560 15104 10566 15116
rect 10689 15113 10701 15116
rect 10735 15113 10747 15147
rect 10689 15107 10747 15113
rect 14090 15104 14096 15156
rect 14148 15144 14154 15156
rect 15010 15144 15016 15156
rect 14148 15116 15016 15144
rect 14148 15104 14154 15116
rect 15010 15104 15016 15116
rect 15068 15104 15074 15156
rect 15378 15144 15384 15156
rect 15339 15116 15384 15144
rect 15378 15104 15384 15116
rect 15436 15104 15442 15156
rect 18690 15144 18696 15156
rect 18651 15116 18696 15144
rect 18690 15104 18696 15116
rect 18748 15104 18754 15156
rect 19978 15104 19984 15156
rect 20036 15144 20042 15156
rect 20441 15147 20499 15153
rect 20441 15144 20453 15147
rect 20036 15116 20453 15144
rect 20036 15104 20042 15116
rect 20441 15113 20453 15116
rect 20487 15113 20499 15147
rect 20441 15107 20499 15113
rect 2501 15079 2559 15085
rect 2501 15045 2513 15079
rect 2547 15076 2559 15079
rect 2866 15076 2872 15088
rect 2547 15048 2872 15076
rect 2547 15045 2559 15048
rect 2501 15039 2559 15045
rect 2866 15036 2872 15048
rect 2924 15036 2930 15088
rect 4985 15079 5043 15085
rect 4985 15045 4997 15079
rect 5031 15076 5043 15079
rect 5442 15076 5448 15088
rect 5031 15048 5448 15076
rect 5031 15045 5043 15048
rect 4985 15039 5043 15045
rect 5442 15036 5448 15048
rect 5500 15076 5506 15088
rect 7469 15079 7527 15085
rect 7469 15076 7481 15079
rect 5500 15048 7481 15076
rect 5500 15036 5506 15048
rect 7469 15045 7481 15048
rect 7515 15045 7527 15079
rect 7469 15039 7527 15045
rect 9490 15036 9496 15088
rect 9548 15076 9554 15088
rect 11011 15079 11069 15085
rect 11011 15076 11023 15079
rect 9548 15048 11023 15076
rect 9548 15036 9554 15048
rect 11011 15045 11023 15048
rect 11057 15045 11069 15079
rect 11011 15039 11069 15045
rect 11425 15079 11483 15085
rect 11425 15045 11437 15079
rect 11471 15076 11483 15079
rect 15102 15076 15108 15088
rect 11471 15048 15108 15076
rect 11471 15045 11483 15048
rect 11425 15039 11483 15045
rect 3467 15011 3525 15017
rect 3467 14977 3479 15011
rect 3513 15008 3525 15011
rect 4433 15011 4491 15017
rect 4433 15008 4445 15011
rect 3513 14980 4445 15008
rect 3513 14977 3525 14980
rect 3467 14971 3525 14977
rect 4433 14977 4445 14980
rect 4479 15008 4491 15011
rect 5353 15011 5411 15017
rect 5353 15008 5365 15011
rect 4479 14980 5365 15008
rect 4479 14977 4491 14980
rect 4433 14971 4491 14977
rect 5353 14977 5365 14980
rect 5399 14977 5411 15011
rect 5353 14971 5411 14977
rect 6917 15011 6975 15017
rect 6917 14977 6929 15011
rect 6963 15008 6975 15011
rect 7374 15008 7380 15020
rect 6963 14980 7380 15008
rect 6963 14977 6975 14980
rect 6917 14971 6975 14977
rect 7374 14968 7380 14980
rect 7432 14968 7438 15020
rect 7926 14968 7932 15020
rect 7984 15008 7990 15020
rect 7984 14980 10983 15008
rect 7984 14968 7990 14980
rect 3050 14900 3056 14952
rect 3108 14940 3114 14952
rect 3364 14943 3422 14949
rect 3364 14940 3376 14943
rect 3108 14912 3376 14940
rect 3108 14900 3114 14912
rect 3364 14909 3376 14912
rect 3410 14940 3422 14943
rect 3789 14943 3847 14949
rect 3789 14940 3801 14943
rect 3410 14912 3801 14940
rect 3410 14909 3422 14912
rect 3364 14903 3422 14909
rect 3528 14884 3556 14912
rect 3789 14909 3801 14912
rect 3835 14909 3847 14943
rect 3789 14903 3847 14909
rect 8754 14900 8760 14952
rect 8812 14940 8818 14952
rect 8884 14943 8942 14949
rect 8884 14940 8896 14943
rect 8812 14912 8896 14940
rect 8812 14900 8818 14912
rect 8884 14909 8896 14912
rect 8930 14940 8942 14943
rect 9306 14940 9312 14952
rect 8930 14912 9312 14940
rect 8930 14909 8942 14912
rect 8884 14903 8942 14909
rect 9306 14900 9312 14912
rect 9364 14900 9370 14952
rect 9928 14943 9986 14949
rect 9928 14909 9940 14943
rect 9974 14940 9986 14943
rect 10410 14940 10416 14952
rect 9974 14912 10416 14940
rect 9974 14909 9986 14912
rect 9928 14903 9986 14909
rect 10410 14900 10416 14912
rect 10468 14900 10474 14952
rect 10955 14949 10983 14980
rect 10940 14943 10998 14949
rect 10940 14909 10952 14943
rect 10986 14940 10998 14943
rect 11440 14940 11468 15039
rect 15102 15036 15108 15048
rect 15160 15036 15166 15088
rect 15194 15036 15200 15088
rect 15252 15076 15258 15088
rect 15657 15079 15715 15085
rect 15657 15076 15669 15079
rect 15252 15048 15669 15076
rect 15252 15036 15258 15048
rect 15657 15045 15669 15048
rect 15703 15045 15715 15079
rect 15657 15039 15715 15045
rect 14550 15008 14556 15020
rect 14511 14980 14556 15008
rect 14550 14968 14556 14980
rect 14608 14968 14614 15020
rect 15010 14968 15016 15020
rect 15068 15008 15074 15020
rect 16209 15011 16267 15017
rect 16209 15008 16221 15011
rect 15068 14980 16221 15008
rect 15068 14968 15074 14980
rect 16209 14977 16221 14980
rect 16255 15008 16267 15011
rect 17129 15011 17187 15017
rect 16255 14980 16896 15008
rect 16255 14977 16267 14980
rect 16209 14971 16267 14977
rect 10986 14912 11468 14940
rect 10986 14909 10998 14912
rect 10940 14903 10998 14909
rect 15562 14900 15568 14952
rect 15620 14940 15626 14952
rect 16390 14940 16396 14952
rect 15620 14912 16396 14940
rect 15620 14900 15626 14912
rect 16390 14900 16396 14912
rect 16448 14900 16454 14952
rect 16868 14949 16896 14980
rect 17129 14977 17141 15011
rect 17175 15008 17187 15011
rect 17310 15008 17316 15020
rect 17175 14980 17316 15008
rect 17175 14977 17187 14980
rect 17129 14971 17187 14977
rect 17310 14968 17316 14980
rect 17368 15008 17374 15020
rect 17773 15011 17831 15017
rect 17773 15008 17785 15011
rect 17368 14980 17785 15008
rect 17368 14968 17374 14980
rect 17773 14977 17785 14980
rect 17819 14977 17831 15011
rect 20456 15008 20484 15107
rect 21266 15036 21272 15088
rect 21324 15076 21330 15088
rect 21324 15048 21404 15076
rect 21324 15036 21330 15048
rect 21376 15017 21404 15048
rect 20717 15011 20775 15017
rect 20717 15008 20729 15011
rect 20456 14980 20729 15008
rect 17773 14971 17831 14977
rect 20717 14977 20729 14980
rect 20763 14977 20775 15011
rect 20717 14971 20775 14977
rect 21361 15011 21419 15017
rect 21361 14977 21373 15011
rect 21407 15008 21419 15011
rect 21450 15008 21456 15020
rect 21407 14980 21456 15008
rect 21407 14977 21419 14980
rect 21361 14971 21419 14977
rect 21450 14968 21456 14980
rect 21508 14968 21514 15020
rect 16853 14943 16911 14949
rect 16853 14909 16865 14943
rect 16899 14909 16911 14943
rect 18877 14943 18935 14949
rect 18877 14940 18889 14943
rect 16853 14903 16911 14909
rect 18340 14912 18889 14940
rect 3510 14832 3516 14884
rect 3568 14832 3574 14884
rect 4522 14872 4528 14884
rect 4483 14844 4528 14872
rect 4522 14832 4528 14844
rect 4580 14832 4586 14884
rect 7006 14872 7012 14884
rect 6967 14844 7012 14872
rect 7006 14832 7012 14844
rect 7064 14832 7070 14884
rect 11885 14875 11943 14881
rect 11885 14841 11897 14875
rect 11931 14872 11943 14875
rect 12526 14872 12532 14884
rect 11931 14844 12532 14872
rect 11931 14841 11943 14844
rect 11885 14835 11943 14841
rect 12526 14832 12532 14844
rect 12584 14832 12590 14884
rect 12621 14875 12679 14881
rect 12621 14841 12633 14875
rect 12667 14841 12679 14875
rect 12621 14835 12679 14841
rect 13173 14875 13231 14881
rect 13173 14841 13185 14875
rect 13219 14872 13231 14875
rect 13354 14872 13360 14884
rect 13219 14844 13360 14872
rect 13219 14841 13231 14844
rect 13173 14835 13231 14841
rect 4154 14764 4160 14816
rect 4212 14804 4218 14816
rect 4212 14776 4257 14804
rect 4212 14764 4218 14776
rect 5994 14764 6000 14816
rect 6052 14804 6058 14816
rect 6181 14807 6239 14813
rect 6181 14804 6193 14807
rect 6052 14776 6193 14804
rect 6052 14764 6058 14776
rect 6181 14773 6193 14776
rect 6227 14773 6239 14807
rect 6181 14767 6239 14773
rect 8021 14807 8079 14813
rect 8021 14773 8033 14807
rect 8067 14804 8079 14807
rect 8110 14804 8116 14816
rect 8067 14776 8116 14804
rect 8067 14773 8079 14776
rect 8021 14767 8079 14773
rect 8110 14764 8116 14776
rect 8168 14764 8174 14816
rect 8294 14804 8300 14816
rect 8255 14776 8300 14804
rect 8294 14764 8300 14776
rect 8352 14764 8358 14816
rect 12158 14804 12164 14816
rect 12119 14776 12164 14804
rect 12158 14764 12164 14776
rect 12216 14804 12222 14816
rect 12636 14804 12664 14835
rect 13354 14832 13360 14844
rect 13412 14832 13418 14884
rect 13725 14875 13783 14881
rect 13725 14841 13737 14875
rect 13771 14872 13783 14875
rect 14090 14872 14096 14884
rect 13771 14844 14096 14872
rect 13771 14841 13783 14844
rect 13725 14835 13783 14841
rect 14090 14832 14096 14844
rect 14148 14832 14154 14884
rect 14277 14875 14335 14881
rect 14277 14841 14289 14875
rect 14323 14841 14335 14875
rect 14277 14835 14335 14841
rect 12216 14776 12664 14804
rect 12216 14764 12222 14776
rect 13814 14764 13820 14816
rect 13872 14804 13878 14816
rect 14001 14807 14059 14813
rect 14001 14804 14013 14807
rect 13872 14776 14013 14804
rect 13872 14764 13878 14776
rect 14001 14773 14013 14776
rect 14047 14773 14059 14807
rect 14292 14804 14320 14835
rect 14366 14832 14372 14884
rect 14424 14872 14430 14884
rect 14424 14844 14469 14872
rect 14424 14832 14430 14844
rect 18340 14816 18368 14912
rect 18877 14909 18889 14912
rect 18923 14909 18935 14943
rect 18877 14903 18935 14909
rect 18966 14832 18972 14884
rect 19024 14872 19030 14884
rect 19198 14875 19256 14881
rect 19198 14872 19210 14875
rect 19024 14844 19210 14872
rect 19024 14832 19030 14844
rect 19198 14841 19210 14844
rect 19244 14841 19256 14875
rect 19198 14835 19256 14841
rect 20809 14875 20867 14881
rect 20809 14841 20821 14875
rect 20855 14841 20867 14875
rect 20809 14835 20867 14841
rect 14458 14804 14464 14816
rect 14292 14776 14464 14804
rect 14001 14767 14059 14773
rect 14458 14764 14464 14776
rect 14516 14764 14522 14816
rect 16298 14764 16304 14816
rect 16356 14804 16362 14816
rect 17402 14804 17408 14816
rect 16356 14776 17408 14804
rect 16356 14764 16362 14776
rect 17402 14764 17408 14776
rect 17460 14764 17466 14816
rect 18322 14804 18328 14816
rect 18283 14776 18328 14804
rect 18322 14764 18328 14776
rect 18380 14764 18386 14816
rect 19797 14807 19855 14813
rect 19797 14773 19809 14807
rect 19843 14804 19855 14807
rect 20622 14804 20628 14816
rect 19843 14776 20628 14804
rect 19843 14773 19855 14776
rect 19797 14767 19855 14773
rect 20622 14764 20628 14776
rect 20680 14804 20686 14816
rect 20824 14804 20852 14835
rect 20680 14776 20852 14804
rect 20680 14764 20686 14776
rect 1104 14714 22816 14736
rect 1104 14662 8982 14714
rect 9034 14662 9046 14714
rect 9098 14662 9110 14714
rect 9162 14662 9174 14714
rect 9226 14662 16982 14714
rect 17034 14662 17046 14714
rect 17098 14662 17110 14714
rect 17162 14662 17174 14714
rect 17226 14662 22816 14714
rect 1104 14640 22816 14662
rect 1118 14560 1124 14612
rect 1176 14600 1182 14612
rect 1581 14603 1639 14609
rect 1581 14600 1593 14603
rect 1176 14572 1593 14600
rect 1176 14560 1182 14572
rect 1581 14569 1593 14572
rect 1627 14569 1639 14603
rect 4522 14600 4528 14612
rect 4483 14572 4528 14600
rect 1581 14563 1639 14569
rect 4522 14560 4528 14572
rect 4580 14560 4586 14612
rect 6963 14603 7021 14609
rect 6963 14569 6975 14603
rect 7009 14600 7021 14603
rect 7374 14600 7380 14612
rect 7009 14572 7380 14600
rect 7009 14569 7021 14572
rect 6963 14563 7021 14569
rect 7374 14560 7380 14572
rect 7432 14560 7438 14612
rect 10042 14600 10048 14612
rect 10003 14572 10048 14600
rect 10042 14560 10048 14572
rect 10100 14560 10106 14612
rect 10502 14560 10508 14612
rect 10560 14600 10566 14612
rect 10597 14603 10655 14609
rect 10597 14600 10609 14603
rect 10560 14572 10609 14600
rect 10560 14560 10566 14572
rect 10597 14569 10609 14572
rect 10643 14569 10655 14603
rect 10870 14600 10876 14612
rect 10831 14572 10876 14600
rect 10597 14563 10655 14569
rect 10870 14560 10876 14572
rect 10928 14600 10934 14612
rect 16666 14600 16672 14612
rect 10928 14572 16672 14600
rect 10928 14560 10934 14572
rect 16666 14560 16672 14572
rect 16724 14600 16730 14612
rect 20622 14600 20628 14612
rect 16724 14572 19012 14600
rect 20583 14572 20628 14600
rect 16724 14560 16730 14572
rect 5994 14532 6000 14544
rect 5955 14504 6000 14532
rect 5994 14492 6000 14504
rect 6052 14492 6058 14544
rect 11606 14492 11612 14544
rect 11664 14532 11670 14544
rect 11746 14535 11804 14541
rect 11746 14532 11758 14535
rect 11664 14504 11758 14532
rect 11664 14492 11670 14504
rect 11746 14501 11758 14504
rect 11792 14501 11804 14535
rect 11746 14495 11804 14501
rect 17865 14535 17923 14541
rect 17865 14501 17877 14535
rect 17911 14532 17923 14535
rect 18322 14532 18328 14544
rect 17911 14504 18328 14532
rect 17911 14501 17923 14504
rect 17865 14495 17923 14501
rect 18322 14492 18328 14504
rect 18380 14492 18386 14544
rect 18984 14476 19012 14572
rect 20622 14560 20628 14572
rect 20680 14560 20686 14612
rect 21085 14603 21143 14609
rect 21085 14569 21097 14603
rect 21131 14600 21143 14603
rect 22278 14600 22284 14612
rect 21131 14572 22284 14600
rect 21131 14569 21143 14572
rect 21085 14563 21143 14569
rect 22278 14560 22284 14572
rect 22336 14560 22342 14612
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14464 1455 14467
rect 2038 14464 2044 14476
rect 1443 14436 2044 14464
rect 1443 14433 1455 14436
rect 1397 14427 1455 14433
rect 2038 14424 2044 14436
rect 2096 14424 2102 14476
rect 4132 14467 4190 14473
rect 4132 14433 4144 14467
rect 4178 14464 4190 14467
rect 5261 14467 5319 14473
rect 4178 14433 4200 14464
rect 4132 14427 4200 14433
rect 5261 14433 5273 14467
rect 5307 14433 5319 14467
rect 5261 14427 5319 14433
rect 4062 14288 4068 14340
rect 4120 14328 4126 14340
rect 4172 14328 4200 14427
rect 5276 14396 5304 14427
rect 5350 14424 5356 14476
rect 5408 14464 5414 14476
rect 5721 14467 5779 14473
rect 5721 14464 5733 14467
rect 5408 14436 5733 14464
rect 5408 14424 5414 14436
rect 5721 14433 5733 14436
rect 5767 14433 5779 14467
rect 5721 14427 5779 14433
rect 6892 14467 6950 14473
rect 6892 14433 6904 14467
rect 6938 14464 6950 14467
rect 7006 14464 7012 14476
rect 6938 14436 7012 14464
rect 6938 14433 6950 14436
rect 6892 14427 6950 14433
rect 7006 14424 7012 14436
rect 7064 14424 7070 14476
rect 7190 14424 7196 14476
rect 7248 14464 7254 14476
rect 7872 14467 7930 14473
rect 7872 14464 7884 14467
rect 7248 14436 7884 14464
rect 7248 14424 7254 14436
rect 7872 14433 7884 14436
rect 7918 14433 7930 14467
rect 7872 14427 7930 14433
rect 13262 14424 13268 14476
rect 13320 14464 13326 14476
rect 13357 14467 13415 14473
rect 13357 14464 13369 14467
rect 13320 14436 13369 14464
rect 13320 14424 13326 14436
rect 13357 14433 13369 14436
rect 13403 14433 13415 14467
rect 13630 14464 13636 14476
rect 13591 14436 13636 14464
rect 13357 14427 13415 14433
rect 5534 14396 5540 14408
rect 5276 14368 5540 14396
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 9674 14396 9680 14408
rect 9635 14368 9680 14396
rect 9674 14356 9680 14368
rect 9732 14356 9738 14408
rect 11425 14399 11483 14405
rect 11425 14365 11437 14399
rect 11471 14396 11483 14399
rect 11974 14396 11980 14408
rect 11471 14368 11980 14396
rect 11471 14365 11483 14368
rect 11425 14359 11483 14365
rect 11974 14356 11980 14368
rect 12032 14356 12038 14408
rect 13372 14396 13400 14427
rect 13630 14424 13636 14436
rect 13688 14424 13694 14476
rect 15194 14424 15200 14476
rect 15252 14464 15258 14476
rect 15562 14464 15568 14476
rect 15252 14436 15568 14464
rect 15252 14424 15258 14436
rect 15562 14424 15568 14436
rect 15620 14424 15626 14476
rect 16025 14467 16083 14473
rect 16025 14433 16037 14467
rect 16071 14464 16083 14467
rect 16390 14464 16396 14476
rect 16071 14436 16396 14464
rect 16071 14433 16083 14436
rect 16025 14427 16083 14433
rect 16390 14424 16396 14436
rect 16448 14424 16454 14476
rect 16850 14424 16856 14476
rect 16908 14464 16914 14476
rect 17129 14467 17187 14473
rect 17129 14464 17141 14467
rect 16908 14436 17141 14464
rect 16908 14424 16914 14436
rect 17129 14433 17141 14436
rect 17175 14464 17187 14467
rect 17310 14464 17316 14476
rect 17175 14436 17316 14464
rect 17175 14433 17187 14436
rect 17129 14427 17187 14433
rect 17310 14424 17316 14436
rect 17368 14424 17374 14476
rect 17586 14464 17592 14476
rect 17547 14436 17592 14464
rect 17586 14424 17592 14436
rect 17644 14424 17650 14476
rect 18966 14464 18972 14476
rect 18927 14436 18972 14464
rect 18966 14424 18972 14436
rect 19024 14424 19030 14476
rect 19058 14424 19064 14476
rect 19116 14464 19122 14476
rect 19153 14467 19211 14473
rect 19153 14464 19165 14467
rect 19116 14436 19165 14464
rect 19116 14424 19122 14436
rect 19153 14433 19165 14436
rect 19199 14433 19211 14467
rect 19153 14427 19211 14433
rect 20806 14424 20812 14476
rect 20864 14464 20870 14476
rect 20901 14467 20959 14473
rect 20901 14464 20913 14467
rect 20864 14436 20913 14464
rect 20864 14424 20870 14436
rect 20901 14433 20913 14436
rect 20947 14433 20959 14467
rect 20901 14427 20959 14433
rect 13722 14396 13728 14408
rect 13372 14368 13492 14396
rect 13683 14368 13728 14396
rect 8386 14328 8392 14340
rect 4120 14300 8392 14328
rect 4120 14288 4126 14300
rect 8386 14288 8392 14300
rect 8444 14288 8450 14340
rect 13464 14328 13492 14368
rect 13722 14356 13728 14368
rect 13780 14356 13786 14408
rect 16114 14396 16120 14408
rect 16075 14368 16120 14396
rect 16114 14356 16120 14368
rect 16172 14356 16178 14408
rect 19242 14396 19248 14408
rect 19203 14368 19248 14396
rect 19242 14356 19248 14368
rect 19300 14356 19306 14408
rect 13998 14328 14004 14340
rect 13464 14300 14004 14328
rect 13998 14288 14004 14300
rect 14056 14288 14062 14340
rect 4203 14263 4261 14269
rect 4203 14229 4215 14263
rect 4249 14260 4261 14263
rect 4338 14260 4344 14272
rect 4249 14232 4344 14260
rect 4249 14229 4261 14232
rect 4203 14223 4261 14229
rect 4338 14220 4344 14232
rect 4396 14220 4402 14272
rect 7469 14263 7527 14269
rect 7469 14229 7481 14263
rect 7515 14260 7527 14263
rect 7558 14260 7564 14272
rect 7515 14232 7564 14260
rect 7515 14229 7527 14232
rect 7469 14223 7527 14229
rect 7558 14220 7564 14232
rect 7616 14220 7622 14272
rect 7650 14220 7656 14272
rect 7708 14260 7714 14272
rect 7975 14263 8033 14269
rect 7975 14260 7987 14263
rect 7708 14232 7987 14260
rect 7708 14220 7714 14232
rect 7975 14229 7987 14232
rect 8021 14229 8033 14263
rect 12342 14260 12348 14272
rect 12303 14232 12348 14260
rect 7975 14223 8033 14229
rect 12342 14220 12348 14232
rect 12400 14220 12406 14272
rect 14274 14260 14280 14272
rect 14235 14232 14280 14260
rect 14274 14220 14280 14232
rect 14332 14220 14338 14272
rect 14458 14220 14464 14272
rect 14516 14260 14522 14272
rect 14553 14263 14611 14269
rect 14553 14260 14565 14263
rect 14516 14232 14565 14260
rect 14516 14220 14522 14232
rect 14553 14229 14565 14232
rect 14599 14229 14611 14263
rect 20162 14260 20168 14272
rect 20123 14232 20168 14260
rect 14553 14223 14611 14229
rect 20162 14220 20168 14232
rect 20220 14220 20226 14272
rect 1104 14170 22816 14192
rect 1104 14118 4982 14170
rect 5034 14118 5046 14170
rect 5098 14118 5110 14170
rect 5162 14118 5174 14170
rect 5226 14118 12982 14170
rect 13034 14118 13046 14170
rect 13098 14118 13110 14170
rect 13162 14118 13174 14170
rect 13226 14118 20982 14170
rect 21034 14118 21046 14170
rect 21098 14118 21110 14170
rect 21162 14118 21174 14170
rect 21226 14118 22816 14170
rect 1104 14096 22816 14118
rect 106 14016 112 14068
rect 164 14056 170 14068
rect 1581 14059 1639 14065
rect 1581 14056 1593 14059
rect 164 14028 1593 14056
rect 164 14016 170 14028
rect 1581 14025 1593 14028
rect 1627 14025 1639 14059
rect 4062 14056 4068 14068
rect 4023 14028 4068 14056
rect 1581 14019 1639 14025
rect 4062 14016 4068 14028
rect 4120 14016 4126 14068
rect 7190 14016 7196 14068
rect 7248 14056 7254 14068
rect 8389 14059 8447 14065
rect 8389 14056 8401 14059
rect 7248 14028 8401 14056
rect 7248 14016 7254 14028
rect 8389 14025 8401 14028
rect 8435 14025 8447 14059
rect 8389 14019 8447 14025
rect 11606 14016 11612 14068
rect 11664 14056 11670 14068
rect 12759 14059 12817 14065
rect 11664 14028 12709 14056
rect 11664 14016 11670 14028
rect 4430 13948 4436 14000
rect 4488 13988 4494 14000
rect 4801 13991 4859 13997
rect 4801 13988 4813 13991
rect 4488 13960 4813 13988
rect 4488 13948 4494 13960
rect 4801 13957 4813 13960
rect 4847 13988 4859 13991
rect 8021 13991 8079 13997
rect 8021 13988 8033 13991
rect 4847 13960 8033 13988
rect 4847 13957 4859 13960
rect 4801 13951 4859 13957
rect 8021 13957 8033 13960
rect 8067 13988 8079 13991
rect 8754 13988 8760 14000
rect 8067 13960 8760 13988
rect 8067 13957 8079 13960
rect 8021 13951 8079 13957
rect 8754 13948 8760 13960
rect 8812 13948 8818 14000
rect 12250 13988 12256 14000
rect 10014 13960 12256 13988
rect 3329 13923 3387 13929
rect 3329 13889 3341 13923
rect 3375 13920 3387 13923
rect 4249 13923 4307 13929
rect 4249 13920 4261 13923
rect 3375 13892 4261 13920
rect 3375 13889 3387 13892
rect 3329 13883 3387 13889
rect 4249 13889 4261 13892
rect 4295 13920 4307 13923
rect 4338 13920 4344 13932
rect 4295 13892 4344 13920
rect 4295 13889 4307 13892
rect 4249 13883 4307 13889
rect 4338 13880 4344 13892
rect 4396 13880 4402 13932
rect 7466 13920 7472 13932
rect 7379 13892 7472 13920
rect 7466 13880 7472 13892
rect 7524 13920 7530 13932
rect 7650 13920 7656 13932
rect 7524 13892 7656 13920
rect 7524 13880 7530 13892
rect 7650 13880 7656 13892
rect 7708 13880 7714 13932
rect 8110 13880 8116 13932
rect 8168 13920 8174 13932
rect 8849 13923 8907 13929
rect 8849 13920 8861 13923
rect 8168 13892 8861 13920
rect 8168 13880 8174 13892
rect 8849 13889 8861 13892
rect 8895 13920 8907 13923
rect 10014 13920 10042 13960
rect 12250 13948 12256 13960
rect 12308 13948 12314 14000
rect 12681 13988 12709 14028
rect 12759 14025 12771 14059
rect 12805 14056 12817 14059
rect 14458 14056 14464 14068
rect 12805 14028 14464 14056
rect 12805 14025 12817 14028
rect 12759 14019 12817 14025
rect 14458 14016 14464 14028
rect 14516 14016 14522 14068
rect 19058 14056 19064 14068
rect 19019 14028 19064 14056
rect 19058 14016 19064 14028
rect 19116 14016 19122 14068
rect 13357 13991 13415 13997
rect 13357 13988 13369 13991
rect 12681 13960 13369 13988
rect 13357 13957 13369 13960
rect 13403 13988 13415 13991
rect 13449 13991 13507 13997
rect 13449 13988 13461 13991
rect 13403 13960 13461 13988
rect 13403 13957 13415 13960
rect 13357 13951 13415 13957
rect 13449 13957 13461 13960
rect 13495 13957 13507 13991
rect 13449 13951 13507 13957
rect 14274 13948 14280 14000
rect 14332 13988 14338 14000
rect 14553 13991 14611 13997
rect 14553 13988 14565 13991
rect 14332 13960 14565 13988
rect 14332 13948 14338 13960
rect 14553 13957 14565 13960
rect 14599 13988 14611 13991
rect 15562 13988 15568 14000
rect 14599 13960 15568 13988
rect 14599 13957 14611 13960
rect 14553 13951 14611 13957
rect 15562 13948 15568 13960
rect 15620 13948 15626 14000
rect 18966 13948 18972 14000
rect 19024 13988 19030 14000
rect 19429 13991 19487 13997
rect 19429 13988 19441 13991
rect 19024 13960 19441 13988
rect 19024 13948 19030 13960
rect 19429 13957 19441 13960
rect 19475 13957 19487 13991
rect 19429 13951 19487 13957
rect 20806 13948 20812 14000
rect 20864 13948 20870 14000
rect 8895 13892 10042 13920
rect 10428 13892 11284 13920
rect 8895 13889 8907 13892
rect 8849 13883 8907 13889
rect 1394 13852 1400 13864
rect 1355 13824 1400 13852
rect 1394 13812 1400 13824
rect 1452 13812 1458 13864
rect 5534 13812 5540 13864
rect 5592 13852 5598 13864
rect 5721 13855 5779 13861
rect 5721 13852 5733 13855
rect 5592 13824 5733 13852
rect 5592 13812 5598 13824
rect 5721 13821 5733 13824
rect 5767 13852 5779 13855
rect 6546 13852 6552 13864
rect 5767 13824 6552 13852
rect 5767 13821 5779 13824
rect 5721 13815 5779 13821
rect 6546 13812 6552 13824
rect 6604 13812 6610 13864
rect 9217 13855 9275 13861
rect 9217 13821 9229 13855
rect 9263 13852 9275 13855
rect 9306 13852 9312 13864
rect 9263 13824 9312 13852
rect 9263 13821 9275 13824
rect 9217 13815 9275 13821
rect 9306 13812 9312 13824
rect 9364 13812 9370 13864
rect 9508 13861 9536 13892
rect 9493 13855 9551 13861
rect 9493 13821 9505 13855
rect 9539 13821 9551 13855
rect 10042 13852 10048 13864
rect 9955 13824 10048 13852
rect 9493 13815 9551 13821
rect 10042 13812 10048 13824
rect 10100 13852 10106 13864
rect 10428 13852 10456 13892
rect 10100 13824 10456 13852
rect 10505 13855 10563 13861
rect 10100 13812 10106 13824
rect 10505 13821 10517 13855
rect 10551 13852 10563 13855
rect 10778 13852 10784 13864
rect 10551 13824 10784 13852
rect 10551 13821 10563 13824
rect 10505 13815 10563 13821
rect 10778 13812 10784 13824
rect 10836 13812 10842 13864
rect 10870 13812 10876 13864
rect 10928 13852 10934 13864
rect 11057 13855 11115 13861
rect 11057 13852 11069 13855
rect 10928 13824 11069 13852
rect 10928 13812 10934 13824
rect 11057 13821 11069 13824
rect 11103 13821 11115 13855
rect 11256 13852 11284 13892
rect 11330 13880 11336 13932
rect 11388 13920 11394 13932
rect 13633 13923 13691 13929
rect 11388 13892 12699 13920
rect 11388 13880 11394 13892
rect 11606 13852 11612 13864
rect 11256 13824 11612 13852
rect 11057 13815 11115 13821
rect 11606 13812 11612 13824
rect 11664 13812 11670 13864
rect 12671 13861 12699 13892
rect 13096 13892 13584 13920
rect 13096 13861 13124 13892
rect 12656 13855 12714 13861
rect 12656 13821 12668 13855
rect 12702 13852 12714 13855
rect 13081 13855 13139 13861
rect 13081 13852 13093 13855
rect 12702 13824 13093 13852
rect 12702 13821 12714 13824
rect 12656 13815 12714 13821
rect 13081 13821 13093 13824
rect 13127 13821 13139 13855
rect 13556 13852 13584 13892
rect 13633 13889 13645 13923
rect 13679 13920 13691 13923
rect 13722 13920 13728 13932
rect 13679 13892 13728 13920
rect 13679 13889 13691 13892
rect 13633 13883 13691 13889
rect 13722 13880 13728 13892
rect 13780 13880 13786 13932
rect 15746 13920 15752 13932
rect 14476 13892 15332 13920
rect 15707 13892 15752 13920
rect 14476 13852 14504 13892
rect 13556 13824 14504 13852
rect 13081 13815 13139 13821
rect 3697 13787 3755 13793
rect 3697 13753 3709 13787
rect 3743 13784 3755 13787
rect 4341 13787 4399 13793
rect 4341 13784 4353 13787
rect 3743 13756 4353 13784
rect 3743 13753 3755 13756
rect 3697 13747 3755 13753
rect 4341 13753 4353 13756
rect 4387 13784 4399 13787
rect 4614 13784 4620 13796
rect 4387 13756 4620 13784
rect 4387 13753 4399 13756
rect 4341 13747 4399 13753
rect 4614 13744 4620 13756
rect 4672 13744 4678 13796
rect 5350 13784 5356 13796
rect 5263 13756 5356 13784
rect 5350 13744 5356 13756
rect 5408 13784 5414 13796
rect 7558 13784 7564 13796
rect 5408 13756 7420 13784
rect 7519 13756 7564 13784
rect 5408 13744 5414 13756
rect 2038 13716 2044 13728
rect 1999 13688 2044 13716
rect 2038 13676 2044 13688
rect 2096 13676 2102 13728
rect 7006 13716 7012 13728
rect 6967 13688 7012 13716
rect 7006 13676 7012 13688
rect 7064 13676 7070 13728
rect 7392 13716 7420 13756
rect 7558 13744 7564 13756
rect 7616 13744 7622 13796
rect 9674 13784 9680 13796
rect 9635 13756 9680 13784
rect 9674 13744 9680 13756
rect 9732 13744 9738 13796
rect 13357 13787 13415 13793
rect 9784 13756 12572 13784
rect 9784 13716 9812 13756
rect 10870 13716 10876 13728
rect 7392 13688 9812 13716
rect 10831 13688 10876 13716
rect 10870 13676 10876 13688
rect 10928 13676 10934 13728
rect 11422 13676 11428 13728
rect 11480 13716 11486 13728
rect 11974 13716 11980 13728
rect 11480 13688 11980 13716
rect 11480 13676 11486 13688
rect 11974 13676 11980 13688
rect 12032 13676 12038 13728
rect 12544 13716 12572 13756
rect 13357 13753 13369 13787
rect 13403 13784 13415 13787
rect 13954 13787 14012 13793
rect 13954 13784 13966 13787
rect 13403 13756 13966 13784
rect 13403 13753 13415 13756
rect 13357 13747 13415 13753
rect 13954 13753 13966 13756
rect 14000 13784 14012 13787
rect 14826 13784 14832 13796
rect 14000 13756 14832 13784
rect 14000 13753 14012 13756
rect 13954 13747 14012 13753
rect 14826 13744 14832 13756
rect 14884 13744 14890 13796
rect 15102 13744 15108 13796
rect 15160 13784 15166 13796
rect 15304 13784 15332 13892
rect 15746 13880 15752 13892
rect 15804 13880 15810 13932
rect 19794 13880 19800 13932
rect 19852 13920 19858 13932
rect 20824 13920 20852 13948
rect 21085 13923 21143 13929
rect 21085 13920 21097 13923
rect 19852 13892 21097 13920
rect 19852 13880 19858 13892
rect 21085 13889 21097 13892
rect 21131 13889 21143 13923
rect 21085 13883 21143 13889
rect 16758 13812 16764 13864
rect 16816 13852 16822 13864
rect 17012 13855 17070 13861
rect 17012 13852 17024 13855
rect 16816 13824 17024 13852
rect 16816 13812 16822 13824
rect 17012 13821 17024 13824
rect 17058 13852 17070 13855
rect 17405 13855 17463 13861
rect 17405 13852 17417 13855
rect 17058 13824 17417 13852
rect 17058 13821 17070 13824
rect 17012 13815 17070 13821
rect 17405 13821 17417 13824
rect 17451 13821 17463 13855
rect 18046 13852 18052 13864
rect 18007 13824 18052 13852
rect 17405 13815 17463 13821
rect 18046 13812 18052 13824
rect 18104 13852 18110 13864
rect 18414 13852 18420 13864
rect 18104 13824 18420 13852
rect 18104 13812 18110 13824
rect 18414 13812 18420 13824
rect 18472 13812 18478 13864
rect 18601 13855 18659 13861
rect 18601 13852 18613 13855
rect 18524 13824 18613 13852
rect 15160 13756 15332 13784
rect 15473 13787 15531 13793
rect 15160 13744 15166 13756
rect 15473 13753 15485 13787
rect 15519 13753 15531 13787
rect 15473 13747 15531 13753
rect 12618 13716 12624 13728
rect 12544 13688 12624 13716
rect 12618 13676 12624 13688
rect 12676 13676 12682 13728
rect 13630 13676 13636 13728
rect 13688 13716 13694 13728
rect 14921 13719 14979 13725
rect 14921 13716 14933 13719
rect 13688 13688 14933 13716
rect 13688 13676 13694 13688
rect 14921 13685 14933 13688
rect 14967 13716 14979 13719
rect 15194 13716 15200 13728
rect 14967 13688 15200 13716
rect 14967 13685 14979 13688
rect 14921 13679 14979 13685
rect 15194 13676 15200 13688
rect 15252 13716 15258 13728
rect 15289 13719 15347 13725
rect 15289 13716 15301 13719
rect 15252 13688 15301 13716
rect 15252 13676 15258 13688
rect 15289 13685 15301 13688
rect 15335 13716 15347 13719
rect 15378 13716 15384 13728
rect 15335 13688 15384 13716
rect 15335 13685 15347 13688
rect 15289 13679 15347 13685
rect 15378 13676 15384 13688
rect 15436 13676 15442 13728
rect 15488 13716 15516 13747
rect 15562 13744 15568 13796
rect 15620 13784 15626 13796
rect 17586 13784 17592 13796
rect 15620 13756 15665 13784
rect 16776 13756 17592 13784
rect 15620 13744 15626 13756
rect 15930 13716 15936 13728
rect 15488 13688 15936 13716
rect 15930 13676 15936 13688
rect 15988 13676 15994 13728
rect 16390 13716 16396 13728
rect 16351 13688 16396 13716
rect 16390 13676 16396 13688
rect 16448 13716 16454 13728
rect 16776 13725 16804 13756
rect 17586 13744 17592 13756
rect 17644 13784 17650 13796
rect 17773 13787 17831 13793
rect 17773 13784 17785 13787
rect 17644 13756 17785 13784
rect 17644 13744 17650 13756
rect 17773 13753 17785 13756
rect 17819 13784 17831 13787
rect 18524 13784 18552 13824
rect 18601 13821 18613 13824
rect 18647 13852 18659 13855
rect 19058 13852 19064 13864
rect 18647 13824 19064 13852
rect 18647 13821 18659 13824
rect 18601 13815 18659 13821
rect 19058 13812 19064 13824
rect 19116 13812 19122 13864
rect 20809 13855 20867 13861
rect 20809 13821 20821 13855
rect 20855 13852 20867 13855
rect 21174 13852 21180 13864
rect 20855 13824 21180 13852
rect 20855 13821 20867 13824
rect 20809 13815 20867 13821
rect 21174 13812 21180 13824
rect 21232 13812 21238 13864
rect 18782 13784 18788 13796
rect 17819 13756 18552 13784
rect 18743 13756 18788 13784
rect 17819 13753 17831 13756
rect 17773 13747 17831 13753
rect 18782 13744 18788 13756
rect 18840 13744 18846 13796
rect 20162 13784 20168 13796
rect 20123 13756 20168 13784
rect 20162 13744 20168 13756
rect 20220 13744 20226 13796
rect 20257 13787 20315 13793
rect 20257 13753 20269 13787
rect 20303 13753 20315 13787
rect 20257 13747 20315 13753
rect 16761 13719 16819 13725
rect 16761 13716 16773 13719
rect 16448 13688 16773 13716
rect 16448 13676 16454 13688
rect 16761 13685 16773 13688
rect 16807 13685 16819 13719
rect 16761 13679 16819 13685
rect 16850 13676 16856 13728
rect 16908 13716 16914 13728
rect 17083 13719 17141 13725
rect 17083 13716 17095 13719
rect 16908 13688 17095 13716
rect 16908 13676 16914 13688
rect 17083 13685 17095 13688
rect 17129 13685 17141 13719
rect 19978 13716 19984 13728
rect 19891 13688 19984 13716
rect 17083 13679 17141 13685
rect 19978 13676 19984 13688
rect 20036 13716 20042 13728
rect 20272 13716 20300 13747
rect 20036 13688 20300 13716
rect 20036 13676 20042 13688
rect 1104 13626 22816 13648
rect 1104 13574 8982 13626
rect 9034 13574 9046 13626
rect 9098 13574 9110 13626
rect 9162 13574 9174 13626
rect 9226 13574 16982 13626
rect 17034 13574 17046 13626
rect 17098 13574 17110 13626
rect 17162 13574 17174 13626
rect 17226 13574 22816 13626
rect 1104 13552 22816 13574
rect 5534 13512 5540 13524
rect 4126 13484 5540 13512
rect 2774 13444 2780 13456
rect 2687 13416 2780 13444
rect 2700 13385 2728 13416
rect 2774 13404 2780 13416
rect 2832 13444 2838 13456
rect 4126 13444 4154 13484
rect 5534 13472 5540 13484
rect 5592 13472 5598 13524
rect 6822 13512 6828 13524
rect 6783 13484 6828 13512
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 7466 13472 7472 13524
rect 7524 13512 7530 13524
rect 7653 13515 7711 13521
rect 7653 13512 7665 13515
rect 7524 13484 7665 13512
rect 7524 13472 7530 13484
rect 7653 13481 7665 13484
rect 7699 13481 7711 13515
rect 7653 13475 7711 13481
rect 9033 13515 9091 13521
rect 9033 13481 9045 13515
rect 9079 13512 9091 13515
rect 9306 13512 9312 13524
rect 9079 13484 9312 13512
rect 9079 13481 9091 13484
rect 9033 13475 9091 13481
rect 9306 13472 9312 13484
rect 9364 13472 9370 13524
rect 9674 13472 9680 13524
rect 9732 13512 9738 13524
rect 9861 13515 9919 13521
rect 9861 13512 9873 13515
rect 9732 13484 9873 13512
rect 9732 13472 9738 13484
rect 9861 13481 9873 13484
rect 9907 13481 9919 13515
rect 9861 13475 9919 13481
rect 10870 13472 10876 13524
rect 10928 13512 10934 13524
rect 11057 13515 11115 13521
rect 11057 13512 11069 13515
rect 10928 13484 11069 13512
rect 10928 13472 10934 13484
rect 11057 13481 11069 13484
rect 11103 13512 11115 13515
rect 11606 13512 11612 13524
rect 11103 13484 11284 13512
rect 11567 13484 11612 13512
rect 11103 13481 11115 13484
rect 11057 13475 11115 13481
rect 2832 13416 4154 13444
rect 2832 13404 2838 13416
rect 4246 13404 4252 13456
rect 4304 13444 4310 13456
rect 4427 13447 4485 13453
rect 4427 13444 4439 13447
rect 4304 13416 4439 13444
rect 4304 13404 4310 13416
rect 4427 13413 4439 13416
rect 4473 13413 4485 13447
rect 4427 13407 4485 13413
rect 7006 13404 7012 13456
rect 7064 13444 7070 13456
rect 9950 13444 9956 13456
rect 7064 13416 9956 13444
rect 7064 13404 7070 13416
rect 9950 13404 9956 13416
rect 10008 13404 10014 13456
rect 2685 13379 2743 13385
rect 2685 13345 2697 13379
rect 2731 13345 2743 13379
rect 2685 13339 2743 13345
rect 2869 13379 2927 13385
rect 2869 13345 2881 13379
rect 2915 13345 2927 13379
rect 2869 13339 2927 13345
rect 7377 13379 7435 13385
rect 7377 13345 7389 13379
rect 7423 13376 7435 13379
rect 7558 13376 7564 13388
rect 7423 13348 7564 13376
rect 7423 13345 7435 13348
rect 7377 13339 7435 13345
rect 2590 13268 2596 13320
rect 2648 13308 2654 13320
rect 2884 13308 2912 13339
rect 7558 13336 7564 13348
rect 7616 13336 7622 13388
rect 8272 13379 8330 13385
rect 8272 13345 8284 13379
rect 8318 13376 8330 13379
rect 8478 13376 8484 13388
rect 8318 13348 8484 13376
rect 8318 13345 8330 13348
rect 8272 13339 8330 13345
rect 8478 13336 8484 13348
rect 8536 13336 8542 13388
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13376 10195 13379
rect 10318 13376 10324 13388
rect 10183 13348 10324 13376
rect 10183 13345 10195 13348
rect 10137 13339 10195 13345
rect 10318 13336 10324 13348
rect 10376 13336 10382 13388
rect 11256 13385 11284 13484
rect 11606 13472 11612 13484
rect 11664 13472 11670 13524
rect 12158 13512 12164 13524
rect 12119 13484 12164 13512
rect 12158 13472 12164 13484
rect 12216 13472 12222 13524
rect 13722 13472 13728 13524
rect 13780 13512 13786 13524
rect 14369 13515 14427 13521
rect 14369 13512 14381 13515
rect 13780 13484 14381 13512
rect 13780 13472 13786 13484
rect 14369 13481 14381 13484
rect 14415 13481 14427 13515
rect 15562 13512 15568 13524
rect 15523 13484 15568 13512
rect 14369 13475 14427 13481
rect 15562 13472 15568 13484
rect 15620 13472 15626 13524
rect 15930 13512 15936 13524
rect 15843 13484 15936 13512
rect 15930 13472 15936 13484
rect 15988 13512 15994 13524
rect 16850 13512 16856 13524
rect 15988 13484 16856 13512
rect 15988 13472 15994 13484
rect 16850 13472 16856 13484
rect 16908 13472 16914 13524
rect 17310 13512 17316 13524
rect 17271 13484 17316 13512
rect 17310 13472 17316 13484
rect 17368 13472 17374 13524
rect 17678 13472 17684 13524
rect 17736 13512 17742 13524
rect 18141 13515 18199 13521
rect 18141 13512 18153 13515
rect 17736 13484 18153 13512
rect 17736 13472 17742 13484
rect 18141 13481 18153 13484
rect 18187 13512 18199 13515
rect 18598 13512 18604 13524
rect 18187 13484 18604 13512
rect 18187 13481 18199 13484
rect 18141 13475 18199 13481
rect 18598 13472 18604 13484
rect 18656 13472 18662 13524
rect 19978 13512 19984 13524
rect 19939 13484 19984 13512
rect 19978 13472 19984 13484
rect 20036 13472 20042 13524
rect 12342 13404 12348 13456
rect 12400 13444 12406 13456
rect 13173 13447 13231 13453
rect 13173 13444 13185 13447
rect 12400 13416 13185 13444
rect 12400 13404 12406 13416
rect 13173 13413 13185 13416
rect 13219 13444 13231 13447
rect 13446 13444 13452 13456
rect 13219 13416 13452 13444
rect 13219 13413 13231 13416
rect 13173 13407 13231 13413
rect 13446 13404 13452 13416
rect 13504 13404 13510 13456
rect 16298 13404 16304 13456
rect 16356 13444 16362 13456
rect 16438 13447 16496 13453
rect 16438 13444 16450 13447
rect 16356 13416 16450 13444
rect 16356 13404 16362 13416
rect 16438 13413 16450 13416
rect 16484 13413 16496 13447
rect 16438 13407 16496 13413
rect 19058 13404 19064 13456
rect 19116 13444 19122 13456
rect 19382 13447 19440 13453
rect 19382 13444 19394 13447
rect 19116 13416 19394 13444
rect 19116 13404 19122 13416
rect 19382 13413 19394 13416
rect 19428 13413 19440 13447
rect 19382 13407 19440 13413
rect 20806 13404 20812 13456
rect 20864 13444 20870 13456
rect 21085 13447 21143 13453
rect 21085 13444 21097 13447
rect 20864 13416 21097 13444
rect 20864 13404 20870 13416
rect 21085 13413 21097 13416
rect 21131 13413 21143 13447
rect 21085 13407 21143 13413
rect 11241 13379 11299 13385
rect 11241 13345 11253 13379
rect 11287 13345 11299 13379
rect 16114 13376 16120 13388
rect 16075 13348 16120 13376
rect 11241 13339 11299 13345
rect 16114 13336 16120 13348
rect 16172 13336 16178 13388
rect 3142 13308 3148 13320
rect 2648 13280 2912 13308
rect 3103 13280 3148 13308
rect 2648 13268 2654 13280
rect 3142 13268 3148 13280
rect 3200 13308 3206 13320
rect 4065 13311 4123 13317
rect 4065 13308 4077 13311
rect 3200 13280 4077 13308
rect 3200 13268 3206 13280
rect 4065 13277 4077 13280
rect 4111 13277 4123 13311
rect 4065 13271 4123 13277
rect 6178 13268 6184 13320
rect 6236 13308 6242 13320
rect 6457 13311 6515 13317
rect 6457 13308 6469 13311
rect 6236 13280 6469 13308
rect 6236 13268 6242 13280
rect 6457 13277 6469 13280
rect 6503 13277 6515 13311
rect 6457 13271 6515 13277
rect 12802 13268 12808 13320
rect 12860 13308 12866 13320
rect 13081 13311 13139 13317
rect 13081 13308 13093 13311
rect 12860 13280 13093 13308
rect 12860 13268 12866 13280
rect 13081 13277 13093 13280
rect 13127 13277 13139 13311
rect 13354 13308 13360 13320
rect 13315 13280 13360 13308
rect 13081 13271 13139 13277
rect 13354 13268 13360 13280
rect 13412 13268 13418 13320
rect 19061 13311 19119 13317
rect 19061 13277 19073 13311
rect 19107 13308 19119 13311
rect 19242 13308 19248 13320
rect 19107 13280 19248 13308
rect 19107 13277 19119 13280
rect 19061 13271 19119 13277
rect 19242 13268 19248 13280
rect 19300 13308 19306 13320
rect 20254 13308 20260 13320
rect 19300 13280 20260 13308
rect 19300 13268 19306 13280
rect 20254 13268 20260 13280
rect 20312 13268 20318 13320
rect 20714 13268 20720 13320
rect 20772 13308 20778 13320
rect 20993 13311 21051 13317
rect 20993 13308 21005 13311
rect 20772 13280 21005 13308
rect 20772 13268 20778 13280
rect 20993 13277 21005 13280
rect 21039 13277 21051 13311
rect 20993 13271 21051 13277
rect 21174 13268 21180 13320
rect 21232 13308 21238 13320
rect 21269 13311 21327 13317
rect 21269 13308 21281 13311
rect 21232 13280 21281 13308
rect 21232 13268 21238 13280
rect 21269 13277 21281 13280
rect 21315 13277 21327 13311
rect 21269 13271 21327 13277
rect 4522 13200 4528 13252
rect 4580 13240 4586 13252
rect 5261 13243 5319 13249
rect 5261 13240 5273 13243
rect 4580 13212 5273 13240
rect 4580 13200 4586 13212
rect 5261 13209 5273 13212
rect 5307 13209 5319 13243
rect 5261 13203 5319 13209
rect 10367 13243 10425 13249
rect 10367 13209 10379 13243
rect 10413 13240 10425 13243
rect 13906 13240 13912 13252
rect 10413 13212 13912 13240
rect 10413 13209 10425 13212
rect 10367 13203 10425 13209
rect 13906 13200 13912 13212
rect 13964 13200 13970 13252
rect 1394 13132 1400 13184
rect 1452 13172 1458 13184
rect 1670 13172 1676 13184
rect 1452 13144 1676 13172
rect 1452 13132 1458 13144
rect 1670 13132 1676 13144
rect 1728 13132 1734 13184
rect 4614 13132 4620 13184
rect 4672 13172 4678 13184
rect 4985 13175 5043 13181
rect 4985 13172 4997 13175
rect 4672 13144 4997 13172
rect 4672 13132 4678 13144
rect 4985 13141 4997 13144
rect 5031 13172 5043 13175
rect 5442 13172 5448 13184
rect 5031 13144 5448 13172
rect 5031 13141 5043 13144
rect 4985 13135 5043 13141
rect 5442 13132 5448 13144
rect 5500 13132 5506 13184
rect 7466 13132 7472 13184
rect 7524 13172 7530 13184
rect 8113 13175 8171 13181
rect 8113 13172 8125 13175
rect 7524 13144 8125 13172
rect 7524 13132 7530 13144
rect 8113 13141 8125 13144
rect 8159 13172 8171 13175
rect 8343 13175 8401 13181
rect 8343 13172 8355 13175
rect 8159 13144 8355 13172
rect 8159 13141 8171 13144
rect 8113 13135 8171 13141
rect 8343 13141 8355 13144
rect 8389 13141 8401 13175
rect 10778 13172 10784 13184
rect 10739 13144 10784 13172
rect 8343 13135 8401 13141
rect 10778 13132 10784 13144
rect 10836 13132 10842 13184
rect 12434 13172 12440 13184
rect 12395 13144 12440 13172
rect 12434 13132 12440 13144
rect 12492 13132 12498 13184
rect 13998 13172 14004 13184
rect 13959 13144 14004 13172
rect 13998 13132 14004 13144
rect 14056 13132 14062 13184
rect 16574 13132 16580 13184
rect 16632 13172 16638 13184
rect 17037 13175 17095 13181
rect 17037 13172 17049 13175
rect 16632 13144 17049 13172
rect 16632 13132 16638 13144
rect 17037 13141 17049 13144
rect 17083 13141 17095 13175
rect 17037 13135 17095 13141
rect 1104 13082 22816 13104
rect 1104 13030 4982 13082
rect 5034 13030 5046 13082
rect 5098 13030 5110 13082
rect 5162 13030 5174 13082
rect 5226 13030 12982 13082
rect 13034 13030 13046 13082
rect 13098 13030 13110 13082
rect 13162 13030 13174 13082
rect 13226 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 22816 13082
rect 1104 13008 22816 13030
rect 2774 12968 2780 12980
rect 2735 12940 2780 12968
rect 2774 12928 2780 12940
rect 2832 12928 2838 12980
rect 3142 12928 3148 12980
rect 3200 12968 3206 12980
rect 3237 12971 3295 12977
rect 3237 12968 3249 12971
rect 3200 12940 3249 12968
rect 3200 12928 3206 12940
rect 3237 12937 3249 12940
rect 3283 12937 3295 12971
rect 5442 12968 5448 12980
rect 5403 12940 5448 12968
rect 3237 12931 3295 12937
rect 5442 12928 5448 12940
rect 5500 12928 5506 12980
rect 7285 12971 7343 12977
rect 7285 12937 7297 12971
rect 7331 12968 7343 12971
rect 7558 12968 7564 12980
rect 7331 12940 7564 12968
rect 7331 12937 7343 12940
rect 7285 12931 7343 12937
rect 7558 12928 7564 12940
rect 7616 12928 7622 12980
rect 13446 12968 13452 12980
rect 13407 12940 13452 12968
rect 13446 12928 13452 12940
rect 13504 12928 13510 12980
rect 13633 12971 13691 12977
rect 13633 12937 13645 12971
rect 13679 12968 13691 12971
rect 13998 12968 14004 12980
rect 13679 12940 14004 12968
rect 13679 12937 13691 12940
rect 13633 12931 13691 12937
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 15841 12971 15899 12977
rect 15841 12937 15853 12971
rect 15887 12968 15899 12971
rect 16114 12968 16120 12980
rect 15887 12940 16120 12968
rect 15887 12937 15899 12940
rect 15841 12931 15899 12937
rect 16114 12928 16120 12940
rect 16172 12928 16178 12980
rect 16298 12928 16304 12980
rect 16356 12968 16362 12980
rect 18877 12971 18935 12977
rect 18877 12968 18889 12971
rect 16356 12940 18889 12968
rect 16356 12928 16362 12940
rect 18877 12937 18889 12940
rect 18923 12968 18935 12971
rect 19058 12968 19064 12980
rect 18923 12940 19064 12968
rect 18923 12937 18935 12940
rect 18877 12931 18935 12937
rect 19058 12928 19064 12940
rect 19116 12928 19122 12980
rect 19981 12971 20039 12977
rect 19981 12937 19993 12971
rect 20027 12968 20039 12971
rect 20806 12968 20812 12980
rect 20027 12940 20812 12968
rect 20027 12937 20039 12940
rect 19981 12931 20039 12937
rect 20806 12928 20812 12940
rect 20864 12928 20870 12980
rect 21085 12971 21143 12977
rect 21085 12937 21097 12971
rect 21131 12968 21143 12971
rect 21358 12968 21364 12980
rect 21131 12940 21364 12968
rect 21131 12937 21143 12940
rect 21085 12931 21143 12937
rect 21358 12928 21364 12940
rect 21416 12928 21422 12980
rect 6362 12860 6368 12912
rect 6420 12900 6426 12912
rect 8570 12900 8576 12912
rect 6420 12872 8576 12900
rect 6420 12860 6426 12872
rect 8570 12860 8576 12872
rect 8628 12900 8634 12912
rect 10502 12900 10508 12912
rect 8628 12872 10508 12900
rect 8628 12860 8634 12872
rect 10502 12860 10508 12872
rect 10560 12860 10566 12912
rect 12526 12860 12532 12912
rect 12584 12900 12590 12912
rect 13081 12903 13139 12909
rect 13081 12900 13093 12903
rect 12584 12872 13093 12900
rect 12584 12860 12590 12872
rect 13081 12869 13093 12872
rect 13127 12900 13139 12903
rect 14645 12903 14703 12909
rect 14645 12900 14657 12903
rect 13127 12872 14657 12900
rect 13127 12869 13139 12872
rect 13081 12863 13139 12869
rect 14645 12869 14657 12872
rect 14691 12900 14703 12903
rect 15746 12900 15752 12912
rect 14691 12872 15752 12900
rect 14691 12869 14703 12872
rect 14645 12863 14703 12869
rect 15746 12860 15752 12872
rect 15804 12860 15810 12912
rect 15930 12860 15936 12912
rect 15988 12900 15994 12912
rect 17310 12900 17316 12912
rect 15988 12872 17316 12900
rect 15988 12860 15994 12872
rect 17310 12860 17316 12872
rect 17368 12860 17374 12912
rect 20254 12900 20260 12912
rect 20215 12872 20260 12900
rect 20254 12860 20260 12872
rect 20312 12860 20318 12912
rect 3559 12835 3617 12841
rect 3559 12801 3571 12835
rect 3605 12832 3617 12835
rect 4522 12832 4528 12844
rect 3605 12804 4528 12832
rect 3605 12801 3617 12804
rect 3559 12795 3617 12801
rect 4522 12792 4528 12804
rect 4580 12792 4586 12844
rect 7466 12832 7472 12844
rect 7427 12804 7472 12832
rect 7466 12792 7472 12804
rect 7524 12792 7530 12844
rect 8754 12792 8760 12844
rect 8812 12832 8818 12844
rect 9309 12835 9367 12841
rect 9309 12832 9321 12835
rect 8812 12804 9321 12832
rect 8812 12792 8818 12804
rect 9309 12801 9321 12804
rect 9355 12801 9367 12835
rect 9309 12795 9367 12801
rect 10778 12792 10784 12844
rect 10836 12832 10842 12844
rect 13633 12835 13691 12841
rect 13633 12832 13645 12835
rect 10836 12804 13645 12832
rect 10836 12792 10842 12804
rect 1670 12724 1676 12776
rect 1728 12764 1734 12776
rect 10980 12773 11008 12804
rect 13633 12801 13645 12804
rect 13679 12801 13691 12835
rect 13633 12795 13691 12801
rect 13906 12792 13912 12844
rect 13964 12832 13970 12844
rect 14093 12835 14151 12841
rect 14093 12832 14105 12835
rect 13964 12804 14105 12832
rect 13964 12792 13970 12804
rect 14093 12801 14105 12804
rect 14139 12832 14151 12835
rect 15013 12835 15071 12841
rect 15013 12832 15025 12835
rect 14139 12804 15025 12832
rect 14139 12801 14151 12804
rect 14093 12795 14151 12801
rect 15013 12801 15025 12804
rect 15059 12801 15071 12835
rect 16482 12832 16488 12844
rect 16395 12804 16488 12832
rect 15013 12795 15071 12801
rect 16482 12792 16488 12804
rect 16540 12832 16546 12844
rect 17405 12835 17463 12841
rect 17405 12832 17417 12835
rect 16540 12804 17417 12832
rect 16540 12792 16546 12804
rect 17405 12801 17417 12804
rect 17451 12801 17463 12835
rect 17405 12795 17463 12801
rect 18782 12792 18788 12844
rect 18840 12832 18846 12844
rect 19061 12835 19119 12841
rect 19061 12832 19073 12835
rect 18840 12804 19073 12832
rect 18840 12792 18846 12804
rect 19061 12801 19073 12804
rect 19107 12801 19119 12835
rect 19061 12795 19119 12801
rect 3472 12767 3530 12773
rect 3472 12764 3484 12767
rect 1728 12736 3484 12764
rect 1728 12724 1734 12736
rect 3472 12733 3484 12736
rect 3518 12764 3530 12767
rect 10965 12767 11023 12773
rect 3518 12736 4016 12764
rect 3518 12733 3530 12736
rect 3472 12727 3530 12733
rect 3988 12640 4016 12736
rect 10965 12733 10977 12767
rect 11011 12733 11023 12767
rect 10965 12727 11023 12733
rect 11241 12767 11299 12773
rect 11241 12733 11253 12767
rect 11287 12733 11299 12767
rect 11422 12764 11428 12776
rect 11383 12736 11428 12764
rect 11241 12727 11299 12733
rect 4614 12696 4620 12708
rect 4575 12668 4620 12696
rect 4614 12656 4620 12668
rect 4672 12656 4678 12708
rect 5166 12696 5172 12708
rect 5127 12668 5172 12696
rect 5166 12656 5172 12668
rect 5224 12656 5230 12708
rect 7558 12696 7564 12708
rect 7519 12668 7564 12696
rect 7558 12656 7564 12668
rect 7616 12656 7622 12708
rect 8113 12699 8171 12705
rect 8113 12665 8125 12699
rect 8159 12696 8171 12699
rect 8202 12696 8208 12708
rect 8159 12668 8208 12696
rect 8159 12665 8171 12668
rect 8113 12659 8171 12665
rect 8202 12656 8208 12668
rect 8260 12656 8266 12708
rect 8846 12656 8852 12708
rect 8904 12696 8910 12708
rect 9033 12699 9091 12705
rect 9033 12696 9045 12699
rect 8904 12668 9045 12696
rect 8904 12656 8910 12668
rect 9033 12665 9045 12668
rect 9079 12665 9091 12699
rect 9033 12659 9091 12665
rect 9125 12699 9183 12705
rect 9125 12665 9137 12699
rect 9171 12665 9183 12699
rect 9125 12659 9183 12665
rect 2501 12631 2559 12637
rect 2501 12597 2513 12631
rect 2547 12628 2559 12631
rect 2590 12628 2596 12640
rect 2547 12600 2596 12628
rect 2547 12597 2559 12600
rect 2501 12591 2559 12597
rect 2590 12588 2596 12600
rect 2648 12588 2654 12640
rect 3970 12628 3976 12640
rect 3931 12600 3976 12628
rect 3970 12588 3976 12600
rect 4028 12588 4034 12640
rect 4341 12631 4399 12637
rect 4341 12597 4353 12631
rect 4387 12628 4399 12631
rect 4522 12628 4528 12640
rect 4387 12600 4528 12628
rect 4387 12597 4399 12600
rect 4341 12591 4399 12597
rect 4522 12588 4528 12600
rect 4580 12588 4586 12640
rect 6178 12628 6184 12640
rect 6139 12600 6184 12628
rect 6178 12588 6184 12600
rect 6236 12588 6242 12640
rect 6549 12631 6607 12637
rect 6549 12597 6561 12631
rect 6595 12628 6607 12631
rect 6822 12628 6828 12640
rect 6595 12600 6828 12628
rect 6595 12597 6607 12600
rect 6549 12591 6607 12597
rect 6822 12588 6828 12600
rect 6880 12628 6886 12640
rect 7466 12628 7472 12640
rect 6880 12600 7472 12628
rect 6880 12588 6886 12600
rect 7466 12588 7472 12600
rect 7524 12588 7530 12640
rect 8478 12628 8484 12640
rect 8439 12600 8484 12628
rect 8478 12588 8484 12600
rect 8536 12588 8542 12640
rect 8754 12628 8760 12640
rect 8667 12600 8760 12628
rect 8754 12588 8760 12600
rect 8812 12628 8818 12640
rect 9140 12628 9168 12659
rect 11054 12656 11060 12708
rect 11112 12696 11118 12708
rect 11256 12696 11284 12727
rect 11422 12724 11428 12736
rect 11480 12724 11486 12776
rect 11790 12764 11796 12776
rect 11618 12736 11796 12764
rect 11618 12696 11646 12736
rect 11790 12724 11796 12736
rect 11848 12724 11854 12776
rect 14826 12724 14832 12776
rect 14884 12764 14890 12776
rect 16117 12767 16175 12773
rect 16117 12764 16129 12767
rect 14884 12736 16129 12764
rect 14884 12724 14890 12736
rect 16117 12733 16129 12736
rect 16163 12764 16175 12767
rect 16298 12764 16304 12776
rect 16163 12736 16304 12764
rect 16163 12733 16175 12736
rect 16117 12727 16175 12733
rect 16298 12724 16304 12736
rect 16356 12724 16362 12776
rect 18084 12767 18142 12773
rect 18084 12764 18096 12767
rect 17788 12736 18096 12764
rect 12526 12696 12532 12708
rect 11112 12668 11646 12696
rect 12487 12668 12532 12696
rect 11112 12656 11118 12668
rect 12526 12656 12532 12668
rect 12584 12656 12590 12708
rect 12621 12699 12679 12705
rect 12621 12665 12633 12699
rect 12667 12665 12679 12699
rect 12621 12659 12679 12665
rect 14185 12699 14243 12705
rect 14185 12665 14197 12699
rect 14231 12665 14243 12699
rect 14185 12659 14243 12665
rect 10318 12628 10324 12640
rect 8812 12600 9168 12628
rect 10279 12600 10324 12628
rect 8812 12588 8818 12600
rect 10318 12588 10324 12600
rect 10376 12588 10382 12640
rect 10686 12588 10692 12640
rect 10744 12628 10750 12640
rect 11606 12628 11612 12640
rect 10744 12600 11612 12628
rect 10744 12588 10750 12600
rect 11606 12588 11612 12600
rect 11664 12628 11670 12640
rect 11701 12631 11759 12637
rect 11701 12628 11713 12631
rect 11664 12600 11713 12628
rect 11664 12588 11670 12600
rect 11701 12597 11713 12600
rect 11747 12597 11759 12631
rect 11701 12591 11759 12597
rect 11790 12588 11796 12640
rect 11848 12628 11854 12640
rect 12253 12631 12311 12637
rect 12253 12628 12265 12631
rect 11848 12600 12265 12628
rect 11848 12588 11854 12600
rect 12253 12597 12265 12600
rect 12299 12628 12311 12631
rect 12636 12628 12664 12659
rect 13906 12628 13912 12640
rect 12299 12600 12664 12628
rect 13867 12600 13912 12628
rect 12299 12597 12311 12600
rect 12253 12591 12311 12597
rect 13906 12588 13912 12600
rect 13964 12628 13970 12640
rect 14200 12628 14228 12659
rect 15102 12656 15108 12708
rect 15160 12696 15166 12708
rect 16574 12696 16580 12708
rect 15160 12668 16481 12696
rect 16535 12668 16580 12696
rect 15160 12656 15166 12668
rect 13964 12600 14228 12628
rect 16453 12628 16481 12668
rect 16574 12656 16580 12668
rect 16632 12656 16638 12708
rect 17129 12699 17187 12705
rect 17129 12665 17141 12699
rect 17175 12696 17187 12699
rect 17310 12696 17316 12708
rect 17175 12668 17316 12696
rect 17175 12665 17187 12668
rect 17129 12659 17187 12665
rect 17310 12656 17316 12668
rect 17368 12656 17374 12708
rect 17788 12628 17816 12736
rect 18084 12733 18096 12736
rect 18130 12764 18142 12767
rect 18509 12767 18567 12773
rect 18509 12764 18521 12767
rect 18130 12736 18521 12764
rect 18130 12733 18142 12736
rect 18084 12727 18142 12733
rect 18509 12733 18521 12736
rect 18555 12764 18567 12767
rect 20901 12767 20959 12773
rect 20901 12764 20913 12767
rect 18555 12736 20913 12764
rect 18555 12733 18567 12736
rect 18509 12727 18567 12733
rect 20901 12733 20913 12736
rect 20947 12764 20959 12767
rect 21453 12767 21511 12773
rect 21453 12764 21465 12767
rect 20947 12736 21465 12764
rect 20947 12733 20959 12736
rect 20901 12727 20959 12733
rect 21453 12733 21465 12736
rect 21499 12764 21511 12767
rect 21542 12764 21548 12776
rect 21499 12736 21548 12764
rect 21499 12733 21511 12736
rect 21453 12727 21511 12733
rect 21542 12724 21548 12736
rect 21600 12724 21606 12776
rect 19058 12656 19064 12708
rect 19116 12696 19122 12708
rect 19382 12699 19440 12705
rect 19382 12696 19394 12699
rect 19116 12668 19394 12696
rect 19116 12656 19122 12668
rect 19382 12665 19394 12668
rect 19428 12665 19440 12699
rect 19382 12659 19440 12665
rect 16453 12600 17816 12628
rect 13964 12588 13970 12600
rect 17862 12588 17868 12640
rect 17920 12628 17926 12640
rect 18187 12631 18245 12637
rect 18187 12628 18199 12631
rect 17920 12600 18199 12628
rect 17920 12588 17926 12600
rect 18187 12597 18199 12600
rect 18233 12597 18245 12631
rect 18187 12591 18245 12597
rect 1104 12538 22816 12560
rect 1104 12486 8982 12538
rect 9034 12486 9046 12538
rect 9098 12486 9110 12538
rect 9162 12486 9174 12538
rect 9226 12486 16982 12538
rect 17034 12486 17046 12538
rect 17098 12486 17110 12538
rect 17162 12486 17174 12538
rect 17226 12486 22816 12538
rect 1104 12464 22816 12486
rect 6178 12424 6184 12436
rect 6139 12396 6184 12424
rect 6178 12384 6184 12396
rect 6236 12384 6242 12436
rect 8846 12384 8852 12436
rect 8904 12424 8910 12436
rect 9033 12427 9091 12433
rect 9033 12424 9045 12427
rect 8904 12396 9045 12424
rect 8904 12384 8910 12396
rect 9033 12393 9045 12396
rect 9079 12424 9091 12427
rect 9815 12427 9873 12433
rect 9815 12424 9827 12427
rect 9079 12396 9827 12424
rect 9079 12393 9091 12396
rect 9033 12387 9091 12393
rect 9815 12393 9827 12396
rect 9861 12393 9873 12427
rect 11054 12424 11060 12436
rect 11015 12396 11060 12424
rect 9815 12387 9873 12393
rect 11054 12384 11060 12396
rect 11112 12384 11118 12436
rect 15427 12427 15485 12433
rect 15427 12393 15439 12427
rect 15473 12424 15485 12427
rect 16482 12424 16488 12436
rect 15473 12396 16488 12424
rect 15473 12393 15485 12396
rect 15427 12387 15485 12393
rect 16482 12384 16488 12396
rect 16540 12384 16546 12436
rect 18782 12384 18788 12436
rect 18840 12424 18846 12436
rect 19797 12427 19855 12433
rect 19797 12424 19809 12427
rect 18840 12396 19809 12424
rect 18840 12384 18846 12396
rect 19797 12393 19809 12396
rect 19843 12393 19855 12427
rect 19797 12387 19855 12393
rect 20714 12384 20720 12436
rect 20772 12424 20778 12436
rect 21085 12427 21143 12433
rect 21085 12424 21097 12427
rect 20772 12396 21097 12424
rect 20772 12384 20778 12396
rect 21085 12393 21097 12396
rect 21131 12393 21143 12427
rect 21085 12387 21143 12393
rect 4522 12356 4528 12368
rect 4483 12328 4528 12356
rect 4522 12316 4528 12328
rect 4580 12316 4586 12368
rect 8205 12359 8263 12365
rect 8205 12325 8217 12359
rect 8251 12356 8263 12359
rect 8754 12356 8760 12368
rect 8251 12328 8760 12356
rect 8251 12325 8263 12328
rect 8205 12319 8263 12325
rect 8754 12316 8760 12328
rect 8812 12316 8818 12368
rect 11790 12356 11796 12368
rect 11751 12328 11796 12356
rect 11790 12316 11796 12328
rect 11848 12316 11854 12368
rect 12345 12359 12403 12365
rect 12345 12325 12357 12359
rect 12391 12356 12403 12359
rect 12802 12356 12808 12368
rect 12391 12328 12808 12356
rect 12391 12325 12403 12328
rect 12345 12319 12403 12325
rect 12802 12316 12808 12328
rect 12860 12356 12866 12368
rect 12989 12359 13047 12365
rect 12989 12356 13001 12359
rect 12860 12328 13001 12356
rect 12860 12316 12866 12328
rect 12989 12325 13001 12328
rect 13035 12325 13047 12359
rect 12989 12319 13047 12325
rect 13817 12359 13875 12365
rect 13817 12325 13829 12359
rect 13863 12356 13875 12359
rect 13906 12356 13912 12368
rect 13863 12328 13912 12356
rect 13863 12325 13875 12328
rect 13817 12319 13875 12325
rect 2498 12288 2504 12300
rect 2459 12260 2504 12288
rect 2498 12248 2504 12260
rect 2556 12248 2562 12300
rect 2590 12248 2596 12300
rect 2648 12288 2654 12300
rect 2869 12291 2927 12297
rect 2869 12288 2881 12291
rect 2648 12260 2881 12288
rect 2648 12248 2654 12260
rect 2869 12257 2881 12260
rect 2915 12257 2927 12291
rect 5902 12288 5908 12300
rect 5863 12260 5908 12288
rect 2869 12251 2927 12257
rect 5902 12248 5908 12260
rect 5960 12248 5966 12300
rect 6454 12288 6460 12300
rect 6415 12260 6460 12288
rect 6454 12248 6460 12260
rect 6512 12248 6518 12300
rect 9744 12291 9802 12297
rect 9744 12257 9756 12291
rect 9790 12288 9802 12291
rect 9950 12288 9956 12300
rect 9790 12260 9956 12288
rect 9790 12257 9802 12260
rect 9744 12251 9802 12257
rect 9950 12248 9956 12260
rect 10008 12248 10014 12300
rect 3142 12220 3148 12232
rect 3103 12192 3148 12220
rect 3142 12180 3148 12192
rect 3200 12180 3206 12232
rect 3878 12180 3884 12232
rect 3936 12220 3942 12232
rect 4430 12220 4436 12232
rect 3936 12192 4436 12220
rect 3936 12180 3942 12192
rect 4430 12180 4436 12192
rect 4488 12180 4494 12232
rect 4706 12220 4712 12232
rect 4667 12192 4712 12220
rect 4706 12180 4712 12192
rect 4764 12180 4770 12232
rect 8110 12220 8116 12232
rect 8071 12192 8116 12220
rect 8110 12180 8116 12192
rect 8168 12180 8174 12232
rect 8202 12180 8208 12232
rect 8260 12220 8266 12232
rect 8389 12223 8447 12229
rect 8389 12220 8401 12223
rect 8260 12192 8401 12220
rect 8260 12180 8266 12192
rect 8389 12189 8401 12192
rect 8435 12189 8447 12223
rect 8389 12183 8447 12189
rect 11701 12223 11759 12229
rect 11701 12189 11713 12223
rect 11747 12220 11759 12223
rect 12158 12220 12164 12232
rect 11747 12192 12164 12220
rect 11747 12189 11759 12192
rect 11701 12183 11759 12189
rect 12158 12180 12164 12192
rect 12216 12180 12222 12232
rect 4798 12112 4804 12164
rect 4856 12152 4862 12164
rect 5166 12152 5172 12164
rect 4856 12124 5172 12152
rect 4856 12112 4862 12124
rect 5166 12112 5172 12124
rect 5224 12152 5230 12164
rect 5445 12155 5503 12161
rect 5445 12152 5457 12155
rect 5224 12124 5457 12152
rect 5224 12112 5230 12124
rect 5445 12121 5457 12124
rect 5491 12152 5503 12155
rect 8220 12152 8248 12180
rect 5491 12124 8248 12152
rect 13004 12152 13032 12319
rect 13906 12316 13912 12328
rect 13964 12356 13970 12368
rect 14366 12356 14372 12368
rect 13964 12328 14372 12356
rect 13964 12316 13970 12328
rect 14366 12316 14372 12328
rect 14424 12316 14430 12368
rect 16393 12359 16451 12365
rect 16393 12325 16405 12359
rect 16439 12356 16451 12359
rect 16574 12356 16580 12368
rect 16439 12328 16580 12356
rect 16439 12325 16451 12328
rect 16393 12319 16451 12325
rect 16574 12316 16580 12328
rect 16632 12356 16638 12368
rect 17221 12359 17279 12365
rect 17221 12356 17233 12359
rect 16632 12328 17233 12356
rect 16632 12316 16638 12328
rect 17221 12325 17233 12328
rect 17267 12356 17279 12359
rect 17402 12356 17408 12368
rect 17267 12328 17408 12356
rect 17267 12325 17279 12328
rect 17221 12319 17279 12325
rect 17402 12316 17408 12328
rect 17460 12316 17466 12368
rect 17773 12359 17831 12365
rect 17773 12325 17785 12359
rect 17819 12356 17831 12359
rect 18598 12356 18604 12368
rect 17819 12328 18604 12356
rect 17819 12325 17831 12328
rect 17773 12319 17831 12325
rect 18598 12316 18604 12328
rect 18656 12356 18662 12368
rect 20732 12356 20760 12384
rect 18656 12328 20760 12356
rect 18656 12316 18662 12328
rect 15194 12248 15200 12300
rect 15252 12288 15258 12300
rect 15324 12291 15382 12297
rect 15324 12288 15336 12291
rect 15252 12260 15336 12288
rect 15252 12248 15258 12260
rect 15324 12257 15336 12260
rect 15370 12288 15382 12291
rect 16758 12288 16764 12300
rect 15370 12260 16764 12288
rect 15370 12257 15382 12260
rect 15324 12251 15382 12257
rect 16758 12248 16764 12260
rect 16816 12248 16822 12300
rect 19058 12288 19064 12300
rect 19019 12260 19064 12288
rect 19058 12248 19064 12260
rect 19116 12248 19122 12300
rect 19245 12291 19303 12297
rect 19245 12257 19257 12291
rect 19291 12288 19303 12291
rect 19334 12288 19340 12300
rect 19291 12260 19340 12288
rect 19291 12257 19303 12260
rect 19245 12251 19303 12257
rect 19334 12248 19340 12260
rect 19392 12248 19398 12300
rect 13722 12220 13728 12232
rect 13683 12192 13728 12220
rect 13722 12180 13728 12192
rect 13780 12180 13786 12232
rect 14369 12223 14427 12229
rect 14369 12189 14381 12223
rect 14415 12220 14427 12223
rect 14550 12220 14556 12232
rect 14415 12192 14556 12220
rect 14415 12189 14427 12192
rect 14369 12183 14427 12189
rect 14384 12152 14412 12183
rect 14550 12180 14556 12192
rect 14608 12180 14614 12232
rect 17129 12223 17187 12229
rect 17129 12189 17141 12223
rect 17175 12220 17187 12223
rect 17862 12220 17868 12232
rect 17175 12192 17868 12220
rect 17175 12189 17187 12192
rect 17129 12183 17187 12189
rect 17862 12180 17868 12192
rect 17920 12180 17926 12232
rect 13004 12124 14412 12152
rect 5491 12121 5503 12124
rect 5445 12115 5503 12121
rect 7742 12084 7748 12096
rect 7703 12056 7748 12084
rect 7742 12044 7748 12056
rect 7800 12044 7806 12096
rect 10686 12084 10692 12096
rect 10647 12056 10692 12084
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 11146 12044 11152 12096
rect 11204 12084 11210 12096
rect 11333 12087 11391 12093
rect 11333 12084 11345 12087
rect 11204 12056 11345 12084
rect 11204 12044 11210 12056
rect 11333 12053 11345 12056
rect 11379 12053 11391 12087
rect 13446 12084 13452 12096
rect 13407 12056 13452 12084
rect 11333 12047 11391 12053
rect 13446 12044 13452 12056
rect 13504 12044 13510 12096
rect 16758 12084 16764 12096
rect 16719 12056 16764 12084
rect 16758 12044 16764 12056
rect 16816 12044 16822 12096
rect 19475 12087 19533 12093
rect 19475 12053 19487 12087
rect 19521 12084 19533 12087
rect 19702 12084 19708 12096
rect 19521 12056 19708 12084
rect 19521 12053 19533 12056
rect 19475 12047 19533 12053
rect 19702 12044 19708 12056
rect 19760 12044 19766 12096
rect 1104 11994 22816 12016
rect 1104 11942 4982 11994
rect 5034 11942 5046 11994
rect 5098 11942 5110 11994
rect 5162 11942 5174 11994
rect 5226 11942 12982 11994
rect 13034 11942 13046 11994
rect 13098 11942 13110 11994
rect 13162 11942 13174 11994
rect 13226 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 22816 11994
rect 1104 11920 22816 11942
rect 4065 11883 4123 11889
rect 4065 11849 4077 11883
rect 4111 11880 4123 11883
rect 4433 11883 4491 11889
rect 4433 11880 4445 11883
rect 4111 11852 4445 11880
rect 4111 11849 4123 11852
rect 4065 11843 4123 11849
rect 4433 11849 4445 11852
rect 4479 11880 4491 11883
rect 4522 11880 4528 11892
rect 4479 11852 4528 11880
rect 4479 11849 4491 11852
rect 4433 11843 4491 11849
rect 4522 11840 4528 11852
rect 4580 11840 4586 11892
rect 5902 11840 5908 11892
rect 5960 11880 5966 11892
rect 6273 11883 6331 11889
rect 6273 11880 6285 11883
rect 5960 11852 6285 11880
rect 5960 11840 5966 11852
rect 6273 11849 6285 11852
rect 6319 11849 6331 11883
rect 6273 11843 6331 11849
rect 8573 11883 8631 11889
rect 8573 11849 8585 11883
rect 8619 11880 8631 11883
rect 8754 11880 8760 11892
rect 8619 11852 8760 11880
rect 8619 11849 8631 11852
rect 8573 11843 8631 11849
rect 8754 11840 8760 11852
rect 8812 11880 8818 11892
rect 8849 11883 8907 11889
rect 8849 11880 8861 11883
rect 8812 11852 8861 11880
rect 8812 11840 8818 11852
rect 8849 11849 8861 11852
rect 8895 11849 8907 11883
rect 8849 11843 8907 11849
rect 10321 11883 10379 11889
rect 10321 11849 10333 11883
rect 10367 11880 10379 11883
rect 10410 11880 10416 11892
rect 10367 11852 10416 11880
rect 10367 11849 10379 11852
rect 10321 11843 10379 11849
rect 3142 11744 3148 11756
rect 3103 11716 3148 11744
rect 3142 11704 3148 11716
rect 3200 11704 3206 11756
rect 4706 11704 4712 11756
rect 4764 11744 4770 11756
rect 5261 11747 5319 11753
rect 5261 11744 5273 11747
rect 4764 11716 5273 11744
rect 4764 11704 4770 11716
rect 5261 11713 5273 11716
rect 5307 11713 5319 11747
rect 5261 11707 5319 11713
rect 2133 11679 2191 11685
rect 2133 11645 2145 11679
rect 2179 11676 2191 11679
rect 2498 11676 2504 11688
rect 2179 11648 2504 11676
rect 2179 11645 2191 11648
rect 2133 11639 2191 11645
rect 2498 11636 2504 11648
rect 2556 11676 2562 11688
rect 3602 11676 3608 11688
rect 2556 11648 3608 11676
rect 2556 11636 2562 11648
rect 3602 11636 3608 11648
rect 3660 11636 3666 11688
rect 7653 11679 7711 11685
rect 7653 11645 7665 11679
rect 7699 11676 7711 11679
rect 7742 11676 7748 11688
rect 7699 11648 7748 11676
rect 7699 11645 7711 11648
rect 7653 11639 7711 11645
rect 7742 11636 7748 11648
rect 7800 11636 7806 11688
rect 9468 11679 9526 11685
rect 9468 11645 9480 11679
rect 9514 11676 9526 11679
rect 10336 11676 10364 11843
rect 10410 11840 10416 11852
rect 10468 11840 10474 11892
rect 11517 11883 11575 11889
rect 11517 11849 11529 11883
rect 11563 11880 11575 11883
rect 11790 11880 11796 11892
rect 11563 11852 11796 11880
rect 11563 11849 11575 11852
rect 11517 11843 11575 11849
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 17402 11880 17408 11892
rect 17363 11852 17408 11880
rect 17402 11840 17408 11852
rect 17460 11840 17466 11892
rect 17862 11880 17868 11892
rect 17823 11852 17868 11880
rect 17862 11840 17868 11852
rect 17920 11840 17926 11892
rect 21634 11880 21640 11892
rect 21595 11852 21640 11880
rect 21634 11840 21640 11852
rect 21692 11840 21698 11892
rect 10502 11772 10508 11824
rect 10560 11812 10566 11824
rect 17037 11815 17095 11821
rect 10560 11784 15459 11812
rect 10560 11772 10566 11784
rect 12575 11747 12633 11753
rect 12575 11713 12587 11747
rect 12621 11744 12633 11747
rect 13722 11744 13728 11756
rect 12621 11716 13728 11744
rect 12621 11713 12633 11716
rect 12575 11707 12633 11713
rect 13722 11704 13728 11716
rect 13780 11704 13786 11756
rect 9514 11648 10364 11676
rect 10597 11679 10655 11685
rect 9514 11645 9526 11648
rect 9468 11639 9526 11645
rect 10597 11645 10609 11679
rect 10643 11676 10655 11679
rect 11146 11676 11152 11688
rect 10643 11648 11152 11676
rect 10643 11645 10655 11648
rect 10597 11639 10655 11645
rect 11146 11636 11152 11648
rect 11204 11636 11210 11688
rect 12488 11679 12546 11685
rect 12488 11645 12500 11679
rect 12534 11676 12546 11679
rect 12710 11676 12716 11688
rect 12534 11648 12716 11676
rect 12534 11645 12546 11648
rect 12488 11639 12546 11645
rect 12710 11636 12716 11648
rect 12768 11676 12774 11688
rect 12897 11679 12955 11685
rect 12897 11676 12909 11679
rect 12768 11648 12909 11676
rect 12768 11636 12774 11648
rect 12897 11645 12909 11648
rect 12943 11645 12955 11679
rect 13446 11676 13452 11688
rect 13407 11648 13452 11676
rect 12897 11639 12955 11645
rect 13446 11636 13452 11648
rect 13504 11636 13510 11688
rect 15431 11685 15459 11784
rect 17037 11781 17049 11815
rect 17083 11812 17095 11815
rect 17310 11812 17316 11824
rect 17083 11784 17316 11812
rect 17083 11781 17095 11784
rect 17037 11775 17095 11781
rect 17310 11772 17316 11784
rect 17368 11812 17374 11824
rect 20162 11812 20168 11824
rect 17368 11784 20168 11812
rect 17368 11772 17374 11784
rect 20162 11772 20168 11784
rect 20220 11772 20226 11824
rect 21269 11815 21327 11821
rect 21269 11781 21281 11815
rect 21315 11812 21327 11815
rect 21358 11812 21364 11824
rect 21315 11784 21364 11812
rect 21315 11781 21327 11784
rect 21269 11775 21327 11781
rect 21358 11772 21364 11784
rect 21416 11772 21422 11824
rect 15519 11747 15577 11753
rect 15519 11713 15531 11747
rect 15565 11744 15577 11747
rect 16485 11747 16543 11753
rect 16485 11744 16497 11747
rect 15565 11716 16497 11744
rect 15565 11713 15577 11716
rect 15519 11707 15577 11713
rect 16485 11713 16497 11716
rect 16531 11744 16543 11747
rect 16758 11744 16764 11756
rect 16531 11716 16764 11744
rect 16531 11713 16543 11716
rect 16485 11707 16543 11713
rect 16758 11704 16764 11716
rect 16816 11704 16822 11756
rect 20257 11747 20315 11753
rect 20257 11713 20269 11747
rect 20303 11744 20315 11747
rect 20714 11744 20720 11756
rect 20303 11716 20720 11744
rect 20303 11713 20315 11716
rect 20257 11707 20315 11713
rect 20714 11704 20720 11716
rect 20772 11704 20778 11756
rect 15416 11679 15474 11685
rect 15416 11645 15428 11679
rect 15462 11676 15474 11679
rect 15841 11679 15899 11685
rect 15841 11676 15853 11679
rect 15462 11648 15853 11676
rect 15462 11645 15474 11648
rect 15416 11639 15474 11645
rect 15841 11645 15853 11648
rect 15887 11645 15899 11679
rect 15841 11639 15899 11645
rect 18116 11679 18174 11685
rect 18116 11645 18128 11679
rect 18162 11676 18174 11679
rect 21085 11679 21143 11685
rect 18162 11648 18644 11676
rect 18162 11645 18174 11648
rect 18116 11639 18174 11645
rect 3466 11611 3524 11617
rect 3466 11577 3478 11611
rect 3512 11577 3524 11611
rect 4982 11608 4988 11620
rect 4943 11580 4988 11608
rect 3466 11571 3524 11577
rect 2501 11543 2559 11549
rect 2501 11509 2513 11543
rect 2547 11540 2559 11543
rect 2590 11540 2596 11552
rect 2547 11512 2596 11540
rect 2547 11509 2559 11512
rect 2501 11503 2559 11509
rect 2590 11500 2596 11512
rect 2648 11500 2654 11552
rect 2682 11500 2688 11552
rect 2740 11540 2746 11552
rect 2961 11543 3019 11549
rect 2961 11540 2973 11543
rect 2740 11512 2973 11540
rect 2740 11500 2746 11512
rect 2961 11509 2973 11512
rect 3007 11540 3019 11543
rect 3481 11540 3509 11571
rect 4982 11568 4988 11580
rect 5040 11568 5046 11620
rect 5077 11611 5135 11617
rect 5077 11577 5089 11611
rect 5123 11577 5135 11611
rect 5994 11608 6000 11620
rect 5907 11580 6000 11608
rect 5077 11571 5135 11577
rect 3007 11512 3509 11540
rect 4801 11543 4859 11549
rect 3007 11509 3019 11512
rect 2961 11503 3019 11509
rect 4801 11509 4813 11543
rect 4847 11540 4859 11543
rect 4890 11540 4896 11552
rect 4847 11512 4896 11540
rect 4847 11509 4859 11512
rect 4801 11503 4859 11509
rect 4890 11500 4896 11512
rect 4948 11540 4954 11552
rect 5092 11540 5120 11571
rect 5994 11568 6000 11580
rect 6052 11608 6058 11620
rect 6454 11608 6460 11620
rect 6052 11580 6460 11608
rect 6052 11568 6058 11580
rect 6454 11568 6460 11580
rect 6512 11608 6518 11620
rect 7558 11608 7564 11620
rect 6512 11580 7564 11608
rect 6512 11568 6518 11580
rect 7558 11568 7564 11580
rect 7616 11568 7622 11620
rect 8015 11611 8073 11617
rect 8015 11608 8027 11611
rect 7668 11580 8027 11608
rect 7466 11540 7472 11552
rect 4948 11512 5120 11540
rect 7379 11512 7472 11540
rect 4948 11500 4954 11512
rect 7466 11500 7472 11512
rect 7524 11540 7530 11552
rect 7668 11540 7696 11580
rect 8015 11577 8027 11580
rect 8061 11608 8073 11611
rect 8570 11608 8576 11620
rect 8061 11580 8576 11608
rect 8061 11577 8073 11580
rect 8015 11571 8073 11577
rect 8570 11568 8576 11580
rect 8628 11608 8634 11620
rect 10686 11608 10692 11620
rect 8628 11580 10692 11608
rect 8628 11568 8634 11580
rect 10686 11568 10692 11580
rect 10744 11608 10750 11620
rect 10918 11611 10976 11617
rect 10918 11608 10930 11611
rect 10744 11580 10930 11608
rect 10744 11568 10750 11580
rect 10918 11577 10930 11580
rect 10964 11608 10976 11611
rect 13265 11611 13323 11617
rect 13265 11608 13277 11611
rect 10964 11580 13277 11608
rect 10964 11577 10976 11580
rect 10918 11571 10976 11577
rect 13265 11577 13277 11580
rect 13311 11608 13323 11611
rect 13770 11611 13828 11617
rect 13770 11608 13782 11611
rect 13311 11580 13782 11608
rect 13311 11577 13323 11580
rect 13265 11571 13323 11577
rect 13770 11577 13782 11580
rect 13816 11577 13828 11611
rect 13770 11571 13828 11577
rect 16301 11611 16359 11617
rect 16301 11577 16313 11611
rect 16347 11608 16359 11611
rect 16574 11608 16580 11620
rect 16347 11580 16580 11608
rect 16347 11577 16359 11580
rect 16301 11571 16359 11577
rect 16574 11568 16580 11580
rect 16632 11568 16638 11620
rect 7524 11512 7696 11540
rect 7524 11500 7530 11512
rect 8110 11500 8116 11552
rect 8168 11540 8174 11552
rect 9539 11543 9597 11549
rect 9539 11540 9551 11543
rect 8168 11512 9551 11540
rect 8168 11500 8174 11512
rect 9539 11509 9551 11512
rect 9585 11509 9597 11543
rect 9950 11540 9956 11552
rect 9911 11512 9956 11540
rect 9539 11503 9597 11509
rect 9950 11500 9956 11512
rect 10008 11500 10014 11552
rect 12158 11540 12164 11552
rect 12119 11512 12164 11540
rect 12158 11500 12164 11512
rect 12216 11500 12222 11552
rect 14366 11540 14372 11552
rect 14327 11512 14372 11540
rect 14366 11500 14372 11512
rect 14424 11500 14430 11552
rect 15194 11540 15200 11552
rect 15155 11512 15200 11540
rect 15194 11500 15200 11512
rect 15252 11500 15258 11552
rect 18046 11500 18052 11552
rect 18104 11540 18110 11552
rect 18616 11549 18644 11648
rect 21085 11645 21097 11679
rect 21131 11676 21143 11679
rect 21634 11676 21640 11688
rect 21131 11648 21640 11676
rect 21131 11645 21143 11648
rect 21085 11639 21143 11645
rect 21634 11636 21640 11648
rect 21692 11636 21698 11688
rect 19061 11611 19119 11617
rect 19061 11577 19073 11611
rect 19107 11608 19119 11611
rect 19610 11608 19616 11620
rect 19107 11580 19466 11608
rect 19571 11580 19616 11608
rect 19107 11577 19119 11580
rect 19061 11571 19119 11577
rect 18187 11543 18245 11549
rect 18187 11540 18199 11543
rect 18104 11512 18199 11540
rect 18104 11500 18110 11512
rect 18187 11509 18199 11512
rect 18233 11509 18245 11543
rect 18187 11503 18245 11509
rect 18601 11543 18659 11549
rect 18601 11509 18613 11543
rect 18647 11540 18659 11543
rect 18782 11540 18788 11552
rect 18647 11512 18788 11540
rect 18647 11509 18659 11512
rect 18601 11503 18659 11509
rect 18782 11500 18788 11512
rect 18840 11500 18846 11552
rect 19334 11540 19340 11552
rect 19295 11512 19340 11540
rect 19334 11500 19340 11512
rect 19392 11500 19398 11552
rect 19438 11540 19466 11580
rect 19610 11568 19616 11580
rect 19668 11568 19674 11620
rect 19705 11611 19763 11617
rect 19705 11577 19717 11611
rect 19751 11577 19763 11611
rect 19705 11571 19763 11577
rect 19518 11540 19524 11552
rect 19438 11512 19524 11540
rect 19518 11500 19524 11512
rect 19576 11540 19582 11552
rect 19720 11540 19748 11571
rect 19576 11512 19748 11540
rect 19576 11500 19582 11512
rect 1104 11450 22816 11472
rect 1104 11398 8982 11450
rect 9034 11398 9046 11450
rect 9098 11398 9110 11450
rect 9162 11398 9174 11450
rect 9226 11398 16982 11450
rect 17034 11398 17046 11450
rect 17098 11398 17110 11450
rect 17162 11398 17174 11450
rect 17226 11398 22816 11450
rect 1104 11376 22816 11398
rect 3142 11336 3148 11348
rect 3103 11308 3148 11336
rect 3142 11296 3148 11308
rect 3200 11296 3206 11348
rect 3878 11336 3884 11348
rect 3839 11308 3884 11336
rect 3878 11296 3884 11308
rect 3936 11296 3942 11348
rect 4890 11296 4896 11348
rect 4948 11336 4954 11348
rect 4985 11339 5043 11345
rect 4985 11336 4997 11339
rect 4948 11308 4997 11336
rect 4948 11296 4954 11308
rect 4985 11305 4997 11308
rect 5031 11305 5043 11339
rect 4985 11299 5043 11305
rect 5353 11339 5411 11345
rect 5353 11305 5365 11339
rect 5399 11336 5411 11339
rect 5442 11336 5448 11348
rect 5399 11308 5448 11336
rect 5399 11305 5411 11308
rect 5353 11299 5411 11305
rect 5442 11296 5448 11308
rect 5500 11336 5506 11348
rect 5902 11336 5908 11348
rect 5500 11308 5908 11336
rect 5500 11296 5506 11308
rect 5902 11296 5908 11308
rect 5960 11296 5966 11348
rect 8110 11336 8116 11348
rect 8071 11308 8116 11336
rect 8110 11296 8116 11308
rect 8168 11296 8174 11348
rect 13817 11339 13875 11345
rect 13817 11305 13829 11339
rect 13863 11336 13875 11339
rect 14366 11336 14372 11348
rect 13863 11308 14372 11336
rect 13863 11305 13875 11308
rect 13817 11299 13875 11305
rect 14366 11296 14372 11308
rect 14424 11296 14430 11348
rect 16574 11296 16580 11348
rect 16632 11336 16638 11348
rect 17037 11339 17095 11345
rect 17037 11336 17049 11339
rect 16632 11308 17049 11336
rect 16632 11296 16638 11308
rect 17037 11305 17049 11308
rect 17083 11336 17095 11339
rect 17770 11336 17776 11348
rect 17083 11308 17776 11336
rect 17083 11305 17095 11308
rect 17037 11299 17095 11305
rect 17770 11296 17776 11308
rect 17828 11296 17834 11348
rect 18046 11336 18052 11348
rect 18007 11308 18052 11336
rect 18046 11296 18052 11308
rect 18104 11296 18110 11348
rect 19058 11336 19064 11348
rect 19019 11308 19064 11336
rect 19058 11296 19064 11308
rect 19116 11296 19122 11348
rect 19610 11296 19616 11348
rect 19668 11336 19674 11348
rect 19889 11339 19947 11345
rect 19889 11336 19901 11339
rect 19668 11308 19901 11336
rect 19668 11296 19674 11308
rect 19889 11305 19901 11308
rect 19935 11336 19947 11339
rect 21039 11339 21097 11345
rect 21039 11336 21051 11339
rect 19935 11308 21051 11336
rect 19935 11305 19947 11308
rect 19889 11299 19947 11305
rect 21039 11305 21051 11308
rect 21085 11305 21097 11339
rect 21039 11299 21097 11305
rect 4427 11271 4485 11277
rect 4427 11237 4439 11271
rect 4473 11268 4485 11271
rect 4614 11268 4620 11280
rect 4473 11240 4620 11268
rect 4473 11237 4485 11240
rect 4427 11231 4485 11237
rect 4614 11228 4620 11240
rect 4672 11228 4678 11280
rect 6270 11268 6276 11280
rect 5895 11240 6276 11268
rect 1464 11203 1522 11209
rect 1464 11169 1476 11203
rect 1510 11200 1522 11203
rect 1670 11200 1676 11212
rect 1510 11172 1676 11200
rect 1510 11169 1522 11172
rect 1464 11163 1522 11169
rect 1670 11160 1676 11172
rect 1728 11160 1734 11212
rect 5895 11209 5923 11240
rect 6270 11228 6276 11240
rect 6328 11268 6334 11280
rect 7190 11268 7196 11280
rect 6328 11240 7196 11268
rect 6328 11228 6334 11240
rect 7190 11228 7196 11240
rect 7248 11228 7254 11280
rect 7742 11268 7748 11280
rect 7703 11240 7748 11268
rect 7742 11228 7748 11240
rect 7800 11228 7806 11280
rect 11146 11268 11152 11280
rect 11107 11240 11152 11268
rect 11146 11228 11152 11240
rect 11204 11228 11210 11280
rect 12621 11271 12679 11277
rect 12621 11237 12633 11271
rect 12667 11268 12679 11271
rect 13446 11268 13452 11280
rect 12667 11240 13216 11268
rect 13407 11240 13452 11268
rect 12667 11237 12679 11240
rect 12621 11231 12679 11237
rect 5880 11203 5938 11209
rect 5880 11169 5892 11203
rect 5926 11169 5938 11203
rect 5880 11163 5938 11169
rect 7101 11203 7159 11209
rect 7101 11169 7113 11203
rect 7147 11169 7159 11203
rect 7558 11200 7564 11212
rect 7519 11172 7564 11200
rect 7101 11163 7159 11169
rect 2406 11132 2412 11144
rect 2367 11104 2412 11132
rect 2406 11092 2412 11104
rect 2464 11092 2470 11144
rect 4065 11135 4123 11141
rect 4065 11101 4077 11135
rect 4111 11132 4123 11135
rect 4246 11132 4252 11144
rect 4111 11104 4252 11132
rect 4111 11101 4123 11104
rect 4065 11095 4123 11101
rect 4246 11092 4252 11104
rect 4304 11092 4310 11144
rect 7116 11076 7144 11163
rect 7558 11160 7564 11172
rect 7616 11160 7622 11212
rect 8640 11203 8698 11209
rect 8640 11169 8652 11203
rect 8686 11200 8698 11203
rect 9306 11200 9312 11212
rect 8686 11172 9312 11200
rect 8686 11169 8698 11172
rect 8640 11163 8698 11169
rect 9306 11160 9312 11172
rect 9364 11160 9370 11212
rect 10686 11200 10692 11212
rect 10647 11172 10692 11200
rect 10686 11160 10692 11172
rect 10744 11160 10750 11212
rect 10965 11203 11023 11209
rect 10965 11169 10977 11203
rect 11011 11200 11023 11203
rect 11238 11200 11244 11212
rect 11011 11172 11244 11200
rect 11011 11169 11023 11172
rect 10965 11163 11023 11169
rect 7742 11132 7748 11144
rect 7392 11104 7748 11132
rect 106 11024 112 11076
rect 164 11064 170 11076
rect 3786 11064 3792 11076
rect 164 11036 3792 11064
rect 164 11024 170 11036
rect 3786 11024 3792 11036
rect 3844 11024 3850 11076
rect 7098 11064 7104 11076
rect 7011 11036 7104 11064
rect 7098 11024 7104 11036
rect 7156 11064 7162 11076
rect 7392 11064 7420 11104
rect 7742 11092 7748 11104
rect 7800 11132 7806 11144
rect 10980 11132 11008 11163
rect 11238 11160 11244 11172
rect 11296 11160 11302 11212
rect 13188 11209 13216 11240
rect 13446 11228 13452 11240
rect 13504 11228 13510 11280
rect 13722 11228 13728 11280
rect 13780 11268 13786 11280
rect 14093 11271 14151 11277
rect 14093 11268 14105 11271
rect 13780 11240 14105 11268
rect 13780 11228 13786 11240
rect 14093 11237 14105 11240
rect 14139 11237 14151 11271
rect 14093 11231 14151 11237
rect 16298 11228 16304 11280
rect 16356 11268 16362 11280
rect 16438 11271 16496 11277
rect 16438 11268 16450 11271
rect 16356 11240 16450 11268
rect 16356 11228 16362 11240
rect 16438 11237 16450 11240
rect 16484 11237 16496 11271
rect 16438 11231 16496 11237
rect 12989 11203 13047 11209
rect 12989 11169 13001 11203
rect 13035 11169 13047 11203
rect 12989 11163 13047 11169
rect 13173 11203 13231 11209
rect 13173 11169 13185 11203
rect 13219 11200 13231 11203
rect 13906 11200 13912 11212
rect 13219 11172 13912 11200
rect 13219 11169 13231 11172
rect 13173 11163 13231 11169
rect 7800 11104 11008 11132
rect 7800 11092 7806 11104
rect 12802 11092 12808 11144
rect 12860 11132 12866 11144
rect 13004 11132 13032 11163
rect 13906 11160 13912 11172
rect 13964 11160 13970 11212
rect 19518 11160 19524 11212
rect 19576 11200 19582 11212
rect 19613 11203 19671 11209
rect 19613 11200 19625 11203
rect 19576 11172 19625 11200
rect 19576 11160 19582 11172
rect 19613 11169 19625 11172
rect 19659 11169 19671 11203
rect 19613 11163 19671 11169
rect 20806 11160 20812 11212
rect 20864 11200 20870 11212
rect 20936 11203 20994 11209
rect 20936 11200 20948 11203
rect 20864 11172 20948 11200
rect 20864 11160 20870 11172
rect 20936 11169 20948 11172
rect 20982 11169 20994 11203
rect 20936 11163 20994 11169
rect 13998 11132 14004 11144
rect 12860 11104 14004 11132
rect 12860 11092 12866 11104
rect 13998 11092 14004 11104
rect 14056 11132 14062 11144
rect 14366 11132 14372 11144
rect 14056 11104 14372 11132
rect 14056 11092 14062 11104
rect 14366 11092 14372 11104
rect 14424 11092 14430 11144
rect 16114 11132 16120 11144
rect 16075 11104 16120 11132
rect 16114 11092 16120 11104
rect 16172 11092 16178 11144
rect 18690 11132 18696 11144
rect 18651 11104 18696 11132
rect 18690 11092 18696 11104
rect 18748 11092 18754 11144
rect 7156 11036 7420 11064
rect 7156 11024 7162 11036
rect 9674 11024 9680 11076
rect 9732 11064 9738 11076
rect 10229 11067 10287 11073
rect 10229 11064 10241 11067
rect 9732 11036 10241 11064
rect 9732 11024 9738 11036
rect 10229 11033 10241 11036
rect 10275 11033 10287 11067
rect 10229 11027 10287 11033
rect 10318 11024 10324 11076
rect 10376 11064 10382 11076
rect 14182 11064 14188 11076
rect 10376 11036 14188 11064
rect 10376 11024 10382 11036
rect 14182 11024 14188 11036
rect 14240 11024 14246 11076
rect 17310 11024 17316 11076
rect 17368 11064 17374 11076
rect 18230 11064 18236 11076
rect 17368 11036 18236 11064
rect 17368 11024 17374 11036
rect 18230 11024 18236 11036
rect 18288 11024 18294 11076
rect 750 10956 756 11008
rect 808 10996 814 11008
rect 1535 10999 1593 11005
rect 1535 10996 1547 10999
rect 808 10968 1547 10996
rect 808 10956 814 10968
rect 1535 10965 1547 10968
rect 1581 10965 1593 10999
rect 1946 10996 1952 11008
rect 1907 10968 1952 10996
rect 1535 10959 1593 10965
rect 1946 10956 1952 10968
rect 2004 10956 2010 11008
rect 5951 10999 6009 11005
rect 5951 10965 5963 10999
rect 5997 10996 6009 10999
rect 6730 10996 6736 11008
rect 5997 10968 6736 10996
rect 5997 10965 6009 10968
rect 5951 10959 6009 10965
rect 6730 10956 6736 10968
rect 6788 10956 6794 11008
rect 6914 10996 6920 11008
rect 6875 10968 6920 10996
rect 6914 10956 6920 10968
rect 6972 10956 6978 11008
rect 8711 10999 8769 11005
rect 8711 10965 8723 10999
rect 8757 10996 8769 10999
rect 9582 10996 9588 11008
rect 8757 10968 9588 10996
rect 8757 10965 8769 10968
rect 8711 10959 8769 10965
rect 9582 10956 9588 10968
rect 9640 10956 9646 11008
rect 9858 10996 9864 11008
rect 9819 10968 9864 10996
rect 9858 10956 9864 10968
rect 9916 10956 9922 11008
rect 1104 10906 22816 10928
rect 1104 10854 4982 10906
rect 5034 10854 5046 10906
rect 5098 10854 5110 10906
rect 5162 10854 5174 10906
rect 5226 10854 12982 10906
rect 13034 10854 13046 10906
rect 13098 10854 13110 10906
rect 13162 10854 13174 10906
rect 13226 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 22816 10906
rect 1104 10832 22816 10854
rect 6270 10792 6276 10804
rect 6231 10764 6276 10792
rect 6270 10752 6276 10764
rect 6328 10752 6334 10804
rect 6641 10795 6699 10801
rect 6641 10761 6653 10795
rect 6687 10792 6699 10795
rect 7098 10792 7104 10804
rect 6687 10764 7104 10792
rect 6687 10761 6699 10764
rect 6641 10755 6699 10761
rect 7098 10752 7104 10764
rect 7156 10752 7162 10804
rect 8938 10792 8944 10804
rect 8899 10764 8944 10792
rect 8938 10752 8944 10764
rect 8996 10752 9002 10804
rect 9306 10792 9312 10804
rect 9219 10764 9312 10792
rect 9306 10752 9312 10764
rect 9364 10792 9370 10804
rect 10318 10792 10324 10804
rect 9364 10764 10324 10792
rect 9364 10752 9370 10764
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 11057 10795 11115 10801
rect 11057 10761 11069 10795
rect 11103 10792 11115 10795
rect 11238 10792 11244 10804
rect 11103 10764 11244 10792
rect 11103 10761 11115 10764
rect 11057 10755 11115 10761
rect 11238 10752 11244 10764
rect 11296 10752 11302 10804
rect 11379 10795 11437 10801
rect 11379 10761 11391 10795
rect 11425 10792 11437 10795
rect 12158 10792 12164 10804
rect 11425 10764 12164 10792
rect 11425 10761 11437 10764
rect 11379 10755 11437 10761
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 14366 10792 14372 10804
rect 14327 10764 14372 10792
rect 14366 10752 14372 10764
rect 14424 10752 14430 10804
rect 16298 10752 16304 10804
rect 16356 10792 16362 10804
rect 16577 10795 16635 10801
rect 16577 10792 16589 10795
rect 16356 10764 16589 10792
rect 16356 10752 16362 10764
rect 16577 10761 16589 10764
rect 16623 10761 16635 10795
rect 17770 10792 17776 10804
rect 17731 10764 17776 10792
rect 16577 10755 16635 10761
rect 17770 10752 17776 10764
rect 17828 10752 17834 10804
rect 19058 10792 19064 10804
rect 19019 10764 19064 10792
rect 19058 10752 19064 10764
rect 19116 10752 19122 10804
rect 19518 10792 19524 10804
rect 19479 10764 19524 10792
rect 19518 10752 19524 10764
rect 19576 10752 19582 10804
rect 1670 10684 1676 10736
rect 1728 10724 1734 10736
rect 2501 10727 2559 10733
rect 2501 10724 2513 10727
rect 1728 10696 2513 10724
rect 1728 10684 1734 10696
rect 2501 10693 2513 10696
rect 2547 10724 2559 10727
rect 4706 10724 4712 10736
rect 2547 10696 4712 10724
rect 2547 10693 2559 10696
rect 2501 10687 2559 10693
rect 4706 10684 4712 10696
rect 4764 10684 4770 10736
rect 7558 10684 7564 10736
rect 7616 10724 7622 10736
rect 7929 10727 7987 10733
rect 7929 10724 7941 10727
rect 7616 10696 7941 10724
rect 7616 10684 7622 10696
rect 7929 10693 7941 10696
rect 7975 10724 7987 10727
rect 10226 10724 10232 10736
rect 7975 10696 10232 10724
rect 7975 10693 7987 10696
rect 7929 10687 7987 10693
rect 10226 10684 10232 10696
rect 10284 10684 10290 10736
rect 10686 10724 10692 10736
rect 10599 10696 10692 10724
rect 10686 10684 10692 10696
rect 10744 10724 10750 10736
rect 12802 10724 12808 10736
rect 10744 10696 12808 10724
rect 10744 10684 10750 10696
rect 12802 10684 12808 10696
rect 12860 10684 12866 10736
rect 13081 10727 13139 10733
rect 13081 10693 13093 10727
rect 13127 10724 13139 10727
rect 13354 10724 13360 10736
rect 13127 10696 13360 10724
rect 13127 10693 13139 10696
rect 13081 10687 13139 10693
rect 13354 10684 13360 10696
rect 13412 10724 13418 10736
rect 14001 10727 14059 10733
rect 14001 10724 14013 10727
rect 13412 10696 14013 10724
rect 13412 10684 13418 10696
rect 14001 10693 14013 10696
rect 14047 10693 14059 10727
rect 14001 10687 14059 10693
rect 18046 10684 18052 10736
rect 18104 10724 18110 10736
rect 18104 10696 18184 10724
rect 18104 10684 18110 10696
rect 1765 10659 1823 10665
rect 1765 10625 1777 10659
rect 1811 10656 1823 10659
rect 1949 10659 2007 10665
rect 1949 10656 1961 10659
rect 1811 10628 1961 10656
rect 1811 10625 1823 10628
rect 1765 10619 1823 10625
rect 1949 10625 1961 10628
rect 1995 10656 2007 10659
rect 2406 10656 2412 10668
rect 1995 10628 2412 10656
rect 1995 10625 2007 10628
rect 1949 10619 2007 10625
rect 2406 10616 2412 10628
rect 2464 10616 2470 10668
rect 2590 10616 2596 10668
rect 2648 10656 2654 10668
rect 3513 10659 3571 10665
rect 3513 10656 3525 10659
rect 2648 10628 3525 10656
rect 2648 10616 2654 10628
rect 3513 10625 3525 10628
rect 3559 10656 3571 10659
rect 4246 10656 4252 10668
rect 3559 10628 4154 10656
rect 4207 10628 4252 10656
rect 3559 10625 3571 10628
rect 3513 10619 3571 10625
rect 4126 10600 4154 10628
rect 4246 10616 4252 10628
rect 4304 10616 4310 10668
rect 5994 10656 6000 10668
rect 4862 10628 6000 10656
rect 3694 10588 3700 10600
rect 3655 10560 3700 10588
rect 3694 10548 3700 10560
rect 3752 10548 3758 10600
rect 4126 10560 4160 10600
rect 4154 10548 4160 10560
rect 4212 10588 4218 10600
rect 4862 10588 4890 10628
rect 5994 10616 6000 10628
rect 6052 10616 6058 10668
rect 6730 10616 6736 10668
rect 6788 10656 6794 10668
rect 6917 10659 6975 10665
rect 6917 10656 6929 10659
rect 6788 10628 6929 10656
rect 6788 10616 6794 10628
rect 6917 10625 6929 10628
rect 6963 10656 6975 10659
rect 8205 10659 8263 10665
rect 8205 10656 8217 10659
rect 6963 10628 8217 10656
rect 6963 10625 6975 10628
rect 6917 10619 6975 10625
rect 8205 10625 8217 10628
rect 8251 10625 8263 10659
rect 8205 10619 8263 10625
rect 8846 10616 8852 10668
rect 8904 10656 8910 10668
rect 8904 10628 13814 10656
rect 8904 10616 8910 10628
rect 5442 10588 5448 10600
rect 4212 10560 4890 10588
rect 5403 10560 5448 10588
rect 4212 10548 4218 10560
rect 5442 10548 5448 10560
rect 5500 10548 5506 10600
rect 5718 10588 5724 10600
rect 5679 10560 5724 10588
rect 5718 10548 5724 10560
rect 5776 10548 5782 10600
rect 8478 10597 8484 10600
rect 8456 10591 8484 10597
rect 8456 10588 8468 10591
rect 8391 10560 8468 10588
rect 8456 10557 8468 10560
rect 8536 10588 8542 10600
rect 8938 10588 8944 10600
rect 8536 10560 8944 10588
rect 8456 10551 8484 10557
rect 8478 10548 8484 10551
rect 8536 10548 8542 10560
rect 8938 10548 8944 10560
rect 8996 10548 9002 10600
rect 11308 10591 11366 10597
rect 11308 10557 11320 10591
rect 11354 10588 11366 10591
rect 12897 10591 12955 10597
rect 11354 10560 11468 10588
rect 11354 10557 11366 10560
rect 11308 10551 11366 10557
rect 1946 10480 1952 10532
rect 2004 10520 2010 10532
rect 2041 10523 2099 10529
rect 2041 10520 2053 10523
rect 2004 10492 2053 10520
rect 2004 10480 2010 10492
rect 2041 10489 2053 10492
rect 2087 10489 2099 10523
rect 2041 10483 2099 10489
rect 4985 10523 5043 10529
rect 4985 10489 4997 10523
rect 5031 10520 5043 10523
rect 5736 10520 5764 10548
rect 5031 10492 5764 10520
rect 5031 10489 5043 10492
rect 4985 10483 5043 10489
rect 6914 10480 6920 10532
rect 6972 10520 6978 10532
rect 7009 10523 7067 10529
rect 7009 10520 7021 10523
rect 6972 10492 7021 10520
rect 6972 10480 6978 10492
rect 7009 10489 7021 10492
rect 7055 10489 7067 10523
rect 7009 10483 7067 10489
rect 7282 10480 7288 10532
rect 7340 10520 7346 10532
rect 7561 10523 7619 10529
rect 7561 10520 7573 10523
rect 7340 10492 7573 10520
rect 7340 10480 7346 10492
rect 7561 10489 7573 10492
rect 7607 10520 7619 10523
rect 9674 10520 9680 10532
rect 7607 10492 9352 10520
rect 9635 10492 9680 10520
rect 7607 10489 7619 10492
rect 7561 10483 7619 10489
rect 3694 10412 3700 10464
rect 3752 10452 3758 10464
rect 4338 10452 4344 10464
rect 3752 10424 4344 10452
rect 3752 10412 3758 10424
rect 4338 10412 4344 10424
rect 4396 10452 4402 10464
rect 4522 10452 4528 10464
rect 4396 10424 4528 10452
rect 4396 10412 4402 10424
rect 4522 10412 4528 10424
rect 4580 10412 4586 10464
rect 4706 10452 4712 10464
rect 4667 10424 4712 10452
rect 4706 10412 4712 10424
rect 4764 10412 4770 10464
rect 5074 10412 5080 10464
rect 5132 10452 5138 10464
rect 5261 10455 5319 10461
rect 5261 10452 5273 10455
rect 5132 10424 5273 10452
rect 5132 10412 5138 10424
rect 5261 10421 5273 10424
rect 5307 10421 5319 10455
rect 5261 10415 5319 10421
rect 7926 10412 7932 10464
rect 7984 10452 7990 10464
rect 8527 10455 8585 10461
rect 8527 10452 8539 10455
rect 7984 10424 8539 10452
rect 7984 10412 7990 10424
rect 8527 10421 8539 10424
rect 8573 10421 8585 10455
rect 9324 10452 9352 10492
rect 9674 10480 9680 10492
rect 9732 10480 9738 10532
rect 9769 10523 9827 10529
rect 9769 10489 9781 10523
rect 9815 10520 9827 10523
rect 9858 10520 9864 10532
rect 9815 10492 9864 10520
rect 9815 10489 9827 10492
rect 9769 10483 9827 10489
rect 9858 10480 9864 10492
rect 9916 10480 9922 10532
rect 10318 10520 10324 10532
rect 10279 10492 10324 10520
rect 10318 10480 10324 10492
rect 10376 10480 10382 10532
rect 10336 10452 10364 10480
rect 11440 10464 11468 10560
rect 12897 10557 12909 10591
rect 12943 10588 12955 10591
rect 12986 10588 12992 10600
rect 12943 10560 12992 10588
rect 12943 10557 12955 10560
rect 12897 10551 12955 10557
rect 12986 10548 12992 10560
rect 13044 10548 13050 10600
rect 13262 10588 13268 10600
rect 13223 10560 13268 10588
rect 13262 10548 13268 10560
rect 13320 10548 13326 10600
rect 13786 10588 13814 10628
rect 16114 10616 16120 10668
rect 16172 10656 16178 10668
rect 18156 10665 18184 10696
rect 16301 10659 16359 10665
rect 16301 10656 16313 10659
rect 16172 10628 16313 10656
rect 16172 10616 16178 10628
rect 16301 10625 16313 10628
rect 16347 10656 16359 10659
rect 16945 10659 17003 10665
rect 16945 10656 16957 10659
rect 16347 10628 16957 10656
rect 16347 10625 16359 10628
rect 16301 10619 16359 10625
rect 16945 10625 16957 10628
rect 16991 10625 17003 10659
rect 16945 10619 17003 10625
rect 18141 10659 18199 10665
rect 18141 10625 18153 10659
rect 18187 10625 18199 10659
rect 18598 10656 18604 10668
rect 18559 10628 18604 10656
rect 18141 10619 18199 10625
rect 18598 10616 18604 10628
rect 18656 10616 18662 10668
rect 19702 10656 19708 10668
rect 19663 10628 19708 10656
rect 19702 10616 19708 10628
rect 19760 10616 19766 10668
rect 20162 10656 20168 10668
rect 20123 10628 20168 10656
rect 20162 10616 20168 10628
rect 20220 10616 20226 10668
rect 14588 10591 14646 10597
rect 14588 10588 14600 10591
rect 13786 10560 14600 10588
rect 14588 10557 14600 10560
rect 14634 10588 14646 10591
rect 15013 10591 15071 10597
rect 15013 10588 15025 10591
rect 14634 10560 15025 10588
rect 14634 10557 14646 10560
rect 14588 10551 14646 10557
rect 15013 10557 15025 10560
rect 15059 10557 15071 10591
rect 15562 10588 15568 10600
rect 15523 10560 15568 10588
rect 15013 10551 15071 10557
rect 15562 10548 15568 10560
rect 15620 10548 15626 10600
rect 16025 10591 16083 10597
rect 16025 10557 16037 10591
rect 16071 10588 16083 10591
rect 16390 10588 16396 10600
rect 16071 10560 16396 10588
rect 16071 10557 16083 10560
rect 16025 10551 16083 10557
rect 12253 10523 12311 10529
rect 12253 10489 12265 10523
rect 12299 10520 12311 10523
rect 12342 10520 12348 10532
rect 12299 10492 12348 10520
rect 12299 10489 12311 10492
rect 12253 10483 12311 10489
rect 12342 10480 12348 10492
rect 12400 10520 12406 10532
rect 13280 10520 13308 10548
rect 16040 10520 16068 10551
rect 16390 10548 16396 10560
rect 16448 10548 16454 10600
rect 12400 10492 13308 10520
rect 15396 10492 16068 10520
rect 12400 10480 12406 10492
rect 15396 10464 15424 10492
rect 17770 10480 17776 10532
rect 17828 10520 17834 10532
rect 18233 10523 18291 10529
rect 18233 10520 18245 10523
rect 17828 10492 18245 10520
rect 17828 10480 17834 10492
rect 18233 10489 18245 10492
rect 18279 10489 18291 10523
rect 18233 10483 18291 10489
rect 19518 10480 19524 10532
rect 19576 10520 19582 10532
rect 19797 10523 19855 10529
rect 19797 10520 19809 10523
rect 19576 10492 19809 10520
rect 19576 10480 19582 10492
rect 19797 10489 19809 10492
rect 19843 10489 19855 10523
rect 19797 10483 19855 10489
rect 9324 10424 10364 10452
rect 8527 10415 8585 10421
rect 11422 10412 11428 10464
rect 11480 10452 11486 10464
rect 11701 10455 11759 10461
rect 11701 10452 11713 10455
rect 11480 10424 11713 10452
rect 11480 10412 11486 10424
rect 11701 10421 11713 10424
rect 11747 10421 11759 10455
rect 11701 10415 11759 10421
rect 11790 10412 11796 10464
rect 11848 10452 11854 10464
rect 13449 10455 13507 10461
rect 13449 10452 13461 10455
rect 11848 10424 13461 10452
rect 11848 10412 11854 10424
rect 13449 10421 13461 10424
rect 13495 10421 13507 10455
rect 13449 10415 13507 10421
rect 14691 10455 14749 10461
rect 14691 10421 14703 10455
rect 14737 10452 14749 10455
rect 15286 10452 15292 10464
rect 14737 10424 15292 10452
rect 14737 10421 14749 10424
rect 14691 10415 14749 10421
rect 15286 10412 15292 10424
rect 15344 10412 15350 10464
rect 15378 10412 15384 10464
rect 15436 10452 15442 10464
rect 15436 10424 15481 10452
rect 15436 10412 15442 10424
rect 20438 10412 20444 10464
rect 20496 10452 20502 10464
rect 20806 10452 20812 10464
rect 20496 10424 20812 10452
rect 20496 10412 20502 10424
rect 20806 10412 20812 10424
rect 20864 10452 20870 10464
rect 20901 10455 20959 10461
rect 20901 10452 20913 10455
rect 20864 10424 20913 10452
rect 20864 10412 20870 10424
rect 20901 10421 20913 10424
rect 20947 10421 20959 10455
rect 20901 10415 20959 10421
rect 1104 10362 22816 10384
rect 1104 10310 8982 10362
rect 9034 10310 9046 10362
rect 9098 10310 9110 10362
rect 9162 10310 9174 10362
rect 9226 10310 16982 10362
rect 17034 10310 17046 10362
rect 17098 10310 17110 10362
rect 17162 10310 17174 10362
rect 17226 10310 22816 10362
rect 1104 10288 22816 10310
rect 1670 10248 1676 10260
rect 1631 10220 1676 10248
rect 1670 10208 1676 10220
rect 1728 10208 1734 10260
rect 1946 10208 1952 10260
rect 2004 10248 2010 10260
rect 2777 10251 2835 10257
rect 2777 10248 2789 10251
rect 2004 10220 2789 10248
rect 2004 10208 2010 10220
rect 2777 10217 2789 10220
rect 2823 10217 2835 10251
rect 3694 10248 3700 10260
rect 3655 10220 3700 10248
rect 2777 10211 2835 10217
rect 3694 10208 3700 10220
rect 3752 10208 3758 10260
rect 4246 10248 4252 10260
rect 4207 10220 4252 10248
rect 4246 10208 4252 10220
rect 4304 10208 4310 10260
rect 5905 10251 5963 10257
rect 5905 10217 5917 10251
rect 5951 10217 5963 10251
rect 5905 10211 5963 10217
rect 2219 10183 2277 10189
rect 2219 10149 2231 10183
rect 2265 10180 2277 10183
rect 2590 10180 2596 10192
rect 2265 10152 2596 10180
rect 2265 10149 2277 10152
rect 2219 10143 2277 10149
rect 2590 10140 2596 10152
rect 2648 10140 2654 10192
rect 4706 10140 4712 10192
rect 4764 10180 4770 10192
rect 5347 10183 5405 10189
rect 5347 10180 5359 10183
rect 4764 10152 5359 10180
rect 4764 10140 4770 10152
rect 5347 10149 5359 10152
rect 5393 10180 5405 10183
rect 5626 10180 5632 10192
rect 5393 10152 5632 10180
rect 5393 10149 5405 10152
rect 5347 10143 5405 10149
rect 5626 10140 5632 10152
rect 5684 10140 5690 10192
rect 5920 10180 5948 10211
rect 12250 10208 12256 10260
rect 12308 10248 12314 10260
rect 12437 10251 12495 10257
rect 12437 10248 12449 10251
rect 12308 10220 12449 10248
rect 12308 10208 12314 10220
rect 12437 10217 12449 10220
rect 12483 10217 12495 10251
rect 12437 10211 12495 10217
rect 13262 10208 13268 10260
rect 13320 10248 13326 10260
rect 13541 10251 13599 10257
rect 13541 10248 13553 10251
rect 13320 10220 13553 10248
rect 13320 10208 13326 10220
rect 13541 10217 13553 10220
rect 13587 10248 13599 10251
rect 14090 10248 14096 10260
rect 13587 10220 13952 10248
rect 14051 10220 14096 10248
rect 13587 10217 13599 10220
rect 13541 10211 13599 10217
rect 6270 10180 6276 10192
rect 5920 10152 6276 10180
rect 6270 10140 6276 10152
rect 6328 10180 6334 10192
rect 6914 10180 6920 10192
rect 6328 10152 6920 10180
rect 6328 10140 6334 10152
rect 6914 10140 6920 10152
rect 6972 10140 6978 10192
rect 9858 10180 9864 10192
rect 9819 10152 9864 10180
rect 9858 10140 9864 10152
rect 9916 10140 9922 10192
rect 11238 10140 11244 10192
rect 11296 10180 11302 10192
rect 13446 10180 13452 10192
rect 11296 10152 13452 10180
rect 11296 10140 11302 10152
rect 13446 10140 13452 10152
rect 13504 10140 13510 10192
rect 4798 10072 4804 10124
rect 4856 10112 4862 10124
rect 4985 10115 5043 10121
rect 4985 10112 4997 10115
rect 4856 10084 4997 10112
rect 4856 10072 4862 10084
rect 4985 10081 4997 10084
rect 5031 10112 5043 10115
rect 5074 10112 5080 10124
rect 5031 10084 5080 10112
rect 5031 10081 5043 10084
rect 4985 10075 5043 10081
rect 5074 10072 5080 10084
rect 5132 10072 5138 10124
rect 8624 10115 8682 10121
rect 8624 10081 8636 10115
rect 8670 10112 8682 10115
rect 8846 10112 8852 10124
rect 8670 10084 8852 10112
rect 8670 10081 8682 10084
rect 8624 10075 8682 10081
rect 8846 10072 8852 10084
rect 8904 10072 8910 10124
rect 11974 10112 11980 10124
rect 11935 10084 11980 10112
rect 11974 10072 11980 10084
rect 12032 10072 12038 10124
rect 12253 10115 12311 10121
rect 12253 10081 12265 10115
rect 12299 10112 12311 10115
rect 12342 10112 12348 10124
rect 12299 10084 12348 10112
rect 12299 10081 12311 10084
rect 12253 10075 12311 10081
rect 1854 10044 1860 10056
rect 1815 10016 1860 10044
rect 1854 10004 1860 10016
rect 1912 10004 1918 10056
rect 4062 10004 4068 10056
rect 4120 10044 4126 10056
rect 5442 10044 5448 10056
rect 4120 10016 5448 10044
rect 4120 10004 4126 10016
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 6638 10004 6644 10056
rect 6696 10044 6702 10056
rect 6825 10047 6883 10053
rect 6825 10044 6837 10047
rect 6696 10016 6837 10044
rect 6696 10004 6702 10016
rect 6825 10013 6837 10016
rect 6871 10044 6883 10047
rect 7926 10044 7932 10056
rect 6871 10016 7932 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 7926 10004 7932 10016
rect 7984 10004 7990 10056
rect 8711 10047 8769 10053
rect 8711 10013 8723 10047
rect 8757 10044 8769 10047
rect 9769 10047 9827 10053
rect 9769 10044 9781 10047
rect 8757 10016 9781 10044
rect 8757 10013 8769 10016
rect 8711 10007 8769 10013
rect 9769 10013 9781 10016
rect 9815 10044 9827 10047
rect 10042 10044 10048 10056
rect 9815 10016 10048 10044
rect 9815 10013 9827 10016
rect 9769 10007 9827 10013
rect 10042 10004 10048 10016
rect 10100 10004 10106 10056
rect 10410 10044 10416 10056
rect 10371 10016 10416 10044
rect 10410 10004 10416 10016
rect 10468 10004 10474 10056
rect 11885 10047 11943 10053
rect 11885 10013 11897 10047
rect 11931 10044 11943 10047
rect 12268 10044 12296 10075
rect 12342 10072 12348 10084
rect 12400 10072 12406 10124
rect 12986 10072 12992 10124
rect 13044 10112 13050 10124
rect 13924 10121 13952 10220
rect 14090 10208 14096 10220
rect 14148 10208 14154 10260
rect 15286 10208 15292 10260
rect 15344 10248 15350 10260
rect 15933 10251 15991 10257
rect 15933 10248 15945 10251
rect 15344 10220 15945 10248
rect 15344 10208 15350 10220
rect 15933 10217 15945 10220
rect 15979 10248 15991 10251
rect 16114 10248 16120 10260
rect 15979 10220 16120 10248
rect 15979 10217 15991 10220
rect 15933 10211 15991 10217
rect 16114 10208 16120 10220
rect 16172 10208 16178 10260
rect 19702 10248 19708 10260
rect 19663 10220 19708 10248
rect 19702 10208 19708 10220
rect 19760 10208 19766 10260
rect 15470 10140 15476 10192
rect 15528 10180 15534 10192
rect 16758 10180 16764 10192
rect 15528 10152 16764 10180
rect 15528 10140 15534 10152
rect 16408 10121 16436 10152
rect 16758 10140 16764 10152
rect 16816 10140 16822 10192
rect 18417 10183 18475 10189
rect 18417 10149 18429 10183
rect 18463 10180 18475 10183
rect 18690 10180 18696 10192
rect 18463 10152 18696 10180
rect 18463 10149 18475 10152
rect 18417 10143 18475 10149
rect 18690 10140 18696 10152
rect 18748 10140 18754 10192
rect 13633 10115 13691 10121
rect 13633 10112 13645 10115
rect 13044 10084 13645 10112
rect 13044 10072 13050 10084
rect 13633 10081 13645 10084
rect 13679 10112 13691 10115
rect 13909 10115 13967 10121
rect 13679 10084 13814 10112
rect 13679 10081 13691 10084
rect 13633 10075 13691 10081
rect 11931 10016 12296 10044
rect 13786 10044 13814 10084
rect 13909 10081 13921 10115
rect 13955 10081 13967 10115
rect 13909 10075 13967 10081
rect 16393 10115 16451 10121
rect 16393 10081 16405 10115
rect 16439 10081 16451 10115
rect 16393 10075 16451 10081
rect 16577 10115 16635 10121
rect 16577 10081 16589 10115
rect 16623 10081 16635 10115
rect 16577 10075 16635 10081
rect 17957 10115 18015 10121
rect 17957 10081 17969 10115
rect 18003 10081 18015 10115
rect 18138 10112 18144 10124
rect 18099 10084 18144 10112
rect 17957 10075 18015 10081
rect 13998 10044 14004 10056
rect 13786 10016 14004 10044
rect 11931 10013 11943 10016
rect 11885 10007 11943 10013
rect 13998 10004 14004 10016
rect 14056 10044 14062 10056
rect 14645 10047 14703 10053
rect 14645 10044 14657 10047
rect 14056 10016 14657 10044
rect 14056 10004 14062 10016
rect 14645 10013 14657 10016
rect 14691 10013 14703 10047
rect 14645 10007 14703 10013
rect 15654 10004 15660 10056
rect 15712 10044 15718 10056
rect 16592 10044 16620 10075
rect 16850 10044 16856 10056
rect 15712 10016 16620 10044
rect 16811 10016 16856 10044
rect 15712 10004 15718 10016
rect 16850 10004 16856 10016
rect 16908 10004 16914 10056
rect 17972 10044 18000 10075
rect 18138 10072 18144 10084
rect 18196 10072 18202 10124
rect 19312 10115 19370 10121
rect 19312 10081 19324 10115
rect 19358 10112 19370 10115
rect 19794 10112 19800 10124
rect 19358 10084 19800 10112
rect 19358 10081 19370 10084
rect 19312 10075 19370 10081
rect 19794 10072 19800 10084
rect 19852 10072 19858 10124
rect 20806 10072 20812 10124
rect 20864 10112 20870 10124
rect 20901 10115 20959 10121
rect 20901 10112 20913 10115
rect 20864 10084 20913 10112
rect 20864 10072 20870 10084
rect 20901 10081 20913 10084
rect 20947 10081 20959 10115
rect 20901 10075 20959 10081
rect 18230 10044 18236 10056
rect 17972 10016 18236 10044
rect 18230 10004 18236 10016
rect 18288 10004 18294 10056
rect 7098 9976 7104 9988
rect 4126 9948 7104 9976
rect 3970 9868 3976 9920
rect 4028 9908 4034 9920
rect 4126 9908 4154 9948
rect 7098 9936 7104 9948
rect 7156 9936 7162 9988
rect 7190 9936 7196 9988
rect 7248 9976 7254 9988
rect 7377 9979 7435 9985
rect 7377 9976 7389 9979
rect 7248 9948 7389 9976
rect 7248 9936 7254 9948
rect 7377 9945 7389 9948
rect 7423 9976 7435 9979
rect 10428 9976 10456 10004
rect 12066 9976 12072 9988
rect 7423 9948 10456 9976
rect 12027 9948 12072 9976
rect 7423 9945 7435 9948
rect 7377 9939 7435 9945
rect 12066 9936 12072 9948
rect 12124 9936 12130 9988
rect 13722 9976 13728 9988
rect 13683 9948 13728 9976
rect 13722 9936 13728 9948
rect 13780 9936 13786 9988
rect 21082 9976 21088 9988
rect 21043 9948 21088 9976
rect 21082 9936 21088 9948
rect 21140 9936 21146 9988
rect 4614 9908 4620 9920
rect 4028 9880 4154 9908
rect 4575 9880 4620 9908
rect 4028 9868 4034 9880
rect 4614 9868 4620 9880
rect 4672 9868 4678 9920
rect 13081 9911 13139 9917
rect 13081 9877 13093 9911
rect 13127 9908 13139 9911
rect 13538 9908 13544 9920
rect 13127 9880 13544 9908
rect 13127 9877 13139 9880
rect 13081 9871 13139 9877
rect 13538 9868 13544 9880
rect 13596 9868 13602 9920
rect 14918 9868 14924 9920
rect 14976 9908 14982 9920
rect 15562 9908 15568 9920
rect 14976 9880 15568 9908
rect 14976 9868 14982 9880
rect 15562 9868 15568 9880
rect 15620 9868 15626 9920
rect 19058 9908 19064 9920
rect 19019 9880 19064 9908
rect 19058 9868 19064 9880
rect 19116 9868 19122 9920
rect 19242 9868 19248 9920
rect 19300 9908 19306 9920
rect 19383 9911 19441 9917
rect 19383 9908 19395 9911
rect 19300 9880 19395 9908
rect 19300 9868 19306 9880
rect 19383 9877 19395 9880
rect 19429 9877 19441 9911
rect 19383 9871 19441 9877
rect 1104 9818 22816 9840
rect 1104 9766 4982 9818
rect 5034 9766 5046 9818
rect 5098 9766 5110 9818
rect 5162 9766 5174 9818
rect 5226 9766 12982 9818
rect 13034 9766 13046 9818
rect 13098 9766 13110 9818
rect 13162 9766 13174 9818
rect 13226 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 22816 9818
rect 1104 9744 22816 9766
rect 6270 9704 6276 9716
rect 6231 9676 6276 9704
rect 6270 9664 6276 9676
rect 6328 9664 6334 9716
rect 7098 9664 7104 9716
rect 7156 9704 7162 9716
rect 8389 9707 8447 9713
rect 8389 9704 8401 9707
rect 7156 9676 8401 9704
rect 7156 9664 7162 9676
rect 8389 9673 8401 9676
rect 8435 9704 8447 9707
rect 8846 9704 8852 9716
rect 8435 9676 8852 9704
rect 8435 9673 8447 9676
rect 8389 9667 8447 9673
rect 8846 9664 8852 9676
rect 8904 9664 8910 9716
rect 9401 9707 9459 9713
rect 9401 9673 9413 9707
rect 9447 9704 9459 9707
rect 9769 9707 9827 9713
rect 9769 9704 9781 9707
rect 9447 9676 9781 9704
rect 9447 9673 9459 9676
rect 9401 9667 9459 9673
rect 9769 9673 9781 9676
rect 9815 9704 9827 9707
rect 9858 9704 9864 9716
rect 9815 9676 9864 9704
rect 9815 9673 9827 9676
rect 9769 9667 9827 9673
rect 9858 9664 9864 9676
rect 9916 9664 9922 9716
rect 10042 9704 10048 9716
rect 10003 9676 10048 9704
rect 10042 9664 10048 9676
rect 10100 9664 10106 9716
rect 11379 9707 11437 9713
rect 11379 9673 11391 9707
rect 11425 9704 11437 9707
rect 12526 9704 12532 9716
rect 11425 9676 12532 9704
rect 11425 9673 11437 9676
rect 11379 9667 11437 9673
rect 12526 9664 12532 9676
rect 12584 9664 12590 9716
rect 15378 9664 15384 9716
rect 15436 9704 15442 9716
rect 17681 9707 17739 9713
rect 17681 9704 17693 9707
rect 15436 9676 17693 9704
rect 15436 9664 15442 9676
rect 17681 9673 17693 9676
rect 17727 9704 17739 9707
rect 18138 9704 18144 9716
rect 17727 9676 18144 9704
rect 17727 9673 17739 9676
rect 17681 9667 17739 9673
rect 18138 9664 18144 9676
rect 18196 9664 18202 9716
rect 12066 9636 12072 9648
rect 12027 9608 12072 9636
rect 12066 9596 12072 9608
rect 12124 9636 12130 9648
rect 12124 9608 12572 9636
rect 12124 9596 12130 9608
rect 1854 9528 1860 9580
rect 1912 9568 1918 9580
rect 2869 9571 2927 9577
rect 2869 9568 2881 9571
rect 1912 9540 2881 9568
rect 1912 9528 1918 9540
rect 2869 9537 2881 9540
rect 2915 9568 2927 9571
rect 3513 9571 3571 9577
rect 3513 9568 3525 9571
rect 2915 9540 3525 9568
rect 2915 9537 2927 9540
rect 2869 9531 2927 9537
rect 3513 9537 3525 9540
rect 3559 9537 3571 9571
rect 3513 9531 3571 9537
rect 5718 9528 5724 9580
rect 5776 9568 5782 9580
rect 6641 9571 6699 9577
rect 6641 9568 6653 9571
rect 5776 9540 6653 9568
rect 5776 9528 5782 9540
rect 6641 9537 6653 9540
rect 6687 9568 6699 9571
rect 8110 9568 8116 9580
rect 6687 9540 8116 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 2130 9500 2136 9512
rect 2091 9472 2136 9500
rect 2130 9460 2136 9472
rect 2188 9460 2194 9512
rect 2222 9460 2228 9512
rect 2280 9500 2286 9512
rect 2685 9503 2743 9509
rect 2685 9500 2697 9503
rect 2280 9472 2697 9500
rect 2280 9460 2286 9472
rect 2685 9469 2697 9472
rect 2731 9500 2743 9503
rect 4154 9500 4160 9512
rect 2731 9472 4160 9500
rect 2731 9469 2743 9472
rect 2685 9463 2743 9469
rect 4154 9460 4160 9472
rect 4212 9460 4218 9512
rect 4614 9500 4620 9512
rect 4575 9472 4620 9500
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 5169 9503 5227 9509
rect 5169 9469 5181 9503
rect 5215 9500 5227 9503
rect 5736 9500 5764 9528
rect 5215 9472 5764 9500
rect 5215 9469 5227 9472
rect 5169 9463 5227 9469
rect 2148 9432 2176 9460
rect 3145 9435 3203 9441
rect 3145 9432 3157 9435
rect 2148 9404 3157 9432
rect 3145 9401 3157 9404
rect 3191 9401 3203 9435
rect 4522 9432 4528 9444
rect 4435 9404 4528 9432
rect 3145 9395 3203 9401
rect 4522 9392 4528 9404
rect 4580 9432 4586 9444
rect 5184 9432 5212 9463
rect 6546 9460 6552 9512
rect 6604 9500 6610 9512
rect 6914 9500 6920 9512
rect 6604 9472 6920 9500
rect 6604 9460 6610 9472
rect 6914 9460 6920 9472
rect 6972 9460 6978 9512
rect 7484 9509 7512 9540
rect 8110 9528 8116 9540
rect 8168 9568 8174 9580
rect 11790 9568 11796 9580
rect 8168 9540 11796 9568
rect 8168 9528 8174 9540
rect 11790 9528 11796 9540
rect 11848 9528 11854 9580
rect 12544 9577 12572 9608
rect 13446 9596 13452 9648
rect 13504 9636 13510 9648
rect 14918 9636 14924 9648
rect 13504 9608 14924 9636
rect 13504 9596 13510 9608
rect 14918 9596 14924 9608
rect 14976 9596 14982 9648
rect 16666 9636 16672 9648
rect 16627 9608 16672 9636
rect 16666 9596 16672 9608
rect 16724 9596 16730 9648
rect 12529 9571 12587 9577
rect 12529 9537 12541 9571
rect 12575 9568 12587 9571
rect 12894 9568 12900 9580
rect 12575 9540 12900 9568
rect 12575 9537 12587 9540
rect 12529 9531 12587 9537
rect 12894 9528 12900 9540
rect 12952 9568 12958 9580
rect 13633 9571 13691 9577
rect 13633 9568 13645 9571
rect 12952 9540 13645 9568
rect 12952 9528 12958 9540
rect 13633 9537 13645 9540
rect 13679 9568 13691 9571
rect 13722 9568 13728 9580
rect 13679 9540 13728 9568
rect 13679 9537 13691 9540
rect 13633 9531 13691 9537
rect 13722 9528 13728 9540
rect 13780 9568 13786 9580
rect 14093 9571 14151 9577
rect 14093 9568 14105 9571
rect 13780 9540 14105 9568
rect 13780 9528 13786 9540
rect 14093 9537 14105 9540
rect 14139 9537 14151 9571
rect 14093 9531 14151 9537
rect 14737 9571 14795 9577
rect 14737 9537 14749 9571
rect 14783 9568 14795 9571
rect 15378 9568 15384 9580
rect 14783 9540 15384 9568
rect 14783 9537 14795 9540
rect 14737 9531 14795 9537
rect 15378 9528 15384 9540
rect 15436 9528 15442 9580
rect 16114 9568 16120 9580
rect 16075 9540 16120 9568
rect 16114 9528 16120 9540
rect 16172 9528 16178 9580
rect 18785 9571 18843 9577
rect 18785 9537 18797 9571
rect 18831 9568 18843 9571
rect 19242 9568 19248 9580
rect 18831 9540 19248 9568
rect 18831 9537 18843 9540
rect 18785 9531 18843 9537
rect 19242 9528 19248 9540
rect 19300 9528 19306 9580
rect 7469 9503 7527 9509
rect 7469 9469 7481 9503
rect 7515 9469 7527 9503
rect 7469 9463 7527 9469
rect 8481 9503 8539 9509
rect 8481 9469 8493 9503
rect 8527 9469 8539 9503
rect 8481 9463 8539 9469
rect 5350 9432 5356 9444
rect 4580 9404 5212 9432
rect 5311 9404 5356 9432
rect 4580 9392 4586 9404
rect 5350 9392 5356 9404
rect 5408 9392 5414 9444
rect 7653 9435 7711 9441
rect 7653 9401 7665 9435
rect 7699 9432 7711 9435
rect 7929 9435 7987 9441
rect 7929 9432 7941 9435
rect 7699 9404 7941 9432
rect 7699 9401 7711 9404
rect 7653 9395 7711 9401
rect 7929 9401 7941 9404
rect 7975 9432 7987 9435
rect 8496 9432 8524 9463
rect 9950 9460 9956 9512
rect 10008 9500 10014 9512
rect 10296 9503 10354 9509
rect 10296 9500 10308 9503
rect 10008 9472 10308 9500
rect 10008 9460 10014 9472
rect 10296 9469 10308 9472
rect 10342 9500 10354 9503
rect 11146 9500 11152 9512
rect 10342 9472 10824 9500
rect 11107 9472 11152 9500
rect 10342 9469 10354 9472
rect 10296 9463 10354 9469
rect 7975 9404 8524 9432
rect 7975 9401 7987 9404
rect 7929 9395 7987 9401
rect 8570 9392 8576 9444
rect 8628 9432 8634 9444
rect 10796 9441 10824 9472
rect 11146 9460 11152 9472
rect 11204 9500 11210 9512
rect 11276 9503 11334 9509
rect 11276 9500 11288 9503
rect 11204 9472 11288 9500
rect 11204 9460 11210 9472
rect 11276 9469 11288 9472
rect 11322 9469 11334 9503
rect 11276 9463 11334 9469
rect 11882 9460 11888 9512
rect 11940 9500 11946 9512
rect 12437 9503 12495 9509
rect 12437 9500 12449 9503
rect 11940 9472 12449 9500
rect 11940 9460 11946 9472
rect 12437 9469 12449 9472
rect 12483 9469 12495 9503
rect 12437 9463 12495 9469
rect 12713 9503 12771 9509
rect 12713 9469 12725 9503
rect 12759 9500 12771 9503
rect 13538 9500 13544 9512
rect 12759 9472 13544 9500
rect 12759 9469 12771 9472
rect 12713 9463 12771 9469
rect 13538 9460 13544 9472
rect 13596 9460 13602 9512
rect 13998 9500 14004 9512
rect 13959 9472 14004 9500
rect 13998 9460 14004 9472
rect 14056 9460 14062 9512
rect 14274 9500 14280 9512
rect 14187 9472 14280 9500
rect 14274 9460 14280 9472
rect 14332 9500 14338 9512
rect 15013 9503 15071 9509
rect 15013 9500 15025 9503
rect 14332 9472 15025 9500
rect 14332 9460 14338 9472
rect 15013 9469 15025 9472
rect 15059 9469 15071 9503
rect 15013 9463 15071 9469
rect 8802 9435 8860 9441
rect 8802 9432 8814 9435
rect 8628 9404 8814 9432
rect 8628 9392 8634 9404
rect 8802 9401 8814 9404
rect 8848 9401 8860 9435
rect 8802 9395 8860 9401
rect 10781 9435 10839 9441
rect 10781 9401 10793 9435
rect 10827 9432 10839 9435
rect 13630 9432 13636 9444
rect 10827 9404 13636 9432
rect 10827 9401 10839 9404
rect 10781 9395 10839 9401
rect 13630 9392 13636 9404
rect 13688 9392 13694 9444
rect 14016 9432 14044 9460
rect 15381 9435 15439 9441
rect 15381 9432 15393 9435
rect 14016 9404 15393 9432
rect 15381 9401 15393 9404
rect 15427 9401 15439 9435
rect 15381 9395 15439 9401
rect 16206 9392 16212 9444
rect 16264 9432 16270 9444
rect 18877 9435 18935 9441
rect 16264 9404 16309 9432
rect 16264 9392 16270 9404
rect 18877 9401 18889 9435
rect 18923 9432 18935 9435
rect 19058 9432 19064 9444
rect 18923 9404 19064 9432
rect 18923 9401 18935 9404
rect 18877 9395 18935 9401
rect 19058 9392 19064 9404
rect 19116 9392 19122 9444
rect 19429 9435 19487 9441
rect 19429 9401 19441 9435
rect 19475 9432 19487 9435
rect 19518 9432 19524 9444
rect 19475 9404 19524 9432
rect 19475 9401 19487 9404
rect 19429 9395 19487 9401
rect 19518 9392 19524 9404
rect 19576 9392 19582 9444
rect 19794 9432 19800 9444
rect 19755 9404 19800 9432
rect 19794 9392 19800 9404
rect 19852 9392 19858 9444
rect 1949 9367 2007 9373
rect 1949 9333 1961 9367
rect 1995 9364 2007 9367
rect 2590 9364 2596 9376
rect 1995 9336 2596 9364
rect 1995 9333 2007 9336
rect 1949 9327 2007 9333
rect 2590 9324 2596 9336
rect 2648 9324 2654 9376
rect 5718 9364 5724 9376
rect 5631 9336 5724 9364
rect 5718 9324 5724 9336
rect 5776 9364 5782 9376
rect 8588 9364 8616 9392
rect 5776 9336 8616 9364
rect 5776 9324 5782 9336
rect 10134 9324 10140 9376
rect 10192 9364 10198 9376
rect 10367 9367 10425 9373
rect 10367 9364 10379 9367
rect 10192 9336 10379 9364
rect 10192 9324 10198 9336
rect 10367 9333 10379 9336
rect 10413 9333 10425 9367
rect 10367 9327 10425 9333
rect 12802 9324 12808 9376
rect 12860 9364 12866 9376
rect 12897 9367 12955 9373
rect 12897 9364 12909 9367
rect 12860 9336 12909 9364
rect 12860 9324 12866 9336
rect 12897 9333 12909 9336
rect 12943 9333 12955 9367
rect 12897 9327 12955 9333
rect 15654 9324 15660 9376
rect 15712 9364 15718 9376
rect 15841 9367 15899 9373
rect 15841 9364 15853 9367
rect 15712 9336 15853 9364
rect 15712 9324 15718 9336
rect 15841 9333 15853 9336
rect 15887 9333 15899 9367
rect 15841 9327 15899 9333
rect 16758 9324 16764 9376
rect 16816 9364 16822 9376
rect 17037 9367 17095 9373
rect 17037 9364 17049 9367
rect 16816 9336 17049 9364
rect 16816 9324 16822 9336
rect 17037 9333 17049 9336
rect 17083 9333 17095 9367
rect 18230 9364 18236 9376
rect 18191 9336 18236 9364
rect 17037 9327 17095 9333
rect 18230 9324 18236 9336
rect 18288 9324 18294 9376
rect 20898 9364 20904 9376
rect 20859 9336 20904 9364
rect 20898 9324 20904 9336
rect 20956 9324 20962 9376
rect 1104 9274 22816 9296
rect 1104 9222 8982 9274
rect 9034 9222 9046 9274
rect 9098 9222 9110 9274
rect 9162 9222 9174 9274
rect 9226 9222 16982 9274
rect 17034 9222 17046 9274
rect 17098 9222 17110 9274
rect 17162 9222 17174 9274
rect 17226 9222 22816 9274
rect 1104 9200 22816 9222
rect 2222 9160 2228 9172
rect 2183 9132 2228 9160
rect 2222 9120 2228 9132
rect 2280 9120 2286 9172
rect 2406 9160 2412 9172
rect 2367 9132 2412 9160
rect 2406 9120 2412 9132
rect 2464 9120 2470 9172
rect 4798 9120 4804 9172
rect 4856 9160 4862 9172
rect 4985 9163 5043 9169
rect 4985 9160 4997 9163
rect 4856 9132 4997 9160
rect 4856 9120 4862 9132
rect 4985 9129 4997 9132
rect 5031 9129 5043 9163
rect 5718 9160 5724 9172
rect 5679 9132 5724 9160
rect 4985 9123 5043 9129
rect 5718 9120 5724 9132
rect 5776 9120 5782 9172
rect 6273 9163 6331 9169
rect 6273 9129 6285 9163
rect 6319 9160 6331 9163
rect 7098 9160 7104 9172
rect 6319 9132 7104 9160
rect 6319 9129 6331 9132
rect 6273 9123 6331 9129
rect 7098 9120 7104 9132
rect 7156 9160 7162 9172
rect 8570 9160 8576 9172
rect 7156 9132 7328 9160
rect 8531 9132 8576 9160
rect 7156 9120 7162 9132
rect 4522 9092 4528 9104
rect 4126 9064 4528 9092
rect 1854 8984 1860 9036
rect 1912 9024 1918 9036
rect 2130 9024 2136 9036
rect 1912 8996 2136 9024
rect 1912 8984 1918 8996
rect 2130 8984 2136 8996
rect 2188 9024 2194 9036
rect 2317 9027 2375 9033
rect 2317 9024 2329 9027
rect 2188 8996 2329 9024
rect 2188 8984 2194 8996
rect 2317 8993 2329 8996
rect 2363 8993 2375 9027
rect 2866 9024 2872 9036
rect 2779 8996 2872 9024
rect 2317 8987 2375 8993
rect 2866 8984 2872 8996
rect 2924 9024 2930 9036
rect 4126 9024 4154 9064
rect 4522 9052 4528 9064
rect 4580 9052 4586 9104
rect 6638 9092 6644 9104
rect 6599 9064 6644 9092
rect 6638 9052 6644 9064
rect 6696 9052 6702 9104
rect 6914 9092 6920 9104
rect 6875 9064 6920 9092
rect 6914 9052 6920 9064
rect 6972 9052 6978 9104
rect 7190 9092 7196 9104
rect 7151 9064 7196 9092
rect 7190 9052 7196 9064
rect 7248 9052 7254 9104
rect 7300 9101 7328 9132
rect 8570 9120 8576 9132
rect 8628 9120 8634 9172
rect 12894 9160 12900 9172
rect 12855 9132 12900 9160
rect 12894 9120 12900 9132
rect 12952 9120 12958 9172
rect 15102 9120 15108 9172
rect 15160 9160 15166 9172
rect 15160 9132 16160 9160
rect 15160 9120 15166 9132
rect 7285 9095 7343 9101
rect 7285 9061 7297 9095
rect 7331 9061 7343 9095
rect 9858 9092 9864 9104
rect 9819 9064 9864 9092
rect 7285 9055 7343 9061
rect 9858 9052 9864 9064
rect 9916 9052 9922 9104
rect 10410 9092 10416 9104
rect 10371 9064 10416 9092
rect 10410 9052 10416 9064
rect 10468 9052 10474 9104
rect 13262 9092 13268 9104
rect 12176 9064 13268 9092
rect 2924 8996 4154 9024
rect 2924 8984 2930 8996
rect 4246 8984 4252 9036
rect 4304 9024 4310 9036
rect 4341 9027 4399 9033
rect 4341 9024 4353 9027
rect 4304 8996 4353 9024
rect 4304 8984 4310 8996
rect 4341 8993 4353 8996
rect 4387 8993 4399 9027
rect 11882 9024 11888 9036
rect 11843 8996 11888 9024
rect 4341 8987 4399 8993
rect 11882 8984 11888 8996
rect 11940 8984 11946 9036
rect 11974 8984 11980 9036
rect 12032 9024 12038 9036
rect 12176 9033 12204 9064
rect 13262 9052 13268 9064
rect 13320 9092 13326 9104
rect 13449 9095 13507 9101
rect 13449 9092 13461 9095
rect 13320 9064 13461 9092
rect 13320 9052 13326 9064
rect 13449 9061 13461 9064
rect 13495 9061 13507 9095
rect 13449 9055 13507 9061
rect 15743 9095 15801 9101
rect 15743 9061 15755 9095
rect 15789 9061 15801 9095
rect 16132 9092 16160 9132
rect 16206 9120 16212 9172
rect 16264 9160 16270 9172
rect 16301 9163 16359 9169
rect 16301 9160 16313 9163
rect 16264 9132 16313 9160
rect 16264 9120 16270 9132
rect 16301 9129 16313 9132
rect 16347 9160 16359 9163
rect 16577 9163 16635 9169
rect 16577 9160 16589 9163
rect 16347 9132 16589 9160
rect 16347 9129 16359 9132
rect 16301 9123 16359 9129
rect 16577 9129 16589 9132
rect 16623 9129 16635 9163
rect 16577 9123 16635 9129
rect 18138 9120 18144 9172
rect 18196 9160 18202 9172
rect 18325 9163 18383 9169
rect 18325 9160 18337 9163
rect 18196 9132 18337 9160
rect 18196 9120 18202 9132
rect 18325 9129 18337 9132
rect 18371 9129 18383 9163
rect 18325 9123 18383 9129
rect 18877 9163 18935 9169
rect 18877 9129 18889 9163
rect 18923 9160 18935 9163
rect 19058 9160 19064 9172
rect 18923 9132 19064 9160
rect 18923 9129 18935 9132
rect 18877 9123 18935 9129
rect 19058 9120 19064 9132
rect 19116 9120 19122 9172
rect 19242 9160 19248 9172
rect 19203 9132 19248 9160
rect 19242 9120 19248 9132
rect 19300 9120 19306 9172
rect 16132 9064 18230 9092
rect 15743 9055 15801 9061
rect 12161 9027 12219 9033
rect 12161 9024 12173 9027
rect 12032 8996 12173 9024
rect 12032 8984 12038 8996
rect 12161 8993 12173 8996
rect 12207 8993 12219 9027
rect 13538 9024 13544 9036
rect 13499 8996 13544 9024
rect 12161 8987 12219 8993
rect 13538 8984 13544 8996
rect 13596 9024 13602 9036
rect 14274 9024 14280 9036
rect 13596 8996 14280 9024
rect 13596 8984 13602 8996
rect 14274 8984 14280 8996
rect 14332 8984 14338 9036
rect 15764 9024 15792 9055
rect 15838 9024 15844 9036
rect 15751 8996 15844 9024
rect 15838 8984 15844 8996
rect 15896 9024 15902 9036
rect 16298 9024 16304 9036
rect 15896 8996 16304 9024
rect 15896 8984 15902 8996
rect 16298 8984 16304 8996
rect 16356 8984 16362 9036
rect 16850 8984 16856 9036
rect 16908 9024 16914 9036
rect 17770 9024 17776 9036
rect 16908 8996 17776 9024
rect 16908 8984 16914 8996
rect 17770 8984 17776 8996
rect 17828 9024 17834 9036
rect 17957 9027 18015 9033
rect 17957 9024 17969 9027
rect 17828 8996 17969 9024
rect 17828 8984 17834 8996
rect 17957 8993 17969 8996
rect 18003 8993 18015 9027
rect 18202 9024 18230 9064
rect 19702 9024 19708 9036
rect 19760 9033 19766 9036
rect 19760 9027 19798 9033
rect 18202 8996 19708 9024
rect 17957 8987 18015 8993
rect 19702 8984 19708 8996
rect 19786 8993 19798 9027
rect 19760 8987 19798 8993
rect 19760 8984 19766 8987
rect 5350 8956 5356 8968
rect 5311 8928 5356 8956
rect 5350 8916 5356 8928
rect 5408 8916 5414 8968
rect 7466 8956 7472 8968
rect 7427 8928 7472 8956
rect 7466 8916 7472 8928
rect 7524 8916 7530 8968
rect 9582 8916 9588 8968
rect 9640 8956 9646 8968
rect 9769 8959 9827 8965
rect 9769 8956 9781 8959
rect 9640 8928 9781 8956
rect 9640 8916 9646 8928
rect 9769 8925 9781 8928
rect 9815 8925 9827 8959
rect 9769 8919 9827 8925
rect 10226 8916 10232 8968
rect 10284 8956 10290 8968
rect 12345 8959 12403 8965
rect 12345 8956 12357 8959
rect 10284 8928 12357 8956
rect 10284 8916 10290 8928
rect 12345 8925 12357 8928
rect 12391 8925 12403 8959
rect 12345 8919 12403 8925
rect 13722 8916 13728 8968
rect 13780 8956 13786 8968
rect 14461 8959 14519 8965
rect 14461 8956 14473 8959
rect 13780 8928 14473 8956
rect 13780 8916 13786 8928
rect 14461 8925 14473 8928
rect 14507 8925 14519 8959
rect 14461 8919 14519 8925
rect 15381 8959 15439 8965
rect 15381 8925 15393 8959
rect 15427 8956 15439 8959
rect 15470 8956 15476 8968
rect 15427 8928 15476 8956
rect 15427 8925 15439 8928
rect 15381 8919 15439 8925
rect 15470 8916 15476 8928
rect 15528 8916 15534 8968
rect 16316 8956 16344 8984
rect 18138 8956 18144 8968
rect 16316 8928 18144 8956
rect 18138 8916 18144 8928
rect 18196 8916 18202 8968
rect 4479 8891 4537 8897
rect 4479 8857 4491 8891
rect 4525 8888 4537 8891
rect 9674 8888 9680 8900
rect 4525 8860 9680 8888
rect 4525 8857 4537 8860
rect 4479 8851 4537 8857
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 11514 8848 11520 8900
rect 11572 8888 11578 8900
rect 11977 8891 12035 8897
rect 11977 8888 11989 8891
rect 11572 8860 11989 8888
rect 11572 8848 11578 8860
rect 11977 8857 11989 8860
rect 12023 8888 12035 8891
rect 13354 8888 13360 8900
rect 12023 8860 13360 8888
rect 12023 8857 12035 8860
rect 11977 8851 12035 8857
rect 13354 8848 13360 8860
rect 13412 8848 13418 8900
rect 11793 8823 11851 8829
rect 11793 8789 11805 8823
rect 11839 8820 11851 8823
rect 11882 8820 11888 8832
rect 11839 8792 11888 8820
rect 11839 8789 11851 8792
rect 11793 8783 11851 8789
rect 11882 8780 11888 8792
rect 11940 8820 11946 8832
rect 13265 8823 13323 8829
rect 13265 8820 13277 8823
rect 11940 8792 13277 8820
rect 11940 8780 11946 8792
rect 13265 8789 13277 8792
rect 13311 8789 13323 8823
rect 13265 8783 13323 8789
rect 18966 8780 18972 8832
rect 19024 8820 19030 8832
rect 19613 8823 19671 8829
rect 19613 8820 19625 8823
rect 19024 8792 19625 8820
rect 19024 8780 19030 8792
rect 19613 8789 19625 8792
rect 19659 8820 19671 8823
rect 19843 8823 19901 8829
rect 19843 8820 19855 8823
rect 19659 8792 19855 8820
rect 19659 8789 19671 8792
rect 19613 8783 19671 8789
rect 19843 8789 19855 8792
rect 19889 8789 19901 8823
rect 19843 8783 19901 8789
rect 1104 8730 22816 8752
rect 1104 8678 4982 8730
rect 5034 8678 5046 8730
rect 5098 8678 5110 8730
rect 5162 8678 5174 8730
rect 5226 8678 12982 8730
rect 13034 8678 13046 8730
rect 13098 8678 13110 8730
rect 13162 8678 13174 8730
rect 13226 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 22816 8730
rect 1104 8656 22816 8678
rect 2225 8619 2283 8625
rect 2225 8585 2237 8619
rect 2271 8616 2283 8619
rect 2866 8616 2872 8628
rect 2271 8588 2872 8616
rect 2271 8585 2283 8588
rect 2225 8579 2283 8585
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 5905 8619 5963 8625
rect 5905 8616 5917 8619
rect 5408 8588 5917 8616
rect 5408 8576 5414 8588
rect 5905 8585 5917 8588
rect 5951 8585 5963 8619
rect 5905 8579 5963 8585
rect 6641 8619 6699 8625
rect 6641 8585 6653 8619
rect 6687 8616 6699 8619
rect 7190 8616 7196 8628
rect 6687 8588 7196 8616
rect 6687 8585 6699 8588
rect 6641 8579 6699 8585
rect 7190 8576 7196 8588
rect 7248 8576 7254 8628
rect 11146 8616 11152 8628
rect 7300 8588 11152 8616
rect 1762 8508 1768 8560
rect 1820 8548 1826 8560
rect 2961 8551 3019 8557
rect 2961 8548 2973 8551
rect 1820 8520 2973 8548
rect 1820 8508 1826 8520
rect 2961 8517 2973 8520
rect 3007 8548 3019 8551
rect 6546 8548 6552 8560
rect 3007 8520 6552 8548
rect 3007 8517 3019 8520
rect 2961 8511 3019 8517
rect 6546 8508 6552 8520
rect 6604 8508 6610 8560
rect 2038 8440 2044 8492
rect 2096 8480 2102 8492
rect 2409 8483 2467 8489
rect 2409 8480 2421 8483
rect 2096 8452 2421 8480
rect 2096 8440 2102 8452
rect 2409 8449 2421 8452
rect 2455 8480 2467 8483
rect 3329 8483 3387 8489
rect 3329 8480 3341 8483
rect 2455 8452 3341 8480
rect 2455 8449 2467 8452
rect 2409 8443 2467 8449
rect 3329 8449 3341 8452
rect 3375 8449 3387 8483
rect 4246 8480 4252 8492
rect 4159 8452 4252 8480
rect 3329 8443 3387 8449
rect 4246 8440 4252 8452
rect 4304 8480 4310 8492
rect 7300 8480 7328 8588
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 11514 8616 11520 8628
rect 11475 8588 11520 8616
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 11885 8619 11943 8625
rect 11885 8585 11897 8619
rect 11931 8616 11943 8619
rect 11974 8616 11980 8628
rect 11931 8588 11980 8616
rect 11931 8585 11943 8588
rect 11885 8579 11943 8585
rect 11974 8576 11980 8588
rect 12032 8576 12038 8628
rect 12066 8576 12072 8628
rect 12124 8616 12130 8628
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 12124 8588 12173 8616
rect 12124 8576 12130 8588
rect 12161 8585 12173 8588
rect 12207 8585 12219 8619
rect 12161 8579 12219 8585
rect 8205 8551 8263 8557
rect 8205 8517 8217 8551
rect 8251 8548 8263 8551
rect 8570 8548 8576 8560
rect 8251 8520 8576 8548
rect 8251 8517 8263 8520
rect 8205 8511 8263 8517
rect 8570 8508 8576 8520
rect 8628 8508 8634 8560
rect 10318 8508 10324 8560
rect 10376 8548 10382 8560
rect 10689 8551 10747 8557
rect 10689 8548 10701 8551
rect 10376 8520 10701 8548
rect 10376 8508 10382 8520
rect 10689 8517 10701 8520
rect 10735 8517 10747 8551
rect 10689 8511 10747 8517
rect 10134 8480 10140 8492
rect 4304 8452 7328 8480
rect 10095 8452 10140 8480
rect 4304 8440 4310 8452
rect 10134 8440 10140 8452
rect 10192 8480 10198 8492
rect 11057 8483 11115 8489
rect 11057 8480 11069 8483
rect 10192 8452 11069 8480
rect 10192 8440 10198 8452
rect 11057 8449 11069 8452
rect 11103 8449 11115 8483
rect 11057 8443 11115 8449
rect 4338 8412 4344 8424
rect 4299 8384 4344 8412
rect 4338 8372 4344 8384
rect 4396 8372 4402 8424
rect 5629 8415 5687 8421
rect 5629 8381 5641 8415
rect 5675 8412 5687 8415
rect 5718 8412 5724 8424
rect 5675 8384 5724 8412
rect 5675 8381 5687 8384
rect 5629 8375 5687 8381
rect 2498 8304 2504 8356
rect 2556 8344 2562 8356
rect 4703 8347 4761 8353
rect 4703 8344 4715 8347
rect 2556 8316 2601 8344
rect 4126 8316 4715 8344
rect 2556 8304 2562 8316
rect 1854 8276 1860 8288
rect 1815 8248 1860 8276
rect 1854 8236 1860 8248
rect 1912 8236 1918 8288
rect 2590 8236 2596 8288
rect 2648 8276 2654 8288
rect 3789 8279 3847 8285
rect 3789 8276 3801 8279
rect 2648 8248 3801 8276
rect 2648 8236 2654 8248
rect 3789 8245 3801 8248
rect 3835 8276 3847 8279
rect 4126 8276 4154 8316
rect 4703 8313 4715 8316
rect 4749 8344 4761 8347
rect 5644 8344 5672 8375
rect 5718 8372 5724 8384
rect 5776 8372 5782 8424
rect 6730 8372 6736 8424
rect 6788 8412 6794 8424
rect 6892 8415 6950 8421
rect 6892 8412 6904 8415
rect 6788 8384 6904 8412
rect 6788 8372 6794 8384
rect 6892 8381 6904 8384
rect 6938 8381 6950 8415
rect 7834 8412 7840 8424
rect 7747 8384 7840 8412
rect 6892 8375 6950 8381
rect 4749 8316 5672 8344
rect 6907 8344 6935 8375
rect 7834 8372 7840 8384
rect 7892 8412 7898 8424
rect 8297 8415 8355 8421
rect 8297 8412 8309 8415
rect 7892 8384 8309 8412
rect 7892 8372 7898 8384
rect 8297 8381 8309 8384
rect 8343 8381 8355 8415
rect 8297 8375 8355 8381
rect 9217 8415 9275 8421
rect 9217 8381 9229 8415
rect 9263 8412 9275 8415
rect 12176 8412 12204 8579
rect 15378 8576 15384 8628
rect 15436 8616 15442 8628
rect 15838 8616 15844 8628
rect 15436 8588 15844 8616
rect 15436 8576 15442 8588
rect 15838 8576 15844 8588
rect 15896 8576 15902 8628
rect 16206 8616 16212 8628
rect 16167 8588 16212 8616
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 17770 8616 17776 8628
rect 17731 8588 17776 8616
rect 17770 8576 17776 8588
rect 17828 8576 17834 8628
rect 18138 8576 18144 8628
rect 18196 8616 18202 8628
rect 18233 8619 18291 8625
rect 18233 8616 18245 8619
rect 18196 8588 18245 8616
rect 18196 8576 18202 8588
rect 18233 8585 18245 8588
rect 18279 8585 18291 8619
rect 19702 8616 19708 8628
rect 19663 8588 19708 8616
rect 18233 8579 18291 8585
rect 19702 8576 19708 8588
rect 19760 8576 19766 8628
rect 16666 8508 16672 8560
rect 16724 8548 16730 8560
rect 16724 8520 19104 8548
rect 16724 8508 16730 8520
rect 13173 8483 13231 8489
rect 13173 8449 13185 8483
rect 13219 8480 13231 8483
rect 13354 8480 13360 8492
rect 13219 8452 13360 8480
rect 13219 8449 13231 8452
rect 13173 8443 13231 8449
rect 13354 8440 13360 8452
rect 13412 8440 13418 8492
rect 16393 8483 16451 8489
rect 16393 8449 16405 8483
rect 16439 8480 16451 8483
rect 16758 8480 16764 8492
rect 16439 8452 16764 8480
rect 16439 8449 16451 8452
rect 16393 8443 16451 8449
rect 16758 8440 16764 8452
rect 16816 8440 16822 8492
rect 18785 8483 18843 8489
rect 18785 8449 18797 8483
rect 18831 8480 18843 8483
rect 18966 8480 18972 8492
rect 18831 8452 18972 8480
rect 18831 8449 18843 8452
rect 18785 8443 18843 8449
rect 18966 8440 18972 8452
rect 19024 8440 19030 8492
rect 19076 8489 19104 8520
rect 19061 8483 19119 8489
rect 19061 8449 19073 8483
rect 19107 8480 19119 8483
rect 19242 8480 19248 8492
rect 19107 8452 19248 8480
rect 19107 8449 19119 8452
rect 19061 8443 19119 8449
rect 19242 8440 19248 8452
rect 19300 8440 19306 8492
rect 12529 8415 12587 8421
rect 12529 8412 12541 8415
rect 9263 8384 9812 8412
rect 12176 8384 12541 8412
rect 9263 8381 9275 8384
rect 9217 8375 9275 8381
rect 7374 8344 7380 8356
rect 6907 8316 7380 8344
rect 4749 8313 4761 8316
rect 4703 8307 4761 8313
rect 7374 8304 7380 8316
rect 7432 8304 7438 8356
rect 9784 8353 9812 8384
rect 12529 8381 12541 8384
rect 12575 8412 12587 8415
rect 12802 8412 12808 8424
rect 12575 8384 12808 8412
rect 12575 8381 12587 8384
rect 12529 8375 12587 8381
rect 12802 8372 12808 8384
rect 12860 8372 12866 8424
rect 14918 8412 14924 8424
rect 14879 8384 14924 8412
rect 14918 8372 14924 8384
rect 14976 8372 14982 8424
rect 15289 8415 15347 8421
rect 15289 8381 15301 8415
rect 15335 8412 15347 8415
rect 15654 8412 15660 8424
rect 15335 8384 15660 8412
rect 15335 8381 15347 8384
rect 15289 8375 15347 8381
rect 9769 8347 9827 8353
rect 9769 8313 9781 8347
rect 9815 8344 9827 8347
rect 9858 8344 9864 8356
rect 9815 8316 9864 8344
rect 9815 8313 9827 8316
rect 9769 8307 9827 8313
rect 9858 8304 9864 8316
rect 9916 8344 9922 8356
rect 10229 8347 10287 8353
rect 10229 8344 10241 8347
rect 9916 8316 10241 8344
rect 9916 8304 9922 8316
rect 10229 8313 10241 8316
rect 10275 8344 10287 8347
rect 10410 8344 10416 8356
rect 10275 8316 10416 8344
rect 10275 8313 10287 8316
rect 10229 8307 10287 8313
rect 10410 8304 10416 8316
rect 10468 8304 10474 8356
rect 14645 8347 14703 8353
rect 14645 8313 14657 8347
rect 14691 8344 14703 8347
rect 15304 8344 15332 8375
rect 15654 8372 15660 8384
rect 15712 8372 15718 8424
rect 15470 8344 15476 8356
rect 14691 8316 15332 8344
rect 15431 8316 15476 8344
rect 14691 8313 14703 8316
rect 14645 8307 14703 8313
rect 15470 8304 15476 8316
rect 15528 8304 15534 8356
rect 16485 8347 16543 8353
rect 16485 8313 16497 8347
rect 16531 8313 16543 8347
rect 16485 8307 16543 8313
rect 5258 8276 5264 8288
rect 3835 8248 4154 8276
rect 5219 8248 5264 8276
rect 3835 8245 3847 8248
rect 3789 8239 3847 8245
rect 5258 8236 5264 8248
rect 5316 8236 5322 8288
rect 6822 8236 6828 8288
rect 6880 8276 6886 8288
rect 6963 8279 7021 8285
rect 6963 8276 6975 8279
rect 6880 8248 6975 8276
rect 6880 8236 6886 8248
rect 6963 8245 6975 8248
rect 7009 8245 7021 8279
rect 6963 8239 7021 8245
rect 8570 8236 8576 8288
rect 8628 8276 8634 8288
rect 8665 8279 8723 8285
rect 8665 8276 8677 8279
rect 8628 8248 8677 8276
rect 8628 8236 8634 8248
rect 8665 8245 8677 8248
rect 8711 8245 8723 8279
rect 8665 8239 8723 8245
rect 13541 8279 13599 8285
rect 13541 8245 13553 8279
rect 13587 8276 13599 8279
rect 13630 8276 13636 8288
rect 13587 8248 13636 8276
rect 13587 8245 13599 8248
rect 13541 8239 13599 8245
rect 13630 8236 13636 8248
rect 13688 8236 13694 8288
rect 16206 8236 16212 8288
rect 16264 8276 16270 8288
rect 16500 8276 16528 8307
rect 16574 8304 16580 8356
rect 16632 8344 16638 8356
rect 17037 8347 17095 8353
rect 17037 8344 17049 8347
rect 16632 8316 17049 8344
rect 16632 8304 16638 8316
rect 17037 8313 17049 8316
rect 17083 8344 17095 8347
rect 18877 8347 18935 8353
rect 17083 8316 18368 8344
rect 17083 8313 17095 8316
rect 17037 8307 17095 8313
rect 16264 8248 16528 8276
rect 18340 8276 18368 8316
rect 18877 8313 18889 8347
rect 18923 8344 18935 8347
rect 19058 8344 19064 8356
rect 18923 8316 19064 8344
rect 18923 8313 18935 8316
rect 18877 8307 18935 8313
rect 19058 8304 19064 8316
rect 19116 8304 19122 8356
rect 19518 8276 19524 8288
rect 18340 8248 19524 8276
rect 16264 8236 16270 8248
rect 19518 8236 19524 8248
rect 19576 8236 19582 8288
rect 1104 8186 22816 8208
rect 1104 8134 8982 8186
rect 9034 8134 9046 8186
rect 9098 8134 9110 8186
rect 9162 8134 9174 8186
rect 9226 8134 16982 8186
rect 17034 8134 17046 8186
rect 17098 8134 17110 8186
rect 17162 8134 17174 8186
rect 17226 8134 22816 8186
rect 1104 8112 22816 8134
rect 1949 8075 2007 8081
rect 1949 8041 1961 8075
rect 1995 8072 2007 8075
rect 2498 8072 2504 8084
rect 1995 8044 2504 8072
rect 1995 8041 2007 8044
rect 1949 8035 2007 8041
rect 2498 8032 2504 8044
rect 2556 8072 2562 8084
rect 2961 8075 3019 8081
rect 2961 8072 2973 8075
rect 2556 8044 2973 8072
rect 2556 8032 2562 8044
rect 2961 8041 2973 8044
rect 3007 8041 3019 8075
rect 4338 8072 4344 8084
rect 4299 8044 4344 8072
rect 2961 8035 3019 8041
rect 4338 8032 4344 8044
rect 4396 8072 4402 8084
rect 5077 8075 5135 8081
rect 5077 8072 5089 8075
rect 4396 8044 5089 8072
rect 4396 8032 4402 8044
rect 5077 8041 5089 8044
rect 5123 8041 5135 8075
rect 7098 8072 7104 8084
rect 7059 8044 7104 8072
rect 5077 8035 5135 8041
rect 7098 8032 7104 8044
rect 7156 8032 7162 8084
rect 7834 8072 7840 8084
rect 7795 8044 7840 8072
rect 7834 8032 7840 8044
rect 7892 8032 7898 8084
rect 9493 8075 9551 8081
rect 9493 8041 9505 8075
rect 9539 8072 9551 8075
rect 9582 8072 9588 8084
rect 9539 8044 9588 8072
rect 9539 8041 9551 8044
rect 9493 8035 9551 8041
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 10410 8072 10416 8084
rect 10371 8044 10416 8072
rect 10410 8032 10416 8044
rect 10468 8032 10474 8084
rect 11974 8032 11980 8084
rect 12032 8072 12038 8084
rect 12345 8075 12403 8081
rect 12345 8072 12357 8075
rect 12032 8044 12357 8072
rect 12032 8032 12038 8044
rect 12345 8041 12357 8044
rect 12391 8041 12403 8075
rect 12345 8035 12403 8041
rect 2403 8007 2461 8013
rect 2403 7973 2415 8007
rect 2449 8004 2461 8007
rect 2590 8004 2596 8016
rect 2449 7976 2596 8004
rect 2449 7973 2461 7976
rect 2403 7967 2461 7973
rect 2590 7964 2596 7976
rect 2648 7964 2654 8016
rect 5258 7964 5264 8016
rect 5316 8004 5322 8016
rect 5902 8004 5908 8016
rect 5316 7976 5908 8004
rect 5316 7964 5322 7976
rect 5902 7964 5908 7976
rect 5960 8004 5966 8016
rect 5997 8007 6055 8013
rect 5997 8004 6009 8007
rect 5960 7976 6009 8004
rect 5960 7964 5966 7976
rect 5997 7973 6009 7976
rect 6043 7973 6055 8007
rect 6546 8004 6552 8016
rect 6459 7976 6552 8004
rect 5997 7967 6055 7973
rect 6546 7964 6552 7976
rect 6604 8004 6610 8016
rect 7466 8004 7472 8016
rect 6604 7976 7472 8004
rect 6604 7964 6610 7976
rect 7466 7964 7472 7976
rect 7524 7964 7530 8016
rect 3694 7896 3700 7948
rect 3752 7936 3758 7948
rect 4065 7939 4123 7945
rect 4065 7936 4077 7939
rect 3752 7908 4077 7936
rect 3752 7896 3758 7908
rect 4065 7905 4077 7908
rect 4111 7905 4123 7939
rect 4522 7936 4528 7948
rect 4483 7908 4528 7936
rect 4065 7899 4123 7905
rect 4522 7896 4528 7908
rect 4580 7896 4586 7948
rect 7742 7936 7748 7948
rect 7703 7908 7748 7936
rect 7742 7896 7748 7908
rect 7800 7896 7806 7948
rect 8110 7936 8116 7948
rect 8071 7908 8116 7936
rect 8110 7896 8116 7908
rect 8168 7896 8174 7948
rect 9950 7936 9956 7948
rect 9911 7908 9956 7936
rect 9950 7896 9956 7908
rect 10008 7896 10014 7948
rect 11124 7939 11182 7945
rect 11124 7905 11136 7939
rect 11170 7936 11182 7939
rect 11330 7936 11336 7948
rect 11170 7908 11336 7936
rect 11170 7905 11182 7908
rect 11124 7899 11182 7905
rect 11330 7896 11336 7908
rect 11388 7896 11394 7948
rect 2041 7871 2099 7877
rect 2041 7837 2053 7871
rect 2087 7868 2099 7871
rect 2406 7868 2412 7880
rect 2087 7840 2412 7868
rect 2087 7837 2099 7840
rect 2041 7831 2099 7837
rect 2406 7828 2412 7840
rect 2464 7828 2470 7880
rect 5905 7871 5963 7877
rect 5905 7837 5917 7871
rect 5951 7868 5963 7871
rect 6270 7868 6276 7880
rect 5951 7840 6276 7868
rect 5951 7837 5963 7840
rect 5905 7831 5963 7837
rect 6270 7828 6276 7840
rect 6328 7868 6334 7880
rect 7282 7868 7288 7880
rect 6328 7840 7288 7868
rect 6328 7828 6334 7840
rect 7282 7828 7288 7840
rect 7340 7828 7346 7880
rect 12360 7868 12388 8035
rect 12618 8032 12624 8084
rect 12676 8072 12682 8084
rect 13173 8075 13231 8081
rect 13173 8072 13185 8075
rect 12676 8044 13185 8072
rect 12676 8032 12682 8044
rect 13173 8041 13185 8044
rect 13219 8041 13231 8075
rect 15470 8072 15476 8084
rect 15431 8044 15476 8072
rect 13173 8035 13231 8041
rect 15470 8032 15476 8044
rect 15528 8032 15534 8084
rect 18785 8075 18843 8081
rect 18785 8041 18797 8075
rect 18831 8072 18843 8075
rect 19058 8072 19064 8084
rect 18831 8044 19064 8072
rect 18831 8041 18843 8044
rect 18785 8035 18843 8041
rect 19058 8032 19064 8044
rect 19116 8032 19122 8084
rect 15838 8004 15844 8016
rect 15799 7976 15844 8004
rect 15838 7964 15844 7976
rect 15896 7964 15902 8016
rect 16393 8007 16451 8013
rect 16393 7973 16405 8007
rect 16439 8004 16451 8007
rect 16574 8004 16580 8016
rect 16439 7976 16580 8004
rect 16439 7973 16451 7976
rect 16393 7967 16451 7973
rect 16574 7964 16580 7976
rect 16632 7964 16638 8016
rect 19150 8004 19156 8016
rect 19111 7976 19156 8004
rect 19150 7964 19156 7976
rect 19208 7964 19214 8016
rect 12529 7939 12587 7945
rect 12529 7905 12541 7939
rect 12575 7936 12587 7939
rect 12618 7936 12624 7948
rect 12575 7908 12624 7936
rect 12575 7905 12587 7908
rect 12529 7899 12587 7905
rect 12618 7896 12624 7908
rect 12676 7896 12682 7948
rect 14093 7939 14151 7945
rect 14093 7905 14105 7939
rect 14139 7936 14151 7939
rect 14182 7936 14188 7948
rect 14139 7908 14188 7936
rect 14139 7905 14151 7908
rect 14093 7899 14151 7905
rect 14182 7896 14188 7908
rect 14240 7896 14246 7948
rect 17678 7936 17684 7948
rect 17639 7908 17684 7936
rect 17678 7896 17684 7908
rect 17736 7896 17742 7948
rect 17865 7939 17923 7945
rect 17865 7905 17877 7939
rect 17911 7905 17923 7939
rect 17865 7899 17923 7905
rect 12897 7871 12955 7877
rect 12897 7868 12909 7871
rect 12360 7840 12909 7868
rect 12897 7837 12909 7840
rect 12943 7837 12955 7871
rect 12897 7831 12955 7837
rect 14323 7871 14381 7877
rect 14323 7837 14335 7871
rect 14369 7868 14381 7871
rect 15749 7871 15807 7877
rect 15749 7868 15761 7871
rect 14369 7840 15761 7868
rect 14369 7837 14381 7840
rect 14323 7831 14381 7837
rect 15749 7837 15761 7840
rect 15795 7868 15807 7871
rect 16482 7868 16488 7880
rect 15795 7840 16488 7868
rect 15795 7837 15807 7840
rect 15749 7831 15807 7837
rect 16482 7828 16488 7840
rect 16540 7828 16546 7880
rect 17586 7828 17592 7880
rect 17644 7868 17650 7880
rect 17880 7868 17908 7899
rect 17644 7840 17908 7868
rect 18141 7871 18199 7877
rect 17644 7828 17650 7840
rect 18141 7837 18153 7871
rect 18187 7868 18199 7871
rect 18414 7868 18420 7880
rect 18187 7840 18420 7868
rect 18187 7837 18199 7840
rect 18141 7831 18199 7837
rect 18414 7828 18420 7840
rect 18472 7828 18478 7880
rect 19061 7871 19119 7877
rect 19061 7837 19073 7871
rect 19107 7868 19119 7871
rect 19518 7868 19524 7880
rect 19107 7840 19524 7868
rect 19107 7837 19119 7840
rect 19061 7831 19119 7837
rect 19518 7828 19524 7840
rect 19576 7828 19582 7880
rect 12694 7803 12752 7809
rect 12694 7769 12706 7803
rect 12740 7800 12752 7803
rect 13354 7800 13360 7812
rect 12740 7772 13360 7800
rect 12740 7769 12752 7772
rect 12694 7763 12752 7769
rect 13354 7760 13360 7772
rect 13412 7800 13418 7812
rect 13909 7803 13967 7809
rect 13909 7800 13921 7803
rect 13412 7772 13921 7800
rect 13412 7760 13418 7772
rect 13909 7769 13921 7772
rect 13955 7769 13967 7803
rect 19610 7800 19616 7812
rect 19571 7772 19616 7800
rect 13909 7763 13967 7769
rect 19610 7760 19616 7772
rect 19668 7760 19674 7812
rect 4798 7692 4804 7744
rect 4856 7732 4862 7744
rect 5445 7735 5503 7741
rect 5445 7732 5457 7735
rect 4856 7704 5457 7732
rect 4856 7692 4862 7704
rect 5445 7701 5457 7704
rect 5491 7701 5503 7735
rect 5445 7695 5503 7701
rect 8478 7692 8484 7744
rect 8536 7732 8542 7744
rect 8573 7735 8631 7741
rect 8573 7732 8585 7735
rect 8536 7704 8585 7732
rect 8536 7692 8542 7704
rect 8573 7701 8585 7704
rect 8619 7701 8631 7735
rect 8573 7695 8631 7701
rect 10091 7735 10149 7741
rect 10091 7701 10103 7735
rect 10137 7732 10149 7735
rect 10318 7732 10324 7744
rect 10137 7704 10324 7732
rect 10137 7701 10149 7704
rect 10091 7695 10149 7701
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 10778 7692 10784 7744
rect 10836 7732 10842 7744
rect 10873 7735 10931 7741
rect 10873 7732 10885 7735
rect 10836 7704 10885 7732
rect 10836 7692 10842 7704
rect 10873 7701 10885 7704
rect 10919 7732 10931 7735
rect 11195 7735 11253 7741
rect 11195 7732 11207 7735
rect 10919 7704 11207 7732
rect 10919 7701 10931 7704
rect 10873 7695 10931 7701
rect 11195 7701 11207 7704
rect 11241 7701 11253 7735
rect 11974 7732 11980 7744
rect 11935 7704 11980 7732
rect 11195 7695 11253 7701
rect 11974 7692 11980 7704
rect 12032 7692 12038 7744
rect 12802 7732 12808 7744
rect 12763 7704 12808 7732
rect 12802 7692 12808 7704
rect 12860 7692 12866 7744
rect 13538 7732 13544 7744
rect 13499 7704 13544 7732
rect 13538 7692 13544 7704
rect 13596 7692 13602 7744
rect 14829 7735 14887 7741
rect 14829 7701 14841 7735
rect 14875 7732 14887 7735
rect 14918 7732 14924 7744
rect 14875 7704 14924 7732
rect 14875 7701 14887 7704
rect 14829 7695 14887 7701
rect 14918 7692 14924 7704
rect 14976 7732 14982 7744
rect 15746 7732 15752 7744
rect 14976 7704 15752 7732
rect 14976 7692 14982 7704
rect 15746 7692 15752 7704
rect 15804 7692 15810 7744
rect 16758 7732 16764 7744
rect 16719 7704 16764 7732
rect 16758 7692 16764 7704
rect 16816 7692 16822 7744
rect 16942 7692 16948 7744
rect 17000 7732 17006 7744
rect 20438 7732 20444 7744
rect 17000 7704 20444 7732
rect 17000 7692 17006 7704
rect 20438 7692 20444 7704
rect 20496 7692 20502 7744
rect 1104 7642 22816 7664
rect 1104 7590 4982 7642
rect 5034 7590 5046 7642
rect 5098 7590 5110 7642
rect 5162 7590 5174 7642
rect 5226 7590 12982 7642
rect 13034 7590 13046 7642
rect 13098 7590 13110 7642
rect 13162 7590 13174 7642
rect 13226 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 22816 7642
rect 1104 7568 22816 7590
rect 2406 7488 2412 7540
rect 2464 7528 2470 7540
rect 2869 7531 2927 7537
rect 2869 7528 2881 7531
rect 2464 7500 2881 7528
rect 2464 7488 2470 7500
rect 2869 7497 2881 7500
rect 2915 7497 2927 7531
rect 4522 7528 4528 7540
rect 4483 7500 4528 7528
rect 2869 7491 2927 7497
rect 4522 7488 4528 7500
rect 4580 7488 4586 7540
rect 5902 7528 5908 7540
rect 5863 7500 5908 7528
rect 5902 7488 5908 7500
rect 5960 7488 5966 7540
rect 6270 7528 6276 7540
rect 6231 7500 6276 7528
rect 6270 7488 6276 7500
rect 6328 7488 6334 7540
rect 8018 7528 8024 7540
rect 7979 7500 8024 7528
rect 8018 7488 8024 7500
rect 8076 7488 8082 7540
rect 8389 7531 8447 7537
rect 8389 7497 8401 7531
rect 8435 7528 8447 7531
rect 8570 7528 8576 7540
rect 8435 7500 8576 7528
rect 8435 7497 8447 7500
rect 8389 7491 8447 7497
rect 8570 7488 8576 7500
rect 8628 7488 8634 7540
rect 11330 7488 11336 7540
rect 11388 7528 11394 7540
rect 11701 7531 11759 7537
rect 11701 7528 11713 7531
rect 11388 7500 11713 7528
rect 11388 7488 11394 7500
rect 11701 7497 11713 7500
rect 11747 7497 11759 7531
rect 11701 7491 11759 7497
rect 12713 7531 12771 7537
rect 12713 7497 12725 7531
rect 12759 7528 12771 7531
rect 12802 7528 12808 7540
rect 12759 7500 12808 7528
rect 12759 7497 12771 7500
rect 12713 7491 12771 7497
rect 12802 7488 12808 7500
rect 12860 7528 12866 7540
rect 13081 7531 13139 7537
rect 13081 7528 13093 7531
rect 12860 7500 13093 7528
rect 12860 7488 12866 7500
rect 13081 7497 13093 7500
rect 13127 7528 13139 7531
rect 13541 7531 13599 7537
rect 13541 7528 13553 7531
rect 13127 7500 13553 7528
rect 13127 7497 13139 7500
rect 13081 7491 13139 7497
rect 13541 7497 13553 7500
rect 13587 7497 13599 7531
rect 13541 7491 13599 7497
rect 7377 7463 7435 7469
rect 7377 7429 7389 7463
rect 7423 7460 7435 7463
rect 8110 7460 8116 7472
rect 7423 7432 8116 7460
rect 7423 7429 7435 7432
rect 7377 7423 7435 7429
rect 8110 7420 8116 7432
rect 8168 7420 8174 7472
rect 13556 7460 13584 7491
rect 13722 7488 13728 7540
rect 13780 7528 13786 7540
rect 15194 7528 15200 7540
rect 13780 7500 15200 7528
rect 13780 7488 13786 7500
rect 15194 7488 15200 7500
rect 15252 7488 15258 7540
rect 15565 7531 15623 7537
rect 15565 7497 15577 7531
rect 15611 7528 15623 7531
rect 16942 7528 16948 7540
rect 15611 7500 16948 7528
rect 15611 7497 15623 7500
rect 15565 7491 15623 7497
rect 14642 7460 14648 7472
rect 13556 7432 14648 7460
rect 14642 7420 14648 7432
rect 14700 7420 14706 7472
rect 15580 7460 15608 7491
rect 16942 7488 16948 7500
rect 17000 7488 17006 7540
rect 17678 7488 17684 7540
rect 17736 7528 17742 7540
rect 17773 7531 17831 7537
rect 17773 7528 17785 7531
rect 17736 7500 17785 7528
rect 17736 7488 17742 7500
rect 17773 7497 17785 7500
rect 17819 7528 17831 7531
rect 17862 7528 17868 7540
rect 17819 7500 17868 7528
rect 17819 7497 17831 7500
rect 17773 7491 17831 7497
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 18969 7531 19027 7537
rect 18969 7497 18981 7531
rect 19015 7528 19027 7531
rect 19150 7528 19156 7540
rect 19015 7500 19156 7528
rect 19015 7497 19027 7500
rect 18969 7491 19027 7497
rect 19150 7488 19156 7500
rect 19208 7488 19214 7540
rect 16666 7460 16672 7472
rect 15079 7432 15608 7460
rect 16627 7432 16672 7460
rect 2038 7392 2044 7404
rect 1999 7364 2044 7392
rect 2038 7352 2044 7364
rect 2096 7352 2102 7404
rect 4798 7392 4804 7404
rect 4759 7364 4804 7392
rect 4798 7352 4804 7364
rect 4856 7352 4862 7404
rect 6454 7352 6460 7404
rect 6512 7392 6518 7404
rect 9950 7392 9956 7404
rect 6512 7364 9956 7392
rect 6512 7352 6518 7364
rect 9950 7352 9956 7364
rect 10008 7352 10014 7404
rect 10778 7392 10784 7404
rect 10739 7364 10784 7392
rect 10778 7352 10784 7364
rect 10836 7352 10842 7404
rect 10962 7352 10968 7404
rect 11020 7392 11026 7404
rect 11057 7395 11115 7401
rect 11057 7392 11069 7395
rect 11020 7364 11069 7392
rect 11020 7352 11026 7364
rect 11057 7361 11069 7364
rect 11103 7361 11115 7395
rect 11057 7355 11115 7361
rect 12894 7352 12900 7404
rect 12952 7392 12958 7404
rect 13354 7392 13360 7404
rect 12952 7364 13360 7392
rect 12952 7352 12958 7364
rect 13354 7352 13360 7364
rect 13412 7401 13418 7404
rect 13412 7395 13470 7401
rect 13412 7361 13424 7395
rect 13458 7361 13470 7395
rect 13630 7392 13636 7404
rect 13591 7364 13636 7392
rect 13412 7355 13470 7361
rect 13412 7352 13418 7355
rect 13630 7352 13636 7364
rect 13688 7352 13694 7404
rect 3786 7333 3792 7336
rect 3764 7327 3792 7333
rect 3764 7324 3776 7327
rect 3699 7296 3776 7324
rect 3764 7293 3776 7296
rect 3844 7324 3850 7336
rect 4157 7327 4215 7333
rect 4157 7324 4169 7327
rect 3844 7296 4169 7324
rect 3764 7287 3792 7293
rect 3786 7284 3792 7287
rect 3844 7284 3850 7296
rect 4157 7293 4169 7296
rect 4203 7293 4215 7327
rect 4157 7287 4215 7293
rect 7520 7327 7578 7333
rect 7520 7293 7532 7327
rect 7566 7324 7578 7327
rect 8018 7324 8024 7336
rect 7566 7296 8024 7324
rect 7566 7293 7578 7296
rect 7520 7287 7578 7293
rect 8018 7284 8024 7296
rect 8076 7284 8082 7336
rect 8478 7324 8484 7336
rect 8439 7296 8484 7324
rect 8478 7284 8484 7296
rect 8536 7284 8542 7336
rect 8570 7284 8576 7336
rect 8628 7324 8634 7336
rect 12253 7327 12311 7333
rect 8628 7296 8845 7324
rect 8628 7284 8634 7296
rect 4893 7259 4951 7265
rect 4893 7225 4905 7259
rect 4939 7256 4951 7259
rect 4982 7256 4988 7268
rect 4939 7228 4988 7256
rect 4939 7225 4951 7228
rect 4893 7219 4951 7225
rect 4982 7216 4988 7228
rect 5040 7216 5046 7268
rect 5445 7259 5503 7265
rect 5445 7225 5457 7259
rect 5491 7256 5503 7259
rect 6546 7256 6552 7268
rect 5491 7228 6552 7256
rect 5491 7225 5503 7228
rect 5445 7219 5503 7225
rect 6546 7216 6552 7228
rect 6604 7216 6610 7268
rect 7607 7259 7665 7265
rect 7607 7225 7619 7259
rect 7653 7256 7665 7259
rect 8662 7256 8668 7268
rect 7653 7228 8668 7256
rect 7653 7225 7665 7228
rect 7607 7219 7665 7225
rect 8662 7216 8668 7228
rect 8720 7216 8726 7268
rect 8817 7265 8845 7296
rect 12253 7293 12265 7327
rect 12299 7324 12311 7327
rect 12618 7324 12624 7336
rect 12299 7296 12624 7324
rect 12299 7293 12311 7296
rect 12253 7287 12311 7293
rect 12618 7284 12624 7296
rect 12676 7324 12682 7336
rect 13265 7327 13323 7333
rect 13265 7324 13277 7327
rect 12676 7296 13277 7324
rect 12676 7284 12682 7296
rect 13265 7293 13277 7296
rect 13311 7324 13323 7327
rect 13538 7324 13544 7336
rect 13311 7296 13544 7324
rect 13311 7293 13323 7296
rect 13265 7287 13323 7293
rect 13538 7284 13544 7296
rect 13596 7284 13602 7336
rect 15079 7333 15107 7432
rect 16666 7420 16672 7432
rect 16724 7420 16730 7472
rect 18506 7420 18512 7472
rect 18564 7460 18570 7472
rect 19610 7460 19616 7472
rect 18564 7432 19616 7460
rect 18564 7420 18570 7432
rect 19610 7420 19616 7432
rect 19668 7460 19674 7472
rect 19705 7463 19763 7469
rect 19705 7460 19717 7463
rect 19668 7432 19717 7460
rect 19668 7420 19674 7432
rect 19705 7429 19717 7432
rect 19751 7429 19763 7463
rect 19705 7423 19763 7429
rect 15151 7395 15209 7401
rect 15151 7361 15163 7395
rect 15197 7392 15209 7395
rect 16117 7395 16175 7401
rect 16117 7392 16129 7395
rect 15197 7364 16129 7392
rect 15197 7361 15209 7364
rect 15151 7355 15209 7361
rect 16117 7361 16129 7364
rect 16163 7392 16175 7395
rect 17037 7395 17095 7401
rect 17037 7392 17049 7395
rect 16163 7364 17049 7392
rect 16163 7361 16175 7364
rect 16117 7355 16175 7361
rect 17037 7361 17049 7364
rect 17083 7361 17095 7395
rect 17037 7355 17095 7361
rect 19153 7395 19211 7401
rect 19153 7361 19165 7395
rect 19199 7392 19211 7395
rect 19242 7392 19248 7404
rect 19199 7364 19248 7392
rect 19199 7361 19211 7364
rect 19153 7355 19211 7361
rect 19242 7352 19248 7364
rect 19300 7392 19306 7404
rect 20073 7395 20131 7401
rect 20073 7392 20085 7395
rect 19300 7364 20085 7392
rect 19300 7352 19306 7364
rect 20073 7361 20085 7364
rect 20119 7361 20131 7395
rect 20073 7355 20131 7361
rect 15064 7327 15122 7333
rect 15064 7324 15076 7327
rect 13786 7296 15076 7324
rect 8802 7259 8860 7265
rect 8802 7225 8814 7259
rect 8848 7225 8860 7259
rect 10505 7259 10563 7265
rect 10505 7256 10517 7259
rect 8802 7219 8860 7225
rect 9692 7228 10517 7256
rect 9692 7200 9720 7228
rect 10505 7225 10517 7228
rect 10551 7256 10563 7259
rect 10873 7259 10931 7265
rect 10873 7256 10885 7259
rect 10551 7228 10885 7256
rect 10551 7225 10563 7228
rect 10505 7219 10563 7225
rect 10873 7225 10885 7228
rect 10919 7225 10931 7259
rect 10873 7219 10931 7225
rect 12710 7216 12716 7268
rect 12768 7256 12774 7268
rect 13786 7256 13814 7296
rect 15064 7293 15076 7296
rect 15110 7293 15122 7327
rect 15064 7287 15122 7293
rect 12768 7228 13814 7256
rect 14001 7259 14059 7265
rect 12768 7216 12774 7228
rect 14001 7225 14013 7259
rect 14047 7256 14059 7259
rect 14090 7256 14096 7268
rect 14047 7228 14096 7256
rect 14047 7225 14059 7228
rect 14001 7219 14059 7225
rect 14090 7216 14096 7228
rect 14148 7216 14154 7268
rect 14921 7259 14979 7265
rect 14921 7225 14933 7259
rect 14967 7256 14979 7259
rect 15838 7256 15844 7268
rect 14967 7228 15844 7256
rect 14967 7225 14979 7228
rect 14921 7219 14979 7225
rect 15838 7216 15844 7228
rect 15896 7256 15902 7268
rect 16206 7256 16212 7268
rect 15896 7228 16212 7256
rect 15896 7216 15902 7228
rect 16206 7216 16212 7228
rect 16264 7216 16270 7268
rect 19245 7259 19303 7265
rect 19245 7225 19257 7259
rect 19291 7225 19303 7259
rect 19245 7219 19303 7225
rect 2590 7188 2596 7200
rect 2503 7160 2596 7188
rect 2590 7148 2596 7160
rect 2648 7188 2654 7200
rect 3142 7188 3148 7200
rect 2648 7160 3148 7188
rect 2648 7148 2654 7160
rect 3142 7148 3148 7160
rect 3200 7148 3206 7200
rect 3605 7191 3663 7197
rect 3605 7157 3617 7191
rect 3651 7188 3663 7191
rect 3694 7188 3700 7200
rect 3651 7160 3700 7188
rect 3651 7157 3663 7160
rect 3605 7151 3663 7157
rect 3694 7148 3700 7160
rect 3752 7148 3758 7200
rect 3835 7191 3893 7197
rect 3835 7157 3847 7191
rect 3881 7188 3893 7191
rect 4430 7188 4436 7200
rect 3881 7160 4436 7188
rect 3881 7157 3893 7160
rect 3835 7151 3893 7157
rect 4430 7148 4436 7160
rect 4488 7148 4494 7200
rect 9401 7191 9459 7197
rect 9401 7157 9413 7191
rect 9447 7188 9459 7191
rect 9674 7188 9680 7200
rect 9447 7160 9680 7188
rect 9447 7157 9459 7160
rect 9401 7151 9459 7157
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 14182 7148 14188 7200
rect 14240 7188 14246 7200
rect 14277 7191 14335 7197
rect 14277 7188 14289 7191
rect 14240 7160 14289 7188
rect 14240 7148 14246 7160
rect 14277 7157 14289 7160
rect 14323 7157 14335 7191
rect 14277 7151 14335 7157
rect 17497 7191 17555 7197
rect 17497 7157 17509 7191
rect 17543 7188 17555 7191
rect 17586 7188 17592 7200
rect 17543 7160 17592 7188
rect 17543 7157 17555 7160
rect 17497 7151 17555 7157
rect 17586 7148 17592 7160
rect 17644 7148 17650 7200
rect 18601 7191 18659 7197
rect 18601 7157 18613 7191
rect 18647 7188 18659 7191
rect 19260 7188 19288 7219
rect 19334 7188 19340 7200
rect 18647 7160 19340 7188
rect 18647 7157 18659 7160
rect 18601 7151 18659 7157
rect 19334 7148 19340 7160
rect 19392 7148 19398 7200
rect 20806 7188 20812 7200
rect 20767 7160 20812 7188
rect 20806 7148 20812 7160
rect 20864 7148 20870 7200
rect 1104 7098 22816 7120
rect 1104 7046 8982 7098
rect 9034 7046 9046 7098
rect 9098 7046 9110 7098
rect 9162 7046 9174 7098
rect 9226 7046 16982 7098
rect 17034 7046 17046 7098
rect 17098 7046 17110 7098
rect 17162 7046 17174 7098
rect 17226 7046 22816 7098
rect 1104 7024 22816 7046
rect 3099 6987 3157 6993
rect 3099 6953 3111 6987
rect 3145 6984 3157 6987
rect 4798 6984 4804 6996
rect 3145 6956 4804 6984
rect 3145 6953 3157 6956
rect 3099 6947 3157 6953
rect 4798 6944 4804 6956
rect 4856 6944 4862 6996
rect 6822 6944 6828 6996
rect 6880 6984 6886 6996
rect 6917 6987 6975 6993
rect 6917 6984 6929 6987
rect 6880 6956 6929 6984
rect 6880 6944 6886 6956
rect 6917 6953 6929 6956
rect 6963 6953 6975 6987
rect 6917 6947 6975 6953
rect 7653 6987 7711 6993
rect 7653 6953 7665 6987
rect 7699 6984 7711 6987
rect 7742 6984 7748 6996
rect 7699 6956 7748 6984
rect 7699 6953 7711 6956
rect 7653 6947 7711 6953
rect 7742 6944 7748 6956
rect 7800 6944 7806 6996
rect 9674 6944 9680 6996
rect 9732 6984 9738 6996
rect 16206 6984 16212 6996
rect 9732 6956 10456 6984
rect 9732 6944 9738 6956
rect 4709 6919 4767 6925
rect 4709 6885 4721 6919
rect 4755 6916 4767 6919
rect 4982 6916 4988 6928
rect 4755 6888 4988 6916
rect 4755 6885 4767 6888
rect 4709 6879 4767 6885
rect 4982 6876 4988 6888
rect 5040 6916 5046 6928
rect 5077 6919 5135 6925
rect 5077 6916 5089 6919
rect 5040 6888 5089 6916
rect 5040 6876 5046 6888
rect 5077 6885 5089 6888
rect 5123 6916 5135 6919
rect 5718 6916 5724 6928
rect 5123 6888 5724 6916
rect 5123 6885 5135 6888
rect 5077 6879 5135 6885
rect 5718 6876 5724 6888
rect 5776 6876 5782 6928
rect 8478 6916 8484 6928
rect 8439 6888 8484 6916
rect 8478 6876 8484 6888
rect 8536 6876 8542 6928
rect 10318 6916 10324 6928
rect 10279 6888 10324 6916
rect 10318 6876 10324 6888
rect 10376 6876 10382 6928
rect 10428 6925 10456 6956
rect 13786 6956 15792 6984
rect 16167 6956 16212 6984
rect 10413 6919 10471 6925
rect 10413 6885 10425 6919
rect 10459 6885 10471 6919
rect 10413 6879 10471 6885
rect 11146 6876 11152 6928
rect 11204 6916 11210 6928
rect 13786 6916 13814 6956
rect 11204 6888 13814 6916
rect 11204 6876 11210 6888
rect 15378 6876 15384 6928
rect 15436 6916 15442 6928
rect 15610 6919 15668 6925
rect 15610 6916 15622 6919
rect 15436 6888 15622 6916
rect 15436 6876 15442 6888
rect 15610 6885 15622 6888
rect 15656 6885 15668 6919
rect 15764 6916 15792 6956
rect 16206 6944 16212 6956
rect 16264 6944 16270 6996
rect 16482 6984 16488 6996
rect 16443 6956 16488 6984
rect 16482 6944 16488 6956
rect 16540 6944 16546 6996
rect 16758 6944 16764 6996
rect 16816 6984 16822 6996
rect 17175 6987 17233 6993
rect 17175 6984 17187 6987
rect 16816 6956 17187 6984
rect 16816 6944 16822 6956
rect 17175 6953 17187 6956
rect 17221 6953 17233 6987
rect 17175 6947 17233 6953
rect 19150 6944 19156 6996
rect 19208 6984 19214 6996
rect 19245 6987 19303 6993
rect 19245 6984 19257 6987
rect 19208 6956 19257 6984
rect 19208 6944 19214 6956
rect 19245 6953 19257 6956
rect 19291 6953 19303 6987
rect 19518 6984 19524 6996
rect 19479 6956 19524 6984
rect 19245 6947 19303 6953
rect 19518 6944 19524 6956
rect 19576 6944 19582 6996
rect 21039 6987 21097 6993
rect 21039 6953 21051 6987
rect 21085 6984 21097 6987
rect 21266 6984 21272 6996
rect 21085 6956 21272 6984
rect 21085 6953 21097 6956
rect 21039 6947 21097 6953
rect 21266 6944 21272 6956
rect 21324 6944 21330 6996
rect 15764 6888 17126 6916
rect 15610 6879 15668 6885
rect 17098 6860 17126 6888
rect 18138 6876 18144 6928
rect 18196 6916 18202 6928
rect 18646 6919 18704 6925
rect 18646 6916 18658 6919
rect 18196 6888 18658 6916
rect 18196 6876 18202 6888
rect 18646 6885 18658 6888
rect 18692 6885 18704 6919
rect 18646 6879 18704 6885
rect 1464 6851 1522 6857
rect 1464 6817 1476 6851
rect 1510 6848 1522 6851
rect 1762 6848 1768 6860
rect 1510 6820 1768 6848
rect 1510 6817 1522 6820
rect 1464 6811 1522 6817
rect 1762 6808 1768 6820
rect 1820 6808 1826 6860
rect 2682 6808 2688 6860
rect 2740 6848 2746 6860
rect 3028 6851 3086 6857
rect 3028 6848 3040 6851
rect 2740 6820 3040 6848
rect 2740 6808 2746 6820
rect 3028 6817 3040 6820
rect 3074 6848 3086 6851
rect 3510 6848 3516 6860
rect 3074 6820 3516 6848
rect 3074 6817 3086 6820
rect 3028 6811 3086 6817
rect 3510 6808 3516 6820
rect 3568 6808 3574 6860
rect 6454 6848 6460 6860
rect 6415 6820 6460 6848
rect 6454 6808 6460 6820
rect 6512 6808 6518 6860
rect 6914 6808 6920 6860
rect 6972 6848 6978 6860
rect 7558 6848 7564 6860
rect 6972 6820 7564 6848
rect 6972 6808 6978 6820
rect 7558 6808 7564 6820
rect 7616 6848 7622 6860
rect 7745 6851 7803 6857
rect 7745 6848 7757 6851
rect 7616 6820 7757 6848
rect 7616 6808 7622 6820
rect 7745 6817 7757 6820
rect 7791 6817 7803 6851
rect 7745 6811 7803 6817
rect 7926 6808 7932 6860
rect 7984 6848 7990 6860
rect 11882 6857 11888 6860
rect 8205 6851 8263 6857
rect 8205 6848 8217 6851
rect 7984 6820 8217 6848
rect 7984 6808 7990 6820
rect 8205 6817 8217 6820
rect 8251 6817 8263 6851
rect 11860 6851 11888 6857
rect 11860 6848 11872 6851
rect 11795 6820 11872 6848
rect 8205 6811 8263 6817
rect 11860 6817 11872 6820
rect 11940 6848 11946 6860
rect 12802 6848 12808 6860
rect 11940 6820 12808 6848
rect 11860 6811 11888 6817
rect 11882 6808 11888 6811
rect 11940 6808 11946 6820
rect 12802 6808 12808 6820
rect 12860 6808 12866 6860
rect 13906 6848 13912 6860
rect 13819 6820 13912 6848
rect 13906 6808 13912 6820
rect 13964 6848 13970 6860
rect 13964 6820 14044 6848
rect 13964 6808 13970 6820
rect 4430 6740 4436 6792
rect 4488 6780 4494 6792
rect 4798 6780 4804 6792
rect 4488 6752 4804 6780
rect 4488 6740 4494 6752
rect 4798 6740 4804 6752
rect 4856 6780 4862 6792
rect 4985 6783 5043 6789
rect 4985 6780 4997 6783
rect 4856 6752 4997 6780
rect 4856 6740 4862 6752
rect 4985 6749 4997 6752
rect 5031 6749 5043 6783
rect 4985 6743 5043 6749
rect 5629 6783 5687 6789
rect 5629 6749 5641 6783
rect 5675 6780 5687 6783
rect 7190 6780 7196 6792
rect 5675 6752 7196 6780
rect 5675 6749 5687 6752
rect 5629 6743 5687 6749
rect 7190 6740 7196 6752
rect 7248 6740 7254 6792
rect 10594 6780 10600 6792
rect 10555 6752 10600 6780
rect 10594 6740 10600 6752
rect 10652 6740 10658 6792
rect 13262 6712 13268 6724
rect 13223 6684 13268 6712
rect 13262 6672 13268 6684
rect 13320 6712 13326 6724
rect 13630 6712 13636 6724
rect 13320 6684 13636 6712
rect 13320 6672 13326 6684
rect 13630 6672 13636 6684
rect 13688 6672 13694 6724
rect 14016 6712 14044 6820
rect 14090 6808 14096 6860
rect 14148 6848 14154 6860
rect 14185 6851 14243 6857
rect 14185 6848 14197 6851
rect 14148 6820 14197 6848
rect 14148 6808 14154 6820
rect 14185 6817 14197 6820
rect 14231 6848 14243 6851
rect 15470 6848 15476 6860
rect 14231 6820 15476 6848
rect 14231 6817 14243 6820
rect 14185 6811 14243 6817
rect 15470 6808 15476 6820
rect 15528 6808 15534 6860
rect 17098 6851 17132 6860
rect 17098 6848 17116 6851
rect 17039 6820 17116 6848
rect 17104 6817 17116 6820
rect 17184 6848 17190 6860
rect 18874 6848 18880 6860
rect 17184 6820 18880 6848
rect 17104 6811 17132 6817
rect 17126 6808 17132 6811
rect 17184 6808 17190 6820
rect 18874 6808 18880 6820
rect 18932 6808 18938 6860
rect 20968 6851 21026 6857
rect 20968 6817 20980 6851
rect 21014 6848 21026 6851
rect 21450 6848 21456 6860
rect 21014 6820 21456 6848
rect 21014 6817 21026 6820
rect 20968 6811 21026 6817
rect 21450 6808 21456 6820
rect 21508 6808 21514 6860
rect 14369 6783 14427 6789
rect 14369 6749 14381 6783
rect 14415 6780 14427 6783
rect 15289 6783 15347 6789
rect 15289 6780 15301 6783
rect 14415 6752 15301 6780
rect 14415 6749 14427 6752
rect 14369 6743 14427 6749
rect 15289 6749 15301 6752
rect 15335 6780 15347 6783
rect 16574 6780 16580 6792
rect 15335 6752 16580 6780
rect 15335 6749 15347 6752
rect 15289 6743 15347 6749
rect 16574 6740 16580 6752
rect 16632 6740 16638 6792
rect 18138 6740 18144 6792
rect 18196 6780 18202 6792
rect 18325 6783 18383 6789
rect 18325 6780 18337 6783
rect 18196 6752 18337 6780
rect 18196 6740 18202 6752
rect 18325 6749 18337 6752
rect 18371 6749 18383 6783
rect 18325 6743 18383 6749
rect 14016 6684 14780 6712
rect 198 6604 204 6656
rect 256 6644 262 6656
rect 1535 6647 1593 6653
rect 1535 6644 1547 6647
rect 256 6616 1547 6644
rect 256 6604 262 6616
rect 1535 6613 1547 6616
rect 1581 6613 1593 6647
rect 1535 6607 1593 6613
rect 2869 6647 2927 6653
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 2958 6644 2964 6656
rect 2915 6616 2964 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 2958 6604 2964 6616
rect 3016 6604 3022 6656
rect 5902 6604 5908 6656
rect 5960 6644 5966 6656
rect 6595 6647 6653 6653
rect 6595 6644 6607 6647
rect 5960 6616 6607 6644
rect 5960 6604 5966 6616
rect 6595 6613 6607 6616
rect 6641 6613 6653 6647
rect 6595 6607 6653 6613
rect 10137 6647 10195 6653
rect 10137 6613 10149 6647
rect 10183 6644 10195 6647
rect 10318 6644 10324 6656
rect 10183 6616 10324 6644
rect 10183 6613 10195 6616
rect 10137 6607 10195 6613
rect 10318 6604 10324 6616
rect 10376 6644 10382 6656
rect 11931 6647 11989 6653
rect 11931 6644 11943 6647
rect 10376 6616 11943 6644
rect 10376 6604 10382 6616
rect 11931 6613 11943 6616
rect 11977 6613 11989 6647
rect 12618 6644 12624 6656
rect 12579 6616 12624 6644
rect 11931 6607 11989 6613
rect 12618 6604 12624 6616
rect 12676 6604 12682 6656
rect 12802 6604 12808 6656
rect 12860 6644 12866 6656
rect 14752 6653 14780 6684
rect 12897 6647 12955 6653
rect 12897 6644 12909 6647
rect 12860 6616 12909 6644
rect 12860 6604 12866 6616
rect 12897 6613 12909 6616
rect 12943 6613 12955 6647
rect 12897 6607 12955 6613
rect 14737 6647 14795 6653
rect 14737 6613 14749 6647
rect 14783 6644 14795 6647
rect 16666 6644 16672 6656
rect 14783 6616 16672 6644
rect 14783 6613 14795 6616
rect 14737 6607 14795 6613
rect 16666 6604 16672 6616
rect 16724 6644 16730 6656
rect 18230 6644 18236 6656
rect 16724 6616 18236 6644
rect 16724 6604 16730 6616
rect 18230 6604 18236 6616
rect 18288 6604 18294 6656
rect 1104 6554 22816 6576
rect 1104 6502 4982 6554
rect 5034 6502 5046 6554
rect 5098 6502 5110 6554
rect 5162 6502 5174 6554
rect 5226 6502 12982 6554
rect 13034 6502 13046 6554
rect 13098 6502 13110 6554
rect 13162 6502 13174 6554
rect 13226 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 22816 6554
rect 1104 6480 22816 6502
rect 1673 6443 1731 6449
rect 1673 6409 1685 6443
rect 1719 6440 1731 6443
rect 1762 6440 1768 6452
rect 1719 6412 1768 6440
rect 1719 6409 1731 6412
rect 1673 6403 1731 6409
rect 1762 6400 1768 6412
rect 1820 6400 1826 6452
rect 2682 6440 2688 6452
rect 2643 6412 2688 6440
rect 2682 6400 2688 6412
rect 2740 6400 2746 6452
rect 3697 6443 3755 6449
rect 3697 6409 3709 6443
rect 3743 6440 3755 6443
rect 5718 6440 5724 6452
rect 3743 6412 5724 6440
rect 3743 6409 3755 6412
rect 3697 6403 3755 6409
rect 5718 6400 5724 6412
rect 5776 6400 5782 6452
rect 8389 6443 8447 6449
rect 8389 6409 8401 6443
rect 8435 6440 8447 6443
rect 8570 6440 8576 6452
rect 8435 6412 8576 6440
rect 8435 6409 8447 6412
rect 8389 6403 8447 6409
rect 8570 6400 8576 6412
rect 8628 6400 8634 6452
rect 9674 6440 9680 6452
rect 9635 6412 9680 6440
rect 9674 6400 9680 6412
rect 9732 6400 9738 6452
rect 11514 6440 11520 6452
rect 11475 6412 11520 6440
rect 11514 6400 11520 6412
rect 11572 6440 11578 6452
rect 11790 6440 11796 6452
rect 11572 6412 11796 6440
rect 11572 6400 11578 6412
rect 11790 6400 11796 6412
rect 11848 6440 11854 6452
rect 12805 6443 12863 6449
rect 12805 6440 12817 6443
rect 11848 6412 12817 6440
rect 11848 6400 11854 6412
rect 12805 6409 12817 6412
rect 12851 6409 12863 6443
rect 12805 6403 12863 6409
rect 13725 6443 13783 6449
rect 13725 6409 13737 6443
rect 13771 6440 13783 6443
rect 14090 6440 14096 6452
rect 13771 6412 14096 6440
rect 13771 6409 13783 6412
rect 13725 6403 13783 6409
rect 14090 6400 14096 6412
rect 14148 6400 14154 6452
rect 15378 6440 15384 6452
rect 15339 6412 15384 6440
rect 15378 6400 15384 6412
rect 15436 6400 15442 6452
rect 16574 6440 16580 6452
rect 16535 6412 16580 6440
rect 16574 6400 16580 6412
rect 16632 6400 16638 6452
rect 17126 6440 17132 6452
rect 17087 6412 17132 6440
rect 17126 6400 17132 6412
rect 17184 6400 17190 6452
rect 17865 6443 17923 6449
rect 17865 6409 17877 6443
rect 17911 6440 17923 6443
rect 18046 6440 18052 6452
rect 17911 6412 18052 6440
rect 17911 6409 17923 6412
rect 17865 6403 17923 6409
rect 18046 6400 18052 6412
rect 18104 6440 18110 6452
rect 18233 6443 18291 6449
rect 18233 6440 18245 6443
rect 18104 6412 18245 6440
rect 18104 6400 18110 6412
rect 18233 6409 18245 6412
rect 18279 6409 18291 6443
rect 19334 6440 19340 6452
rect 19295 6412 19340 6440
rect 18233 6403 18291 6409
rect 4706 6332 4712 6384
rect 4764 6372 4770 6384
rect 6454 6372 6460 6384
rect 4764 6344 6460 6372
rect 4764 6332 4770 6344
rect 6454 6332 6460 6344
rect 6512 6332 6518 6384
rect 6822 6332 6828 6384
rect 6880 6372 6886 6384
rect 11882 6372 11888 6384
rect 6880 6344 6960 6372
rect 11843 6344 11888 6372
rect 6880 6332 6886 6344
rect 6932 6313 6960 6344
rect 11882 6332 11888 6344
rect 11940 6332 11946 6384
rect 12710 6381 12716 6384
rect 12694 6375 12716 6381
rect 12694 6341 12706 6375
rect 12694 6335 12716 6341
rect 12710 6332 12716 6335
rect 12768 6332 12774 6384
rect 6917 6307 6975 6313
rect 6917 6273 6929 6307
rect 6963 6273 6975 6307
rect 7190 6304 7196 6316
rect 7151 6276 7196 6304
rect 6917 6267 6975 6273
rect 7190 6264 7196 6276
rect 7248 6264 7254 6316
rect 10318 6304 10324 6316
rect 10279 6276 10324 6304
rect 10318 6264 10324 6276
rect 10376 6264 10382 6316
rect 10962 6304 10968 6316
rect 10923 6276 10968 6304
rect 10962 6264 10968 6276
rect 11020 6264 11026 6316
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 12176 6276 12909 6304
rect 2777 6239 2835 6245
rect 2777 6205 2789 6239
rect 2823 6236 2835 6239
rect 2958 6236 2964 6248
rect 2823 6208 2964 6236
rect 2823 6205 2835 6208
rect 2777 6199 2835 6205
rect 2958 6196 2964 6208
rect 3016 6196 3022 6248
rect 4065 6239 4123 6245
rect 4065 6205 4077 6239
rect 4111 6236 4123 6239
rect 4522 6236 4528 6248
rect 4111 6208 4528 6236
rect 4111 6205 4123 6208
rect 4065 6199 4123 6205
rect 4522 6196 4528 6208
rect 4580 6196 4586 6248
rect 5445 6239 5503 6245
rect 5445 6205 5457 6239
rect 5491 6236 5503 6239
rect 5994 6236 6000 6248
rect 5491 6208 6000 6236
rect 5491 6205 5503 6208
rect 5445 6199 5503 6205
rect 5994 6196 6000 6208
rect 6052 6196 6058 6248
rect 8478 6236 8484 6248
rect 8439 6208 8484 6236
rect 8478 6196 8484 6208
rect 8536 6196 8542 6248
rect 9401 6239 9459 6245
rect 9401 6205 9413 6239
rect 9447 6236 9459 6239
rect 10042 6236 10048 6248
rect 9447 6208 10048 6236
rect 9447 6205 9459 6208
rect 9401 6199 9459 6205
rect 10042 6196 10048 6208
rect 10100 6196 10106 6248
rect 6012 6168 6040 6196
rect 7009 6171 7067 6177
rect 7009 6168 7021 6171
rect 6012 6140 7021 6168
rect 7009 6137 7021 6140
rect 7055 6137 7067 6171
rect 7009 6131 7067 6137
rect 8570 6128 8576 6180
rect 8628 6168 8634 6180
rect 8802 6171 8860 6177
rect 8802 6168 8814 6171
rect 8628 6140 8814 6168
rect 8628 6128 8634 6140
rect 8802 6137 8814 6140
rect 8848 6137 8860 6171
rect 10060 6168 10088 6196
rect 10413 6171 10471 6177
rect 10413 6168 10425 6171
rect 10060 6140 10425 6168
rect 8802 6131 8860 6137
rect 10413 6137 10425 6140
rect 10459 6137 10471 6171
rect 10413 6131 10471 6137
rect 11698 6128 11704 6180
rect 11756 6168 11762 6180
rect 12176 6177 12204 6276
rect 12897 6273 12909 6276
rect 12943 6304 12955 6307
rect 13262 6304 13268 6316
rect 12943 6276 13268 6304
rect 12943 6273 12955 6276
rect 12897 6267 12955 6273
rect 13262 6264 13268 6276
rect 13320 6264 13326 6316
rect 14553 6307 14611 6313
rect 14553 6304 14565 6307
rect 13786 6276 14565 6304
rect 12529 6239 12587 6245
rect 12529 6205 12541 6239
rect 12575 6236 12587 6239
rect 12618 6236 12624 6248
rect 12575 6208 12624 6236
rect 12575 6205 12587 6208
rect 12529 6199 12587 6205
rect 12618 6196 12624 6208
rect 12676 6236 12682 6248
rect 13786 6236 13814 6276
rect 14553 6273 14565 6276
rect 14599 6273 14611 6307
rect 16114 6304 16120 6316
rect 16075 6276 16120 6304
rect 14553 6267 14611 6273
rect 16114 6264 16120 6276
rect 16172 6264 16178 6316
rect 14093 6239 14151 6245
rect 14093 6236 14105 6239
rect 12676 6208 13814 6236
rect 13924 6208 14105 6236
rect 12676 6196 12682 6208
rect 12161 6171 12219 6177
rect 12161 6168 12173 6171
rect 11756 6140 12173 6168
rect 11756 6128 11762 6140
rect 12161 6137 12173 6140
rect 12207 6137 12219 6171
rect 13262 6168 13268 6180
rect 13223 6140 13268 6168
rect 12161 6131 12219 6137
rect 13262 6128 13268 6140
rect 13320 6128 13326 6180
rect 13354 6128 13360 6180
rect 13412 6168 13418 6180
rect 13924 6168 13952 6208
rect 14093 6205 14105 6208
rect 14139 6236 14151 6239
rect 14277 6239 14335 6245
rect 14139 6208 14228 6236
rect 14139 6205 14151 6208
rect 14093 6199 14151 6205
rect 13412 6140 13952 6168
rect 14200 6168 14228 6208
rect 14277 6205 14289 6239
rect 14323 6236 14335 6239
rect 14366 6236 14372 6248
rect 14323 6208 14372 6236
rect 14323 6205 14335 6208
rect 14277 6199 14335 6205
rect 14366 6196 14372 6208
rect 14424 6196 14430 6248
rect 15841 6239 15899 6245
rect 15841 6205 15853 6239
rect 15887 6236 15899 6239
rect 15930 6236 15936 6248
rect 15887 6208 15936 6236
rect 15887 6205 15899 6208
rect 15841 6199 15899 6205
rect 15930 6196 15936 6208
rect 15988 6196 15994 6248
rect 16025 6239 16083 6245
rect 16025 6205 16037 6239
rect 16071 6236 16083 6239
rect 17586 6236 17592 6248
rect 16071 6208 17592 6236
rect 16071 6205 16083 6208
rect 16025 6199 16083 6205
rect 14200 6140 14964 6168
rect 13412 6128 13418 6140
rect 14936 6112 14964 6140
rect 15654 6128 15660 6180
rect 15712 6168 15718 6180
rect 16040 6168 16068 6199
rect 17586 6196 17592 6208
rect 17644 6196 17650 6248
rect 15712 6140 16068 6168
rect 17497 6171 17555 6177
rect 15712 6128 15718 6140
rect 17497 6137 17509 6171
rect 17543 6168 17555 6171
rect 18138 6168 18144 6180
rect 17543 6140 18144 6168
rect 17543 6137 17555 6140
rect 17497 6131 17555 6137
rect 18138 6128 18144 6140
rect 18196 6128 18202 6180
rect 18248 6168 18276 6403
rect 19334 6400 19340 6412
rect 19392 6400 19398 6452
rect 21450 6440 21456 6452
rect 21411 6412 21456 6440
rect 21450 6400 21456 6412
rect 21508 6400 21514 6452
rect 18414 6304 18420 6316
rect 18375 6276 18420 6304
rect 18414 6264 18420 6276
rect 18472 6264 18478 6316
rect 20533 6239 20591 6245
rect 20533 6205 20545 6239
rect 20579 6205 20591 6239
rect 20533 6199 20591 6205
rect 18598 6168 18604 6180
rect 18248 6140 18604 6168
rect 18598 6128 18604 6140
rect 18656 6168 18662 6180
rect 18738 6171 18796 6177
rect 18738 6168 18750 6171
rect 18656 6140 18750 6168
rect 18656 6128 18662 6140
rect 18738 6137 18750 6140
rect 18784 6137 18796 6171
rect 18738 6131 18796 6137
rect 3142 6100 3148 6112
rect 3103 6072 3148 6100
rect 3142 6060 3148 6072
rect 3200 6100 3206 6112
rect 4433 6103 4491 6109
rect 4433 6100 4445 6103
rect 3200 6072 4445 6100
rect 3200 6060 3206 6072
rect 4433 6069 4445 6072
rect 4479 6100 4491 6103
rect 4893 6103 4951 6109
rect 4893 6100 4905 6103
rect 4479 6072 4905 6100
rect 4479 6069 4491 6072
rect 4433 6063 4491 6069
rect 4893 6069 4905 6072
rect 4939 6069 4951 6103
rect 7926 6100 7932 6112
rect 7887 6072 7932 6100
rect 4893 6063 4951 6069
rect 7926 6060 7932 6072
rect 7984 6060 7990 6112
rect 14918 6100 14924 6112
rect 14879 6072 14924 6100
rect 14918 6060 14924 6072
rect 14976 6060 14982 6112
rect 20349 6103 20407 6109
rect 20349 6069 20361 6103
rect 20395 6100 20407 6103
rect 20548 6100 20576 6199
rect 21174 6168 21180 6180
rect 21135 6140 21180 6168
rect 21174 6128 21180 6140
rect 21232 6128 21238 6180
rect 20714 6100 20720 6112
rect 20395 6072 20720 6100
rect 20395 6069 20407 6072
rect 20349 6063 20407 6069
rect 20714 6060 20720 6072
rect 20772 6060 20778 6112
rect 1104 6010 22816 6032
rect 1104 5958 8982 6010
rect 9034 5958 9046 6010
rect 9098 5958 9110 6010
rect 9162 5958 9174 6010
rect 9226 5958 16982 6010
rect 17034 5958 17046 6010
rect 17098 5958 17110 6010
rect 17162 5958 17174 6010
rect 17226 5958 22816 6010
rect 1104 5936 22816 5958
rect 4341 5899 4399 5905
rect 4341 5865 4353 5899
rect 4387 5896 4399 5899
rect 4522 5896 4528 5908
rect 4387 5868 4528 5896
rect 4387 5865 4399 5868
rect 4341 5859 4399 5865
rect 4522 5856 4528 5868
rect 4580 5856 4586 5908
rect 4798 5856 4804 5908
rect 4856 5896 4862 5908
rect 5077 5899 5135 5905
rect 5077 5896 5089 5899
rect 4856 5868 5089 5896
rect 4856 5856 4862 5868
rect 5077 5865 5089 5868
rect 5123 5865 5135 5899
rect 7558 5896 7564 5908
rect 5077 5859 5135 5865
rect 5184 5868 7564 5896
rect 5184 5828 5212 5868
rect 7558 5856 7564 5868
rect 7616 5856 7622 5908
rect 10410 5856 10416 5908
rect 10468 5896 10474 5908
rect 10873 5899 10931 5905
rect 10873 5896 10885 5899
rect 10468 5868 10885 5896
rect 10468 5856 10474 5868
rect 10873 5865 10885 5868
rect 10919 5865 10931 5899
rect 12069 5899 12127 5905
rect 12069 5896 12081 5899
rect 10873 5859 10931 5865
rect 11618 5868 12081 5896
rect 5902 5828 5908 5840
rect 4356 5800 5212 5828
rect 5863 5800 5908 5828
rect 4154 5720 4160 5772
rect 4212 5760 4218 5772
rect 4356 5769 4384 5800
rect 5902 5788 5908 5800
rect 5960 5788 5966 5840
rect 5994 5788 6000 5840
rect 6052 5828 6058 5840
rect 6825 5831 6883 5837
rect 6825 5828 6837 5831
rect 6052 5800 6837 5828
rect 6052 5788 6058 5800
rect 6825 5797 6837 5800
rect 6871 5797 6883 5831
rect 8478 5828 8484 5840
rect 8391 5800 8484 5828
rect 6825 5791 6883 5797
rect 8478 5788 8484 5800
rect 8536 5828 8542 5840
rect 8757 5831 8815 5837
rect 8757 5828 8769 5831
rect 8536 5800 8769 5828
rect 8536 5788 8542 5800
rect 8757 5797 8769 5800
rect 8803 5797 8815 5831
rect 10042 5828 10048 5840
rect 10003 5800 10048 5828
rect 8757 5791 8815 5797
rect 10042 5788 10048 5800
rect 10100 5788 10106 5840
rect 10594 5828 10600 5840
rect 10555 5800 10600 5828
rect 10594 5788 10600 5800
rect 10652 5788 10658 5840
rect 11618 5828 11646 5868
rect 12069 5865 12081 5868
rect 12115 5865 12127 5899
rect 15654 5896 15660 5908
rect 15615 5868 15660 5896
rect 12069 5859 12127 5865
rect 15654 5856 15660 5868
rect 15712 5856 15718 5908
rect 15930 5896 15936 5908
rect 15891 5868 15936 5896
rect 15930 5856 15936 5868
rect 15988 5896 15994 5908
rect 16298 5896 16304 5908
rect 15988 5868 16304 5896
rect 15988 5856 15994 5868
rect 16298 5856 16304 5868
rect 16356 5856 16362 5908
rect 18414 5856 18420 5908
rect 18472 5896 18478 5908
rect 18877 5899 18935 5905
rect 18877 5896 18889 5899
rect 18472 5868 18889 5896
rect 18472 5856 18478 5868
rect 18877 5865 18889 5868
rect 18923 5865 18935 5899
rect 18877 5859 18935 5865
rect 10704 5800 11646 5828
rect 12713 5831 12771 5837
rect 4341 5763 4399 5769
rect 4341 5760 4353 5763
rect 4212 5732 4353 5760
rect 4212 5720 4218 5732
rect 4341 5729 4353 5732
rect 4387 5729 4399 5763
rect 4341 5723 4399 5729
rect 4522 5720 4528 5772
rect 4580 5760 4586 5772
rect 4617 5763 4675 5769
rect 4617 5760 4629 5763
rect 4580 5732 4629 5760
rect 4580 5720 4586 5732
rect 4617 5729 4629 5732
rect 4663 5760 4675 5763
rect 4893 5763 4951 5769
rect 4893 5760 4905 5763
rect 4663 5732 4905 5760
rect 4663 5729 4675 5732
rect 4617 5723 4675 5729
rect 4893 5729 4905 5732
rect 4939 5729 4951 5763
rect 4893 5723 4951 5729
rect 6546 5720 6552 5772
rect 6604 5760 6610 5772
rect 7745 5763 7803 5769
rect 6604 5732 6649 5760
rect 6604 5720 6610 5732
rect 7745 5729 7757 5763
rect 7791 5729 7803 5763
rect 7745 5723 7803 5729
rect 7760 5692 7788 5723
rect 7926 5720 7932 5772
rect 7984 5760 7990 5772
rect 8297 5763 8355 5769
rect 8297 5760 8309 5763
rect 7984 5732 8309 5760
rect 7984 5720 7990 5732
rect 8297 5729 8309 5732
rect 8343 5729 8355 5763
rect 8297 5723 8355 5729
rect 7834 5692 7840 5704
rect 4126 5664 7840 5692
rect 4126 5568 4154 5664
rect 7834 5652 7840 5664
rect 7892 5652 7898 5704
rect 8312 5692 8340 5723
rect 8478 5692 8484 5704
rect 8312 5664 8484 5692
rect 8478 5652 8484 5664
rect 8536 5652 8542 5704
rect 8662 5652 8668 5704
rect 8720 5692 8726 5704
rect 9398 5692 9404 5704
rect 8720 5664 9404 5692
rect 8720 5652 8726 5664
rect 9398 5652 9404 5664
rect 9456 5692 9462 5704
rect 9953 5695 10011 5701
rect 9953 5692 9965 5695
rect 9456 5664 9965 5692
rect 9456 5652 9462 5664
rect 9953 5661 9965 5664
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 4893 5627 4951 5633
rect 4893 5593 4905 5627
rect 4939 5624 4951 5627
rect 9490 5624 9496 5636
rect 4939 5596 9496 5624
rect 4939 5593 4951 5596
rect 4893 5587 4951 5593
rect 9490 5584 9496 5596
rect 9548 5624 9554 5636
rect 10704 5624 10732 5800
rect 12713 5797 12725 5831
rect 12759 5828 12771 5831
rect 12802 5828 12808 5840
rect 12759 5800 12808 5828
rect 12759 5797 12771 5800
rect 12713 5791 12771 5797
rect 12802 5788 12808 5800
rect 12860 5828 12866 5840
rect 13265 5831 13323 5837
rect 13265 5828 13277 5831
rect 12860 5800 13277 5828
rect 12860 5788 12866 5800
rect 13265 5797 13277 5800
rect 13311 5828 13323 5831
rect 13311 5800 13676 5828
rect 13311 5797 13323 5800
rect 13265 5791 13323 5797
rect 13648 5772 13676 5800
rect 15378 5788 15384 5840
rect 15436 5828 15442 5840
rect 16438 5831 16496 5837
rect 16438 5828 16450 5831
rect 15436 5800 16450 5828
rect 15436 5788 15442 5800
rect 16438 5797 16450 5800
rect 16484 5797 16496 5831
rect 18046 5828 18052 5840
rect 16438 5791 16496 5797
rect 17052 5800 18052 5828
rect 11609 5763 11667 5769
rect 11609 5729 11621 5763
rect 11655 5729 11667 5763
rect 11609 5723 11667 5729
rect 9548 5596 10732 5624
rect 9548 5584 9554 5596
rect 2869 5559 2927 5565
rect 2869 5525 2881 5559
rect 2915 5556 2927 5559
rect 3142 5556 3148 5568
rect 2915 5528 3148 5556
rect 2915 5525 2927 5528
rect 2869 5519 2927 5525
rect 3142 5516 3148 5528
rect 3200 5516 3206 5568
rect 4062 5516 4068 5568
rect 4120 5528 4154 5568
rect 7190 5556 7196 5568
rect 7151 5528 7196 5556
rect 4120 5516 4126 5528
rect 7190 5516 7196 5528
rect 7248 5516 7254 5568
rect 11517 5559 11575 5565
rect 11517 5525 11529 5559
rect 11563 5556 11575 5559
rect 11624 5556 11652 5723
rect 11698 5720 11704 5772
rect 11756 5760 11762 5772
rect 11885 5763 11943 5769
rect 11885 5760 11897 5763
rect 11756 5732 11897 5760
rect 11756 5720 11762 5732
rect 11885 5729 11897 5732
rect 11931 5729 11943 5763
rect 13354 5760 13360 5772
rect 13315 5732 13360 5760
rect 11885 5723 11943 5729
rect 13354 5720 13360 5732
rect 13412 5720 13418 5772
rect 13630 5760 13636 5772
rect 13591 5732 13636 5760
rect 13630 5720 13636 5732
rect 13688 5720 13694 5772
rect 16114 5760 16120 5772
rect 16075 5732 16120 5760
rect 16114 5720 16120 5732
rect 16172 5720 16178 5772
rect 17052 5769 17080 5800
rect 18046 5788 18052 5800
rect 18104 5788 18110 5840
rect 20806 5788 20812 5840
rect 20864 5828 20870 5840
rect 20993 5831 21051 5837
rect 20993 5828 21005 5831
rect 20864 5800 21005 5828
rect 20864 5788 20870 5800
rect 20993 5797 21005 5800
rect 21039 5797 21051 5831
rect 20993 5791 21051 5797
rect 21085 5831 21143 5837
rect 21085 5797 21097 5831
rect 21131 5828 21143 5831
rect 21174 5828 21180 5840
rect 21131 5800 21180 5828
rect 21131 5797 21143 5800
rect 21085 5791 21143 5797
rect 21174 5788 21180 5800
rect 21232 5788 21238 5840
rect 17037 5763 17095 5769
rect 17037 5729 17049 5763
rect 17083 5729 17095 5763
rect 17037 5723 17095 5729
rect 13998 5692 14004 5704
rect 13959 5664 14004 5692
rect 13998 5652 14004 5664
rect 14056 5652 14062 5704
rect 17494 5652 17500 5704
rect 17552 5692 17558 5704
rect 17957 5695 18015 5701
rect 17957 5692 17969 5695
rect 17552 5664 17969 5692
rect 17552 5652 17558 5664
rect 17957 5661 17969 5664
rect 18003 5692 18015 5695
rect 19429 5695 19487 5701
rect 19429 5692 19441 5695
rect 18003 5664 19441 5692
rect 18003 5661 18015 5664
rect 17957 5655 18015 5661
rect 19429 5661 19441 5664
rect 19475 5661 19487 5695
rect 21450 5692 21456 5704
rect 21411 5664 21456 5692
rect 19429 5655 19487 5661
rect 21450 5652 21456 5664
rect 21508 5652 21514 5704
rect 11701 5627 11759 5633
rect 11701 5593 11713 5627
rect 11747 5624 11759 5627
rect 11790 5624 11796 5636
rect 11747 5596 11796 5624
rect 11747 5593 11759 5596
rect 11701 5587 11759 5593
rect 11790 5584 11796 5596
rect 11848 5584 11854 5636
rect 13449 5627 13507 5633
rect 13449 5593 13461 5627
rect 13495 5624 13507 5627
rect 13538 5624 13544 5636
rect 13495 5596 13544 5624
rect 13495 5593 13507 5596
rect 13449 5587 13507 5593
rect 13538 5584 13544 5596
rect 13596 5624 13602 5636
rect 14274 5624 14280 5636
rect 13596 5596 14280 5624
rect 13596 5584 13602 5596
rect 14274 5584 14280 5596
rect 14332 5584 14338 5636
rect 18506 5624 18512 5636
rect 18467 5596 18512 5624
rect 18506 5584 18512 5596
rect 18564 5584 18570 5636
rect 11974 5556 11980 5568
rect 11563 5528 11980 5556
rect 11563 5525 11575 5528
rect 11517 5519 11575 5525
rect 11974 5516 11980 5528
rect 12032 5556 12038 5568
rect 12526 5556 12532 5568
rect 12032 5528 12532 5556
rect 12032 5516 12038 5528
rect 12526 5516 12532 5528
rect 12584 5516 12590 5568
rect 14366 5556 14372 5568
rect 14327 5528 14372 5556
rect 14366 5516 14372 5528
rect 14424 5516 14430 5568
rect 20346 5516 20352 5568
rect 20404 5556 20410 5568
rect 20533 5559 20591 5565
rect 20533 5556 20545 5559
rect 20404 5528 20545 5556
rect 20404 5516 20410 5528
rect 20533 5525 20545 5528
rect 20579 5525 20591 5559
rect 20533 5519 20591 5525
rect 1104 5466 22816 5488
rect 1104 5414 4982 5466
rect 5034 5414 5046 5466
rect 5098 5414 5110 5466
rect 5162 5414 5174 5466
rect 5226 5414 12982 5466
rect 13034 5414 13046 5466
rect 13098 5414 13110 5466
rect 13162 5414 13174 5466
rect 13226 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 22816 5466
rect 1104 5392 22816 5414
rect 4154 5312 4160 5364
rect 4212 5352 4218 5364
rect 4522 5352 4528 5364
rect 4212 5324 4257 5352
rect 4483 5324 4528 5352
rect 4212 5312 4218 5324
rect 4522 5312 4528 5324
rect 4580 5312 4586 5364
rect 5629 5355 5687 5361
rect 5629 5321 5641 5355
rect 5675 5352 5687 5355
rect 5994 5352 6000 5364
rect 5675 5324 6000 5352
rect 5675 5321 5687 5324
rect 5629 5315 5687 5321
rect 5994 5312 6000 5324
rect 6052 5312 6058 5364
rect 6273 5355 6331 5361
rect 6273 5321 6285 5355
rect 6319 5352 6331 5355
rect 6362 5352 6368 5364
rect 6319 5324 6368 5352
rect 6319 5321 6331 5324
rect 6273 5315 6331 5321
rect 6362 5312 6368 5324
rect 6420 5312 6426 5364
rect 6546 5312 6552 5364
rect 6604 5352 6610 5364
rect 7374 5352 7380 5364
rect 6604 5324 7380 5352
rect 6604 5312 6610 5324
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 9769 5355 9827 5361
rect 9769 5321 9781 5355
rect 9815 5352 9827 5355
rect 10042 5352 10048 5364
rect 9815 5324 10048 5352
rect 9815 5321 9827 5324
rect 9769 5315 9827 5321
rect 10042 5312 10048 5324
rect 10100 5312 10106 5364
rect 11333 5355 11391 5361
rect 11333 5321 11345 5355
rect 11379 5352 11391 5355
rect 11790 5352 11796 5364
rect 11379 5324 11796 5352
rect 11379 5321 11391 5324
rect 11333 5315 11391 5321
rect 11790 5312 11796 5324
rect 11848 5352 11854 5364
rect 12250 5352 12256 5364
rect 11848 5324 12256 5352
rect 11848 5312 11854 5324
rect 12250 5312 12256 5324
rect 12308 5312 12314 5364
rect 12526 5352 12532 5364
rect 12487 5324 12532 5352
rect 12526 5312 12532 5324
rect 12584 5312 12590 5364
rect 15378 5312 15384 5364
rect 15436 5352 15442 5364
rect 15473 5355 15531 5361
rect 15473 5352 15485 5355
rect 15436 5324 15485 5352
rect 15436 5312 15442 5324
rect 15473 5321 15485 5324
rect 15519 5321 15531 5355
rect 17494 5352 17500 5364
rect 17455 5324 17500 5352
rect 15473 5315 15531 5321
rect 17494 5312 17500 5324
rect 17552 5312 17558 5364
rect 18046 5312 18052 5364
rect 18104 5352 18110 5364
rect 19061 5355 19119 5361
rect 19061 5352 19073 5355
rect 18104 5324 19073 5352
rect 18104 5312 18110 5324
rect 19061 5321 19073 5324
rect 19107 5321 19119 5355
rect 19061 5315 19119 5321
rect 20441 5355 20499 5361
rect 20441 5321 20453 5355
rect 20487 5352 20499 5355
rect 20806 5352 20812 5364
rect 20487 5324 20812 5352
rect 20487 5321 20499 5324
rect 20441 5315 20499 5321
rect 20806 5312 20812 5324
rect 20864 5312 20870 5364
rect 21266 5312 21272 5364
rect 21324 5352 21330 5364
rect 21545 5355 21603 5361
rect 21545 5352 21557 5355
rect 21324 5324 21557 5352
rect 21324 5312 21330 5324
rect 21545 5321 21557 5324
rect 21591 5321 21603 5355
rect 21545 5315 21603 5321
rect 106 5244 112 5296
rect 164 5284 170 5296
rect 1535 5287 1593 5293
rect 1535 5284 1547 5287
rect 164 5256 1547 5284
rect 164 5244 170 5256
rect 1535 5253 1547 5256
rect 1581 5253 1593 5287
rect 1535 5247 1593 5253
rect 5859 5287 5917 5293
rect 5859 5253 5871 5287
rect 5905 5284 5917 5287
rect 11238 5284 11244 5296
rect 5905 5256 11244 5284
rect 5905 5253 5917 5256
rect 5859 5247 5917 5253
rect 11238 5244 11244 5256
rect 11296 5244 11302 5296
rect 14274 5244 14280 5296
rect 14332 5284 14338 5296
rect 14369 5287 14427 5293
rect 14369 5284 14381 5287
rect 14332 5256 14381 5284
rect 14332 5244 14338 5256
rect 14369 5253 14381 5256
rect 14415 5284 14427 5287
rect 21358 5284 21364 5296
rect 14415 5256 21364 5284
rect 14415 5253 14427 5256
rect 14369 5247 14427 5253
rect 21358 5244 21364 5256
rect 21416 5244 21422 5296
rect 2961 5219 3019 5225
rect 2961 5185 2973 5219
rect 3007 5216 3019 5219
rect 4062 5216 4068 5228
rect 3007 5188 4068 5216
rect 3007 5185 3019 5188
rect 2961 5179 3019 5185
rect 1464 5151 1522 5157
rect 1464 5117 1476 5151
rect 1510 5148 1522 5151
rect 1946 5148 1952 5160
rect 1510 5120 1952 5148
rect 1510 5117 1522 5120
rect 1464 5111 1522 5117
rect 1946 5108 1952 5120
rect 2004 5108 2010 5160
rect 3344 5157 3372 5188
rect 4062 5176 4068 5188
rect 4120 5176 4126 5228
rect 5626 5176 5632 5228
rect 5684 5216 5690 5228
rect 6917 5219 6975 5225
rect 6917 5216 6929 5219
rect 5684 5188 6929 5216
rect 5684 5176 5690 5188
rect 6917 5185 6929 5188
rect 6963 5216 6975 5219
rect 7190 5216 7196 5228
rect 6963 5188 7196 5216
rect 6963 5185 6975 5188
rect 6917 5179 6975 5185
rect 7190 5176 7196 5188
rect 7248 5176 7254 5228
rect 7374 5216 7380 5228
rect 7335 5188 7380 5216
rect 7374 5176 7380 5188
rect 7432 5176 7438 5228
rect 10962 5216 10968 5228
rect 10923 5188 10968 5216
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 12253 5219 12311 5225
rect 12253 5185 12265 5219
rect 12299 5216 12311 5219
rect 13354 5216 13360 5228
rect 12299 5188 13360 5216
rect 12299 5185 12311 5188
rect 12253 5179 12311 5185
rect 3329 5151 3387 5157
rect 3329 5117 3341 5151
rect 3375 5117 3387 5151
rect 3329 5111 3387 5117
rect 3513 5151 3571 5157
rect 3513 5117 3525 5151
rect 3559 5148 3571 5151
rect 4522 5148 4528 5160
rect 3559 5120 4528 5148
rect 3559 5117 3571 5120
rect 3513 5111 3571 5117
rect 2593 5083 2651 5089
rect 2593 5049 2605 5083
rect 2639 5080 2651 5083
rect 3418 5080 3424 5092
rect 2639 5052 3424 5080
rect 2639 5049 2651 5052
rect 2593 5043 2651 5049
rect 3418 5040 3424 5052
rect 3476 5080 3482 5092
rect 3528 5080 3556 5111
rect 4522 5108 4528 5120
rect 4580 5108 4586 5160
rect 4760 5151 4818 5157
rect 4760 5117 4772 5151
rect 4806 5148 4818 5151
rect 5169 5151 5227 5157
rect 5169 5148 5181 5151
rect 4806 5120 5181 5148
rect 4806 5117 4818 5120
rect 4760 5111 4818 5117
rect 5169 5117 5181 5120
rect 5215 5148 5227 5151
rect 5534 5148 5540 5160
rect 5215 5120 5540 5148
rect 5215 5117 5227 5120
rect 5169 5111 5227 5117
rect 5534 5108 5540 5120
rect 5592 5108 5598 5160
rect 5810 5157 5816 5160
rect 5788 5151 5816 5157
rect 5788 5117 5800 5151
rect 5868 5148 5874 5160
rect 6362 5148 6368 5160
rect 5868 5120 6368 5148
rect 5788 5111 5816 5117
rect 5810 5108 5816 5111
rect 5868 5108 5874 5120
rect 6362 5108 6368 5120
rect 6420 5108 6426 5160
rect 7742 5108 7748 5160
rect 7800 5148 7806 5160
rect 8386 5148 8392 5160
rect 7800 5120 8392 5148
rect 7800 5108 7806 5120
rect 8386 5108 8392 5120
rect 8444 5108 8450 5160
rect 12728 5157 12756 5188
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 13630 5176 13636 5228
rect 13688 5216 13694 5228
rect 14461 5219 14519 5225
rect 14461 5216 14473 5219
rect 13688 5188 14473 5216
rect 13688 5176 13694 5188
rect 14461 5185 14473 5188
rect 14507 5185 14519 5219
rect 14461 5179 14519 5185
rect 16761 5219 16819 5225
rect 16761 5185 16773 5219
rect 16807 5216 16819 5219
rect 16850 5216 16856 5228
rect 16807 5188 16856 5216
rect 16807 5185 16819 5188
rect 16761 5179 16819 5185
rect 16850 5176 16856 5188
rect 16908 5176 16914 5228
rect 17586 5176 17592 5228
rect 17644 5216 17650 5228
rect 17865 5219 17923 5225
rect 17865 5216 17877 5219
rect 17644 5188 17877 5216
rect 17644 5176 17650 5188
rect 17865 5185 17877 5188
rect 17911 5216 17923 5219
rect 21269 5219 21327 5225
rect 17911 5188 18276 5216
rect 17911 5185 17923 5188
rect 17865 5179 17923 5185
rect 8849 5151 8907 5157
rect 8849 5148 8861 5151
rect 8496 5120 8861 5148
rect 3476 5052 3556 5080
rect 4847 5083 4905 5089
rect 3476 5040 3482 5052
rect 4847 5049 4859 5083
rect 4893 5080 4905 5083
rect 6730 5080 6736 5092
rect 4893 5052 6736 5080
rect 4893 5049 4905 5052
rect 4847 5043 4905 5049
rect 6730 5040 6736 5052
rect 6788 5040 6794 5092
rect 7006 5040 7012 5092
rect 7064 5080 7070 5092
rect 7064 5052 7109 5080
rect 7064 5040 7070 5052
rect 1946 5012 1952 5024
rect 1907 4984 1952 5012
rect 1946 4972 1952 4984
rect 2004 4972 2010 5024
rect 2958 4972 2964 5024
rect 3016 5012 3022 5024
rect 3145 5015 3203 5021
rect 3145 5012 3157 5015
rect 3016 4984 3157 5012
rect 3016 4972 3022 4984
rect 3145 4981 3157 4984
rect 3191 4981 3203 5015
rect 3145 4975 3203 4981
rect 6641 5015 6699 5021
rect 6641 4981 6653 5015
rect 6687 5012 6699 5015
rect 7024 5012 7052 5040
rect 8496 5024 8524 5120
rect 8849 5117 8861 5120
rect 8895 5117 8907 5151
rect 8849 5111 8907 5117
rect 12713 5151 12771 5157
rect 12713 5117 12725 5151
rect 12759 5117 12771 5151
rect 12894 5148 12900 5160
rect 12855 5120 12900 5148
rect 12713 5111 12771 5117
rect 12894 5108 12900 5120
rect 12952 5108 12958 5160
rect 13173 5151 13231 5157
rect 13173 5148 13185 5151
rect 13004 5120 13185 5148
rect 9125 5083 9183 5089
rect 9125 5049 9137 5083
rect 9171 5080 9183 5083
rect 9582 5080 9588 5092
rect 9171 5052 9588 5080
rect 9171 5049 9183 5052
rect 9125 5043 9183 5049
rect 9582 5040 9588 5052
rect 9640 5040 9646 5092
rect 10318 5080 10324 5092
rect 10279 5052 10324 5080
rect 10318 5040 10324 5052
rect 10376 5040 10382 5092
rect 10413 5083 10471 5089
rect 10413 5049 10425 5083
rect 10459 5049 10471 5083
rect 10413 5043 10471 5049
rect 6687 4984 7052 5012
rect 7929 5015 7987 5021
rect 6687 4981 6699 4984
rect 6641 4975 6699 4981
rect 7929 4981 7941 5015
rect 7975 5012 7987 5015
rect 8297 5015 8355 5021
rect 8297 5012 8309 5015
rect 7975 4984 8309 5012
rect 7975 4981 7987 4984
rect 7929 4975 7987 4981
rect 8297 4981 8309 4984
rect 8343 5012 8355 5015
rect 8478 5012 8484 5024
rect 8343 4984 8484 5012
rect 8343 4981 8355 4984
rect 8297 4975 8355 4981
rect 8478 4972 8484 4984
rect 8536 4972 8542 5024
rect 10137 5015 10195 5021
rect 10137 4981 10149 5015
rect 10183 5012 10195 5015
rect 10428 5012 10456 5043
rect 10594 5012 10600 5024
rect 10183 4984 10600 5012
rect 10183 4981 10195 4984
rect 10137 4975 10195 4981
rect 10594 4972 10600 4984
rect 10652 4972 10658 5024
rect 11606 5012 11612 5024
rect 11567 4984 11612 5012
rect 11606 4972 11612 4984
rect 11664 4972 11670 5024
rect 12434 4972 12440 5024
rect 12492 5012 12498 5024
rect 13004 5012 13032 5120
rect 13173 5117 13185 5120
rect 13219 5148 13231 5151
rect 14550 5148 14556 5160
rect 13219 5120 14556 5148
rect 13219 5117 13231 5120
rect 13173 5111 13231 5117
rect 14550 5108 14556 5120
rect 14608 5108 14614 5160
rect 16025 5151 16083 5157
rect 16025 5148 16037 5151
rect 15856 5120 16037 5148
rect 12492 4984 13032 5012
rect 14001 5015 14059 5021
rect 12492 4972 12498 4984
rect 14001 4981 14013 5015
rect 14047 5012 14059 5015
rect 14090 5012 14096 5024
rect 14047 4984 14096 5012
rect 14047 4981 14059 4984
rect 14001 4975 14059 4981
rect 14090 4972 14096 4984
rect 14148 4972 14154 5024
rect 15654 4972 15660 5024
rect 15712 5012 15718 5024
rect 15856 5021 15884 5120
rect 16025 5117 16037 5120
rect 16071 5117 16083 5151
rect 16025 5111 16083 5117
rect 16114 5108 16120 5160
rect 16172 5148 16178 5160
rect 16301 5151 16359 5157
rect 16172 5120 16217 5148
rect 16172 5108 16178 5120
rect 16301 5117 16313 5151
rect 16347 5148 16359 5151
rect 18046 5148 18052 5160
rect 16347 5120 17172 5148
rect 18007 5120 18052 5148
rect 16347 5117 16359 5120
rect 16301 5111 16359 5117
rect 17144 5021 17172 5120
rect 18046 5108 18052 5120
rect 18104 5108 18110 5160
rect 18248 5148 18276 5188
rect 21269 5185 21281 5219
rect 21315 5216 21327 5219
rect 21450 5216 21456 5228
rect 21315 5188 21456 5216
rect 21315 5185 21327 5188
rect 21269 5179 21327 5185
rect 21450 5176 21456 5188
rect 21508 5176 21514 5228
rect 18509 5151 18567 5157
rect 18509 5148 18521 5151
rect 18248 5120 18521 5148
rect 18509 5117 18521 5120
rect 18555 5117 18567 5151
rect 18509 5111 18567 5117
rect 20346 5040 20352 5092
rect 20404 5080 20410 5092
rect 20625 5083 20683 5089
rect 20625 5080 20637 5083
rect 20404 5052 20637 5080
rect 20404 5040 20410 5052
rect 20625 5049 20637 5052
rect 20671 5049 20683 5083
rect 20625 5043 20683 5049
rect 20714 5040 20720 5092
rect 20772 5080 20778 5092
rect 20772 5052 20817 5080
rect 20772 5040 20778 5052
rect 15841 5015 15899 5021
rect 15841 5012 15853 5015
rect 15712 4984 15853 5012
rect 15712 4972 15718 4984
rect 15841 4981 15853 4984
rect 15887 4981 15899 5015
rect 15841 4975 15899 4981
rect 17129 5015 17187 5021
rect 17129 4981 17141 5015
rect 17175 5012 17187 5015
rect 17310 5012 17316 5024
rect 17175 4984 17316 5012
rect 17175 4981 17187 4984
rect 17129 4975 17187 4981
rect 17310 4972 17316 4984
rect 17368 4972 17374 5024
rect 18138 5012 18144 5024
rect 18099 4984 18144 5012
rect 18138 4972 18144 4984
rect 18196 4972 18202 5024
rect 1104 4922 22816 4944
rect 1104 4870 8982 4922
rect 9034 4870 9046 4922
rect 9098 4870 9110 4922
rect 9162 4870 9174 4922
rect 9226 4870 16982 4922
rect 17034 4870 17046 4922
rect 17098 4870 17110 4922
rect 17162 4870 17174 4922
rect 17226 4870 22816 4922
rect 1104 4848 22816 4870
rect 3099 4811 3157 4817
rect 3099 4777 3111 4811
rect 3145 4808 3157 4811
rect 5626 4808 5632 4820
rect 3145 4780 5632 4808
rect 3145 4777 3157 4780
rect 3099 4771 3157 4777
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 5902 4808 5908 4820
rect 5863 4780 5908 4808
rect 5902 4768 5908 4780
rect 5960 4768 5966 4820
rect 6730 4808 6736 4820
rect 6691 4780 6736 4808
rect 6730 4768 6736 4780
rect 6788 4768 6794 4820
rect 7834 4768 7840 4820
rect 7892 4808 7898 4820
rect 7929 4811 7987 4817
rect 7929 4808 7941 4811
rect 7892 4780 7941 4808
rect 7892 4768 7898 4780
rect 7929 4777 7941 4780
rect 7975 4777 7987 4811
rect 8386 4808 8392 4820
rect 8347 4780 8392 4808
rect 7929 4771 7987 4777
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 8711 4811 8769 4817
rect 8711 4777 8723 4811
rect 8757 4808 8769 4811
rect 10318 4808 10324 4820
rect 8757 4780 10324 4808
rect 8757 4777 8769 4780
rect 8711 4771 8769 4777
rect 10318 4768 10324 4780
rect 10376 4808 10382 4820
rect 10873 4811 10931 4817
rect 10873 4808 10885 4811
rect 10376 4780 10885 4808
rect 10376 4768 10382 4780
rect 10873 4777 10885 4780
rect 10919 4777 10931 4811
rect 11238 4808 11244 4820
rect 11199 4780 11244 4808
rect 10873 4771 10931 4777
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 12894 4808 12900 4820
rect 12855 4780 12900 4808
rect 12894 4768 12900 4780
rect 12952 4808 12958 4820
rect 14550 4808 14556 4820
rect 12952 4780 13032 4808
rect 14511 4780 14556 4808
rect 12952 4768 12958 4780
rect 4798 4700 4804 4752
rect 4856 4740 4862 4752
rect 5077 4743 5135 4749
rect 5077 4740 5089 4743
rect 4856 4712 5089 4740
rect 4856 4700 4862 4712
rect 5077 4709 5089 4712
rect 5123 4709 5135 4743
rect 5077 4703 5135 4709
rect 7006 4700 7012 4752
rect 7064 4740 7070 4752
rect 7101 4743 7159 4749
rect 7101 4740 7113 4743
rect 7064 4712 7113 4740
rect 7064 4700 7070 4712
rect 7101 4709 7113 4712
rect 7147 4740 7159 4743
rect 7742 4740 7748 4752
rect 7147 4712 7748 4740
rect 7147 4709 7159 4712
rect 7101 4703 7159 4709
rect 7742 4700 7748 4712
rect 7800 4700 7806 4752
rect 9398 4740 9404 4752
rect 9359 4712 9404 4740
rect 9398 4700 9404 4712
rect 9456 4700 9462 4752
rect 9766 4700 9772 4752
rect 9824 4740 9830 4752
rect 9998 4743 10056 4749
rect 9998 4740 10010 4743
rect 9824 4712 10010 4740
rect 9824 4700 9830 4712
rect 9998 4709 10010 4712
rect 10044 4709 10056 4743
rect 11609 4743 11667 4749
rect 11609 4740 11621 4743
rect 9998 4703 10056 4709
rect 10612 4712 11621 4740
rect 10612 4684 10640 4712
rect 11609 4709 11621 4712
rect 11655 4740 11667 4743
rect 11698 4740 11704 4752
rect 11655 4712 11704 4740
rect 11655 4709 11667 4712
rect 11609 4703 11667 4709
rect 11698 4700 11704 4712
rect 11756 4700 11762 4752
rect 13004 4749 13032 4780
rect 14550 4768 14556 4780
rect 14608 4768 14614 4820
rect 15749 4811 15807 4817
rect 15749 4777 15761 4811
rect 15795 4808 15807 4811
rect 16022 4808 16028 4820
rect 15795 4780 16028 4808
rect 15795 4777 15807 4780
rect 15749 4771 15807 4777
rect 16022 4768 16028 4780
rect 16080 4768 16086 4820
rect 16666 4808 16672 4820
rect 16627 4780 16672 4808
rect 16666 4768 16672 4780
rect 16724 4768 16730 4820
rect 18046 4808 18052 4820
rect 18007 4780 18052 4808
rect 18046 4768 18052 4780
rect 18104 4768 18110 4820
rect 18598 4808 18604 4820
rect 18559 4780 18604 4808
rect 18598 4768 18604 4780
rect 18656 4768 18662 4820
rect 19153 4811 19211 4817
rect 19153 4777 19165 4811
rect 19199 4808 19211 4811
rect 20533 4811 20591 4817
rect 20533 4808 20545 4811
rect 19199 4780 20545 4808
rect 19199 4777 19211 4780
rect 19153 4771 19211 4777
rect 20533 4777 20545 4780
rect 20579 4808 20591 4811
rect 20714 4808 20720 4820
rect 20579 4780 20720 4808
rect 20579 4777 20591 4780
rect 20533 4771 20591 4777
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 12989 4743 13047 4749
rect 12989 4709 13001 4743
rect 13035 4740 13047 4743
rect 14366 4740 14372 4752
rect 13035 4712 14372 4740
rect 13035 4709 13047 4712
rect 12989 4703 13047 4709
rect 14366 4700 14372 4712
rect 14424 4700 14430 4752
rect 2866 4672 2872 4684
rect 2827 4644 2872 4672
rect 2866 4632 2872 4644
rect 2924 4632 2930 4684
rect 8386 4672 8392 4684
rect 7944 4644 8392 4672
rect 4985 4607 5043 4613
rect 4985 4573 4997 4607
rect 5031 4573 5043 4607
rect 5626 4604 5632 4616
rect 5587 4576 5632 4604
rect 4985 4567 5043 4573
rect 5000 4536 5028 4567
rect 5626 4564 5632 4576
rect 5684 4564 5690 4616
rect 6546 4604 6552 4616
rect 5736 4576 6552 4604
rect 5350 4536 5356 4548
rect 5000 4508 5356 4536
rect 5350 4496 5356 4508
rect 5408 4536 5414 4548
rect 5736 4536 5764 4576
rect 6546 4564 6552 4576
rect 6604 4564 6610 4616
rect 6730 4564 6736 4616
rect 6788 4604 6794 4616
rect 7009 4607 7067 4613
rect 7009 4604 7021 4607
rect 6788 4576 7021 4604
rect 6788 4564 6794 4576
rect 7009 4573 7021 4576
rect 7055 4573 7067 4607
rect 7282 4604 7288 4616
rect 7243 4576 7288 4604
rect 7009 4567 7067 4573
rect 7282 4564 7288 4576
rect 7340 4564 7346 4616
rect 5408 4508 5764 4536
rect 5408 4496 5414 4508
rect 6362 4496 6368 4548
rect 6420 4536 6426 4548
rect 7300 4536 7328 4564
rect 6420 4508 7328 4536
rect 6420 4496 6426 4508
rect 3602 4468 3608 4480
rect 3563 4440 3608 4468
rect 3602 4428 3608 4440
rect 3660 4428 3666 4480
rect 5534 4428 5540 4480
rect 5592 4468 5598 4480
rect 7944 4468 7972 4644
rect 8386 4632 8392 4644
rect 8444 4672 8450 4684
rect 8608 4675 8666 4681
rect 8608 4672 8620 4675
rect 8444 4644 8620 4672
rect 8444 4632 8450 4644
rect 8608 4641 8620 4644
rect 8654 4641 8666 4675
rect 8608 4635 8666 4641
rect 9582 4632 9588 4684
rect 9640 4672 9646 4684
rect 9677 4675 9735 4681
rect 9677 4672 9689 4675
rect 9640 4644 9689 4672
rect 9640 4632 9646 4644
rect 9677 4641 9689 4644
rect 9723 4641 9735 4675
rect 10594 4672 10600 4684
rect 10555 4644 10600 4672
rect 9677 4635 9735 4641
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 13538 4672 13544 4684
rect 13499 4644 13544 4672
rect 13538 4632 13544 4644
rect 13596 4632 13602 4684
rect 15378 4632 15384 4684
rect 15436 4672 15442 4684
rect 16209 4675 16267 4681
rect 16209 4672 16221 4675
rect 15436 4644 16221 4672
rect 15436 4632 15442 4644
rect 16209 4641 16221 4644
rect 16255 4641 16267 4675
rect 16482 4672 16488 4684
rect 16443 4644 16488 4672
rect 16209 4635 16267 4641
rect 16482 4632 16488 4644
rect 16540 4632 16546 4684
rect 20622 4632 20628 4684
rect 20680 4672 20686 4684
rect 20936 4675 20994 4681
rect 20936 4672 20948 4675
rect 20680 4644 20948 4672
rect 20680 4632 20686 4644
rect 20936 4641 20948 4644
rect 20982 4641 20994 4675
rect 20936 4635 20994 4641
rect 11238 4564 11244 4616
rect 11296 4604 11302 4616
rect 11517 4607 11575 4613
rect 11517 4604 11529 4607
rect 11296 4576 11529 4604
rect 11296 4564 11302 4576
rect 11517 4573 11529 4576
rect 11563 4573 11575 4607
rect 11517 4567 11575 4573
rect 11793 4607 11851 4613
rect 11793 4573 11805 4607
rect 11839 4573 11851 4607
rect 11793 4567 11851 4573
rect 10502 4496 10508 4548
rect 10560 4536 10566 4548
rect 11808 4536 11836 4567
rect 17402 4564 17408 4616
rect 17460 4604 17466 4616
rect 18233 4607 18291 4613
rect 18233 4604 18245 4607
rect 17460 4576 18245 4604
rect 17460 4564 17466 4576
rect 18233 4573 18245 4576
rect 18279 4573 18291 4607
rect 18233 4567 18291 4573
rect 10560 4508 11836 4536
rect 16301 4539 16359 4545
rect 10560 4496 10566 4508
rect 16301 4505 16313 4539
rect 16347 4505 16359 4539
rect 20162 4536 20168 4548
rect 20075 4508 20168 4536
rect 16301 4499 16359 4505
rect 12434 4468 12440 4480
rect 5592 4440 7972 4468
rect 12395 4440 12440 4468
rect 5592 4428 5598 4440
rect 12434 4428 12440 4440
rect 12492 4428 12498 4480
rect 13998 4468 14004 4480
rect 13959 4440 14004 4468
rect 13998 4428 14004 4440
rect 14056 4428 14062 4480
rect 16114 4468 16120 4480
rect 16075 4440 16120 4468
rect 16114 4428 16120 4440
rect 16172 4468 16178 4480
rect 16316 4468 16344 4499
rect 20162 4496 20168 4508
rect 20220 4536 20226 4548
rect 21039 4539 21097 4545
rect 21039 4536 21051 4539
rect 20220 4508 21051 4536
rect 20220 4496 20226 4508
rect 21039 4505 21051 4508
rect 21085 4505 21097 4539
rect 21039 4499 21097 4505
rect 16172 4440 16344 4468
rect 16172 4428 16178 4440
rect 1104 4378 22816 4400
rect 1104 4326 4982 4378
rect 5034 4326 5046 4378
rect 5098 4326 5110 4378
rect 5162 4326 5174 4378
rect 5226 4326 12982 4378
rect 13034 4326 13046 4378
rect 13098 4326 13110 4378
rect 13162 4326 13174 4378
rect 13226 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 22816 4378
rect 1104 4304 22816 4326
rect 4525 4267 4583 4273
rect 4525 4233 4537 4267
rect 4571 4264 4583 4267
rect 4798 4264 4804 4276
rect 4571 4236 4804 4264
rect 4571 4233 4583 4236
rect 4525 4227 4583 4233
rect 4798 4224 4804 4236
rect 4856 4264 4862 4276
rect 4893 4267 4951 4273
rect 4893 4264 4905 4267
rect 4856 4236 4905 4264
rect 4856 4224 4862 4236
rect 4893 4233 4905 4236
rect 4939 4233 4951 4267
rect 5350 4264 5356 4276
rect 5311 4236 5356 4264
rect 4893 4227 4951 4233
rect 5350 4224 5356 4236
rect 5408 4224 5414 4276
rect 6273 4267 6331 4273
rect 6273 4233 6285 4267
rect 6319 4264 6331 4267
rect 7742 4264 7748 4276
rect 6319 4236 7748 4264
rect 6319 4233 6331 4236
rect 6273 4227 6331 4233
rect 7742 4224 7748 4236
rect 7800 4224 7806 4276
rect 8386 4264 8392 4276
rect 8347 4236 8392 4264
rect 8386 4224 8392 4236
rect 8444 4264 8450 4276
rect 9306 4264 9312 4276
rect 8444 4236 9312 4264
rect 8444 4224 8450 4236
rect 9306 4224 9312 4236
rect 9364 4224 9370 4276
rect 9582 4224 9588 4276
rect 9640 4264 9646 4276
rect 10045 4267 10103 4273
rect 10045 4264 10057 4267
rect 9640 4236 10057 4264
rect 9640 4224 9646 4236
rect 10045 4233 10057 4236
rect 10091 4233 10103 4267
rect 11698 4264 11704 4276
rect 11659 4236 11704 4264
rect 10045 4227 10103 4233
rect 11698 4224 11704 4236
rect 11756 4224 11762 4276
rect 18782 4264 18788 4276
rect 15304 4236 18788 4264
rect 2866 4156 2872 4208
rect 2924 4196 2930 4208
rect 3145 4199 3203 4205
rect 3145 4196 3157 4199
rect 2924 4168 3157 4196
rect 2924 4156 2930 4168
rect 3145 4165 3157 4168
rect 3191 4196 3203 4199
rect 5810 4196 5816 4208
rect 3191 4168 5816 4196
rect 3191 4165 3203 4168
rect 3145 4159 3203 4165
rect 5810 4156 5816 4168
rect 5868 4156 5874 4208
rect 8113 4199 8171 4205
rect 8113 4165 8125 4199
rect 8159 4196 8171 4199
rect 8294 4196 8300 4208
rect 8159 4168 8300 4196
rect 8159 4165 8171 4168
rect 8113 4159 8171 4165
rect 8294 4156 8300 4168
rect 8352 4156 8358 4208
rect 9674 4196 9680 4208
rect 9646 4156 9680 4196
rect 9732 4156 9738 4208
rect 11974 4156 11980 4208
rect 12032 4196 12038 4208
rect 12621 4199 12679 4205
rect 12032 4168 12296 4196
rect 12032 4156 12038 4168
rect 3418 4128 3424 4140
rect 2608 4100 3424 4128
rect 2608 4069 2636 4100
rect 3418 4088 3424 4100
rect 3476 4088 3482 4140
rect 9490 4128 9496 4140
rect 6748 4100 7189 4128
rect 2317 4063 2375 4069
rect 2317 4029 2329 4063
rect 2363 4029 2375 4063
rect 2317 4023 2375 4029
rect 2593 4063 2651 4069
rect 2593 4029 2605 4063
rect 2639 4029 2651 4063
rect 2593 4023 2651 4029
rect 2777 4063 2835 4069
rect 2777 4029 2789 4063
rect 2823 4060 2835 4063
rect 3602 4060 3608 4072
rect 2823 4032 3608 4060
rect 2823 4029 2835 4032
rect 2777 4023 2835 4029
rect 1949 3995 2007 4001
rect 1949 3961 1961 3995
rect 1995 3992 2007 3995
rect 2332 3992 2360 4023
rect 3602 4020 3608 4032
rect 3660 4020 3666 4072
rect 5537 4063 5595 4069
rect 5537 4029 5549 4063
rect 5583 4060 5595 4063
rect 5626 4060 5632 4072
rect 5583 4032 5632 4060
rect 5583 4029 5595 4032
rect 5537 4023 5595 4029
rect 5626 4020 5632 4032
rect 5684 4020 5690 4072
rect 3694 3992 3700 4004
rect 1995 3964 3700 3992
rect 1995 3961 2007 3964
rect 1949 3955 2007 3961
rect 3694 3952 3700 3964
rect 3752 3952 3758 4004
rect 3926 3995 3984 4001
rect 3926 3961 3938 3995
rect 3972 3961 3984 3995
rect 3926 3955 3984 3961
rect 5767 3995 5825 4001
rect 5767 3961 5779 3995
rect 5813 3992 5825 3995
rect 6638 3992 6644 4004
rect 5813 3964 6644 3992
rect 5813 3961 5825 3964
rect 5767 3955 5825 3961
rect 3142 3884 3148 3936
rect 3200 3924 3206 3936
rect 3421 3927 3479 3933
rect 3421 3924 3433 3927
rect 3200 3896 3433 3924
rect 3200 3884 3206 3896
rect 3421 3893 3433 3896
rect 3467 3924 3479 3927
rect 3941 3924 3969 3955
rect 6638 3952 6644 3964
rect 6696 3952 6702 4004
rect 3467 3896 3969 3924
rect 3467 3893 3479 3896
rect 3421 3887 3479 3893
rect 5534 3884 5540 3936
rect 5592 3924 5598 3936
rect 6549 3927 6607 3933
rect 6549 3924 6561 3927
rect 5592 3896 6561 3924
rect 5592 3884 5598 3896
rect 6549 3893 6561 3896
rect 6595 3924 6607 3927
rect 6748 3924 6776 4100
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 6595 3896 6776 3924
rect 6840 3924 6868 4023
rect 7161 4001 7189 4100
rect 9140 4100 9496 4128
rect 8294 4020 8300 4072
rect 8352 4060 8358 4072
rect 9140 4069 9168 4100
rect 9490 4088 9496 4100
rect 9548 4088 9554 4140
rect 8573 4063 8631 4069
rect 8573 4060 8585 4063
rect 8352 4032 8585 4060
rect 8352 4020 8358 4032
rect 8573 4029 8585 4032
rect 8619 4029 8631 4063
rect 8573 4023 8631 4029
rect 9125 4063 9183 4069
rect 9125 4029 9137 4063
rect 9171 4029 9183 4063
rect 9125 4023 9183 4029
rect 9306 4020 9312 4072
rect 9364 4060 9370 4072
rect 9646 4060 9674 4156
rect 10594 4088 10600 4140
rect 10652 4128 10658 4140
rect 12268 4137 12296 4168
rect 12621 4165 12633 4199
rect 12667 4196 12679 4199
rect 15010 4196 15016 4208
rect 12667 4168 15016 4196
rect 12667 4165 12679 4168
rect 12621 4159 12679 4165
rect 15010 4156 15016 4168
rect 15068 4156 15074 4208
rect 10781 4131 10839 4137
rect 10781 4128 10793 4131
rect 10652 4100 10793 4128
rect 10652 4088 10658 4100
rect 10781 4097 10793 4100
rect 10827 4097 10839 4131
rect 12253 4131 12311 4137
rect 12253 4128 12265 4131
rect 12163 4100 12265 4128
rect 10781 4091 10839 4097
rect 12253 4097 12265 4100
rect 12299 4128 12311 4131
rect 15304 4128 15332 4236
rect 18782 4224 18788 4236
rect 18840 4224 18846 4276
rect 20622 4224 20628 4276
rect 20680 4264 20686 4276
rect 21085 4267 21143 4273
rect 21085 4264 21097 4267
rect 20680 4236 21097 4264
rect 20680 4224 20686 4236
rect 21085 4233 21097 4236
rect 21131 4233 21143 4267
rect 21085 4227 21143 4233
rect 18230 4156 18236 4208
rect 18288 4196 18294 4208
rect 18325 4199 18383 4205
rect 18325 4196 18337 4199
rect 18288 4168 18337 4196
rect 18288 4156 18294 4168
rect 18325 4165 18337 4168
rect 18371 4196 18383 4199
rect 18598 4196 18604 4208
rect 18371 4168 18604 4196
rect 18371 4165 18383 4168
rect 18325 4159 18383 4165
rect 18598 4156 18604 4168
rect 18656 4156 18662 4208
rect 12299 4100 15332 4128
rect 16945 4131 17003 4137
rect 12299 4097 12311 4100
rect 12253 4091 12311 4097
rect 12452 4069 12480 4100
rect 16945 4097 16957 4131
rect 16991 4128 17003 4131
rect 17310 4128 17316 4140
rect 16991 4100 17316 4128
rect 16991 4097 17003 4100
rect 16945 4091 17003 4097
rect 17310 4088 17316 4100
rect 17368 4088 17374 4140
rect 20162 4128 20168 4140
rect 20123 4100 20168 4128
rect 20162 4088 20168 4100
rect 20220 4088 20226 4140
rect 20346 4088 20352 4140
rect 20404 4128 20410 4140
rect 20441 4131 20499 4137
rect 20441 4128 20453 4131
rect 20404 4100 20453 4128
rect 20404 4088 20410 4100
rect 20441 4097 20453 4100
rect 20487 4097 20499 4131
rect 20441 4091 20499 4097
rect 12437 4063 12495 4069
rect 12437 4060 12449 4063
rect 9364 4032 9674 4060
rect 12415 4032 12449 4060
rect 9364 4020 9370 4032
rect 12437 4029 12449 4032
rect 12483 4029 12495 4063
rect 13541 4063 13599 4069
rect 13541 4060 13553 4063
rect 12437 4023 12495 4029
rect 13004 4032 13553 4060
rect 7146 3995 7204 4001
rect 7146 3961 7158 3995
rect 7192 3992 7204 3995
rect 7466 3992 7472 4004
rect 7192 3964 7472 3992
rect 7192 3961 7204 3964
rect 7146 3955 7204 3961
rect 7466 3952 7472 3964
rect 7524 3992 7530 4004
rect 9398 3992 9404 4004
rect 7524 3964 9404 3992
rect 7524 3952 7530 3964
rect 9398 3952 9404 3964
rect 9456 3992 9462 4004
rect 9677 3995 9735 4001
rect 9677 3992 9689 3995
rect 9456 3964 9689 3992
rect 9456 3952 9462 3964
rect 9677 3961 9689 3964
rect 9723 3992 9735 3995
rect 9766 3992 9772 4004
rect 9723 3964 9772 3992
rect 9723 3961 9735 3964
rect 9677 3955 9735 3961
rect 9766 3952 9772 3964
rect 9824 3952 9830 4004
rect 10597 3995 10655 4001
rect 10597 3961 10609 3995
rect 10643 3992 10655 3995
rect 10870 3992 10876 4004
rect 10643 3964 10876 3992
rect 10643 3961 10655 3964
rect 10597 3955 10655 3961
rect 10870 3952 10876 3964
rect 10928 3952 10934 4004
rect 11425 3995 11483 4001
rect 11425 3961 11437 3995
rect 11471 3992 11483 3995
rect 11698 3992 11704 4004
rect 11471 3964 11704 3992
rect 11471 3961 11483 3964
rect 11425 3955 11483 3961
rect 11698 3952 11704 3964
rect 11756 3952 11762 4004
rect 7374 3924 7380 3936
rect 6840 3896 7380 3924
rect 6595 3893 6607 3896
rect 6549 3887 6607 3893
rect 7374 3884 7380 3896
rect 7432 3924 7438 3936
rect 8665 3927 8723 3933
rect 8665 3924 8677 3927
rect 7432 3896 8677 3924
rect 7432 3884 7438 3896
rect 8665 3893 8677 3896
rect 8711 3893 8723 3927
rect 8665 3887 8723 3893
rect 11606 3884 11612 3936
rect 11664 3924 11670 3936
rect 13004 3933 13032 4032
rect 13541 4029 13553 4032
rect 13587 4060 13599 4063
rect 13630 4060 13636 4072
rect 13587 4032 13636 4060
rect 13587 4029 13599 4032
rect 13541 4023 13599 4029
rect 13630 4020 13636 4032
rect 13688 4020 13694 4072
rect 13906 4020 13912 4072
rect 13964 4060 13970 4072
rect 14001 4063 14059 4069
rect 14001 4060 14013 4063
rect 13964 4032 14013 4060
rect 13964 4020 13970 4032
rect 14001 4029 14013 4032
rect 14047 4029 14059 4063
rect 14001 4023 14059 4029
rect 14090 4020 14096 4072
rect 14148 4060 14154 4072
rect 14366 4060 14372 4072
rect 14148 4032 14372 4060
rect 14148 4020 14154 4032
rect 14366 4020 14372 4032
rect 14424 4020 14430 4072
rect 14737 4063 14795 4069
rect 14737 4060 14749 4063
rect 14476 4032 14749 4060
rect 14476 3992 14504 4032
rect 14737 4029 14749 4032
rect 14783 4029 14795 4063
rect 14737 4023 14795 4029
rect 16206 4020 16212 4072
rect 16264 4060 16270 4072
rect 16301 4063 16359 4069
rect 16301 4060 16313 4063
rect 16264 4032 16313 4060
rect 16264 4020 16270 4032
rect 16301 4029 16313 4032
rect 16347 4060 16359 4063
rect 16482 4060 16488 4072
rect 16347 4032 16488 4060
rect 16347 4029 16359 4032
rect 16301 4023 16359 4029
rect 16482 4020 16488 4032
rect 16540 4020 16546 4072
rect 17865 4063 17923 4069
rect 17865 4029 17877 4063
rect 17911 4060 17923 4063
rect 18601 4063 18659 4069
rect 18601 4060 18613 4063
rect 17911 4032 18613 4060
rect 17911 4029 17923 4032
rect 17865 4023 17923 4029
rect 18601 4029 18613 4032
rect 18647 4060 18659 4063
rect 19334 4060 19340 4072
rect 18647 4032 19340 4060
rect 18647 4029 18659 4032
rect 18601 4023 18659 4029
rect 19334 4020 19340 4032
rect 19392 4020 19398 4072
rect 13786 3964 14504 3992
rect 15013 3995 15071 4001
rect 12989 3927 13047 3933
rect 12989 3924 13001 3927
rect 11664 3896 13001 3924
rect 11664 3884 11670 3896
rect 12989 3893 13001 3896
rect 13035 3893 13047 3927
rect 13446 3924 13452 3936
rect 13407 3896 13452 3924
rect 12989 3887 13047 3893
rect 13446 3884 13452 3896
rect 13504 3924 13510 3936
rect 13786 3924 13814 3964
rect 15013 3961 15025 3995
rect 15059 3992 15071 3995
rect 17678 3992 17684 4004
rect 15059 3964 17684 3992
rect 15059 3961 15071 3964
rect 15013 3955 15071 3961
rect 17678 3952 17684 3964
rect 17736 3952 17742 4004
rect 19245 3995 19303 4001
rect 19245 3961 19257 3995
rect 19291 3992 19303 3995
rect 19889 3995 19947 4001
rect 19889 3992 19901 3995
rect 19291 3964 19901 3992
rect 19291 3961 19303 3964
rect 19245 3955 19303 3961
rect 19889 3961 19901 3964
rect 19935 3992 19947 3995
rect 20257 3995 20315 4001
rect 20257 3992 20269 3995
rect 19935 3964 20269 3992
rect 19935 3961 19947 3964
rect 19889 3955 19947 3961
rect 20257 3961 20269 3964
rect 20303 3961 20315 3995
rect 20257 3955 20315 3961
rect 15378 3924 15384 3936
rect 13504 3896 13814 3924
rect 15339 3896 15384 3924
rect 13504 3884 13510 3896
rect 15378 3884 15384 3896
rect 15436 3884 15442 3936
rect 15746 3924 15752 3936
rect 15707 3896 15752 3924
rect 15746 3884 15752 3896
rect 15804 3924 15810 3936
rect 16025 3927 16083 3933
rect 16025 3924 16037 3927
rect 15804 3896 16037 3924
rect 15804 3884 15810 3896
rect 16025 3893 16037 3896
rect 16071 3893 16083 3927
rect 16025 3887 16083 3893
rect 16758 3884 16764 3936
rect 16816 3924 16822 3936
rect 17402 3924 17408 3936
rect 16816 3896 17408 3924
rect 16816 3884 16822 3896
rect 17402 3884 17408 3896
rect 17460 3884 17466 3936
rect 1104 3834 22816 3856
rect 1104 3782 8982 3834
rect 9034 3782 9046 3834
rect 9098 3782 9110 3834
rect 9162 3782 9174 3834
rect 9226 3782 16982 3834
rect 17034 3782 17046 3834
rect 17098 3782 17110 3834
rect 17162 3782 17174 3834
rect 17226 3782 22816 3834
rect 1104 3760 22816 3782
rect 2133 3723 2191 3729
rect 2133 3689 2145 3723
rect 2179 3720 2191 3723
rect 3418 3720 3424 3732
rect 2179 3692 3424 3720
rect 2179 3689 2191 3692
rect 2133 3683 2191 3689
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 5445 3723 5503 3729
rect 5445 3689 5457 3723
rect 5491 3720 5503 3723
rect 6270 3720 6276 3732
rect 5491 3692 6276 3720
rect 5491 3689 5503 3692
rect 5445 3683 5503 3689
rect 6270 3680 6276 3692
rect 6328 3720 6334 3732
rect 7374 3720 7380 3732
rect 6328 3692 6500 3720
rect 7335 3692 7380 3720
rect 6328 3680 6334 3692
rect 4430 3612 4436 3664
rect 4488 3652 4494 3664
rect 4846 3655 4904 3661
rect 4846 3652 4858 3655
rect 4488 3624 4858 3652
rect 4488 3612 4494 3624
rect 4846 3621 4858 3624
rect 4892 3652 4904 3655
rect 5534 3652 5540 3664
rect 4892 3624 5540 3652
rect 4892 3621 4904 3624
rect 4846 3615 4904 3621
rect 5534 3612 5540 3624
rect 5592 3612 5598 3664
rect 5626 3612 5632 3664
rect 5684 3652 5690 3664
rect 6472 3661 6500 3692
rect 7374 3680 7380 3692
rect 7432 3680 7438 3732
rect 7650 3680 7656 3732
rect 7708 3720 7714 3732
rect 7929 3723 7987 3729
rect 7929 3720 7941 3723
rect 7708 3692 7941 3720
rect 7708 3680 7714 3692
rect 7929 3689 7941 3692
rect 7975 3689 7987 3723
rect 7929 3683 7987 3689
rect 8941 3723 8999 3729
rect 8941 3689 8953 3723
rect 8987 3720 8999 3723
rect 9490 3720 9496 3732
rect 8987 3692 9496 3720
rect 8987 3689 8999 3692
rect 8941 3683 8999 3689
rect 9490 3680 9496 3692
rect 9548 3680 9554 3732
rect 9950 3720 9956 3732
rect 9911 3692 9956 3720
rect 9950 3680 9956 3692
rect 10008 3680 10014 3732
rect 10594 3680 10600 3732
rect 10652 3720 10658 3732
rect 10689 3723 10747 3729
rect 10689 3720 10701 3723
rect 10652 3692 10701 3720
rect 10652 3680 10658 3692
rect 10689 3689 10701 3692
rect 10735 3689 10747 3723
rect 10689 3683 10747 3689
rect 10962 3680 10968 3732
rect 11020 3720 11026 3732
rect 11149 3723 11207 3729
rect 11149 3720 11161 3723
rect 11020 3692 11161 3720
rect 11020 3680 11026 3692
rect 11149 3689 11161 3692
rect 11195 3689 11207 3723
rect 11149 3683 11207 3689
rect 5721 3655 5779 3661
rect 5721 3652 5733 3655
rect 5684 3624 5733 3652
rect 5684 3612 5690 3624
rect 5721 3621 5733 3624
rect 5767 3621 5779 3655
rect 5721 3615 5779 3621
rect 6457 3655 6515 3661
rect 6457 3621 6469 3655
rect 6503 3621 6515 3655
rect 6457 3615 6515 3621
rect 8110 3584 8116 3596
rect 8071 3556 8116 3584
rect 8110 3544 8116 3556
rect 8168 3544 8174 3596
rect 8389 3587 8447 3593
rect 8389 3553 8401 3587
rect 8435 3584 8447 3587
rect 8478 3584 8484 3596
rect 8435 3556 8484 3584
rect 8435 3553 8447 3556
rect 8389 3547 8447 3553
rect 8478 3544 8484 3556
rect 8536 3544 8542 3596
rect 9677 3587 9735 3593
rect 9677 3553 9689 3587
rect 9723 3553 9735 3587
rect 10226 3584 10232 3596
rect 10139 3556 10232 3584
rect 9677 3547 9735 3553
rect 4522 3516 4528 3528
rect 4483 3488 4528 3516
rect 4522 3476 4528 3488
rect 4580 3476 4586 3528
rect 6362 3516 6368 3528
rect 6323 3488 6368 3516
rect 6362 3476 6368 3488
rect 6420 3476 6426 3528
rect 6641 3519 6699 3525
rect 6641 3485 6653 3519
rect 6687 3485 6699 3519
rect 6641 3479 6699 3485
rect 5626 3408 5632 3460
rect 5684 3448 5690 3460
rect 6656 3448 6684 3479
rect 9582 3476 9588 3528
rect 9640 3516 9646 3528
rect 9692 3516 9720 3547
rect 10226 3544 10232 3556
rect 10284 3584 10290 3596
rect 10505 3587 10563 3593
rect 10505 3584 10517 3587
rect 10284 3556 10517 3584
rect 10284 3544 10290 3556
rect 10505 3553 10517 3556
rect 10551 3553 10563 3587
rect 10505 3547 10563 3553
rect 9640 3488 9720 3516
rect 11164 3516 11192 3683
rect 12250 3680 12256 3732
rect 12308 3720 12314 3732
rect 12621 3723 12679 3729
rect 12621 3720 12633 3723
rect 12308 3692 12633 3720
rect 12308 3680 12314 3692
rect 12621 3689 12633 3692
rect 12667 3689 12679 3723
rect 12621 3683 12679 3689
rect 13081 3723 13139 3729
rect 13081 3689 13093 3723
rect 13127 3720 13139 3723
rect 13538 3720 13544 3732
rect 13127 3692 13544 3720
rect 13127 3689 13139 3692
rect 13081 3683 13139 3689
rect 11514 3652 11520 3664
rect 11475 3624 11520 3652
rect 11514 3612 11520 3624
rect 11572 3612 11578 3664
rect 12636 3652 12664 3683
rect 13538 3680 13544 3692
rect 13596 3680 13602 3732
rect 16022 3720 16028 3732
rect 15983 3692 16028 3720
rect 16022 3680 16028 3692
rect 16080 3680 16086 3732
rect 17678 3720 17684 3732
rect 17639 3692 17684 3720
rect 17678 3680 17684 3692
rect 17736 3680 17742 3732
rect 19334 3720 19340 3732
rect 19295 3692 19340 3720
rect 19334 3680 19340 3692
rect 19392 3720 19398 3732
rect 19797 3723 19855 3729
rect 19797 3720 19809 3723
rect 19392 3692 19809 3720
rect 19392 3680 19398 3692
rect 19797 3689 19809 3692
rect 19843 3720 19855 3723
rect 19978 3720 19984 3732
rect 19843 3692 19984 3720
rect 19843 3689 19855 3692
rect 19797 3683 19855 3689
rect 19978 3680 19984 3692
rect 20036 3680 20042 3732
rect 13906 3652 13912 3664
rect 12636 3624 13912 3652
rect 13906 3612 13912 3624
rect 13964 3612 13970 3664
rect 13446 3544 13452 3596
rect 13504 3584 13510 3596
rect 13725 3587 13783 3593
rect 13725 3584 13737 3587
rect 13504 3556 13737 3584
rect 13504 3544 13510 3556
rect 13725 3553 13737 3556
rect 13771 3584 13783 3587
rect 15565 3587 15623 3593
rect 15565 3584 15577 3587
rect 13771 3556 15577 3584
rect 13771 3553 13783 3556
rect 13725 3547 13783 3553
rect 15565 3553 15577 3556
rect 15611 3584 15623 3587
rect 15654 3584 15660 3596
rect 15611 3556 15660 3584
rect 15611 3553 15623 3556
rect 15565 3547 15623 3553
rect 15654 3544 15660 3556
rect 15712 3544 15718 3596
rect 15746 3544 15752 3596
rect 15804 3584 15810 3596
rect 15841 3587 15899 3593
rect 15841 3584 15853 3587
rect 15804 3556 15853 3584
rect 15804 3544 15810 3556
rect 15841 3553 15853 3556
rect 15887 3584 15899 3587
rect 16206 3584 16212 3596
rect 15887 3556 16212 3584
rect 15887 3553 15899 3556
rect 15841 3547 15899 3553
rect 16206 3544 16212 3556
rect 16264 3544 16270 3596
rect 16850 3544 16856 3596
rect 16908 3584 16914 3596
rect 17129 3587 17187 3593
rect 17129 3584 17141 3587
rect 16908 3556 17141 3584
rect 16908 3544 16914 3556
rect 17129 3553 17141 3556
rect 17175 3553 17187 3587
rect 17696 3584 17724 3680
rect 18230 3612 18236 3664
rect 18288 3652 18294 3664
rect 18738 3655 18796 3661
rect 18738 3652 18750 3655
rect 18288 3624 18750 3652
rect 18288 3612 18294 3624
rect 18738 3621 18750 3624
rect 18784 3652 18796 3655
rect 19058 3652 19064 3664
rect 18784 3624 19064 3652
rect 18784 3621 18796 3624
rect 18738 3615 18796 3621
rect 19058 3612 19064 3624
rect 19116 3612 19122 3664
rect 18417 3587 18475 3593
rect 18417 3584 18429 3587
rect 17696 3556 18429 3584
rect 17129 3547 17187 3553
rect 18417 3553 18429 3556
rect 18463 3553 18475 3587
rect 18417 3547 18475 3553
rect 20936 3587 20994 3593
rect 20936 3553 20948 3587
rect 20982 3553 20994 3587
rect 20936 3547 20994 3553
rect 11425 3519 11483 3525
rect 11425 3516 11437 3519
rect 11164 3488 11437 3516
rect 9640 3476 9646 3488
rect 11425 3485 11437 3488
rect 11471 3485 11483 3519
rect 11698 3516 11704 3528
rect 11659 3488 11704 3516
rect 11425 3479 11483 3485
rect 11698 3476 11704 3488
rect 11756 3476 11762 3528
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3516 13599 3519
rect 14369 3519 14427 3525
rect 14369 3516 14381 3519
rect 13587 3488 14381 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 14369 3485 14381 3488
rect 14415 3516 14427 3519
rect 15378 3516 15384 3528
rect 14415 3488 15384 3516
rect 14415 3485 14427 3488
rect 14369 3479 14427 3485
rect 15378 3476 15384 3488
rect 15436 3476 15442 3528
rect 17770 3476 17776 3528
rect 17828 3516 17834 3528
rect 20806 3516 20812 3528
rect 17828 3488 20812 3516
rect 17828 3476 17834 3488
rect 20806 3476 20812 3488
rect 20864 3516 20870 3528
rect 20951 3516 20979 3547
rect 20864 3488 20979 3516
rect 20864 3476 20870 3488
rect 5684 3420 6684 3448
rect 9493 3451 9551 3457
rect 5684 3408 5690 3420
rect 9493 3417 9505 3451
rect 9539 3448 9551 3451
rect 9674 3448 9680 3460
rect 9539 3420 9680 3448
rect 9539 3417 9551 3420
rect 9493 3411 9551 3417
rect 9674 3408 9680 3420
rect 9732 3448 9738 3460
rect 11716 3448 11744 3476
rect 13262 3448 13268 3460
rect 9732 3420 11744 3448
rect 12452 3420 13268 3448
rect 9732 3408 9738 3420
rect 7745 3383 7803 3389
rect 7745 3349 7757 3383
rect 7791 3380 7803 3383
rect 8386 3380 8392 3392
rect 7791 3352 8392 3380
rect 7791 3349 7803 3352
rect 7745 3343 7803 3349
rect 8386 3340 8392 3352
rect 8444 3340 8450 3392
rect 10505 3383 10563 3389
rect 10505 3349 10517 3383
rect 10551 3380 10563 3383
rect 12452 3380 12480 3420
rect 13262 3408 13268 3420
rect 13320 3408 13326 3460
rect 13354 3408 13360 3460
rect 13412 3448 13418 3460
rect 15470 3448 15476 3460
rect 13412 3420 15476 3448
rect 13412 3408 13418 3420
rect 15470 3408 15476 3420
rect 15528 3408 15534 3460
rect 15657 3451 15715 3457
rect 15657 3417 15669 3451
rect 15703 3448 15715 3451
rect 16114 3448 16120 3460
rect 15703 3420 16120 3448
rect 15703 3417 15715 3420
rect 15657 3411 15715 3417
rect 16114 3408 16120 3420
rect 16172 3448 16178 3460
rect 16172 3420 16712 3448
rect 16172 3408 16178 3420
rect 16684 3392 16712 3420
rect 10551 3352 12480 3380
rect 15105 3383 15163 3389
rect 10551 3349 10563 3352
rect 10505 3343 10563 3349
rect 15105 3349 15117 3383
rect 15151 3380 15163 3383
rect 15930 3380 15936 3392
rect 15151 3352 15936 3380
rect 15151 3349 15163 3352
rect 15105 3343 15163 3349
rect 15930 3340 15936 3352
rect 15988 3340 15994 3392
rect 16666 3380 16672 3392
rect 16627 3352 16672 3380
rect 16666 3340 16672 3352
rect 16724 3340 16730 3392
rect 17310 3380 17316 3392
rect 17271 3352 17316 3380
rect 17310 3340 17316 3352
rect 17368 3340 17374 3392
rect 18046 3380 18052 3392
rect 18007 3352 18052 3380
rect 18046 3340 18052 3352
rect 18104 3340 18110 3392
rect 19886 3340 19892 3392
rect 19944 3380 19950 3392
rect 20257 3383 20315 3389
rect 20257 3380 20269 3383
rect 19944 3352 20269 3380
rect 19944 3340 19950 3352
rect 20257 3349 20269 3352
rect 20303 3380 20315 3383
rect 21039 3383 21097 3389
rect 21039 3380 21051 3383
rect 20303 3352 21051 3380
rect 20303 3349 20315 3352
rect 20257 3343 20315 3349
rect 21039 3349 21051 3352
rect 21085 3349 21097 3383
rect 21039 3343 21097 3349
rect 1104 3290 22816 3312
rect 1104 3238 4982 3290
rect 5034 3238 5046 3290
rect 5098 3238 5110 3290
rect 5162 3238 5174 3290
rect 5226 3238 12982 3290
rect 13034 3238 13046 3290
rect 13098 3238 13110 3290
rect 13162 3238 13174 3290
rect 13226 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 22816 3290
rect 1104 3216 22816 3238
rect 4522 3136 4528 3188
rect 4580 3176 4586 3188
rect 5905 3179 5963 3185
rect 5905 3176 5917 3179
rect 4580 3148 5917 3176
rect 4580 3136 4586 3148
rect 5905 3145 5917 3148
rect 5951 3145 5963 3179
rect 6270 3176 6276 3188
rect 6231 3148 6276 3176
rect 5905 3139 5963 3145
rect 6270 3136 6276 3148
rect 6328 3136 6334 3188
rect 7929 3179 7987 3185
rect 7929 3145 7941 3179
rect 7975 3176 7987 3179
rect 8478 3176 8484 3188
rect 7975 3148 8484 3176
rect 7975 3145 7987 3148
rect 7929 3139 7987 3145
rect 8478 3136 8484 3148
rect 8536 3176 8542 3188
rect 9493 3179 9551 3185
rect 9493 3176 9505 3179
rect 8536 3148 9505 3176
rect 8536 3136 8542 3148
rect 9493 3145 9505 3148
rect 9539 3176 9551 3179
rect 10226 3176 10232 3188
rect 9539 3148 10232 3176
rect 9539 3145 9551 3148
rect 9493 3139 9551 3145
rect 10226 3136 10232 3148
rect 10284 3136 10290 3188
rect 10870 3176 10876 3188
rect 10831 3148 10876 3176
rect 10870 3136 10876 3148
rect 10928 3136 10934 3188
rect 11514 3176 11520 3188
rect 11475 3148 11520 3176
rect 11514 3136 11520 3148
rect 11572 3136 11578 3188
rect 12250 3176 12256 3188
rect 12211 3148 12256 3176
rect 12250 3136 12256 3148
rect 12308 3136 12314 3188
rect 19058 3176 19064 3188
rect 19019 3148 19064 3176
rect 19058 3136 19064 3148
rect 19116 3136 19122 3188
rect 20806 3136 20812 3188
rect 20864 3176 20870 3188
rect 20901 3179 20959 3185
rect 20901 3176 20913 3179
rect 20864 3148 20913 3176
rect 20864 3136 20870 3148
rect 20901 3145 20913 3148
rect 20947 3145 20959 3179
rect 20901 3139 20959 3145
rect 4540 3108 4568 3136
rect 3988 3080 4568 3108
rect 3418 3000 3424 3052
rect 3476 3040 3482 3052
rect 3988 3049 4016 3080
rect 9398 3068 9404 3120
rect 9456 3108 9462 3120
rect 9769 3111 9827 3117
rect 9769 3108 9781 3111
rect 9456 3080 9781 3108
rect 9456 3068 9462 3080
rect 9769 3077 9781 3080
rect 9815 3077 9827 3111
rect 9769 3071 9827 3077
rect 3973 3043 4031 3049
rect 3476 3012 3832 3040
rect 3476 3000 3482 3012
rect 3804 2981 3832 3012
rect 3973 3009 3985 3043
rect 4019 3009 4031 3043
rect 5626 3040 5632 3052
rect 5587 3012 5632 3040
rect 3973 3003 4031 3009
rect 5626 3000 5632 3012
rect 5684 3000 5690 3052
rect 8941 3043 8999 3049
rect 8941 3009 8953 3043
rect 8987 3040 8999 3043
rect 9674 3040 9680 3052
rect 8987 3012 9680 3040
rect 8987 3009 8999 3012
rect 8941 3003 8999 3009
rect 9674 3000 9680 3012
rect 9732 3000 9738 3052
rect 3605 2975 3663 2981
rect 3605 2941 3617 2975
rect 3651 2941 3663 2975
rect 3605 2935 3663 2941
rect 3789 2975 3847 2981
rect 3789 2941 3801 2975
rect 3835 2941 3847 2975
rect 7098 2972 7104 2984
rect 7011 2944 7104 2972
rect 3789 2935 3847 2941
rect 3237 2907 3295 2913
rect 3237 2873 3249 2907
rect 3283 2904 3295 2907
rect 3620 2904 3648 2935
rect 7098 2932 7104 2944
rect 7156 2972 7162 2984
rect 8110 2972 8116 2984
rect 7156 2944 8116 2972
rect 7156 2932 7162 2944
rect 8110 2932 8116 2944
rect 8168 2932 8174 2984
rect 4614 2904 4620 2916
rect 3283 2876 4620 2904
rect 3283 2873 3295 2876
rect 3237 2867 3295 2873
rect 4614 2864 4620 2876
rect 4672 2864 4678 2916
rect 4982 2904 4988 2916
rect 4943 2876 4988 2904
rect 4982 2864 4988 2876
rect 5040 2864 5046 2916
rect 5074 2864 5080 2916
rect 5132 2904 5138 2916
rect 7193 2907 7251 2913
rect 5132 2876 5177 2904
rect 5132 2864 5138 2876
rect 7193 2873 7205 2907
rect 7239 2904 7251 2907
rect 8294 2904 8300 2916
rect 7239 2876 8300 2904
rect 7239 2873 7251 2876
rect 7193 2867 7251 2873
rect 8294 2864 8300 2876
rect 8352 2864 8358 2916
rect 8386 2864 8392 2916
rect 8444 2904 8450 2916
rect 9784 2904 9812 3071
rect 11054 3068 11060 3120
rect 11112 3108 11118 3120
rect 12621 3111 12679 3117
rect 12621 3108 12633 3111
rect 11112 3080 12633 3108
rect 11112 3068 11118 3080
rect 12621 3077 12633 3080
rect 12667 3077 12679 3111
rect 12621 3071 12679 3077
rect 15013 3111 15071 3117
rect 15013 3077 15025 3111
rect 15059 3108 15071 3111
rect 16758 3108 16764 3120
rect 15059 3080 16764 3108
rect 15059 3077 15071 3080
rect 15013 3071 15071 3077
rect 16758 3068 16764 3080
rect 16816 3068 16822 3120
rect 17037 3111 17095 3117
rect 17037 3077 17049 3111
rect 17083 3108 17095 3111
rect 17313 3111 17371 3117
rect 17313 3108 17325 3111
rect 17083 3080 17325 3108
rect 17083 3077 17095 3080
rect 17037 3071 17095 3077
rect 17313 3077 17325 3080
rect 17359 3108 17371 3111
rect 17865 3111 17923 3117
rect 17865 3108 17877 3111
rect 17359 3080 17877 3108
rect 17359 3077 17371 3080
rect 17313 3071 17371 3077
rect 17865 3077 17877 3080
rect 17911 3108 17923 3111
rect 18230 3108 18236 3120
rect 17911 3080 18236 3108
rect 17911 3077 17923 3080
rect 17865 3071 17923 3077
rect 9950 3040 9956 3052
rect 9911 3012 9956 3040
rect 9950 3000 9956 3012
rect 10008 3040 10014 3052
rect 11149 3043 11207 3049
rect 11149 3040 11161 3043
rect 10008 3012 11161 3040
rect 10008 3000 10014 3012
rect 11149 3009 11161 3012
rect 11195 3009 11207 3043
rect 15930 3040 15936 3052
rect 15891 3012 15936 3040
rect 11149 3003 11207 3009
rect 15930 3000 15936 3012
rect 15988 3000 15994 3052
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2972 12495 2975
rect 13078 2972 13084 2984
rect 12483 2944 13084 2972
rect 12483 2941 12495 2944
rect 12437 2935 12495 2941
rect 13078 2932 13084 2944
rect 13136 2932 13142 2984
rect 13630 2972 13636 2984
rect 13591 2944 13636 2972
rect 13630 2932 13636 2944
rect 13688 2932 13694 2984
rect 13906 2932 13912 2984
rect 13964 2972 13970 2984
rect 14093 2975 14151 2981
rect 14093 2972 14105 2975
rect 13964 2944 14105 2972
rect 13964 2932 13970 2944
rect 14093 2941 14105 2944
rect 14139 2941 14151 2975
rect 14093 2935 14151 2941
rect 14366 2932 14372 2984
rect 14424 2972 14430 2984
rect 14461 2975 14519 2981
rect 14461 2972 14473 2975
rect 14424 2944 14473 2972
rect 14424 2932 14430 2944
rect 14461 2941 14473 2944
rect 14507 2941 14519 2975
rect 14461 2935 14519 2941
rect 15013 2975 15071 2981
rect 15013 2941 15025 2975
rect 15059 2972 15071 2975
rect 15378 2972 15384 2984
rect 15059 2944 15384 2972
rect 15059 2941 15071 2944
rect 15013 2935 15071 2941
rect 15378 2932 15384 2944
rect 15436 2972 15442 2984
rect 16022 2972 16028 2984
rect 15436 2944 16028 2972
rect 15436 2932 15442 2944
rect 16022 2932 16028 2944
rect 16080 2932 16086 2984
rect 16577 2975 16635 2981
rect 16577 2941 16589 2975
rect 16623 2972 16635 2975
rect 16666 2972 16672 2984
rect 16623 2944 16672 2972
rect 16623 2941 16635 2944
rect 16577 2935 16635 2941
rect 16666 2932 16672 2944
rect 16724 2972 16730 2984
rect 17052 2972 17080 3071
rect 18230 3068 18236 3080
rect 18288 3068 18294 3120
rect 17402 3000 17408 3052
rect 17460 3040 17466 3052
rect 19429 3043 19487 3049
rect 19429 3040 19441 3043
rect 17460 3012 19441 3040
rect 17460 3000 17466 3012
rect 18046 2972 18052 2984
rect 16724 2944 17080 2972
rect 18007 2944 18052 2972
rect 16724 2932 16730 2944
rect 18046 2932 18052 2944
rect 18104 2932 18110 2984
rect 18141 2975 18199 2981
rect 18141 2941 18153 2975
rect 18187 2972 18199 2975
rect 18230 2972 18236 2984
rect 18187 2944 18236 2972
rect 18187 2941 18199 2944
rect 18141 2935 18199 2941
rect 18230 2932 18236 2944
rect 18288 2932 18294 2984
rect 18340 2981 18368 3012
rect 19429 3009 19441 3012
rect 19475 3009 19487 3043
rect 19886 3040 19892 3052
rect 19847 3012 19892 3040
rect 19429 3003 19487 3009
rect 19886 3000 19892 3012
rect 19944 3000 19950 3052
rect 20346 3040 20352 3052
rect 20307 3012 20352 3040
rect 20346 3000 20352 3012
rect 20404 3000 20410 3052
rect 18325 2975 18383 2981
rect 18325 2941 18337 2975
rect 18371 2941 18383 2975
rect 18325 2935 18383 2941
rect 10274 2907 10332 2913
rect 10274 2904 10286 2907
rect 8444 2876 8489 2904
rect 9784 2876 10286 2904
rect 8444 2864 8450 2876
rect 10274 2873 10286 2876
rect 10320 2904 10332 2907
rect 10594 2904 10600 2916
rect 10320 2876 10600 2904
rect 10320 2873 10332 2876
rect 10274 2867 10332 2873
rect 10594 2864 10600 2876
rect 10652 2864 10658 2916
rect 15470 2864 15476 2916
rect 15528 2904 15534 2916
rect 19978 2904 19984 2916
rect 15528 2876 18552 2904
rect 19939 2876 19984 2904
rect 15528 2864 15534 2876
rect 18156 2848 18184 2876
rect 4522 2836 4528 2848
rect 4483 2808 4528 2836
rect 4522 2796 4528 2808
rect 4580 2796 4586 2848
rect 13446 2836 13452 2848
rect 13407 2808 13452 2836
rect 13446 2796 13452 2808
rect 13504 2796 13510 2848
rect 15654 2836 15660 2848
rect 15615 2808 15660 2836
rect 15654 2796 15660 2808
rect 15712 2796 15718 2848
rect 16022 2796 16028 2848
rect 16080 2836 16086 2848
rect 18046 2836 18052 2848
rect 16080 2808 18052 2836
rect 16080 2796 16086 2808
rect 18046 2796 18052 2808
rect 18104 2796 18110 2848
rect 18138 2796 18144 2848
rect 18196 2796 18202 2848
rect 18524 2845 18552 2876
rect 19978 2864 19984 2876
rect 20036 2864 20042 2916
rect 18509 2839 18567 2845
rect 18509 2805 18521 2839
rect 18555 2805 18567 2839
rect 18509 2799 18567 2805
rect 1104 2746 22816 2768
rect 1104 2694 8982 2746
rect 9034 2694 9046 2746
rect 9098 2694 9110 2746
rect 9162 2694 9174 2746
rect 9226 2694 16982 2746
rect 17034 2694 17046 2746
rect 17098 2694 17110 2746
rect 17162 2694 17174 2746
rect 17226 2694 22816 2746
rect 1104 2672 22816 2694
rect 1854 2592 1860 2644
rect 1912 2632 1918 2644
rect 2133 2635 2191 2641
rect 2133 2632 2145 2635
rect 1912 2604 2145 2632
rect 1912 2592 1918 2604
rect 2133 2601 2145 2604
rect 2179 2632 2191 2635
rect 2225 2635 2283 2641
rect 2225 2632 2237 2635
rect 2179 2604 2237 2632
rect 2179 2601 2191 2604
rect 2133 2595 2191 2601
rect 2225 2601 2237 2604
rect 2271 2601 2283 2635
rect 2225 2595 2283 2601
rect 4982 2592 4988 2644
rect 5040 2632 5046 2644
rect 5261 2635 5319 2641
rect 5261 2632 5273 2635
rect 5040 2604 5273 2632
rect 5040 2592 5046 2604
rect 5261 2601 5273 2604
rect 5307 2632 5319 2635
rect 5813 2635 5871 2641
rect 5813 2632 5825 2635
rect 5307 2604 5825 2632
rect 5307 2601 5319 2604
rect 5261 2595 5319 2601
rect 5813 2601 5825 2604
rect 5859 2601 5871 2635
rect 6362 2632 6368 2644
rect 6323 2604 6368 2632
rect 5813 2595 5871 2601
rect 6362 2592 6368 2604
rect 6420 2592 6426 2644
rect 7466 2632 7472 2644
rect 7427 2604 7472 2632
rect 7466 2592 7472 2604
rect 7524 2592 7530 2644
rect 8386 2592 8392 2644
rect 8444 2632 8450 2644
rect 8573 2635 8631 2641
rect 8573 2632 8585 2635
rect 8444 2604 8585 2632
rect 8444 2592 8450 2604
rect 8573 2601 8585 2604
rect 8619 2601 8631 2635
rect 8573 2595 8631 2601
rect 9582 2592 9588 2644
rect 9640 2632 9646 2644
rect 10229 2635 10287 2641
rect 10229 2632 10241 2635
rect 9640 2604 10241 2632
rect 9640 2592 9646 2604
rect 10229 2601 10241 2604
rect 10275 2601 10287 2635
rect 10594 2632 10600 2644
rect 10555 2604 10600 2632
rect 10229 2595 10287 2601
rect 10594 2592 10600 2604
rect 10652 2632 10658 2644
rect 10652 2604 11145 2632
rect 10652 2592 10658 2604
rect 1949 2567 2007 2573
rect 1949 2533 1961 2567
rect 1995 2564 2007 2567
rect 3418 2564 3424 2576
rect 1995 2536 3424 2564
rect 1995 2533 2007 2536
rect 1949 2527 2007 2533
rect 2976 2505 3004 2536
rect 3418 2524 3424 2536
rect 3476 2524 3482 2576
rect 3697 2567 3755 2573
rect 3697 2533 3709 2567
rect 3743 2564 3755 2567
rect 4386 2567 4444 2573
rect 4386 2564 4398 2567
rect 3743 2536 4398 2564
rect 3743 2533 3755 2536
rect 3697 2527 3755 2533
rect 4386 2533 4398 2536
rect 4432 2564 4444 2567
rect 4522 2564 4528 2576
rect 4432 2536 4528 2564
rect 4432 2533 4444 2536
rect 4386 2527 4444 2533
rect 4522 2524 4528 2536
rect 4580 2524 4586 2576
rect 7484 2564 7512 2592
rect 7974 2567 8032 2573
rect 7974 2564 7986 2567
rect 7484 2536 7986 2564
rect 7974 2533 7986 2536
rect 8020 2533 8032 2567
rect 7974 2527 8032 2533
rect 8294 2524 8300 2576
rect 8352 2564 8358 2576
rect 11117 2573 11145 2604
rect 11514 2592 11520 2644
rect 11572 2632 11578 2644
rect 11701 2635 11759 2641
rect 11701 2632 11713 2635
rect 11572 2604 11713 2632
rect 11572 2592 11578 2604
rect 11701 2601 11713 2604
rect 11747 2601 11759 2635
rect 12713 2635 12771 2641
rect 12713 2632 12725 2635
rect 11701 2595 11759 2601
rect 11808 2604 12725 2632
rect 8849 2567 8907 2573
rect 8849 2564 8861 2567
rect 8352 2536 8861 2564
rect 8352 2524 8358 2536
rect 8849 2533 8861 2536
rect 8895 2533 8907 2567
rect 8849 2527 8907 2533
rect 11102 2567 11160 2573
rect 11102 2533 11114 2567
rect 11148 2533 11160 2567
rect 11102 2527 11160 2533
rect 2133 2499 2191 2505
rect 2133 2465 2145 2499
rect 2179 2496 2191 2499
rect 2409 2499 2467 2505
rect 2409 2496 2421 2499
rect 2179 2468 2421 2496
rect 2179 2465 2191 2468
rect 2133 2459 2191 2465
rect 2409 2465 2421 2468
rect 2455 2465 2467 2499
rect 2409 2459 2467 2465
rect 2961 2499 3019 2505
rect 2961 2465 2973 2499
rect 3007 2465 3019 2499
rect 2961 2459 3019 2465
rect 4985 2499 5043 2505
rect 4985 2465 4997 2499
rect 5031 2496 5043 2499
rect 5074 2496 5080 2508
rect 5031 2468 5080 2496
rect 5031 2465 5043 2468
rect 4985 2459 5043 2465
rect 2424 2360 2452 2459
rect 5074 2456 5080 2468
rect 5132 2496 5138 2508
rect 5629 2499 5687 2505
rect 5629 2496 5641 2499
rect 5132 2468 5641 2496
rect 5132 2456 5138 2468
rect 5629 2465 5641 2468
rect 5675 2465 5687 2499
rect 5629 2459 5687 2465
rect 7193 2499 7251 2505
rect 7193 2465 7205 2499
rect 7239 2496 7251 2499
rect 7650 2496 7656 2508
rect 7239 2468 7656 2496
rect 7239 2465 7251 2468
rect 7193 2459 7251 2465
rect 7650 2456 7656 2468
rect 7708 2456 7714 2508
rect 9674 2496 9680 2508
rect 9635 2468 9680 2496
rect 9674 2456 9680 2468
rect 9732 2456 9738 2508
rect 10781 2499 10839 2505
rect 10781 2465 10793 2499
rect 10827 2496 10839 2499
rect 11808 2496 11836 2604
rect 12713 2601 12725 2604
rect 12759 2601 12771 2635
rect 13630 2632 13636 2644
rect 13591 2604 13636 2632
rect 12713 2595 12771 2601
rect 13630 2592 13636 2604
rect 13688 2592 13694 2644
rect 14093 2635 14151 2641
rect 14093 2601 14105 2635
rect 14139 2632 14151 2635
rect 14366 2632 14372 2644
rect 14139 2604 14372 2632
rect 14139 2601 14151 2604
rect 14093 2595 14151 2601
rect 14366 2592 14372 2604
rect 14424 2592 14430 2644
rect 16390 2632 16396 2644
rect 16351 2604 16396 2632
rect 16390 2592 16396 2604
rect 16448 2592 16454 2644
rect 18046 2592 18052 2644
rect 18104 2632 18110 2644
rect 19337 2635 19395 2641
rect 19337 2632 19349 2635
rect 18104 2604 19349 2632
rect 18104 2592 18110 2604
rect 19337 2601 19349 2604
rect 19383 2601 19395 2635
rect 19337 2595 19395 2601
rect 20533 2635 20591 2641
rect 20533 2601 20545 2635
rect 20579 2632 20591 2635
rect 20806 2632 20812 2644
rect 20579 2604 20812 2632
rect 20579 2601 20591 2604
rect 20533 2595 20591 2601
rect 12437 2567 12495 2573
rect 12437 2533 12449 2567
rect 12483 2564 12495 2567
rect 12483 2536 13216 2564
rect 12483 2533 12495 2536
rect 12437 2527 12495 2533
rect 13188 2505 13216 2536
rect 15654 2524 15660 2576
rect 15712 2564 15718 2576
rect 20548 2564 20576 2595
rect 20806 2592 20812 2604
rect 20864 2592 20870 2644
rect 15712 2536 18184 2564
rect 15712 2524 15718 2536
rect 10827 2468 11836 2496
rect 12897 2499 12955 2505
rect 10827 2465 10839 2468
rect 10781 2459 10839 2465
rect 12897 2465 12909 2499
rect 12943 2465 12955 2499
rect 12897 2459 12955 2465
rect 13173 2499 13231 2505
rect 13173 2465 13185 2499
rect 13219 2496 13231 2499
rect 13262 2496 13268 2508
rect 13219 2468 13268 2496
rect 13219 2465 13231 2468
rect 13173 2459 13231 2465
rect 3145 2431 3203 2437
rect 3145 2397 3157 2431
rect 3191 2428 3203 2431
rect 3421 2431 3479 2437
rect 3421 2428 3433 2431
rect 3191 2400 3433 2428
rect 3191 2397 3203 2400
rect 3145 2391 3203 2397
rect 3421 2397 3433 2400
rect 3467 2428 3479 2431
rect 4065 2431 4123 2437
rect 4065 2428 4077 2431
rect 3467 2400 4077 2428
rect 3467 2397 3479 2400
rect 3421 2391 3479 2397
rect 4065 2397 4077 2400
rect 4111 2397 4123 2431
rect 4065 2391 4123 2397
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2428 9643 2431
rect 10796 2428 10824 2459
rect 9631 2400 10824 2428
rect 12069 2431 12127 2437
rect 9631 2397 9643 2400
rect 9585 2391 9643 2397
rect 12069 2397 12081 2431
rect 12115 2428 12127 2431
rect 12912 2428 12940 2459
rect 13262 2456 13268 2468
rect 13320 2456 13326 2508
rect 14182 2496 14188 2508
rect 14143 2468 14188 2496
rect 14182 2456 14188 2468
rect 14240 2496 14246 2508
rect 14737 2499 14795 2505
rect 14737 2496 14749 2499
rect 14240 2468 14749 2496
rect 14240 2456 14246 2468
rect 14737 2465 14749 2468
rect 14783 2465 14795 2499
rect 14737 2459 14795 2465
rect 15933 2499 15991 2505
rect 15933 2465 15945 2499
rect 15979 2496 15991 2499
rect 16022 2496 16028 2508
rect 15979 2468 16028 2496
rect 15979 2465 15991 2468
rect 15933 2459 15991 2465
rect 16022 2456 16028 2468
rect 16080 2456 16086 2508
rect 16206 2496 16212 2508
rect 16167 2468 16212 2496
rect 16206 2456 16212 2468
rect 16264 2456 16270 2508
rect 16850 2456 16856 2508
rect 16908 2496 16914 2508
rect 17126 2496 17132 2508
rect 16908 2468 17132 2496
rect 16908 2456 16914 2468
rect 17126 2456 17132 2468
rect 17184 2456 17190 2508
rect 18156 2505 18184 2536
rect 19904 2536 20576 2564
rect 18141 2499 18199 2505
rect 18141 2465 18153 2499
rect 18187 2496 18199 2499
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 18187 2468 18337 2496
rect 18187 2465 18199 2468
rect 18141 2459 18199 2465
rect 18325 2465 18337 2468
rect 18371 2465 18383 2499
rect 18598 2496 18604 2508
rect 18559 2468 18604 2496
rect 18325 2459 18383 2465
rect 18598 2456 18604 2468
rect 18656 2456 18662 2508
rect 19904 2505 19932 2536
rect 19889 2499 19947 2505
rect 19889 2465 19901 2499
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 20438 2456 20444 2508
rect 20496 2496 20502 2508
rect 21177 2499 21235 2505
rect 21177 2496 21189 2499
rect 20496 2468 21189 2496
rect 20496 2456 20502 2468
rect 21177 2465 21189 2468
rect 21223 2496 21235 2499
rect 21729 2499 21787 2505
rect 21729 2496 21741 2499
rect 21223 2468 21741 2496
rect 21223 2465 21235 2468
rect 21177 2459 21235 2465
rect 21729 2465 21741 2468
rect 21775 2465 21787 2499
rect 21729 2459 21787 2465
rect 13722 2428 13728 2440
rect 12115 2400 13728 2428
rect 12115 2397 12127 2400
rect 12069 2391 12127 2397
rect 13722 2388 13728 2400
rect 13780 2388 13786 2440
rect 17862 2428 17868 2440
rect 15120 2400 17868 2428
rect 7098 2360 7104 2372
rect 2424 2332 7104 2360
rect 7098 2320 7104 2332
rect 7156 2320 7162 2372
rect 9214 2320 9220 2372
rect 9272 2360 9278 2372
rect 9907 2363 9965 2369
rect 9907 2360 9919 2363
rect 9272 2332 9919 2360
rect 9272 2320 9278 2332
rect 9907 2329 9919 2332
rect 9953 2329 9965 2363
rect 9907 2323 9965 2329
rect 13262 2320 13268 2372
rect 13320 2360 13326 2372
rect 14369 2363 14427 2369
rect 14369 2360 14381 2363
rect 13320 2332 14381 2360
rect 13320 2320 13326 2332
rect 14369 2329 14381 2332
rect 14415 2329 14427 2363
rect 14369 2323 14427 2329
rect 3142 2252 3148 2304
rect 3200 2292 3206 2304
rect 3697 2295 3755 2301
rect 3697 2292 3709 2295
rect 3200 2264 3709 2292
rect 3200 2252 3206 2264
rect 3697 2261 3709 2264
rect 3743 2292 3755 2295
rect 3789 2295 3847 2301
rect 3789 2292 3801 2295
rect 3743 2264 3801 2292
rect 3743 2261 3755 2264
rect 3697 2255 3755 2261
rect 3789 2261 3801 2264
rect 3835 2261 3847 2295
rect 3789 2255 3847 2261
rect 13722 2252 13728 2304
rect 13780 2292 13786 2304
rect 15120 2292 15148 2400
rect 17862 2388 17868 2400
rect 17920 2428 17926 2440
rect 18785 2431 18843 2437
rect 18785 2428 18797 2431
rect 17920 2400 18797 2428
rect 17920 2388 17926 2400
rect 18785 2397 18797 2400
rect 18831 2397 18843 2431
rect 18785 2391 18843 2397
rect 15930 2320 15936 2372
rect 15988 2360 15994 2372
rect 16025 2363 16083 2369
rect 16025 2360 16037 2363
rect 15988 2332 16037 2360
rect 15988 2320 15994 2332
rect 16025 2329 16037 2332
rect 16071 2360 16083 2363
rect 18417 2363 18475 2369
rect 18417 2360 18429 2363
rect 16071 2332 18429 2360
rect 16071 2329 16083 2332
rect 16025 2323 16083 2329
rect 18417 2329 18429 2332
rect 18463 2360 18475 2363
rect 19705 2363 19763 2369
rect 19705 2360 19717 2363
rect 18463 2332 19717 2360
rect 18463 2329 18475 2332
rect 18417 2323 18475 2329
rect 19705 2329 19717 2332
rect 19751 2329 19763 2363
rect 19705 2323 19763 2329
rect 20073 2363 20131 2369
rect 20073 2329 20085 2363
rect 20119 2360 20131 2363
rect 20622 2360 20628 2372
rect 20119 2332 20628 2360
rect 20119 2329 20131 2332
rect 20073 2323 20131 2329
rect 20622 2320 20628 2332
rect 20680 2320 20686 2372
rect 21361 2363 21419 2369
rect 21361 2329 21373 2363
rect 21407 2360 21419 2363
rect 22646 2360 22652 2372
rect 21407 2332 22652 2360
rect 21407 2329 21419 2332
rect 21361 2323 21419 2329
rect 22646 2320 22652 2332
rect 22704 2320 22710 2372
rect 13780 2264 15148 2292
rect 15289 2295 15347 2301
rect 13780 2252 13786 2264
rect 15289 2261 15301 2295
rect 15335 2292 15347 2295
rect 15749 2295 15807 2301
rect 15749 2292 15761 2295
rect 15335 2264 15761 2292
rect 15335 2261 15347 2264
rect 15289 2255 15347 2261
rect 15749 2261 15761 2264
rect 15795 2292 15807 2295
rect 16206 2292 16212 2304
rect 15795 2264 16212 2292
rect 15795 2261 15807 2264
rect 15749 2255 15807 2261
rect 16206 2252 16212 2264
rect 16264 2292 16270 2304
rect 17773 2295 17831 2301
rect 17773 2292 17785 2295
rect 16264 2264 17785 2292
rect 16264 2252 16270 2264
rect 17773 2261 17785 2264
rect 17819 2292 17831 2295
rect 18598 2292 18604 2304
rect 17819 2264 18604 2292
rect 17819 2261 17831 2264
rect 17773 2255 17831 2261
rect 18598 2252 18604 2264
rect 18656 2252 18662 2304
rect 1104 2202 22816 2224
rect 1104 2150 4982 2202
rect 5034 2150 5046 2202
rect 5098 2150 5110 2202
rect 5162 2150 5174 2202
rect 5226 2150 12982 2202
rect 13034 2150 13046 2202
rect 13098 2150 13110 2202
rect 13162 2150 13174 2202
rect 13226 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 22816 2202
rect 1104 2128 22816 2150
rect 5166 1980 5172 2032
rect 5224 2020 5230 2032
rect 11606 2020 11612 2032
rect 5224 1992 11612 2020
rect 5224 1980 5230 1992
rect 11606 1980 11612 1992
rect 11664 1980 11670 2032
<< via1 >>
rect 13820 23536 13872 23588
rect 14648 23536 14700 23588
rect 4982 21734 5034 21786
rect 5046 21734 5098 21786
rect 5110 21734 5162 21786
rect 5174 21734 5226 21786
rect 12982 21734 13034 21786
rect 13046 21734 13098 21786
rect 13110 21734 13162 21786
rect 13174 21734 13226 21786
rect 20982 21734 21034 21786
rect 21046 21734 21098 21786
rect 21110 21734 21162 21786
rect 21174 21734 21226 21786
rect 8982 21190 9034 21242
rect 9046 21190 9098 21242
rect 9110 21190 9162 21242
rect 9174 21190 9226 21242
rect 16982 21190 17034 21242
rect 17046 21190 17098 21242
rect 17110 21190 17162 21242
rect 17174 21190 17226 21242
rect 8208 20927 8260 20936
rect 8208 20893 8217 20927
rect 8217 20893 8251 20927
rect 8251 20893 8260 20927
rect 8208 20884 8260 20893
rect 18420 20884 18472 20936
rect 4982 20646 5034 20698
rect 5046 20646 5098 20698
rect 5110 20646 5162 20698
rect 5174 20646 5226 20698
rect 12982 20646 13034 20698
rect 13046 20646 13098 20698
rect 13110 20646 13162 20698
rect 13174 20646 13226 20698
rect 20982 20646 21034 20698
rect 21046 20646 21098 20698
rect 21110 20646 21162 20698
rect 21174 20646 21226 20698
rect 1584 20587 1636 20596
rect 1584 20553 1593 20587
rect 1593 20553 1627 20587
rect 1627 20553 1636 20587
rect 1584 20544 1636 20553
rect 6368 20544 6420 20596
rect 8208 20544 8260 20596
rect 8576 20544 8628 20596
rect 11612 20544 11664 20596
rect 19708 20544 19760 20596
rect 20352 20587 20404 20596
rect 20352 20553 20361 20587
rect 20361 20553 20395 20587
rect 20395 20553 20404 20587
rect 20352 20544 20404 20553
rect 4160 20476 4212 20528
rect 9404 20476 9456 20528
rect 8576 20451 8628 20460
rect 8576 20417 8585 20451
rect 8585 20417 8619 20451
rect 8619 20417 8628 20451
rect 8576 20408 8628 20417
rect 5540 20340 5592 20392
rect 10968 20383 11020 20392
rect 10968 20349 10977 20383
rect 10977 20349 11011 20383
rect 11011 20349 11020 20383
rect 10968 20340 11020 20349
rect 8760 20272 8812 20324
rect 11336 20272 11388 20324
rect 11612 20204 11664 20256
rect 18880 20340 18932 20392
rect 19248 20340 19300 20392
rect 13360 20204 13412 20256
rect 8982 20102 9034 20154
rect 9046 20102 9098 20154
rect 9110 20102 9162 20154
rect 9174 20102 9226 20154
rect 16982 20102 17034 20154
rect 17046 20102 17098 20154
rect 17110 20102 17162 20154
rect 17174 20102 17226 20154
rect 8760 20043 8812 20052
rect 8760 20009 8769 20043
rect 8769 20009 8803 20043
rect 8803 20009 8812 20043
rect 8760 20000 8812 20009
rect 5356 19932 5408 19984
rect 8668 19932 8720 19984
rect 10784 19975 10836 19984
rect 10784 19941 10793 19975
rect 10793 19941 10827 19975
rect 10827 19941 10836 19975
rect 10784 19932 10836 19941
rect 18420 19975 18472 19984
rect 18420 19941 18429 19975
rect 18429 19941 18463 19975
rect 18463 19941 18472 19975
rect 18420 19932 18472 19941
rect 18512 19975 18564 19984
rect 18512 19941 18521 19975
rect 18521 19941 18555 19975
rect 18555 19941 18564 19975
rect 18512 19932 18564 19941
rect 4804 19796 4856 19848
rect 5540 19839 5592 19848
rect 5540 19805 5549 19839
rect 5549 19805 5583 19839
rect 5583 19805 5592 19839
rect 5540 19796 5592 19805
rect 7840 19839 7892 19848
rect 7840 19805 7849 19839
rect 7849 19805 7883 19839
rect 7883 19805 7892 19839
rect 7840 19796 7892 19805
rect 11336 19839 11388 19848
rect 10600 19728 10652 19780
rect 11336 19805 11345 19839
rect 11345 19805 11379 19839
rect 11379 19805 11388 19839
rect 11336 19796 11388 19805
rect 11704 19796 11756 19848
rect 19248 19796 19300 19848
rect 9956 19703 10008 19712
rect 9956 19669 9965 19703
rect 9965 19669 9999 19703
rect 9999 19669 10008 19703
rect 9956 19660 10008 19669
rect 18052 19703 18104 19712
rect 18052 19669 18061 19703
rect 18061 19669 18095 19703
rect 18095 19669 18104 19703
rect 18052 19660 18104 19669
rect 4982 19558 5034 19610
rect 5046 19558 5098 19610
rect 5110 19558 5162 19610
rect 5174 19558 5226 19610
rect 12982 19558 13034 19610
rect 13046 19558 13098 19610
rect 13110 19558 13162 19610
rect 13174 19558 13226 19610
rect 20982 19558 21034 19610
rect 21046 19558 21098 19610
rect 21110 19558 21162 19610
rect 21174 19558 21226 19610
rect 4804 19456 4856 19508
rect 10784 19456 10836 19508
rect 18512 19456 18564 19508
rect 21272 19456 21324 19508
rect 5356 19388 5408 19440
rect 9956 19363 10008 19372
rect 7656 19295 7708 19304
rect 7656 19261 7665 19295
rect 7665 19261 7699 19295
rect 7699 19261 7708 19295
rect 7656 19252 7708 19261
rect 9956 19329 9965 19363
rect 9965 19329 9999 19363
rect 9999 19329 10008 19363
rect 9956 19320 10008 19329
rect 8576 19252 8628 19304
rect 16672 19295 16724 19304
rect 16672 19261 16681 19295
rect 16681 19261 16715 19295
rect 16715 19261 16724 19295
rect 16672 19252 16724 19261
rect 3608 19159 3660 19168
rect 3608 19125 3617 19159
rect 3617 19125 3651 19159
rect 3651 19125 3660 19159
rect 3608 19116 3660 19125
rect 4160 19116 4212 19168
rect 7840 19116 7892 19168
rect 8668 19159 8720 19168
rect 8668 19125 8677 19159
rect 8677 19125 8711 19159
rect 8711 19125 8720 19159
rect 17316 19252 17368 19304
rect 18052 19295 18104 19304
rect 18052 19261 18061 19295
rect 18061 19261 18095 19295
rect 18095 19261 18104 19295
rect 18052 19252 18104 19261
rect 21456 19252 21508 19304
rect 17408 19184 17460 19236
rect 8668 19116 8720 19125
rect 10600 19116 10652 19168
rect 16212 19159 16264 19168
rect 16212 19125 16221 19159
rect 16221 19125 16255 19159
rect 16255 19125 16264 19159
rect 16212 19116 16264 19125
rect 17776 19159 17828 19168
rect 17776 19125 17785 19159
rect 17785 19125 17819 19159
rect 17819 19125 17828 19159
rect 17776 19116 17828 19125
rect 8982 19014 9034 19066
rect 9046 19014 9098 19066
rect 9110 19014 9162 19066
rect 9174 19014 9226 19066
rect 16982 19014 17034 19066
rect 17046 19014 17098 19066
rect 17110 19014 17162 19066
rect 17174 19014 17226 19066
rect 1584 18955 1636 18964
rect 1584 18921 1593 18955
rect 1593 18921 1627 18955
rect 1627 18921 1636 18955
rect 1584 18912 1636 18921
rect 6460 18955 6512 18964
rect 6460 18921 6469 18955
rect 6469 18921 6503 18955
rect 6503 18921 6512 18955
rect 6460 18912 6512 18921
rect 9956 18955 10008 18964
rect 9956 18921 9965 18955
rect 9965 18921 9999 18955
rect 9999 18921 10008 18955
rect 9956 18912 10008 18921
rect 18420 18955 18472 18964
rect 18420 18921 18429 18955
rect 18429 18921 18463 18955
rect 18463 18921 18472 18955
rect 18420 18912 18472 18921
rect 4712 18844 4764 18896
rect 11520 18887 11572 18896
rect 11520 18853 11529 18887
rect 11529 18853 11563 18887
rect 11563 18853 11572 18887
rect 11520 18844 11572 18853
rect 17316 18887 17368 18896
rect 17316 18853 17325 18887
rect 17325 18853 17359 18887
rect 17359 18853 17368 18887
rect 17316 18844 17368 18853
rect 18788 18887 18840 18896
rect 18788 18853 18797 18887
rect 18797 18853 18831 18887
rect 18831 18853 18840 18887
rect 18788 18844 18840 18853
rect 1400 18819 1452 18828
rect 1400 18785 1409 18819
rect 1409 18785 1443 18819
rect 1443 18785 1452 18819
rect 1400 18776 1452 18785
rect 5540 18751 5592 18760
rect 5540 18717 5549 18751
rect 5549 18717 5583 18751
rect 5583 18717 5592 18751
rect 5540 18708 5592 18717
rect 6092 18708 6144 18760
rect 6736 18776 6788 18828
rect 8300 18819 8352 18828
rect 8300 18785 8309 18819
rect 8309 18785 8343 18819
rect 8343 18785 8352 18819
rect 8300 18776 8352 18785
rect 8576 18819 8628 18828
rect 8576 18785 8585 18819
rect 8585 18785 8619 18819
rect 8619 18785 8628 18819
rect 8576 18776 8628 18785
rect 10140 18819 10192 18828
rect 8760 18751 8812 18760
rect 8760 18717 8769 18751
rect 8769 18717 8803 18751
rect 8803 18717 8812 18751
rect 8760 18708 8812 18717
rect 10140 18785 10149 18819
rect 10149 18785 10183 18819
rect 10183 18785 10192 18819
rect 10140 18776 10192 18785
rect 15200 18819 15252 18828
rect 15200 18785 15209 18819
rect 15209 18785 15243 18819
rect 15243 18785 15252 18819
rect 15200 18776 15252 18785
rect 16856 18819 16908 18828
rect 16856 18785 16865 18819
rect 16865 18785 16899 18819
rect 16899 18785 16908 18819
rect 16856 18776 16908 18785
rect 17040 18819 17092 18828
rect 17040 18785 17049 18819
rect 17049 18785 17083 18819
rect 17083 18785 17092 18819
rect 17040 18776 17092 18785
rect 10416 18708 10468 18760
rect 11428 18751 11480 18760
rect 11428 18717 11437 18751
rect 11437 18717 11471 18751
rect 11471 18717 11480 18751
rect 11428 18708 11480 18717
rect 11704 18751 11756 18760
rect 11704 18717 11713 18751
rect 11713 18717 11747 18751
rect 11747 18717 11756 18751
rect 11704 18708 11756 18717
rect 18696 18751 18748 18760
rect 18696 18717 18705 18751
rect 18705 18717 18739 18751
rect 18739 18717 18748 18751
rect 18696 18708 18748 18717
rect 5448 18640 5500 18692
rect 19248 18683 19300 18692
rect 19248 18649 19257 18683
rect 19257 18649 19291 18683
rect 19291 18649 19300 18683
rect 19248 18640 19300 18649
rect 3516 18572 3568 18624
rect 7656 18615 7708 18624
rect 7656 18581 7665 18615
rect 7665 18581 7699 18615
rect 7699 18581 7708 18615
rect 7656 18572 7708 18581
rect 10784 18615 10836 18624
rect 10784 18581 10793 18615
rect 10793 18581 10827 18615
rect 10827 18581 10836 18615
rect 10784 18572 10836 18581
rect 12532 18615 12584 18624
rect 12532 18581 12541 18615
rect 12541 18581 12575 18615
rect 12575 18581 12584 18615
rect 12532 18572 12584 18581
rect 15568 18572 15620 18624
rect 16672 18572 16724 18624
rect 4982 18470 5034 18522
rect 5046 18470 5098 18522
rect 5110 18470 5162 18522
rect 5174 18470 5226 18522
rect 12982 18470 13034 18522
rect 13046 18470 13098 18522
rect 13110 18470 13162 18522
rect 13174 18470 13226 18522
rect 20982 18470 21034 18522
rect 21046 18470 21098 18522
rect 21110 18470 21162 18522
rect 21174 18470 21226 18522
rect 1400 18368 1452 18420
rect 4712 18411 4764 18420
rect 4712 18377 4721 18411
rect 4721 18377 4755 18411
rect 4755 18377 4764 18411
rect 4712 18368 4764 18377
rect 6092 18411 6144 18420
rect 5540 18343 5592 18352
rect 5540 18309 5549 18343
rect 5549 18309 5583 18343
rect 5583 18309 5592 18343
rect 5540 18300 5592 18309
rect 6092 18377 6101 18411
rect 6101 18377 6135 18411
rect 6135 18377 6144 18411
rect 6092 18368 6144 18377
rect 17408 18411 17460 18420
rect 17408 18377 17417 18411
rect 17417 18377 17451 18411
rect 17451 18377 17460 18411
rect 17408 18368 17460 18377
rect 18788 18368 18840 18420
rect 8208 18300 8260 18352
rect 10048 18300 10100 18352
rect 10784 18300 10836 18352
rect 11520 18300 11572 18352
rect 14188 18300 14240 18352
rect 16212 18300 16264 18352
rect 17040 18300 17092 18352
rect 3516 18207 3568 18216
rect 3516 18173 3525 18207
rect 3525 18173 3559 18207
rect 3559 18173 3568 18207
rect 3516 18164 3568 18173
rect 6736 18232 6788 18284
rect 7012 18232 7064 18284
rect 8760 18232 8812 18284
rect 11428 18232 11480 18284
rect 11796 18232 11848 18284
rect 15200 18232 15252 18284
rect 4988 18139 5040 18148
rect 2872 18028 2924 18080
rect 4988 18105 4997 18139
rect 4997 18105 5031 18139
rect 5031 18105 5040 18139
rect 4988 18096 5040 18105
rect 6920 18139 6972 18148
rect 3608 18071 3660 18080
rect 3608 18037 3617 18071
rect 3617 18037 3651 18071
rect 3651 18037 3660 18071
rect 3608 18028 3660 18037
rect 4804 18028 4856 18080
rect 6920 18105 6929 18139
rect 6929 18105 6963 18139
rect 6963 18105 6972 18139
rect 6920 18096 6972 18105
rect 7104 18096 7156 18148
rect 8576 18164 8628 18216
rect 10140 18164 10192 18216
rect 12532 18164 12584 18216
rect 19800 18207 19852 18216
rect 10692 18139 10744 18148
rect 10692 18105 10701 18139
rect 10701 18105 10735 18139
rect 10735 18105 10744 18139
rect 10692 18096 10744 18105
rect 10784 18139 10836 18148
rect 10784 18105 10793 18139
rect 10793 18105 10827 18139
rect 10827 18105 10836 18139
rect 15016 18139 15068 18148
rect 10784 18096 10836 18105
rect 15016 18105 15025 18139
rect 15025 18105 15059 18139
rect 15059 18105 15068 18139
rect 15016 18096 15068 18105
rect 8116 18071 8168 18080
rect 8116 18037 8125 18071
rect 8125 18037 8159 18071
rect 8159 18037 8168 18071
rect 8116 18028 8168 18037
rect 8668 18071 8720 18080
rect 8668 18037 8677 18071
rect 8677 18037 8711 18071
rect 8711 18037 8720 18071
rect 8668 18028 8720 18037
rect 10416 18071 10468 18080
rect 10416 18037 10425 18071
rect 10425 18037 10459 18071
rect 10459 18037 10468 18071
rect 10416 18028 10468 18037
rect 12624 18028 12676 18080
rect 12808 18071 12860 18080
rect 12808 18037 12817 18071
rect 12817 18037 12851 18071
rect 12851 18037 12860 18071
rect 12808 18028 12860 18037
rect 16028 18096 16080 18148
rect 19800 18173 19809 18207
rect 19809 18173 19843 18207
rect 19843 18173 19852 18207
rect 19800 18164 19852 18173
rect 15752 18028 15804 18080
rect 16212 18028 16264 18080
rect 16856 18028 16908 18080
rect 17776 18071 17828 18080
rect 17776 18037 17785 18071
rect 17785 18037 17819 18071
rect 17819 18037 17828 18071
rect 17776 18028 17828 18037
rect 18512 18028 18564 18080
rect 19892 18071 19944 18080
rect 19892 18037 19901 18071
rect 19901 18037 19935 18071
rect 19935 18037 19944 18071
rect 19892 18028 19944 18037
rect 8982 17926 9034 17978
rect 9046 17926 9098 17978
rect 9110 17926 9162 17978
rect 9174 17926 9226 17978
rect 16982 17926 17034 17978
rect 17046 17926 17098 17978
rect 17110 17926 17162 17978
rect 17174 17926 17226 17978
rect 4712 17824 4764 17876
rect 6920 17824 6972 17876
rect 8760 17824 8812 17876
rect 11428 17867 11480 17876
rect 11428 17833 11437 17867
rect 11437 17833 11471 17867
rect 11471 17833 11480 17867
rect 11428 17824 11480 17833
rect 15016 17867 15068 17876
rect 15016 17833 15025 17867
rect 15025 17833 15059 17867
rect 15059 17833 15068 17867
rect 15016 17824 15068 17833
rect 16212 17867 16264 17876
rect 16212 17833 16221 17867
rect 16221 17833 16255 17867
rect 16255 17833 16264 17867
rect 16212 17824 16264 17833
rect 18696 17824 18748 17876
rect 21272 17824 21324 17876
rect 4160 17756 4212 17808
rect 6736 17799 6788 17808
rect 6736 17765 6745 17799
rect 6745 17765 6779 17799
rect 6779 17765 6788 17799
rect 6736 17756 6788 17765
rect 8668 17756 8720 17808
rect 10048 17799 10100 17808
rect 10048 17765 10057 17799
rect 10057 17765 10091 17799
rect 10091 17765 10100 17799
rect 10048 17756 10100 17765
rect 12532 17799 12584 17808
rect 12532 17765 12541 17799
rect 12541 17765 12575 17799
rect 12575 17765 12584 17799
rect 12532 17756 12584 17765
rect 15292 17756 15344 17808
rect 17776 17756 17828 17808
rect 18512 17756 18564 17808
rect 2596 17731 2648 17740
rect 2596 17697 2605 17731
rect 2605 17697 2639 17731
rect 2639 17697 2648 17731
rect 2596 17688 2648 17697
rect 2872 17731 2924 17740
rect 2872 17697 2881 17731
rect 2881 17697 2915 17731
rect 2915 17697 2924 17731
rect 2872 17688 2924 17697
rect 4712 17688 4764 17740
rect 4988 17688 5040 17740
rect 6460 17731 6512 17740
rect 6460 17697 6469 17731
rect 6469 17697 6503 17731
rect 6503 17697 6512 17731
rect 6460 17688 6512 17697
rect 8484 17688 8536 17740
rect 11888 17731 11940 17740
rect 11888 17697 11897 17731
rect 11897 17697 11931 17731
rect 11931 17697 11940 17731
rect 11888 17688 11940 17697
rect 12256 17731 12308 17740
rect 12256 17697 12265 17731
rect 12265 17697 12299 17731
rect 12299 17697 12308 17731
rect 12256 17688 12308 17697
rect 14004 17688 14056 17740
rect 14188 17731 14240 17740
rect 14188 17697 14197 17731
rect 14197 17697 14231 17731
rect 14231 17697 14240 17731
rect 14188 17688 14240 17697
rect 17132 17688 17184 17740
rect 17868 17688 17920 17740
rect 19892 17688 19944 17740
rect 20720 17688 20772 17740
rect 3148 17663 3200 17672
rect 3148 17629 3157 17663
rect 3157 17629 3191 17663
rect 3191 17629 3200 17663
rect 3148 17620 3200 17629
rect 11152 17620 11204 17672
rect 10600 17552 10652 17604
rect 13268 17595 13320 17604
rect 13268 17561 13277 17595
rect 13277 17561 13311 17595
rect 13311 17561 13320 17595
rect 13268 17552 13320 17561
rect 16488 17620 16540 17672
rect 18052 17552 18104 17604
rect 19800 17595 19852 17604
rect 19800 17561 19809 17595
rect 19809 17561 19843 17595
rect 19843 17561 19852 17595
rect 19800 17552 19852 17561
rect 5448 17484 5500 17536
rect 7012 17484 7064 17536
rect 7104 17484 7156 17536
rect 8300 17484 8352 17536
rect 9588 17484 9640 17536
rect 10692 17484 10744 17536
rect 12808 17527 12860 17536
rect 12808 17493 12817 17527
rect 12817 17493 12851 17527
rect 12851 17493 12860 17527
rect 12808 17484 12860 17493
rect 16580 17484 16632 17536
rect 19064 17527 19116 17536
rect 19064 17493 19073 17527
rect 19073 17493 19107 17527
rect 19107 17493 19116 17527
rect 19064 17484 19116 17493
rect 4982 17382 5034 17434
rect 5046 17382 5098 17434
rect 5110 17382 5162 17434
rect 5174 17382 5226 17434
rect 12982 17382 13034 17434
rect 13046 17382 13098 17434
rect 13110 17382 13162 17434
rect 13174 17382 13226 17434
rect 20982 17382 21034 17434
rect 21046 17382 21098 17434
rect 21110 17382 21162 17434
rect 21174 17382 21226 17434
rect 3148 17323 3200 17332
rect 3148 17289 3157 17323
rect 3157 17289 3191 17323
rect 3191 17289 3200 17323
rect 3148 17280 3200 17289
rect 4804 17280 4856 17332
rect 6460 17280 6512 17332
rect 8208 17323 8260 17332
rect 8208 17289 8217 17323
rect 8217 17289 8251 17323
rect 8251 17289 8260 17323
rect 8208 17280 8260 17289
rect 8484 17280 8536 17332
rect 9588 17280 9640 17332
rect 10048 17280 10100 17332
rect 11152 17323 11204 17332
rect 11152 17289 11161 17323
rect 11161 17289 11195 17323
rect 11195 17289 11204 17323
rect 11152 17280 11204 17289
rect 15016 17280 15068 17332
rect 16488 17323 16540 17332
rect 16488 17289 16497 17323
rect 16497 17289 16531 17323
rect 16531 17289 16540 17323
rect 16488 17280 16540 17289
rect 17868 17323 17920 17332
rect 17868 17289 17877 17323
rect 17877 17289 17911 17323
rect 17911 17289 17920 17323
rect 17868 17280 17920 17289
rect 21272 17280 21324 17332
rect 2596 17212 2648 17264
rect 10416 17212 10468 17264
rect 10876 17212 10928 17264
rect 10968 17212 11020 17264
rect 13360 17255 13412 17264
rect 7748 17144 7800 17196
rect 9956 17144 10008 17196
rect 13360 17221 13369 17255
rect 13369 17221 13403 17255
rect 13403 17221 13412 17255
rect 13360 17212 13412 17221
rect 15108 17212 15160 17264
rect 17132 17255 17184 17264
rect 17132 17221 17141 17255
rect 17141 17221 17175 17255
rect 17175 17221 17184 17255
rect 17132 17212 17184 17221
rect 20536 17212 20588 17264
rect 15568 17187 15620 17196
rect 2872 17008 2924 17060
rect 9312 17076 9364 17128
rect 11796 17119 11848 17128
rect 11796 17085 11805 17119
rect 11805 17085 11839 17119
rect 11839 17085 11848 17119
rect 11796 17076 11848 17085
rect 15568 17153 15577 17187
rect 15577 17153 15611 17187
rect 15611 17153 15620 17187
rect 15568 17144 15620 17153
rect 17776 17144 17828 17196
rect 18972 17144 19024 17196
rect 19248 17187 19300 17196
rect 19248 17153 19257 17187
rect 19257 17153 19291 17187
rect 19291 17153 19300 17187
rect 19248 17144 19300 17153
rect 19524 17076 19576 17128
rect 7104 17008 7156 17060
rect 7288 17008 7340 17060
rect 9496 17008 9548 17060
rect 2596 16940 2648 16992
rect 4160 16940 4212 16992
rect 5264 16983 5316 16992
rect 5264 16949 5273 16983
rect 5273 16949 5307 16983
rect 5307 16949 5316 16983
rect 5264 16940 5316 16949
rect 5816 16940 5868 16992
rect 6736 16940 6788 16992
rect 9312 16983 9364 16992
rect 9312 16949 9321 16983
rect 9321 16949 9355 16983
rect 9355 16949 9364 16983
rect 9312 16940 9364 16949
rect 10600 17008 10652 17060
rect 12440 17008 12492 17060
rect 12808 17051 12860 17060
rect 12808 17017 12817 17051
rect 12817 17017 12851 17051
rect 12851 17017 12860 17051
rect 12808 17008 12860 17017
rect 13268 17008 13320 17060
rect 14004 17008 14056 17060
rect 14188 17008 14240 17060
rect 15752 17008 15804 17060
rect 16212 17051 16264 17060
rect 16212 17017 16221 17051
rect 16221 17017 16255 17051
rect 16255 17017 16264 17051
rect 16212 17008 16264 17017
rect 10140 16940 10192 16992
rect 12256 16983 12308 16992
rect 12256 16949 12265 16983
rect 12265 16949 12299 16983
rect 12299 16949 12308 16983
rect 12256 16940 12308 16949
rect 14096 16983 14148 16992
rect 14096 16949 14105 16983
rect 14105 16949 14139 16983
rect 14139 16949 14148 16983
rect 14096 16940 14148 16949
rect 15292 16983 15344 16992
rect 15292 16949 15301 16983
rect 15301 16949 15335 16983
rect 15335 16949 15344 16983
rect 15292 16940 15344 16949
rect 19064 17008 19116 17060
rect 20720 16983 20772 16992
rect 20720 16949 20729 16983
rect 20729 16949 20763 16983
rect 20763 16949 20772 16983
rect 20720 16940 20772 16949
rect 8982 16838 9034 16890
rect 9046 16838 9098 16890
rect 9110 16838 9162 16890
rect 9174 16838 9226 16890
rect 16982 16838 17034 16890
rect 17046 16838 17098 16890
rect 17110 16838 17162 16890
rect 17174 16838 17226 16890
rect 7104 16779 7156 16788
rect 7104 16745 7113 16779
rect 7113 16745 7147 16779
rect 7147 16745 7156 16779
rect 7104 16736 7156 16745
rect 12716 16779 12768 16788
rect 12716 16745 12725 16779
rect 12725 16745 12759 16779
rect 12759 16745 12768 16779
rect 12716 16736 12768 16745
rect 13268 16779 13320 16788
rect 13268 16745 13277 16779
rect 13277 16745 13311 16779
rect 13311 16745 13320 16779
rect 13268 16736 13320 16745
rect 15568 16736 15620 16788
rect 5264 16668 5316 16720
rect 7748 16668 7800 16720
rect 10140 16711 10192 16720
rect 10140 16677 10149 16711
rect 10149 16677 10183 16711
rect 10183 16677 10192 16711
rect 10140 16668 10192 16677
rect 10968 16668 11020 16720
rect 11428 16668 11480 16720
rect 15844 16711 15896 16720
rect 15844 16677 15853 16711
rect 15853 16677 15887 16711
rect 15887 16677 15896 16711
rect 15844 16668 15896 16677
rect 18328 16711 18380 16720
rect 18328 16677 18337 16711
rect 18337 16677 18371 16711
rect 18371 16677 18380 16711
rect 18328 16668 18380 16677
rect 4252 16643 4304 16652
rect 4252 16609 4261 16643
rect 4261 16609 4295 16643
rect 4295 16609 4304 16643
rect 4252 16600 4304 16609
rect 4620 16643 4672 16652
rect 4620 16609 4629 16643
rect 4629 16609 4663 16643
rect 4663 16609 4672 16643
rect 4620 16600 4672 16609
rect 7932 16600 7984 16652
rect 8392 16600 8444 16652
rect 13912 16600 13964 16652
rect 6368 16575 6420 16584
rect 6368 16541 6377 16575
rect 6377 16541 6411 16575
rect 6411 16541 6420 16575
rect 6368 16532 6420 16541
rect 10048 16575 10100 16584
rect 10048 16541 10057 16575
rect 10057 16541 10091 16575
rect 10091 16541 10100 16575
rect 10048 16532 10100 16541
rect 12348 16575 12400 16584
rect 12348 16541 12357 16575
rect 12357 16541 12391 16575
rect 12391 16541 12400 16575
rect 12348 16532 12400 16541
rect 16580 16532 16632 16584
rect 18236 16575 18288 16584
rect 18236 16541 18245 16575
rect 18245 16541 18279 16575
rect 18279 16541 18288 16575
rect 18236 16532 18288 16541
rect 16212 16464 16264 16516
rect 18696 16464 18748 16516
rect 4436 16396 4488 16448
rect 6184 16396 6236 16448
rect 9036 16439 9088 16448
rect 9036 16405 9045 16439
rect 9045 16405 9079 16439
rect 9079 16405 9088 16439
rect 9036 16396 9088 16405
rect 9496 16439 9548 16448
rect 9496 16405 9505 16439
rect 9505 16405 9539 16439
rect 9539 16405 9548 16439
rect 9496 16396 9548 16405
rect 10508 16396 10560 16448
rect 11796 16439 11848 16448
rect 11796 16405 11805 16439
rect 11805 16405 11839 16439
rect 11839 16405 11848 16439
rect 11796 16396 11848 16405
rect 15200 16396 15252 16448
rect 15752 16396 15804 16448
rect 16028 16396 16080 16448
rect 18972 16464 19024 16516
rect 4982 16294 5034 16346
rect 5046 16294 5098 16346
rect 5110 16294 5162 16346
rect 5174 16294 5226 16346
rect 12982 16294 13034 16346
rect 13046 16294 13098 16346
rect 13110 16294 13162 16346
rect 13174 16294 13226 16346
rect 20982 16294 21034 16346
rect 21046 16294 21098 16346
rect 21110 16294 21162 16346
rect 21174 16294 21226 16346
rect 6184 16235 6236 16244
rect 6184 16201 6193 16235
rect 6193 16201 6227 16235
rect 6227 16201 6236 16235
rect 6184 16192 6236 16201
rect 6368 16192 6420 16244
rect 6736 16192 6788 16244
rect 9312 16192 9364 16244
rect 10140 16192 10192 16244
rect 10324 16192 10376 16244
rect 13820 16192 13872 16244
rect 13912 16192 13964 16244
rect 16580 16192 16632 16244
rect 18236 16192 18288 16244
rect 19248 16192 19300 16244
rect 2872 16124 2924 16176
rect 4620 16124 4672 16176
rect 5356 16124 5408 16176
rect 4436 16099 4488 16108
rect 4436 16065 4445 16099
rect 4445 16065 4479 16099
rect 4479 16065 4488 16099
rect 4436 16056 4488 16065
rect 4712 16099 4764 16108
rect 4712 16065 4721 16099
rect 4721 16065 4755 16099
rect 4755 16065 4764 16099
rect 7288 16124 7340 16176
rect 7656 16124 7708 16176
rect 10968 16167 11020 16176
rect 4712 16056 4764 16065
rect 3792 15988 3844 16040
rect 8668 16056 8720 16108
rect 9036 16056 9088 16108
rect 10968 16133 10977 16167
rect 10977 16133 11011 16167
rect 11011 16133 11020 16167
rect 10968 16124 11020 16133
rect 18696 16167 18748 16176
rect 18696 16133 18705 16167
rect 18705 16133 18739 16167
rect 18739 16133 18748 16167
rect 18696 16124 18748 16133
rect 12716 16056 12768 16108
rect 12532 15988 12584 16040
rect 13268 15988 13320 16040
rect 4252 15920 4304 15972
rect 4528 15963 4580 15972
rect 4528 15929 4537 15963
rect 4537 15929 4571 15963
rect 4571 15929 4580 15963
rect 4528 15920 4580 15929
rect 7012 15963 7064 15972
rect 7012 15929 7021 15963
rect 7021 15929 7055 15963
rect 7055 15929 7064 15963
rect 7012 15920 7064 15929
rect 8760 15920 8812 15972
rect 10416 15963 10468 15972
rect 10416 15929 10425 15963
rect 10425 15929 10459 15963
rect 10459 15929 10468 15963
rect 10416 15920 10468 15929
rect 10508 15963 10560 15972
rect 10508 15929 10517 15963
rect 10517 15929 10551 15963
rect 10551 15929 10560 15963
rect 10508 15920 10560 15929
rect 14832 16031 14884 16040
rect 14832 15997 14841 16031
rect 14841 15997 14875 16031
rect 14875 15997 14884 16031
rect 14832 15988 14884 15997
rect 15292 15920 15344 15972
rect 3792 15895 3844 15904
rect 3792 15861 3801 15895
rect 3801 15861 3835 15895
rect 3835 15861 3844 15895
rect 3792 15852 3844 15861
rect 4988 15852 5040 15904
rect 7932 15895 7984 15904
rect 7932 15861 7941 15895
rect 7941 15861 7975 15895
rect 7975 15861 7984 15895
rect 7932 15852 7984 15861
rect 8392 15895 8444 15904
rect 8392 15861 8401 15895
rect 8401 15861 8435 15895
rect 8435 15861 8444 15895
rect 8392 15852 8444 15861
rect 11612 15852 11664 15904
rect 12348 15852 12400 15904
rect 15384 15852 15436 15904
rect 15844 15852 15896 15904
rect 18328 15920 18380 15972
rect 18144 15852 18196 15904
rect 19524 15852 19576 15904
rect 19984 15895 20036 15904
rect 19984 15861 19993 15895
rect 19993 15861 20027 15895
rect 20027 15861 20036 15895
rect 19984 15852 20036 15861
rect 8982 15750 9034 15802
rect 9046 15750 9098 15802
rect 9110 15750 9162 15802
rect 9174 15750 9226 15802
rect 16982 15750 17034 15802
rect 17046 15750 17098 15802
rect 17110 15750 17162 15802
rect 17174 15750 17226 15802
rect 4160 15648 4212 15700
rect 2780 15580 2832 15632
rect 4528 15648 4580 15700
rect 4988 15691 5040 15700
rect 4988 15657 4997 15691
rect 4997 15657 5031 15691
rect 5031 15657 5040 15691
rect 4988 15648 5040 15657
rect 7012 15691 7064 15700
rect 7012 15657 7021 15691
rect 7021 15657 7055 15691
rect 7055 15657 7064 15691
rect 7012 15648 7064 15657
rect 8760 15648 8812 15700
rect 10048 15691 10100 15700
rect 2872 15555 2924 15564
rect 2872 15521 2881 15555
rect 2881 15521 2915 15555
rect 2915 15521 2924 15555
rect 2872 15512 2924 15521
rect 5816 15580 5868 15632
rect 8668 15623 8720 15632
rect 8668 15589 8677 15623
rect 8677 15589 8711 15623
rect 8711 15589 8720 15623
rect 8668 15580 8720 15589
rect 5908 15512 5960 15564
rect 8300 15512 8352 15564
rect 10048 15657 10057 15691
rect 10057 15657 10091 15691
rect 10091 15657 10100 15691
rect 10048 15648 10100 15657
rect 12440 15691 12492 15700
rect 12440 15657 12449 15691
rect 12449 15657 12483 15691
rect 12483 15657 12492 15691
rect 12440 15648 12492 15657
rect 18328 15648 18380 15700
rect 10508 15580 10560 15632
rect 14832 15623 14884 15632
rect 14832 15589 14841 15623
rect 14841 15589 14875 15623
rect 14875 15589 14884 15623
rect 14832 15580 14884 15589
rect 15384 15580 15436 15632
rect 16028 15623 16080 15632
rect 16028 15589 16037 15623
rect 16037 15589 16071 15623
rect 16071 15589 16080 15623
rect 16028 15580 16080 15589
rect 17408 15580 17460 15632
rect 18972 15580 19024 15632
rect 19248 15623 19300 15632
rect 19248 15589 19257 15623
rect 19257 15589 19291 15623
rect 19291 15589 19300 15623
rect 19248 15580 19300 15589
rect 3148 15487 3200 15496
rect 3148 15453 3157 15487
rect 3157 15453 3191 15487
rect 3191 15453 3200 15487
rect 3148 15444 3200 15453
rect 6000 15444 6052 15496
rect 8116 15444 8168 15496
rect 10048 15512 10100 15564
rect 13820 15555 13872 15564
rect 13820 15521 13829 15555
rect 13829 15521 13863 15555
rect 13863 15521 13872 15555
rect 14096 15555 14148 15564
rect 13820 15512 13872 15521
rect 14096 15521 14105 15555
rect 14105 15521 14139 15555
rect 14139 15521 14148 15555
rect 14096 15512 14148 15521
rect 18696 15512 18748 15564
rect 21640 15512 21692 15564
rect 23572 15512 23624 15564
rect 9772 15444 9824 15496
rect 10600 15487 10652 15496
rect 10600 15453 10609 15487
rect 10609 15453 10643 15487
rect 10643 15453 10652 15487
rect 10600 15444 10652 15453
rect 15200 15444 15252 15496
rect 17316 15487 17368 15496
rect 17316 15453 17325 15487
rect 17325 15453 17359 15487
rect 17359 15453 17368 15487
rect 17316 15444 17368 15453
rect 13268 15376 13320 15428
rect 7380 15351 7432 15360
rect 7380 15317 7389 15351
rect 7389 15317 7423 15351
rect 7423 15317 7432 15351
rect 7380 15308 7432 15317
rect 10416 15308 10468 15360
rect 16396 15351 16448 15360
rect 16396 15317 16405 15351
rect 16405 15317 16439 15351
rect 16439 15317 16448 15351
rect 16396 15308 16448 15317
rect 4982 15206 5034 15258
rect 5046 15206 5098 15258
rect 5110 15206 5162 15258
rect 5174 15206 5226 15258
rect 12982 15206 13034 15258
rect 13046 15206 13098 15258
rect 13110 15206 13162 15258
rect 13174 15206 13226 15258
rect 20982 15206 21034 15258
rect 21046 15206 21098 15258
rect 21110 15206 21162 15258
rect 21174 15206 21226 15258
rect 2780 15147 2832 15156
rect 2780 15113 2789 15147
rect 2789 15113 2823 15147
rect 2823 15113 2832 15147
rect 2780 15104 2832 15113
rect 3148 15147 3200 15156
rect 3148 15113 3157 15147
rect 3157 15113 3191 15147
rect 3191 15113 3200 15147
rect 3148 15104 3200 15113
rect 4160 15104 4212 15156
rect 5816 15147 5868 15156
rect 5816 15113 5825 15147
rect 5825 15113 5859 15147
rect 5859 15113 5868 15147
rect 5816 15104 5868 15113
rect 7012 15104 7064 15156
rect 9772 15147 9824 15156
rect 9772 15113 9781 15147
rect 9781 15113 9815 15147
rect 9815 15113 9824 15147
rect 9772 15104 9824 15113
rect 10416 15104 10468 15156
rect 10508 15104 10560 15156
rect 14096 15104 14148 15156
rect 15016 15104 15068 15156
rect 15384 15147 15436 15156
rect 15384 15113 15393 15147
rect 15393 15113 15427 15147
rect 15427 15113 15436 15147
rect 15384 15104 15436 15113
rect 18696 15147 18748 15156
rect 18696 15113 18705 15147
rect 18705 15113 18739 15147
rect 18739 15113 18748 15147
rect 18696 15104 18748 15113
rect 19984 15104 20036 15156
rect 2872 15036 2924 15088
rect 5448 15036 5500 15088
rect 9496 15036 9548 15088
rect 7380 14968 7432 15020
rect 7932 14968 7984 15020
rect 3056 14900 3108 14952
rect 8760 14900 8812 14952
rect 9312 14943 9364 14952
rect 9312 14909 9321 14943
rect 9321 14909 9355 14943
rect 9355 14909 9364 14943
rect 9312 14900 9364 14909
rect 10416 14943 10468 14952
rect 10416 14909 10425 14943
rect 10425 14909 10459 14943
rect 10459 14909 10468 14943
rect 10416 14900 10468 14909
rect 15108 15036 15160 15088
rect 15200 15036 15252 15088
rect 14556 15011 14608 15020
rect 14556 14977 14565 15011
rect 14565 14977 14599 15011
rect 14599 14977 14608 15011
rect 14556 14968 14608 14977
rect 15016 14968 15068 15020
rect 15568 14900 15620 14952
rect 16396 14943 16448 14952
rect 16396 14909 16405 14943
rect 16405 14909 16439 14943
rect 16439 14909 16448 14943
rect 16396 14900 16448 14909
rect 17316 14968 17368 15020
rect 21272 15036 21324 15088
rect 21456 14968 21508 15020
rect 3516 14832 3568 14884
rect 4528 14875 4580 14884
rect 4528 14841 4537 14875
rect 4537 14841 4571 14875
rect 4571 14841 4580 14875
rect 4528 14832 4580 14841
rect 7012 14875 7064 14884
rect 7012 14841 7021 14875
rect 7021 14841 7055 14875
rect 7055 14841 7064 14875
rect 7012 14832 7064 14841
rect 12532 14875 12584 14884
rect 12532 14841 12541 14875
rect 12541 14841 12575 14875
rect 12575 14841 12584 14875
rect 12532 14832 12584 14841
rect 4160 14807 4212 14816
rect 4160 14773 4169 14807
rect 4169 14773 4203 14807
rect 4203 14773 4212 14807
rect 4160 14764 4212 14773
rect 6000 14764 6052 14816
rect 8116 14764 8168 14816
rect 8300 14807 8352 14816
rect 8300 14773 8309 14807
rect 8309 14773 8343 14807
rect 8343 14773 8352 14807
rect 8300 14764 8352 14773
rect 12164 14807 12216 14816
rect 12164 14773 12173 14807
rect 12173 14773 12207 14807
rect 12207 14773 12216 14807
rect 13360 14832 13412 14884
rect 14096 14832 14148 14884
rect 12164 14764 12216 14773
rect 13820 14764 13872 14816
rect 14372 14875 14424 14884
rect 14372 14841 14381 14875
rect 14381 14841 14415 14875
rect 14415 14841 14424 14875
rect 14372 14832 14424 14841
rect 18972 14832 19024 14884
rect 14464 14764 14516 14816
rect 16304 14764 16356 14816
rect 17408 14807 17460 14816
rect 17408 14773 17417 14807
rect 17417 14773 17451 14807
rect 17451 14773 17460 14807
rect 17408 14764 17460 14773
rect 18328 14807 18380 14816
rect 18328 14773 18337 14807
rect 18337 14773 18371 14807
rect 18371 14773 18380 14807
rect 18328 14764 18380 14773
rect 20628 14764 20680 14816
rect 8982 14662 9034 14714
rect 9046 14662 9098 14714
rect 9110 14662 9162 14714
rect 9174 14662 9226 14714
rect 16982 14662 17034 14714
rect 17046 14662 17098 14714
rect 17110 14662 17162 14714
rect 17174 14662 17226 14714
rect 1124 14560 1176 14612
rect 4528 14603 4580 14612
rect 4528 14569 4537 14603
rect 4537 14569 4571 14603
rect 4571 14569 4580 14603
rect 4528 14560 4580 14569
rect 7380 14560 7432 14612
rect 10048 14603 10100 14612
rect 10048 14569 10057 14603
rect 10057 14569 10091 14603
rect 10091 14569 10100 14603
rect 10048 14560 10100 14569
rect 10508 14560 10560 14612
rect 10876 14603 10928 14612
rect 10876 14569 10885 14603
rect 10885 14569 10919 14603
rect 10919 14569 10928 14603
rect 10876 14560 10928 14569
rect 16672 14560 16724 14612
rect 20628 14603 20680 14612
rect 6000 14535 6052 14544
rect 6000 14501 6009 14535
rect 6009 14501 6043 14535
rect 6043 14501 6052 14535
rect 6000 14492 6052 14501
rect 11612 14492 11664 14544
rect 18328 14492 18380 14544
rect 20628 14569 20637 14603
rect 20637 14569 20671 14603
rect 20671 14569 20680 14603
rect 20628 14560 20680 14569
rect 22284 14560 22336 14612
rect 2044 14424 2096 14476
rect 4068 14288 4120 14340
rect 5356 14424 5408 14476
rect 7012 14424 7064 14476
rect 7196 14424 7248 14476
rect 13268 14424 13320 14476
rect 13636 14467 13688 14476
rect 5540 14356 5592 14408
rect 9680 14399 9732 14408
rect 9680 14365 9689 14399
rect 9689 14365 9723 14399
rect 9723 14365 9732 14399
rect 9680 14356 9732 14365
rect 11980 14356 12032 14408
rect 13636 14433 13645 14467
rect 13645 14433 13679 14467
rect 13679 14433 13688 14467
rect 13636 14424 13688 14433
rect 15200 14424 15252 14476
rect 15568 14467 15620 14476
rect 15568 14433 15577 14467
rect 15577 14433 15611 14467
rect 15611 14433 15620 14467
rect 15568 14424 15620 14433
rect 16396 14424 16448 14476
rect 16856 14424 16908 14476
rect 17316 14424 17368 14476
rect 17592 14467 17644 14476
rect 17592 14433 17601 14467
rect 17601 14433 17635 14467
rect 17635 14433 17644 14467
rect 17592 14424 17644 14433
rect 18972 14467 19024 14476
rect 18972 14433 18981 14467
rect 18981 14433 19015 14467
rect 19015 14433 19024 14467
rect 18972 14424 19024 14433
rect 19064 14424 19116 14476
rect 20812 14424 20864 14476
rect 13728 14399 13780 14408
rect 8392 14288 8444 14340
rect 13728 14365 13737 14399
rect 13737 14365 13771 14399
rect 13771 14365 13780 14399
rect 13728 14356 13780 14365
rect 16120 14399 16172 14408
rect 16120 14365 16129 14399
rect 16129 14365 16163 14399
rect 16163 14365 16172 14399
rect 16120 14356 16172 14365
rect 19248 14399 19300 14408
rect 19248 14365 19257 14399
rect 19257 14365 19291 14399
rect 19291 14365 19300 14399
rect 19248 14356 19300 14365
rect 14004 14288 14056 14340
rect 4344 14220 4396 14272
rect 7564 14220 7616 14272
rect 7656 14220 7708 14272
rect 12348 14263 12400 14272
rect 12348 14229 12357 14263
rect 12357 14229 12391 14263
rect 12391 14229 12400 14263
rect 12348 14220 12400 14229
rect 14280 14263 14332 14272
rect 14280 14229 14289 14263
rect 14289 14229 14323 14263
rect 14323 14229 14332 14263
rect 14280 14220 14332 14229
rect 14464 14220 14516 14272
rect 20168 14263 20220 14272
rect 20168 14229 20177 14263
rect 20177 14229 20211 14263
rect 20211 14229 20220 14263
rect 20168 14220 20220 14229
rect 4982 14118 5034 14170
rect 5046 14118 5098 14170
rect 5110 14118 5162 14170
rect 5174 14118 5226 14170
rect 12982 14118 13034 14170
rect 13046 14118 13098 14170
rect 13110 14118 13162 14170
rect 13174 14118 13226 14170
rect 20982 14118 21034 14170
rect 21046 14118 21098 14170
rect 21110 14118 21162 14170
rect 21174 14118 21226 14170
rect 112 14016 164 14068
rect 4068 14059 4120 14068
rect 4068 14025 4077 14059
rect 4077 14025 4111 14059
rect 4111 14025 4120 14059
rect 4068 14016 4120 14025
rect 7196 14016 7248 14068
rect 11612 14016 11664 14068
rect 4436 13948 4488 14000
rect 8760 13948 8812 14000
rect 4344 13880 4396 13932
rect 7472 13923 7524 13932
rect 7472 13889 7481 13923
rect 7481 13889 7515 13923
rect 7515 13889 7524 13923
rect 7472 13880 7524 13889
rect 7656 13880 7708 13932
rect 8116 13880 8168 13932
rect 12256 13948 12308 14000
rect 14464 14016 14516 14068
rect 19064 14059 19116 14068
rect 19064 14025 19073 14059
rect 19073 14025 19107 14059
rect 19107 14025 19116 14059
rect 19064 14016 19116 14025
rect 14280 13948 14332 14000
rect 15568 13948 15620 14000
rect 18972 13948 19024 14000
rect 20812 13948 20864 14000
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 5540 13812 5592 13864
rect 6552 13812 6604 13864
rect 9312 13812 9364 13864
rect 10048 13855 10100 13864
rect 10048 13821 10057 13855
rect 10057 13821 10091 13855
rect 10091 13821 10100 13855
rect 10048 13812 10100 13821
rect 10784 13855 10836 13864
rect 10784 13821 10793 13855
rect 10793 13821 10827 13855
rect 10827 13821 10836 13855
rect 10784 13812 10836 13821
rect 10876 13812 10928 13864
rect 11336 13880 11388 13932
rect 11612 13855 11664 13864
rect 11612 13821 11621 13855
rect 11621 13821 11655 13855
rect 11655 13821 11664 13855
rect 11612 13812 11664 13821
rect 13728 13880 13780 13932
rect 15752 13923 15804 13932
rect 4620 13744 4672 13796
rect 5356 13787 5408 13796
rect 5356 13753 5365 13787
rect 5365 13753 5399 13787
rect 5399 13753 5408 13787
rect 7564 13787 7616 13796
rect 5356 13744 5408 13753
rect 2044 13719 2096 13728
rect 2044 13685 2053 13719
rect 2053 13685 2087 13719
rect 2087 13685 2096 13719
rect 2044 13676 2096 13685
rect 7012 13719 7064 13728
rect 7012 13685 7021 13719
rect 7021 13685 7055 13719
rect 7055 13685 7064 13719
rect 7012 13676 7064 13685
rect 7564 13753 7573 13787
rect 7573 13753 7607 13787
rect 7607 13753 7616 13787
rect 7564 13744 7616 13753
rect 9680 13787 9732 13796
rect 9680 13753 9689 13787
rect 9689 13753 9723 13787
rect 9723 13753 9732 13787
rect 9680 13744 9732 13753
rect 10876 13719 10928 13728
rect 10876 13685 10885 13719
rect 10885 13685 10919 13719
rect 10919 13685 10928 13719
rect 10876 13676 10928 13685
rect 11428 13676 11480 13728
rect 11980 13719 12032 13728
rect 11980 13685 11989 13719
rect 11989 13685 12023 13719
rect 12023 13685 12032 13719
rect 11980 13676 12032 13685
rect 14832 13744 14884 13796
rect 15108 13744 15160 13796
rect 15752 13889 15761 13923
rect 15761 13889 15795 13923
rect 15795 13889 15804 13923
rect 15752 13880 15804 13889
rect 19800 13880 19852 13932
rect 16764 13812 16816 13864
rect 18052 13855 18104 13864
rect 18052 13821 18061 13855
rect 18061 13821 18095 13855
rect 18095 13821 18104 13855
rect 18052 13812 18104 13821
rect 18420 13812 18472 13864
rect 12624 13676 12676 13728
rect 13636 13676 13688 13728
rect 15200 13676 15252 13728
rect 15384 13676 15436 13728
rect 15568 13787 15620 13796
rect 15568 13753 15577 13787
rect 15577 13753 15611 13787
rect 15611 13753 15620 13787
rect 15568 13744 15620 13753
rect 15936 13676 15988 13728
rect 16396 13719 16448 13728
rect 16396 13685 16405 13719
rect 16405 13685 16439 13719
rect 16439 13685 16448 13719
rect 17592 13744 17644 13796
rect 19064 13812 19116 13864
rect 21180 13812 21232 13864
rect 18788 13787 18840 13796
rect 18788 13753 18797 13787
rect 18797 13753 18831 13787
rect 18831 13753 18840 13787
rect 18788 13744 18840 13753
rect 20168 13787 20220 13796
rect 20168 13753 20177 13787
rect 20177 13753 20211 13787
rect 20211 13753 20220 13787
rect 20168 13744 20220 13753
rect 16396 13676 16448 13685
rect 16856 13676 16908 13728
rect 19984 13719 20036 13728
rect 19984 13685 19993 13719
rect 19993 13685 20027 13719
rect 20027 13685 20036 13719
rect 19984 13676 20036 13685
rect 8982 13574 9034 13626
rect 9046 13574 9098 13626
rect 9110 13574 9162 13626
rect 9174 13574 9226 13626
rect 16982 13574 17034 13626
rect 17046 13574 17098 13626
rect 17110 13574 17162 13626
rect 17174 13574 17226 13626
rect 2780 13404 2832 13456
rect 5540 13472 5592 13524
rect 6828 13515 6880 13524
rect 6828 13481 6837 13515
rect 6837 13481 6871 13515
rect 6871 13481 6880 13515
rect 6828 13472 6880 13481
rect 7472 13472 7524 13524
rect 9312 13472 9364 13524
rect 9680 13472 9732 13524
rect 10876 13472 10928 13524
rect 11612 13515 11664 13524
rect 4252 13404 4304 13456
rect 7012 13404 7064 13456
rect 9956 13404 10008 13456
rect 2596 13268 2648 13320
rect 7564 13336 7616 13388
rect 8484 13336 8536 13388
rect 10324 13336 10376 13388
rect 11612 13481 11621 13515
rect 11621 13481 11655 13515
rect 11655 13481 11664 13515
rect 11612 13472 11664 13481
rect 12164 13515 12216 13524
rect 12164 13481 12173 13515
rect 12173 13481 12207 13515
rect 12207 13481 12216 13515
rect 12164 13472 12216 13481
rect 13728 13472 13780 13524
rect 15568 13515 15620 13524
rect 15568 13481 15577 13515
rect 15577 13481 15611 13515
rect 15611 13481 15620 13515
rect 15568 13472 15620 13481
rect 15936 13515 15988 13524
rect 15936 13481 15945 13515
rect 15945 13481 15979 13515
rect 15979 13481 15988 13515
rect 15936 13472 15988 13481
rect 16856 13472 16908 13524
rect 17316 13515 17368 13524
rect 17316 13481 17325 13515
rect 17325 13481 17359 13515
rect 17359 13481 17368 13515
rect 17316 13472 17368 13481
rect 17684 13472 17736 13524
rect 18604 13472 18656 13524
rect 19984 13515 20036 13524
rect 19984 13481 19993 13515
rect 19993 13481 20027 13515
rect 20027 13481 20036 13515
rect 19984 13472 20036 13481
rect 12348 13404 12400 13456
rect 13452 13404 13504 13456
rect 16304 13404 16356 13456
rect 19064 13404 19116 13456
rect 20812 13404 20864 13456
rect 16120 13379 16172 13388
rect 16120 13345 16129 13379
rect 16129 13345 16163 13379
rect 16163 13345 16172 13379
rect 16120 13336 16172 13345
rect 3148 13311 3200 13320
rect 3148 13277 3157 13311
rect 3157 13277 3191 13311
rect 3191 13277 3200 13311
rect 3148 13268 3200 13277
rect 6184 13268 6236 13320
rect 12808 13268 12860 13320
rect 13360 13311 13412 13320
rect 13360 13277 13369 13311
rect 13369 13277 13403 13311
rect 13403 13277 13412 13311
rect 13360 13268 13412 13277
rect 19248 13268 19300 13320
rect 20260 13268 20312 13320
rect 20720 13268 20772 13320
rect 21180 13268 21232 13320
rect 4528 13200 4580 13252
rect 13912 13200 13964 13252
rect 1400 13132 1452 13184
rect 1676 13175 1728 13184
rect 1676 13141 1685 13175
rect 1685 13141 1719 13175
rect 1719 13141 1728 13175
rect 1676 13132 1728 13141
rect 4620 13132 4672 13184
rect 5448 13132 5500 13184
rect 7472 13132 7524 13184
rect 10784 13175 10836 13184
rect 10784 13141 10793 13175
rect 10793 13141 10827 13175
rect 10827 13141 10836 13175
rect 10784 13132 10836 13141
rect 12440 13175 12492 13184
rect 12440 13141 12449 13175
rect 12449 13141 12483 13175
rect 12483 13141 12492 13175
rect 12440 13132 12492 13141
rect 14004 13175 14056 13184
rect 14004 13141 14013 13175
rect 14013 13141 14047 13175
rect 14047 13141 14056 13175
rect 14004 13132 14056 13141
rect 16580 13132 16632 13184
rect 4982 13030 5034 13082
rect 5046 13030 5098 13082
rect 5110 13030 5162 13082
rect 5174 13030 5226 13082
rect 12982 13030 13034 13082
rect 13046 13030 13098 13082
rect 13110 13030 13162 13082
rect 13174 13030 13226 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 2780 12971 2832 12980
rect 2780 12937 2789 12971
rect 2789 12937 2823 12971
rect 2823 12937 2832 12971
rect 2780 12928 2832 12937
rect 3148 12928 3200 12980
rect 5448 12971 5500 12980
rect 5448 12937 5457 12971
rect 5457 12937 5491 12971
rect 5491 12937 5500 12971
rect 5448 12928 5500 12937
rect 7564 12928 7616 12980
rect 13452 12971 13504 12980
rect 13452 12937 13461 12971
rect 13461 12937 13495 12971
rect 13495 12937 13504 12971
rect 13452 12928 13504 12937
rect 14004 12928 14056 12980
rect 16120 12928 16172 12980
rect 16304 12928 16356 12980
rect 19064 12928 19116 12980
rect 20812 12971 20864 12980
rect 20812 12937 20821 12971
rect 20821 12937 20855 12971
rect 20855 12937 20864 12971
rect 20812 12928 20864 12937
rect 21364 12928 21416 12980
rect 6368 12860 6420 12912
rect 8576 12860 8628 12912
rect 10508 12860 10560 12912
rect 12532 12860 12584 12912
rect 15752 12860 15804 12912
rect 15936 12860 15988 12912
rect 17316 12860 17368 12912
rect 20260 12903 20312 12912
rect 20260 12869 20269 12903
rect 20269 12869 20303 12903
rect 20303 12869 20312 12903
rect 20260 12860 20312 12869
rect 4528 12835 4580 12844
rect 4528 12801 4537 12835
rect 4537 12801 4571 12835
rect 4571 12801 4580 12835
rect 4528 12792 4580 12801
rect 7472 12835 7524 12844
rect 7472 12801 7481 12835
rect 7481 12801 7515 12835
rect 7515 12801 7524 12835
rect 7472 12792 7524 12801
rect 8760 12792 8812 12844
rect 10784 12792 10836 12844
rect 1676 12724 1728 12776
rect 13912 12792 13964 12844
rect 16488 12835 16540 12844
rect 16488 12801 16497 12835
rect 16497 12801 16531 12835
rect 16531 12801 16540 12835
rect 16488 12792 16540 12801
rect 18788 12792 18840 12844
rect 11428 12767 11480 12776
rect 4620 12699 4672 12708
rect 4620 12665 4629 12699
rect 4629 12665 4663 12699
rect 4663 12665 4672 12699
rect 4620 12656 4672 12665
rect 5172 12699 5224 12708
rect 5172 12665 5181 12699
rect 5181 12665 5215 12699
rect 5215 12665 5224 12699
rect 5172 12656 5224 12665
rect 7564 12699 7616 12708
rect 7564 12665 7573 12699
rect 7573 12665 7607 12699
rect 7607 12665 7616 12699
rect 7564 12656 7616 12665
rect 8208 12656 8260 12708
rect 8852 12656 8904 12708
rect 2596 12588 2648 12640
rect 3976 12631 4028 12640
rect 3976 12597 3985 12631
rect 3985 12597 4019 12631
rect 4019 12597 4028 12631
rect 3976 12588 4028 12597
rect 4528 12588 4580 12640
rect 6184 12631 6236 12640
rect 6184 12597 6193 12631
rect 6193 12597 6227 12631
rect 6227 12597 6236 12631
rect 6184 12588 6236 12597
rect 6828 12588 6880 12640
rect 7472 12588 7524 12640
rect 8484 12631 8536 12640
rect 8484 12597 8493 12631
rect 8493 12597 8527 12631
rect 8527 12597 8536 12631
rect 8484 12588 8536 12597
rect 8760 12631 8812 12640
rect 8760 12597 8769 12631
rect 8769 12597 8803 12631
rect 8803 12597 8812 12631
rect 11060 12656 11112 12708
rect 11428 12733 11437 12767
rect 11437 12733 11471 12767
rect 11471 12733 11480 12767
rect 11428 12724 11480 12733
rect 11796 12724 11848 12776
rect 14832 12724 14884 12776
rect 16304 12724 16356 12776
rect 12532 12699 12584 12708
rect 12532 12665 12541 12699
rect 12541 12665 12575 12699
rect 12575 12665 12584 12699
rect 12532 12656 12584 12665
rect 10324 12631 10376 12640
rect 8760 12588 8812 12597
rect 10324 12597 10333 12631
rect 10333 12597 10367 12631
rect 10367 12597 10376 12631
rect 10324 12588 10376 12597
rect 10692 12588 10744 12640
rect 11612 12588 11664 12640
rect 11796 12588 11848 12640
rect 13912 12631 13964 12640
rect 13912 12597 13921 12631
rect 13921 12597 13955 12631
rect 13955 12597 13964 12631
rect 15108 12656 15160 12708
rect 16580 12699 16632 12708
rect 16580 12665 16589 12699
rect 16589 12665 16623 12699
rect 16623 12665 16632 12699
rect 16580 12656 16632 12665
rect 17316 12656 17368 12708
rect 21548 12724 21600 12776
rect 19064 12656 19116 12708
rect 13912 12588 13964 12597
rect 17868 12588 17920 12640
rect 8982 12486 9034 12538
rect 9046 12486 9098 12538
rect 9110 12486 9162 12538
rect 9174 12486 9226 12538
rect 16982 12486 17034 12538
rect 17046 12486 17098 12538
rect 17110 12486 17162 12538
rect 17174 12486 17226 12538
rect 6184 12427 6236 12436
rect 6184 12393 6193 12427
rect 6193 12393 6227 12427
rect 6227 12393 6236 12427
rect 6184 12384 6236 12393
rect 8852 12384 8904 12436
rect 11060 12427 11112 12436
rect 11060 12393 11069 12427
rect 11069 12393 11103 12427
rect 11103 12393 11112 12427
rect 11060 12384 11112 12393
rect 16488 12384 16540 12436
rect 18788 12384 18840 12436
rect 20720 12384 20772 12436
rect 4528 12359 4580 12368
rect 4528 12325 4537 12359
rect 4537 12325 4571 12359
rect 4571 12325 4580 12359
rect 4528 12316 4580 12325
rect 8760 12316 8812 12368
rect 11796 12359 11848 12368
rect 11796 12325 11805 12359
rect 11805 12325 11839 12359
rect 11839 12325 11848 12359
rect 11796 12316 11848 12325
rect 12808 12316 12860 12368
rect 2504 12291 2556 12300
rect 2504 12257 2513 12291
rect 2513 12257 2547 12291
rect 2547 12257 2556 12291
rect 2504 12248 2556 12257
rect 2596 12248 2648 12300
rect 5908 12291 5960 12300
rect 5908 12257 5917 12291
rect 5917 12257 5951 12291
rect 5951 12257 5960 12291
rect 5908 12248 5960 12257
rect 6460 12291 6512 12300
rect 6460 12257 6469 12291
rect 6469 12257 6503 12291
rect 6503 12257 6512 12291
rect 6460 12248 6512 12257
rect 9956 12248 10008 12300
rect 3148 12223 3200 12232
rect 3148 12189 3157 12223
rect 3157 12189 3191 12223
rect 3191 12189 3200 12223
rect 3148 12180 3200 12189
rect 3884 12180 3936 12232
rect 4436 12223 4488 12232
rect 4436 12189 4445 12223
rect 4445 12189 4479 12223
rect 4479 12189 4488 12223
rect 4436 12180 4488 12189
rect 4712 12223 4764 12232
rect 4712 12189 4721 12223
rect 4721 12189 4755 12223
rect 4755 12189 4764 12223
rect 4712 12180 4764 12189
rect 8116 12223 8168 12232
rect 8116 12189 8125 12223
rect 8125 12189 8159 12223
rect 8159 12189 8168 12223
rect 8116 12180 8168 12189
rect 8208 12180 8260 12232
rect 12164 12180 12216 12232
rect 4804 12112 4856 12164
rect 5172 12112 5224 12164
rect 13912 12316 13964 12368
rect 14372 12316 14424 12368
rect 16580 12316 16632 12368
rect 17408 12316 17460 12368
rect 18604 12316 18656 12368
rect 15200 12248 15252 12300
rect 16764 12248 16816 12300
rect 19064 12291 19116 12300
rect 19064 12257 19073 12291
rect 19073 12257 19107 12291
rect 19107 12257 19116 12291
rect 19064 12248 19116 12257
rect 19340 12248 19392 12300
rect 13728 12223 13780 12232
rect 13728 12189 13737 12223
rect 13737 12189 13771 12223
rect 13771 12189 13780 12223
rect 13728 12180 13780 12189
rect 14556 12180 14608 12232
rect 17868 12180 17920 12232
rect 7748 12087 7800 12096
rect 7748 12053 7757 12087
rect 7757 12053 7791 12087
rect 7791 12053 7800 12087
rect 7748 12044 7800 12053
rect 10692 12087 10744 12096
rect 10692 12053 10701 12087
rect 10701 12053 10735 12087
rect 10735 12053 10744 12087
rect 10692 12044 10744 12053
rect 11152 12044 11204 12096
rect 13452 12087 13504 12096
rect 13452 12053 13461 12087
rect 13461 12053 13495 12087
rect 13495 12053 13504 12087
rect 13452 12044 13504 12053
rect 16764 12087 16816 12096
rect 16764 12053 16773 12087
rect 16773 12053 16807 12087
rect 16807 12053 16816 12087
rect 16764 12044 16816 12053
rect 19708 12044 19760 12096
rect 4982 11942 5034 11994
rect 5046 11942 5098 11994
rect 5110 11942 5162 11994
rect 5174 11942 5226 11994
rect 12982 11942 13034 11994
rect 13046 11942 13098 11994
rect 13110 11942 13162 11994
rect 13174 11942 13226 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 4528 11840 4580 11892
rect 5908 11840 5960 11892
rect 8760 11840 8812 11892
rect 3148 11747 3200 11756
rect 3148 11713 3157 11747
rect 3157 11713 3191 11747
rect 3191 11713 3200 11747
rect 3148 11704 3200 11713
rect 4712 11704 4764 11756
rect 2504 11636 2556 11688
rect 3608 11636 3660 11688
rect 7748 11636 7800 11688
rect 10416 11840 10468 11892
rect 11796 11883 11848 11892
rect 11796 11849 11805 11883
rect 11805 11849 11839 11883
rect 11839 11849 11848 11883
rect 11796 11840 11848 11849
rect 17408 11883 17460 11892
rect 17408 11849 17417 11883
rect 17417 11849 17451 11883
rect 17451 11849 17460 11883
rect 17408 11840 17460 11849
rect 17868 11883 17920 11892
rect 17868 11849 17877 11883
rect 17877 11849 17911 11883
rect 17911 11849 17920 11883
rect 17868 11840 17920 11849
rect 21640 11883 21692 11892
rect 21640 11849 21649 11883
rect 21649 11849 21683 11883
rect 21683 11849 21692 11883
rect 21640 11840 21692 11849
rect 10508 11772 10560 11824
rect 13728 11704 13780 11756
rect 11152 11636 11204 11688
rect 12716 11636 12768 11688
rect 13452 11679 13504 11688
rect 13452 11645 13461 11679
rect 13461 11645 13495 11679
rect 13495 11645 13504 11679
rect 13452 11636 13504 11645
rect 17316 11772 17368 11824
rect 20168 11772 20220 11824
rect 21364 11772 21416 11824
rect 16764 11704 16816 11756
rect 20720 11704 20772 11756
rect 4988 11611 5040 11620
rect 2596 11500 2648 11552
rect 2688 11500 2740 11552
rect 4988 11577 4997 11611
rect 4997 11577 5031 11611
rect 5031 11577 5040 11611
rect 4988 11568 5040 11577
rect 6000 11611 6052 11620
rect 4896 11500 4948 11552
rect 6000 11577 6009 11611
rect 6009 11577 6043 11611
rect 6043 11577 6052 11611
rect 6000 11568 6052 11577
rect 6460 11568 6512 11620
rect 7564 11568 7616 11620
rect 7472 11543 7524 11552
rect 7472 11509 7481 11543
rect 7481 11509 7515 11543
rect 7515 11509 7524 11543
rect 8576 11568 8628 11620
rect 10692 11568 10744 11620
rect 16580 11611 16632 11620
rect 16580 11577 16589 11611
rect 16589 11577 16623 11611
rect 16623 11577 16632 11611
rect 16580 11568 16632 11577
rect 7472 11500 7524 11509
rect 8116 11500 8168 11552
rect 9956 11543 10008 11552
rect 9956 11509 9965 11543
rect 9965 11509 9999 11543
rect 9999 11509 10008 11543
rect 9956 11500 10008 11509
rect 12164 11543 12216 11552
rect 12164 11509 12173 11543
rect 12173 11509 12207 11543
rect 12207 11509 12216 11543
rect 12164 11500 12216 11509
rect 14372 11543 14424 11552
rect 14372 11509 14381 11543
rect 14381 11509 14415 11543
rect 14415 11509 14424 11543
rect 14372 11500 14424 11509
rect 15200 11543 15252 11552
rect 15200 11509 15209 11543
rect 15209 11509 15243 11543
rect 15243 11509 15252 11543
rect 15200 11500 15252 11509
rect 18052 11500 18104 11552
rect 21640 11636 21692 11688
rect 19616 11611 19668 11620
rect 18788 11500 18840 11552
rect 19340 11543 19392 11552
rect 19340 11509 19349 11543
rect 19349 11509 19383 11543
rect 19383 11509 19392 11543
rect 19340 11500 19392 11509
rect 19616 11577 19625 11611
rect 19625 11577 19659 11611
rect 19659 11577 19668 11611
rect 19616 11568 19668 11577
rect 19524 11500 19576 11552
rect 8982 11398 9034 11450
rect 9046 11398 9098 11450
rect 9110 11398 9162 11450
rect 9174 11398 9226 11450
rect 16982 11398 17034 11450
rect 17046 11398 17098 11450
rect 17110 11398 17162 11450
rect 17174 11398 17226 11450
rect 3148 11339 3200 11348
rect 3148 11305 3157 11339
rect 3157 11305 3191 11339
rect 3191 11305 3200 11339
rect 3148 11296 3200 11305
rect 3884 11339 3936 11348
rect 3884 11305 3893 11339
rect 3893 11305 3927 11339
rect 3927 11305 3936 11339
rect 3884 11296 3936 11305
rect 4896 11296 4948 11348
rect 5448 11296 5500 11348
rect 5908 11296 5960 11348
rect 8116 11339 8168 11348
rect 8116 11305 8125 11339
rect 8125 11305 8159 11339
rect 8159 11305 8168 11339
rect 8116 11296 8168 11305
rect 14372 11296 14424 11348
rect 16580 11296 16632 11348
rect 17776 11296 17828 11348
rect 18052 11339 18104 11348
rect 18052 11305 18061 11339
rect 18061 11305 18095 11339
rect 18095 11305 18104 11339
rect 18052 11296 18104 11305
rect 19064 11339 19116 11348
rect 19064 11305 19073 11339
rect 19073 11305 19107 11339
rect 19107 11305 19116 11339
rect 19064 11296 19116 11305
rect 19616 11296 19668 11348
rect 4620 11228 4672 11280
rect 1676 11160 1728 11212
rect 6276 11228 6328 11280
rect 7196 11228 7248 11280
rect 7748 11271 7800 11280
rect 7748 11237 7757 11271
rect 7757 11237 7791 11271
rect 7791 11237 7800 11271
rect 7748 11228 7800 11237
rect 11152 11271 11204 11280
rect 11152 11237 11161 11271
rect 11161 11237 11195 11271
rect 11195 11237 11204 11271
rect 11152 11228 11204 11237
rect 13452 11271 13504 11280
rect 7564 11203 7616 11212
rect 2412 11135 2464 11144
rect 2412 11101 2421 11135
rect 2421 11101 2455 11135
rect 2455 11101 2464 11135
rect 2412 11092 2464 11101
rect 4252 11092 4304 11144
rect 7564 11169 7573 11203
rect 7573 11169 7607 11203
rect 7607 11169 7616 11203
rect 7564 11160 7616 11169
rect 9312 11160 9364 11212
rect 10692 11203 10744 11212
rect 10692 11169 10701 11203
rect 10701 11169 10735 11203
rect 10735 11169 10744 11203
rect 10692 11160 10744 11169
rect 112 11024 164 11076
rect 3792 11024 3844 11076
rect 7104 11024 7156 11076
rect 7748 11092 7800 11144
rect 11244 11160 11296 11212
rect 13452 11237 13461 11271
rect 13461 11237 13495 11271
rect 13495 11237 13504 11271
rect 13452 11228 13504 11237
rect 13728 11228 13780 11280
rect 16304 11228 16356 11280
rect 12808 11092 12860 11144
rect 13912 11160 13964 11212
rect 19524 11160 19576 11212
rect 20812 11160 20864 11212
rect 14004 11092 14056 11144
rect 14372 11092 14424 11144
rect 16120 11135 16172 11144
rect 16120 11101 16129 11135
rect 16129 11101 16163 11135
rect 16163 11101 16172 11135
rect 16120 11092 16172 11101
rect 18696 11135 18748 11144
rect 18696 11101 18705 11135
rect 18705 11101 18739 11135
rect 18739 11101 18748 11135
rect 18696 11092 18748 11101
rect 9680 11024 9732 11076
rect 10324 11024 10376 11076
rect 14188 11024 14240 11076
rect 17316 11024 17368 11076
rect 18236 11024 18288 11076
rect 756 10956 808 11008
rect 1952 10999 2004 11008
rect 1952 10965 1961 10999
rect 1961 10965 1995 10999
rect 1995 10965 2004 10999
rect 1952 10956 2004 10965
rect 6736 10956 6788 11008
rect 6920 10999 6972 11008
rect 6920 10965 6929 10999
rect 6929 10965 6963 10999
rect 6963 10965 6972 10999
rect 6920 10956 6972 10965
rect 9588 10956 9640 11008
rect 9864 10999 9916 11008
rect 9864 10965 9873 10999
rect 9873 10965 9907 10999
rect 9907 10965 9916 10999
rect 9864 10956 9916 10965
rect 4982 10854 5034 10906
rect 5046 10854 5098 10906
rect 5110 10854 5162 10906
rect 5174 10854 5226 10906
rect 12982 10854 13034 10906
rect 13046 10854 13098 10906
rect 13110 10854 13162 10906
rect 13174 10854 13226 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 6276 10795 6328 10804
rect 6276 10761 6285 10795
rect 6285 10761 6319 10795
rect 6319 10761 6328 10795
rect 6276 10752 6328 10761
rect 7104 10752 7156 10804
rect 8944 10795 8996 10804
rect 8944 10761 8953 10795
rect 8953 10761 8987 10795
rect 8987 10761 8996 10795
rect 8944 10752 8996 10761
rect 9312 10795 9364 10804
rect 9312 10761 9321 10795
rect 9321 10761 9355 10795
rect 9355 10761 9364 10795
rect 9312 10752 9364 10761
rect 10324 10752 10376 10804
rect 11244 10752 11296 10804
rect 12164 10752 12216 10804
rect 14372 10795 14424 10804
rect 14372 10761 14381 10795
rect 14381 10761 14415 10795
rect 14415 10761 14424 10795
rect 14372 10752 14424 10761
rect 16304 10752 16356 10804
rect 17776 10795 17828 10804
rect 17776 10761 17785 10795
rect 17785 10761 17819 10795
rect 17819 10761 17828 10795
rect 17776 10752 17828 10761
rect 19064 10795 19116 10804
rect 19064 10761 19073 10795
rect 19073 10761 19107 10795
rect 19107 10761 19116 10795
rect 19064 10752 19116 10761
rect 19524 10795 19576 10804
rect 19524 10761 19533 10795
rect 19533 10761 19567 10795
rect 19567 10761 19576 10795
rect 19524 10752 19576 10761
rect 1676 10684 1728 10736
rect 4712 10684 4764 10736
rect 7564 10684 7616 10736
rect 10232 10684 10284 10736
rect 10692 10727 10744 10736
rect 10692 10693 10701 10727
rect 10701 10693 10735 10727
rect 10735 10693 10744 10727
rect 10692 10684 10744 10693
rect 12808 10684 12860 10736
rect 13360 10684 13412 10736
rect 18052 10684 18104 10736
rect 2412 10616 2464 10668
rect 2596 10616 2648 10668
rect 4252 10659 4304 10668
rect 4252 10625 4261 10659
rect 4261 10625 4295 10659
rect 4295 10625 4304 10659
rect 4252 10616 4304 10625
rect 3700 10591 3752 10600
rect 3700 10557 3709 10591
rect 3709 10557 3743 10591
rect 3743 10557 3752 10591
rect 3700 10548 3752 10557
rect 4160 10591 4212 10600
rect 4160 10557 4169 10591
rect 4169 10557 4203 10591
rect 4203 10557 4212 10591
rect 6000 10616 6052 10668
rect 6736 10616 6788 10668
rect 8852 10616 8904 10668
rect 5448 10591 5500 10600
rect 4160 10548 4212 10557
rect 5448 10557 5457 10591
rect 5457 10557 5491 10591
rect 5491 10557 5500 10591
rect 5448 10548 5500 10557
rect 5724 10591 5776 10600
rect 5724 10557 5733 10591
rect 5733 10557 5767 10591
rect 5767 10557 5776 10591
rect 5724 10548 5776 10557
rect 8484 10591 8536 10600
rect 8484 10557 8502 10591
rect 8502 10557 8536 10591
rect 8484 10548 8536 10557
rect 8944 10548 8996 10600
rect 1952 10480 2004 10532
rect 6920 10480 6972 10532
rect 7288 10480 7340 10532
rect 9680 10523 9732 10532
rect 3700 10412 3752 10464
rect 4344 10412 4396 10464
rect 4528 10412 4580 10464
rect 4712 10455 4764 10464
rect 4712 10421 4721 10455
rect 4721 10421 4755 10455
rect 4755 10421 4764 10455
rect 4712 10412 4764 10421
rect 5080 10412 5132 10464
rect 7932 10412 7984 10464
rect 9680 10489 9689 10523
rect 9689 10489 9723 10523
rect 9723 10489 9732 10523
rect 9680 10480 9732 10489
rect 9864 10480 9916 10532
rect 10324 10523 10376 10532
rect 10324 10489 10333 10523
rect 10333 10489 10367 10523
rect 10367 10489 10376 10523
rect 10324 10480 10376 10489
rect 12992 10591 13044 10600
rect 12992 10557 13001 10591
rect 13001 10557 13035 10591
rect 13035 10557 13044 10591
rect 12992 10548 13044 10557
rect 13268 10591 13320 10600
rect 13268 10557 13277 10591
rect 13277 10557 13311 10591
rect 13311 10557 13320 10591
rect 13268 10548 13320 10557
rect 16120 10616 16172 10668
rect 18604 10659 18656 10668
rect 18604 10625 18613 10659
rect 18613 10625 18647 10659
rect 18647 10625 18656 10659
rect 18604 10616 18656 10625
rect 19708 10659 19760 10668
rect 19708 10625 19717 10659
rect 19717 10625 19751 10659
rect 19751 10625 19760 10659
rect 19708 10616 19760 10625
rect 20168 10659 20220 10668
rect 20168 10625 20177 10659
rect 20177 10625 20211 10659
rect 20211 10625 20220 10659
rect 20168 10616 20220 10625
rect 15568 10591 15620 10600
rect 15568 10557 15577 10591
rect 15577 10557 15611 10591
rect 15611 10557 15620 10591
rect 15568 10548 15620 10557
rect 12348 10480 12400 10532
rect 16396 10548 16448 10600
rect 17776 10480 17828 10532
rect 19524 10480 19576 10532
rect 11428 10412 11480 10464
rect 11796 10412 11848 10464
rect 15292 10412 15344 10464
rect 15384 10455 15436 10464
rect 15384 10421 15393 10455
rect 15393 10421 15427 10455
rect 15427 10421 15436 10455
rect 15384 10412 15436 10421
rect 20444 10412 20496 10464
rect 20812 10412 20864 10464
rect 8982 10310 9034 10362
rect 9046 10310 9098 10362
rect 9110 10310 9162 10362
rect 9174 10310 9226 10362
rect 16982 10310 17034 10362
rect 17046 10310 17098 10362
rect 17110 10310 17162 10362
rect 17174 10310 17226 10362
rect 1676 10251 1728 10260
rect 1676 10217 1685 10251
rect 1685 10217 1719 10251
rect 1719 10217 1728 10251
rect 1676 10208 1728 10217
rect 1952 10208 2004 10260
rect 3700 10251 3752 10260
rect 3700 10217 3709 10251
rect 3709 10217 3743 10251
rect 3743 10217 3752 10251
rect 3700 10208 3752 10217
rect 4252 10251 4304 10260
rect 4252 10217 4261 10251
rect 4261 10217 4295 10251
rect 4295 10217 4304 10251
rect 4252 10208 4304 10217
rect 2596 10140 2648 10192
rect 4712 10140 4764 10192
rect 5632 10140 5684 10192
rect 12256 10208 12308 10260
rect 13268 10208 13320 10260
rect 14096 10251 14148 10260
rect 6276 10140 6328 10192
rect 6920 10183 6972 10192
rect 6920 10149 6929 10183
rect 6929 10149 6963 10183
rect 6963 10149 6972 10183
rect 6920 10140 6972 10149
rect 9864 10183 9916 10192
rect 9864 10149 9873 10183
rect 9873 10149 9907 10183
rect 9907 10149 9916 10183
rect 9864 10140 9916 10149
rect 11244 10140 11296 10192
rect 13452 10140 13504 10192
rect 4804 10072 4856 10124
rect 5080 10072 5132 10124
rect 8852 10072 8904 10124
rect 11980 10115 12032 10124
rect 11980 10081 11989 10115
rect 11989 10081 12023 10115
rect 12023 10081 12032 10115
rect 11980 10072 12032 10081
rect 1860 10047 1912 10056
rect 1860 10013 1869 10047
rect 1869 10013 1903 10047
rect 1903 10013 1912 10047
rect 1860 10004 1912 10013
rect 4068 10004 4120 10056
rect 5448 10004 5500 10056
rect 6644 10004 6696 10056
rect 7932 10004 7984 10056
rect 10048 10004 10100 10056
rect 10416 10047 10468 10056
rect 10416 10013 10425 10047
rect 10425 10013 10459 10047
rect 10459 10013 10468 10047
rect 10416 10004 10468 10013
rect 12348 10072 12400 10124
rect 12992 10072 13044 10124
rect 14096 10217 14105 10251
rect 14105 10217 14139 10251
rect 14139 10217 14148 10251
rect 14096 10208 14148 10217
rect 15292 10208 15344 10260
rect 16120 10208 16172 10260
rect 19708 10251 19760 10260
rect 19708 10217 19717 10251
rect 19717 10217 19751 10251
rect 19751 10217 19760 10251
rect 19708 10208 19760 10217
rect 15476 10140 15528 10192
rect 16764 10140 16816 10192
rect 18696 10183 18748 10192
rect 18696 10149 18705 10183
rect 18705 10149 18739 10183
rect 18739 10149 18748 10183
rect 18696 10140 18748 10149
rect 18144 10115 18196 10124
rect 14004 10004 14056 10056
rect 15660 10004 15712 10056
rect 16856 10047 16908 10056
rect 16856 10013 16865 10047
rect 16865 10013 16899 10047
rect 16899 10013 16908 10047
rect 16856 10004 16908 10013
rect 18144 10081 18153 10115
rect 18153 10081 18187 10115
rect 18187 10081 18196 10115
rect 18144 10072 18196 10081
rect 19800 10072 19852 10124
rect 20812 10072 20864 10124
rect 18236 10004 18288 10056
rect 3976 9868 4028 9920
rect 7104 9936 7156 9988
rect 7196 9936 7248 9988
rect 12072 9979 12124 9988
rect 12072 9945 12081 9979
rect 12081 9945 12115 9979
rect 12115 9945 12124 9979
rect 12072 9936 12124 9945
rect 13728 9979 13780 9988
rect 13728 9945 13737 9979
rect 13737 9945 13771 9979
rect 13771 9945 13780 9979
rect 13728 9936 13780 9945
rect 21088 9979 21140 9988
rect 21088 9945 21097 9979
rect 21097 9945 21131 9979
rect 21131 9945 21140 9979
rect 21088 9936 21140 9945
rect 4620 9911 4672 9920
rect 4620 9877 4629 9911
rect 4629 9877 4663 9911
rect 4663 9877 4672 9911
rect 4620 9868 4672 9877
rect 13544 9868 13596 9920
rect 14924 9868 14976 9920
rect 15568 9911 15620 9920
rect 15568 9877 15577 9911
rect 15577 9877 15611 9911
rect 15611 9877 15620 9911
rect 15568 9868 15620 9877
rect 19064 9911 19116 9920
rect 19064 9877 19073 9911
rect 19073 9877 19107 9911
rect 19107 9877 19116 9911
rect 19064 9868 19116 9877
rect 19248 9868 19300 9920
rect 4982 9766 5034 9818
rect 5046 9766 5098 9818
rect 5110 9766 5162 9818
rect 5174 9766 5226 9818
rect 12982 9766 13034 9818
rect 13046 9766 13098 9818
rect 13110 9766 13162 9818
rect 13174 9766 13226 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 6276 9707 6328 9716
rect 6276 9673 6285 9707
rect 6285 9673 6319 9707
rect 6319 9673 6328 9707
rect 6276 9664 6328 9673
rect 7104 9664 7156 9716
rect 8852 9664 8904 9716
rect 9864 9664 9916 9716
rect 10048 9707 10100 9716
rect 10048 9673 10057 9707
rect 10057 9673 10091 9707
rect 10091 9673 10100 9707
rect 10048 9664 10100 9673
rect 12532 9664 12584 9716
rect 15384 9664 15436 9716
rect 18144 9664 18196 9716
rect 12072 9639 12124 9648
rect 12072 9605 12081 9639
rect 12081 9605 12115 9639
rect 12115 9605 12124 9639
rect 12072 9596 12124 9605
rect 1860 9528 1912 9580
rect 5724 9528 5776 9580
rect 2136 9503 2188 9512
rect 2136 9469 2145 9503
rect 2145 9469 2179 9503
rect 2179 9469 2188 9503
rect 2136 9460 2188 9469
rect 2228 9460 2280 9512
rect 4160 9460 4212 9512
rect 4620 9503 4672 9512
rect 4620 9469 4629 9503
rect 4629 9469 4663 9503
rect 4663 9469 4672 9503
rect 4620 9460 4672 9469
rect 4528 9435 4580 9444
rect 4528 9401 4537 9435
rect 4537 9401 4571 9435
rect 4571 9401 4580 9435
rect 6552 9460 6604 9512
rect 6920 9503 6972 9512
rect 6920 9469 6929 9503
rect 6929 9469 6963 9503
rect 6963 9469 6972 9503
rect 6920 9460 6972 9469
rect 8116 9528 8168 9580
rect 11796 9528 11848 9580
rect 13452 9596 13504 9648
rect 14924 9596 14976 9648
rect 16672 9639 16724 9648
rect 16672 9605 16681 9639
rect 16681 9605 16715 9639
rect 16715 9605 16724 9639
rect 16672 9596 16724 9605
rect 12900 9528 12952 9580
rect 13728 9528 13780 9580
rect 15384 9528 15436 9580
rect 16120 9571 16172 9580
rect 16120 9537 16129 9571
rect 16129 9537 16163 9571
rect 16163 9537 16172 9571
rect 16120 9528 16172 9537
rect 19248 9528 19300 9580
rect 5356 9435 5408 9444
rect 4528 9392 4580 9401
rect 5356 9401 5365 9435
rect 5365 9401 5399 9435
rect 5399 9401 5408 9435
rect 5356 9392 5408 9401
rect 9956 9460 10008 9512
rect 11152 9503 11204 9512
rect 8576 9392 8628 9444
rect 11152 9469 11161 9503
rect 11161 9469 11195 9503
rect 11195 9469 11204 9503
rect 11152 9460 11204 9469
rect 11888 9460 11940 9512
rect 13544 9460 13596 9512
rect 14004 9503 14056 9512
rect 14004 9469 14013 9503
rect 14013 9469 14047 9503
rect 14047 9469 14056 9503
rect 14004 9460 14056 9469
rect 14280 9503 14332 9512
rect 14280 9469 14289 9503
rect 14289 9469 14323 9503
rect 14323 9469 14332 9503
rect 14280 9460 14332 9469
rect 13636 9392 13688 9444
rect 16212 9435 16264 9444
rect 16212 9401 16221 9435
rect 16221 9401 16255 9435
rect 16255 9401 16264 9435
rect 16212 9392 16264 9401
rect 19064 9392 19116 9444
rect 19524 9392 19576 9444
rect 19800 9435 19852 9444
rect 19800 9401 19809 9435
rect 19809 9401 19843 9435
rect 19843 9401 19852 9435
rect 19800 9392 19852 9401
rect 2596 9324 2648 9376
rect 5724 9367 5776 9376
rect 5724 9333 5733 9367
rect 5733 9333 5767 9367
rect 5767 9333 5776 9367
rect 5724 9324 5776 9333
rect 10140 9324 10192 9376
rect 12808 9324 12860 9376
rect 15660 9324 15712 9376
rect 16764 9324 16816 9376
rect 18236 9367 18288 9376
rect 18236 9333 18245 9367
rect 18245 9333 18279 9367
rect 18279 9333 18288 9367
rect 18236 9324 18288 9333
rect 20904 9367 20956 9376
rect 20904 9333 20913 9367
rect 20913 9333 20947 9367
rect 20947 9333 20956 9367
rect 20904 9324 20956 9333
rect 8982 9222 9034 9274
rect 9046 9222 9098 9274
rect 9110 9222 9162 9274
rect 9174 9222 9226 9274
rect 16982 9222 17034 9274
rect 17046 9222 17098 9274
rect 17110 9222 17162 9274
rect 17174 9222 17226 9274
rect 2228 9163 2280 9172
rect 2228 9129 2237 9163
rect 2237 9129 2271 9163
rect 2271 9129 2280 9163
rect 2228 9120 2280 9129
rect 2412 9163 2464 9172
rect 2412 9129 2421 9163
rect 2421 9129 2455 9163
rect 2455 9129 2464 9163
rect 2412 9120 2464 9129
rect 4804 9120 4856 9172
rect 5724 9163 5776 9172
rect 5724 9129 5733 9163
rect 5733 9129 5767 9163
rect 5767 9129 5776 9163
rect 5724 9120 5776 9129
rect 7104 9120 7156 9172
rect 8576 9163 8628 9172
rect 1860 8984 1912 9036
rect 2136 8984 2188 9036
rect 2872 9027 2924 9036
rect 2872 8993 2881 9027
rect 2881 8993 2915 9027
rect 2915 8993 2924 9027
rect 4528 9052 4580 9104
rect 6644 9095 6696 9104
rect 6644 9061 6653 9095
rect 6653 9061 6687 9095
rect 6687 9061 6696 9095
rect 6644 9052 6696 9061
rect 6920 9095 6972 9104
rect 6920 9061 6929 9095
rect 6929 9061 6963 9095
rect 6963 9061 6972 9095
rect 6920 9052 6972 9061
rect 7196 9095 7248 9104
rect 7196 9061 7205 9095
rect 7205 9061 7239 9095
rect 7239 9061 7248 9095
rect 7196 9052 7248 9061
rect 8576 9129 8585 9163
rect 8585 9129 8619 9163
rect 8619 9129 8628 9163
rect 8576 9120 8628 9129
rect 12900 9163 12952 9172
rect 12900 9129 12909 9163
rect 12909 9129 12943 9163
rect 12943 9129 12952 9163
rect 12900 9120 12952 9129
rect 15108 9120 15160 9172
rect 9864 9095 9916 9104
rect 9864 9061 9873 9095
rect 9873 9061 9907 9095
rect 9907 9061 9916 9095
rect 9864 9052 9916 9061
rect 10416 9095 10468 9104
rect 10416 9061 10425 9095
rect 10425 9061 10459 9095
rect 10459 9061 10468 9095
rect 10416 9052 10468 9061
rect 2872 8984 2924 8993
rect 4252 8984 4304 9036
rect 11888 9027 11940 9036
rect 11888 8993 11897 9027
rect 11897 8993 11931 9027
rect 11931 8993 11940 9027
rect 11888 8984 11940 8993
rect 11980 8984 12032 9036
rect 13268 9052 13320 9104
rect 16212 9120 16264 9172
rect 18144 9120 18196 9172
rect 19064 9120 19116 9172
rect 19248 9163 19300 9172
rect 19248 9129 19257 9163
rect 19257 9129 19291 9163
rect 19291 9129 19300 9163
rect 19248 9120 19300 9129
rect 13544 9027 13596 9036
rect 13544 8993 13553 9027
rect 13553 8993 13587 9027
rect 13587 8993 13596 9027
rect 13544 8984 13596 8993
rect 14280 8984 14332 9036
rect 15844 8984 15896 9036
rect 16304 8984 16356 9036
rect 16856 8984 16908 9036
rect 17776 8984 17828 9036
rect 19708 9027 19760 9036
rect 19708 8993 19752 9027
rect 19752 8993 19760 9027
rect 19708 8984 19760 8993
rect 5356 8959 5408 8968
rect 5356 8925 5365 8959
rect 5365 8925 5399 8959
rect 5399 8925 5408 8959
rect 5356 8916 5408 8925
rect 7472 8959 7524 8968
rect 7472 8925 7481 8959
rect 7481 8925 7515 8959
rect 7515 8925 7524 8959
rect 7472 8916 7524 8925
rect 9588 8916 9640 8968
rect 10232 8916 10284 8968
rect 13728 8916 13780 8968
rect 15476 8916 15528 8968
rect 18144 8916 18196 8968
rect 9680 8848 9732 8900
rect 11520 8848 11572 8900
rect 13360 8848 13412 8900
rect 11888 8780 11940 8832
rect 18972 8780 19024 8832
rect 4982 8678 5034 8730
rect 5046 8678 5098 8730
rect 5110 8678 5162 8730
rect 5174 8678 5226 8730
rect 12982 8678 13034 8730
rect 13046 8678 13098 8730
rect 13110 8678 13162 8730
rect 13174 8678 13226 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 2872 8576 2924 8628
rect 5356 8576 5408 8628
rect 7196 8576 7248 8628
rect 1768 8508 1820 8560
rect 6552 8508 6604 8560
rect 2044 8440 2096 8492
rect 4252 8483 4304 8492
rect 4252 8449 4261 8483
rect 4261 8449 4295 8483
rect 4295 8449 4304 8483
rect 11152 8576 11204 8628
rect 11520 8619 11572 8628
rect 11520 8585 11529 8619
rect 11529 8585 11563 8619
rect 11563 8585 11572 8619
rect 11520 8576 11572 8585
rect 11980 8576 12032 8628
rect 12072 8576 12124 8628
rect 8576 8508 8628 8560
rect 10324 8508 10376 8560
rect 10140 8483 10192 8492
rect 4252 8440 4304 8449
rect 10140 8449 10149 8483
rect 10149 8449 10183 8483
rect 10183 8449 10192 8483
rect 10140 8440 10192 8449
rect 4344 8415 4396 8424
rect 4344 8381 4353 8415
rect 4353 8381 4387 8415
rect 4387 8381 4396 8415
rect 4344 8372 4396 8381
rect 2504 8347 2556 8356
rect 2504 8313 2513 8347
rect 2513 8313 2547 8347
rect 2547 8313 2556 8347
rect 2504 8304 2556 8313
rect 1860 8279 1912 8288
rect 1860 8245 1869 8279
rect 1869 8245 1903 8279
rect 1903 8245 1912 8279
rect 1860 8236 1912 8245
rect 2596 8236 2648 8288
rect 5724 8372 5776 8424
rect 6736 8372 6788 8424
rect 7840 8415 7892 8424
rect 7840 8381 7849 8415
rect 7849 8381 7883 8415
rect 7883 8381 7892 8415
rect 7840 8372 7892 8381
rect 15384 8576 15436 8628
rect 15844 8619 15896 8628
rect 15844 8585 15853 8619
rect 15853 8585 15887 8619
rect 15887 8585 15896 8619
rect 15844 8576 15896 8585
rect 16212 8619 16264 8628
rect 16212 8585 16221 8619
rect 16221 8585 16255 8619
rect 16255 8585 16264 8619
rect 16212 8576 16264 8585
rect 17776 8619 17828 8628
rect 17776 8585 17785 8619
rect 17785 8585 17819 8619
rect 17819 8585 17828 8619
rect 17776 8576 17828 8585
rect 18144 8576 18196 8628
rect 19708 8619 19760 8628
rect 19708 8585 19717 8619
rect 19717 8585 19751 8619
rect 19751 8585 19760 8619
rect 19708 8576 19760 8585
rect 16672 8508 16724 8560
rect 13360 8440 13412 8492
rect 16764 8440 16816 8492
rect 18972 8440 19024 8492
rect 19248 8440 19300 8492
rect 7380 8347 7432 8356
rect 7380 8313 7389 8347
rect 7389 8313 7423 8347
rect 7423 8313 7432 8347
rect 7380 8304 7432 8313
rect 12808 8372 12860 8424
rect 14924 8415 14976 8424
rect 14924 8381 14933 8415
rect 14933 8381 14967 8415
rect 14967 8381 14976 8415
rect 14924 8372 14976 8381
rect 9864 8304 9916 8356
rect 10416 8304 10468 8356
rect 15660 8372 15712 8424
rect 15476 8347 15528 8356
rect 15476 8313 15485 8347
rect 15485 8313 15519 8347
rect 15519 8313 15528 8347
rect 15476 8304 15528 8313
rect 5264 8279 5316 8288
rect 5264 8245 5273 8279
rect 5273 8245 5307 8279
rect 5307 8245 5316 8279
rect 5264 8236 5316 8245
rect 6828 8236 6880 8288
rect 8576 8236 8628 8288
rect 13636 8236 13688 8288
rect 16212 8236 16264 8288
rect 16580 8304 16632 8356
rect 19064 8304 19116 8356
rect 19524 8236 19576 8288
rect 8982 8134 9034 8186
rect 9046 8134 9098 8186
rect 9110 8134 9162 8186
rect 9174 8134 9226 8186
rect 16982 8134 17034 8186
rect 17046 8134 17098 8186
rect 17110 8134 17162 8186
rect 17174 8134 17226 8186
rect 2504 8032 2556 8084
rect 4344 8075 4396 8084
rect 4344 8041 4353 8075
rect 4353 8041 4387 8075
rect 4387 8041 4396 8075
rect 4344 8032 4396 8041
rect 7104 8075 7156 8084
rect 7104 8041 7113 8075
rect 7113 8041 7147 8075
rect 7147 8041 7156 8075
rect 7104 8032 7156 8041
rect 7840 8075 7892 8084
rect 7840 8041 7849 8075
rect 7849 8041 7883 8075
rect 7883 8041 7892 8075
rect 7840 8032 7892 8041
rect 9588 8032 9640 8084
rect 10416 8075 10468 8084
rect 10416 8041 10425 8075
rect 10425 8041 10459 8075
rect 10459 8041 10468 8075
rect 10416 8032 10468 8041
rect 11980 8032 12032 8084
rect 2596 7964 2648 8016
rect 5264 7964 5316 8016
rect 5908 7964 5960 8016
rect 6552 8007 6604 8016
rect 6552 7973 6561 8007
rect 6561 7973 6595 8007
rect 6595 7973 6604 8007
rect 6552 7964 6604 7973
rect 7472 7964 7524 8016
rect 3700 7896 3752 7948
rect 4528 7939 4580 7948
rect 4528 7905 4537 7939
rect 4537 7905 4571 7939
rect 4571 7905 4580 7939
rect 4528 7896 4580 7905
rect 7748 7939 7800 7948
rect 7748 7905 7757 7939
rect 7757 7905 7791 7939
rect 7791 7905 7800 7939
rect 7748 7896 7800 7905
rect 8116 7939 8168 7948
rect 8116 7905 8125 7939
rect 8125 7905 8159 7939
rect 8159 7905 8168 7939
rect 8116 7896 8168 7905
rect 9956 7939 10008 7948
rect 9956 7905 9965 7939
rect 9965 7905 9999 7939
rect 9999 7905 10008 7939
rect 9956 7896 10008 7905
rect 11336 7896 11388 7948
rect 2412 7828 2464 7880
rect 6276 7828 6328 7880
rect 7288 7828 7340 7880
rect 12624 8032 12676 8084
rect 15476 8075 15528 8084
rect 15476 8041 15485 8075
rect 15485 8041 15519 8075
rect 15519 8041 15528 8075
rect 15476 8032 15528 8041
rect 19064 8032 19116 8084
rect 15844 8007 15896 8016
rect 15844 7973 15853 8007
rect 15853 7973 15887 8007
rect 15887 7973 15896 8007
rect 15844 7964 15896 7973
rect 16580 7964 16632 8016
rect 19156 8007 19208 8016
rect 19156 7973 19165 8007
rect 19165 7973 19199 8007
rect 19199 7973 19208 8007
rect 19156 7964 19208 7973
rect 12624 7896 12676 7948
rect 14188 7896 14240 7948
rect 17684 7939 17736 7948
rect 17684 7905 17693 7939
rect 17693 7905 17727 7939
rect 17727 7905 17736 7939
rect 17684 7896 17736 7905
rect 16488 7828 16540 7880
rect 17592 7828 17644 7880
rect 18420 7828 18472 7880
rect 19524 7828 19576 7880
rect 13360 7760 13412 7812
rect 19616 7803 19668 7812
rect 19616 7769 19625 7803
rect 19625 7769 19659 7803
rect 19659 7769 19668 7803
rect 19616 7760 19668 7769
rect 4804 7692 4856 7744
rect 8484 7692 8536 7744
rect 10324 7692 10376 7744
rect 10784 7692 10836 7744
rect 11980 7735 12032 7744
rect 11980 7701 11989 7735
rect 11989 7701 12023 7735
rect 12023 7701 12032 7735
rect 11980 7692 12032 7701
rect 12808 7735 12860 7744
rect 12808 7701 12817 7735
rect 12817 7701 12851 7735
rect 12851 7701 12860 7735
rect 12808 7692 12860 7701
rect 13544 7735 13596 7744
rect 13544 7701 13553 7735
rect 13553 7701 13587 7735
rect 13587 7701 13596 7735
rect 13544 7692 13596 7701
rect 14924 7692 14976 7744
rect 15752 7692 15804 7744
rect 16764 7735 16816 7744
rect 16764 7701 16773 7735
rect 16773 7701 16807 7735
rect 16807 7701 16816 7735
rect 16764 7692 16816 7701
rect 16948 7692 17000 7744
rect 20444 7692 20496 7744
rect 4982 7590 5034 7642
rect 5046 7590 5098 7642
rect 5110 7590 5162 7642
rect 5174 7590 5226 7642
rect 12982 7590 13034 7642
rect 13046 7590 13098 7642
rect 13110 7590 13162 7642
rect 13174 7590 13226 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 2412 7488 2464 7540
rect 4528 7531 4580 7540
rect 4528 7497 4537 7531
rect 4537 7497 4571 7531
rect 4571 7497 4580 7531
rect 4528 7488 4580 7497
rect 5908 7531 5960 7540
rect 5908 7497 5917 7531
rect 5917 7497 5951 7531
rect 5951 7497 5960 7531
rect 5908 7488 5960 7497
rect 6276 7531 6328 7540
rect 6276 7497 6285 7531
rect 6285 7497 6319 7531
rect 6319 7497 6328 7531
rect 6276 7488 6328 7497
rect 8024 7531 8076 7540
rect 8024 7497 8033 7531
rect 8033 7497 8067 7531
rect 8067 7497 8076 7531
rect 8024 7488 8076 7497
rect 8576 7488 8628 7540
rect 11336 7488 11388 7540
rect 12808 7488 12860 7540
rect 8116 7420 8168 7472
rect 13728 7488 13780 7540
rect 15200 7488 15252 7540
rect 14648 7420 14700 7472
rect 16948 7488 17000 7540
rect 17684 7488 17736 7540
rect 17868 7488 17920 7540
rect 19156 7488 19208 7540
rect 16672 7463 16724 7472
rect 2044 7395 2096 7404
rect 2044 7361 2053 7395
rect 2053 7361 2087 7395
rect 2087 7361 2096 7395
rect 2044 7352 2096 7361
rect 4804 7395 4856 7404
rect 4804 7361 4813 7395
rect 4813 7361 4847 7395
rect 4847 7361 4856 7395
rect 4804 7352 4856 7361
rect 6460 7352 6512 7404
rect 9956 7395 10008 7404
rect 9956 7361 9965 7395
rect 9965 7361 9999 7395
rect 9999 7361 10008 7395
rect 9956 7352 10008 7361
rect 10784 7395 10836 7404
rect 10784 7361 10793 7395
rect 10793 7361 10827 7395
rect 10827 7361 10836 7395
rect 10784 7352 10836 7361
rect 10968 7352 11020 7404
rect 12900 7352 12952 7404
rect 13360 7352 13412 7404
rect 13636 7395 13688 7404
rect 13636 7361 13645 7395
rect 13645 7361 13679 7395
rect 13679 7361 13688 7395
rect 13636 7352 13688 7361
rect 3792 7327 3844 7336
rect 3792 7293 3810 7327
rect 3810 7293 3844 7327
rect 3792 7284 3844 7293
rect 8024 7284 8076 7336
rect 8484 7327 8536 7336
rect 8484 7293 8493 7327
rect 8493 7293 8527 7327
rect 8527 7293 8536 7327
rect 8484 7284 8536 7293
rect 8576 7284 8628 7336
rect 4988 7216 5040 7268
rect 6552 7216 6604 7268
rect 8668 7216 8720 7268
rect 12624 7284 12676 7336
rect 13544 7284 13596 7336
rect 16672 7429 16681 7463
rect 16681 7429 16715 7463
rect 16715 7429 16724 7463
rect 16672 7420 16724 7429
rect 18512 7420 18564 7472
rect 19616 7420 19668 7472
rect 19248 7352 19300 7404
rect 12716 7216 12768 7268
rect 14096 7216 14148 7268
rect 15844 7259 15896 7268
rect 15844 7225 15853 7259
rect 15853 7225 15887 7259
rect 15887 7225 15896 7259
rect 16212 7259 16264 7268
rect 15844 7216 15896 7225
rect 16212 7225 16221 7259
rect 16221 7225 16255 7259
rect 16255 7225 16264 7259
rect 16212 7216 16264 7225
rect 2596 7191 2648 7200
rect 2596 7157 2605 7191
rect 2605 7157 2639 7191
rect 2639 7157 2648 7191
rect 2596 7148 2648 7157
rect 3148 7148 3200 7200
rect 3700 7148 3752 7200
rect 4436 7148 4488 7200
rect 9680 7148 9732 7200
rect 14188 7148 14240 7200
rect 17592 7148 17644 7200
rect 19340 7148 19392 7200
rect 20812 7191 20864 7200
rect 20812 7157 20821 7191
rect 20821 7157 20855 7191
rect 20855 7157 20864 7191
rect 20812 7148 20864 7157
rect 8982 7046 9034 7098
rect 9046 7046 9098 7098
rect 9110 7046 9162 7098
rect 9174 7046 9226 7098
rect 16982 7046 17034 7098
rect 17046 7046 17098 7098
rect 17110 7046 17162 7098
rect 17174 7046 17226 7098
rect 4804 6944 4856 6996
rect 6828 6944 6880 6996
rect 7748 6944 7800 6996
rect 9680 6944 9732 6996
rect 16212 6987 16264 6996
rect 4988 6876 5040 6928
rect 5724 6876 5776 6928
rect 8484 6919 8536 6928
rect 8484 6885 8493 6919
rect 8493 6885 8527 6919
rect 8527 6885 8536 6919
rect 8484 6876 8536 6885
rect 10324 6919 10376 6928
rect 10324 6885 10333 6919
rect 10333 6885 10367 6919
rect 10367 6885 10376 6919
rect 10324 6876 10376 6885
rect 11152 6876 11204 6928
rect 15384 6876 15436 6928
rect 16212 6953 16221 6987
rect 16221 6953 16255 6987
rect 16255 6953 16264 6987
rect 16212 6944 16264 6953
rect 16488 6987 16540 6996
rect 16488 6953 16497 6987
rect 16497 6953 16531 6987
rect 16531 6953 16540 6987
rect 16488 6944 16540 6953
rect 16764 6944 16816 6996
rect 19156 6944 19208 6996
rect 19524 6987 19576 6996
rect 19524 6953 19533 6987
rect 19533 6953 19567 6987
rect 19567 6953 19576 6987
rect 19524 6944 19576 6953
rect 21272 6944 21324 6996
rect 18144 6876 18196 6928
rect 1768 6808 1820 6860
rect 2688 6808 2740 6860
rect 3516 6808 3568 6860
rect 6460 6851 6512 6860
rect 6460 6817 6469 6851
rect 6469 6817 6503 6851
rect 6503 6817 6512 6851
rect 6460 6808 6512 6817
rect 6920 6808 6972 6860
rect 7564 6808 7616 6860
rect 7932 6808 7984 6860
rect 11888 6851 11940 6860
rect 11888 6817 11906 6851
rect 11906 6817 11940 6851
rect 11888 6808 11940 6817
rect 12808 6808 12860 6860
rect 13912 6851 13964 6860
rect 13912 6817 13921 6851
rect 13921 6817 13955 6851
rect 13955 6817 13964 6851
rect 13912 6808 13964 6817
rect 4436 6740 4488 6792
rect 4804 6740 4856 6792
rect 7196 6740 7248 6792
rect 10600 6783 10652 6792
rect 10600 6749 10609 6783
rect 10609 6749 10643 6783
rect 10643 6749 10652 6783
rect 10600 6740 10652 6749
rect 13268 6715 13320 6724
rect 13268 6681 13277 6715
rect 13277 6681 13311 6715
rect 13311 6681 13320 6715
rect 13268 6672 13320 6681
rect 13636 6672 13688 6724
rect 14096 6808 14148 6860
rect 15476 6808 15528 6860
rect 17132 6851 17184 6860
rect 17132 6817 17150 6851
rect 17150 6817 17184 6851
rect 17132 6808 17184 6817
rect 18880 6808 18932 6860
rect 21456 6808 21508 6860
rect 16580 6740 16632 6792
rect 18144 6740 18196 6792
rect 204 6604 256 6656
rect 2964 6604 3016 6656
rect 5908 6604 5960 6656
rect 10324 6604 10376 6656
rect 12624 6647 12676 6656
rect 12624 6613 12633 6647
rect 12633 6613 12667 6647
rect 12667 6613 12676 6647
rect 12624 6604 12676 6613
rect 12808 6604 12860 6656
rect 16672 6604 16724 6656
rect 18236 6604 18288 6656
rect 4982 6502 5034 6554
rect 5046 6502 5098 6554
rect 5110 6502 5162 6554
rect 5174 6502 5226 6554
rect 12982 6502 13034 6554
rect 13046 6502 13098 6554
rect 13110 6502 13162 6554
rect 13174 6502 13226 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 1768 6400 1820 6452
rect 2688 6443 2740 6452
rect 2688 6409 2697 6443
rect 2697 6409 2731 6443
rect 2731 6409 2740 6443
rect 2688 6400 2740 6409
rect 5724 6443 5776 6452
rect 5724 6409 5733 6443
rect 5733 6409 5767 6443
rect 5767 6409 5776 6443
rect 5724 6400 5776 6409
rect 8576 6400 8628 6452
rect 9680 6443 9732 6452
rect 9680 6409 9689 6443
rect 9689 6409 9723 6443
rect 9723 6409 9732 6443
rect 9680 6400 9732 6409
rect 11520 6443 11572 6452
rect 11520 6409 11529 6443
rect 11529 6409 11563 6443
rect 11563 6409 11572 6443
rect 11520 6400 11572 6409
rect 11796 6400 11848 6452
rect 14096 6400 14148 6452
rect 15384 6443 15436 6452
rect 15384 6409 15393 6443
rect 15393 6409 15427 6443
rect 15427 6409 15436 6443
rect 15384 6400 15436 6409
rect 16580 6443 16632 6452
rect 16580 6409 16589 6443
rect 16589 6409 16623 6443
rect 16623 6409 16632 6443
rect 16580 6400 16632 6409
rect 17132 6443 17184 6452
rect 17132 6409 17141 6443
rect 17141 6409 17175 6443
rect 17175 6409 17184 6443
rect 17132 6400 17184 6409
rect 18052 6400 18104 6452
rect 19340 6443 19392 6452
rect 4712 6332 4764 6384
rect 6460 6375 6512 6384
rect 6460 6341 6469 6375
rect 6469 6341 6503 6375
rect 6503 6341 6512 6375
rect 6460 6332 6512 6341
rect 6828 6332 6880 6384
rect 11888 6375 11940 6384
rect 11888 6341 11897 6375
rect 11897 6341 11931 6375
rect 11931 6341 11940 6375
rect 11888 6332 11940 6341
rect 12716 6375 12768 6384
rect 12716 6341 12740 6375
rect 12740 6341 12768 6375
rect 12716 6332 12768 6341
rect 7196 6307 7248 6316
rect 7196 6273 7205 6307
rect 7205 6273 7239 6307
rect 7239 6273 7248 6307
rect 7196 6264 7248 6273
rect 10324 6307 10376 6316
rect 10324 6273 10333 6307
rect 10333 6273 10367 6307
rect 10367 6273 10376 6307
rect 10324 6264 10376 6273
rect 10968 6307 11020 6316
rect 10968 6273 10977 6307
rect 10977 6273 11011 6307
rect 11011 6273 11020 6307
rect 10968 6264 11020 6273
rect 2964 6196 3016 6248
rect 4528 6239 4580 6248
rect 4528 6205 4537 6239
rect 4537 6205 4571 6239
rect 4571 6205 4580 6239
rect 4528 6196 4580 6205
rect 6000 6196 6052 6248
rect 8484 6239 8536 6248
rect 8484 6205 8493 6239
rect 8493 6205 8527 6239
rect 8527 6205 8536 6239
rect 8484 6196 8536 6205
rect 10048 6239 10100 6248
rect 10048 6205 10057 6239
rect 10057 6205 10091 6239
rect 10091 6205 10100 6239
rect 10048 6196 10100 6205
rect 8576 6128 8628 6180
rect 11704 6128 11756 6180
rect 13268 6264 13320 6316
rect 12624 6196 12676 6248
rect 16120 6307 16172 6316
rect 16120 6273 16129 6307
rect 16129 6273 16163 6307
rect 16163 6273 16172 6307
rect 16120 6264 16172 6273
rect 13268 6171 13320 6180
rect 13268 6137 13277 6171
rect 13277 6137 13311 6171
rect 13311 6137 13320 6171
rect 13268 6128 13320 6137
rect 13360 6128 13412 6180
rect 14372 6196 14424 6248
rect 15936 6196 15988 6248
rect 15660 6128 15712 6180
rect 17592 6196 17644 6248
rect 18144 6128 18196 6180
rect 19340 6409 19349 6443
rect 19349 6409 19383 6443
rect 19383 6409 19392 6443
rect 19340 6400 19392 6409
rect 21456 6443 21508 6452
rect 21456 6409 21465 6443
rect 21465 6409 21499 6443
rect 21499 6409 21508 6443
rect 21456 6400 21508 6409
rect 18420 6307 18472 6316
rect 18420 6273 18429 6307
rect 18429 6273 18463 6307
rect 18463 6273 18472 6307
rect 18420 6264 18472 6273
rect 18604 6128 18656 6180
rect 3148 6103 3200 6112
rect 3148 6069 3157 6103
rect 3157 6069 3191 6103
rect 3191 6069 3200 6103
rect 3148 6060 3200 6069
rect 7932 6103 7984 6112
rect 7932 6069 7941 6103
rect 7941 6069 7975 6103
rect 7975 6069 7984 6103
rect 7932 6060 7984 6069
rect 14924 6103 14976 6112
rect 14924 6069 14933 6103
rect 14933 6069 14967 6103
rect 14967 6069 14976 6103
rect 14924 6060 14976 6069
rect 21180 6171 21232 6180
rect 21180 6137 21189 6171
rect 21189 6137 21223 6171
rect 21223 6137 21232 6171
rect 21180 6128 21232 6137
rect 20720 6060 20772 6112
rect 8982 5958 9034 6010
rect 9046 5958 9098 6010
rect 9110 5958 9162 6010
rect 9174 5958 9226 6010
rect 16982 5958 17034 6010
rect 17046 5958 17098 6010
rect 17110 5958 17162 6010
rect 17174 5958 17226 6010
rect 4528 5856 4580 5908
rect 4804 5856 4856 5908
rect 7564 5899 7616 5908
rect 7564 5865 7573 5899
rect 7573 5865 7607 5899
rect 7607 5865 7616 5899
rect 7564 5856 7616 5865
rect 10416 5856 10468 5908
rect 5908 5831 5960 5840
rect 4160 5720 4212 5772
rect 5908 5797 5917 5831
rect 5917 5797 5951 5831
rect 5951 5797 5960 5831
rect 5908 5788 5960 5797
rect 6000 5831 6052 5840
rect 6000 5797 6009 5831
rect 6009 5797 6043 5831
rect 6043 5797 6052 5831
rect 6000 5788 6052 5797
rect 8484 5831 8536 5840
rect 8484 5797 8493 5831
rect 8493 5797 8527 5831
rect 8527 5797 8536 5831
rect 8484 5788 8536 5797
rect 10048 5831 10100 5840
rect 10048 5797 10057 5831
rect 10057 5797 10091 5831
rect 10091 5797 10100 5831
rect 10048 5788 10100 5797
rect 10600 5831 10652 5840
rect 10600 5797 10609 5831
rect 10609 5797 10643 5831
rect 10643 5797 10652 5831
rect 10600 5788 10652 5797
rect 15660 5899 15712 5908
rect 15660 5865 15669 5899
rect 15669 5865 15703 5899
rect 15703 5865 15712 5899
rect 15660 5856 15712 5865
rect 15936 5899 15988 5908
rect 15936 5865 15945 5899
rect 15945 5865 15979 5899
rect 15979 5865 15988 5899
rect 15936 5856 15988 5865
rect 16304 5856 16356 5908
rect 18420 5856 18472 5908
rect 4528 5720 4580 5772
rect 6552 5763 6604 5772
rect 6552 5729 6561 5763
rect 6561 5729 6595 5763
rect 6595 5729 6604 5763
rect 6552 5720 6604 5729
rect 7932 5720 7984 5772
rect 7840 5652 7892 5704
rect 8484 5652 8536 5704
rect 8668 5652 8720 5704
rect 9404 5652 9456 5704
rect 9496 5584 9548 5636
rect 12808 5788 12860 5840
rect 15384 5788 15436 5840
rect 18052 5831 18104 5840
rect 3148 5516 3200 5568
rect 4068 5516 4120 5568
rect 7196 5559 7248 5568
rect 7196 5525 7205 5559
rect 7205 5525 7239 5559
rect 7239 5525 7248 5559
rect 7196 5516 7248 5525
rect 11704 5720 11756 5772
rect 13360 5763 13412 5772
rect 13360 5729 13369 5763
rect 13369 5729 13403 5763
rect 13403 5729 13412 5763
rect 13360 5720 13412 5729
rect 13636 5763 13688 5772
rect 13636 5729 13645 5763
rect 13645 5729 13679 5763
rect 13679 5729 13688 5763
rect 13636 5720 13688 5729
rect 16120 5763 16172 5772
rect 16120 5729 16129 5763
rect 16129 5729 16163 5763
rect 16163 5729 16172 5763
rect 16120 5720 16172 5729
rect 18052 5797 18061 5831
rect 18061 5797 18095 5831
rect 18095 5797 18104 5831
rect 18052 5788 18104 5797
rect 20812 5788 20864 5840
rect 21180 5788 21232 5840
rect 14004 5695 14056 5704
rect 14004 5661 14013 5695
rect 14013 5661 14047 5695
rect 14047 5661 14056 5695
rect 14004 5652 14056 5661
rect 17500 5652 17552 5704
rect 21456 5695 21508 5704
rect 21456 5661 21465 5695
rect 21465 5661 21499 5695
rect 21499 5661 21508 5695
rect 21456 5652 21508 5661
rect 11796 5584 11848 5636
rect 13544 5584 13596 5636
rect 14280 5584 14332 5636
rect 18512 5627 18564 5636
rect 18512 5593 18521 5627
rect 18521 5593 18555 5627
rect 18555 5593 18564 5627
rect 18512 5584 18564 5593
rect 11980 5516 12032 5568
rect 12532 5516 12584 5568
rect 14372 5559 14424 5568
rect 14372 5525 14381 5559
rect 14381 5525 14415 5559
rect 14415 5525 14424 5559
rect 14372 5516 14424 5525
rect 20352 5516 20404 5568
rect 4982 5414 5034 5466
rect 5046 5414 5098 5466
rect 5110 5414 5162 5466
rect 5174 5414 5226 5466
rect 12982 5414 13034 5466
rect 13046 5414 13098 5466
rect 13110 5414 13162 5466
rect 13174 5414 13226 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 4160 5355 4212 5364
rect 4160 5321 4169 5355
rect 4169 5321 4203 5355
rect 4203 5321 4212 5355
rect 4528 5355 4580 5364
rect 4160 5312 4212 5321
rect 4528 5321 4537 5355
rect 4537 5321 4571 5355
rect 4571 5321 4580 5355
rect 4528 5312 4580 5321
rect 6000 5312 6052 5364
rect 6368 5312 6420 5364
rect 6552 5312 6604 5364
rect 7380 5312 7432 5364
rect 10048 5312 10100 5364
rect 11796 5312 11848 5364
rect 12256 5312 12308 5364
rect 12532 5355 12584 5364
rect 12532 5321 12541 5355
rect 12541 5321 12575 5355
rect 12575 5321 12584 5355
rect 12532 5312 12584 5321
rect 15384 5312 15436 5364
rect 17500 5355 17552 5364
rect 17500 5321 17509 5355
rect 17509 5321 17543 5355
rect 17543 5321 17552 5355
rect 17500 5312 17552 5321
rect 18052 5312 18104 5364
rect 20812 5312 20864 5364
rect 21272 5312 21324 5364
rect 112 5244 164 5296
rect 11244 5244 11296 5296
rect 14280 5244 14332 5296
rect 21364 5244 21416 5296
rect 1952 5108 2004 5160
rect 4068 5176 4120 5228
rect 5632 5176 5684 5228
rect 7196 5176 7248 5228
rect 7380 5219 7432 5228
rect 7380 5185 7389 5219
rect 7389 5185 7423 5219
rect 7423 5185 7432 5219
rect 7380 5176 7432 5185
rect 10968 5219 11020 5228
rect 10968 5185 10977 5219
rect 10977 5185 11011 5219
rect 11011 5185 11020 5219
rect 10968 5176 11020 5185
rect 3424 5040 3476 5092
rect 4528 5108 4580 5160
rect 5540 5108 5592 5160
rect 5816 5151 5868 5160
rect 5816 5117 5834 5151
rect 5834 5117 5868 5151
rect 5816 5108 5868 5117
rect 6368 5108 6420 5160
rect 7748 5108 7800 5160
rect 8392 5151 8444 5160
rect 8392 5117 8401 5151
rect 8401 5117 8435 5151
rect 8435 5117 8444 5151
rect 8392 5108 8444 5117
rect 13360 5176 13412 5228
rect 13636 5176 13688 5228
rect 16856 5176 16908 5228
rect 17592 5176 17644 5228
rect 6736 5040 6788 5092
rect 7012 5083 7064 5092
rect 7012 5049 7021 5083
rect 7021 5049 7055 5083
rect 7055 5049 7064 5083
rect 7012 5040 7064 5049
rect 1952 5015 2004 5024
rect 1952 4981 1961 5015
rect 1961 4981 1995 5015
rect 1995 4981 2004 5015
rect 1952 4972 2004 4981
rect 2964 4972 3016 5024
rect 12900 5151 12952 5160
rect 12900 5117 12909 5151
rect 12909 5117 12943 5151
rect 12943 5117 12952 5151
rect 12900 5108 12952 5117
rect 9588 5040 9640 5092
rect 10324 5083 10376 5092
rect 10324 5049 10333 5083
rect 10333 5049 10367 5083
rect 10367 5049 10376 5083
rect 10324 5040 10376 5049
rect 8484 4972 8536 5024
rect 10600 4972 10652 5024
rect 11612 5015 11664 5024
rect 11612 4981 11621 5015
rect 11621 4981 11655 5015
rect 11655 4981 11664 5015
rect 11612 4972 11664 4981
rect 12440 4972 12492 5024
rect 14556 5151 14608 5160
rect 14556 5117 14565 5151
rect 14565 5117 14599 5151
rect 14599 5117 14608 5151
rect 14556 5108 14608 5117
rect 14096 4972 14148 5024
rect 15660 4972 15712 5024
rect 16120 5151 16172 5160
rect 16120 5117 16129 5151
rect 16129 5117 16163 5151
rect 16163 5117 16172 5151
rect 16120 5108 16172 5117
rect 18052 5151 18104 5160
rect 18052 5117 18061 5151
rect 18061 5117 18095 5151
rect 18095 5117 18104 5151
rect 18052 5108 18104 5117
rect 21456 5176 21508 5228
rect 20352 5040 20404 5092
rect 20720 5083 20772 5092
rect 20720 5049 20729 5083
rect 20729 5049 20763 5083
rect 20763 5049 20772 5083
rect 20720 5040 20772 5049
rect 17316 4972 17368 5024
rect 18144 5015 18196 5024
rect 18144 4981 18153 5015
rect 18153 4981 18187 5015
rect 18187 4981 18196 5015
rect 18144 4972 18196 4981
rect 8982 4870 9034 4922
rect 9046 4870 9098 4922
rect 9110 4870 9162 4922
rect 9174 4870 9226 4922
rect 16982 4870 17034 4922
rect 17046 4870 17098 4922
rect 17110 4870 17162 4922
rect 17174 4870 17226 4922
rect 5632 4768 5684 4820
rect 5908 4811 5960 4820
rect 5908 4777 5917 4811
rect 5917 4777 5951 4811
rect 5951 4777 5960 4811
rect 5908 4768 5960 4777
rect 6736 4811 6788 4820
rect 6736 4777 6745 4811
rect 6745 4777 6779 4811
rect 6779 4777 6788 4811
rect 6736 4768 6788 4777
rect 7840 4768 7892 4820
rect 8392 4811 8444 4820
rect 8392 4777 8401 4811
rect 8401 4777 8435 4811
rect 8435 4777 8444 4811
rect 8392 4768 8444 4777
rect 10324 4768 10376 4820
rect 11244 4811 11296 4820
rect 11244 4777 11253 4811
rect 11253 4777 11287 4811
rect 11287 4777 11296 4811
rect 11244 4768 11296 4777
rect 12900 4811 12952 4820
rect 12900 4777 12909 4811
rect 12909 4777 12943 4811
rect 12943 4777 12952 4811
rect 14556 4811 14608 4820
rect 12900 4768 12952 4777
rect 4804 4700 4856 4752
rect 7012 4700 7064 4752
rect 7748 4700 7800 4752
rect 9404 4743 9456 4752
rect 9404 4709 9413 4743
rect 9413 4709 9447 4743
rect 9447 4709 9456 4743
rect 9404 4700 9456 4709
rect 9772 4700 9824 4752
rect 11704 4700 11756 4752
rect 14556 4777 14565 4811
rect 14565 4777 14599 4811
rect 14599 4777 14608 4811
rect 14556 4768 14608 4777
rect 16028 4768 16080 4820
rect 16672 4811 16724 4820
rect 16672 4777 16681 4811
rect 16681 4777 16715 4811
rect 16715 4777 16724 4811
rect 16672 4768 16724 4777
rect 18052 4811 18104 4820
rect 18052 4777 18061 4811
rect 18061 4777 18095 4811
rect 18095 4777 18104 4811
rect 18052 4768 18104 4777
rect 18604 4811 18656 4820
rect 18604 4777 18613 4811
rect 18613 4777 18647 4811
rect 18647 4777 18656 4811
rect 18604 4768 18656 4777
rect 20720 4768 20772 4820
rect 14372 4700 14424 4752
rect 2872 4675 2924 4684
rect 2872 4641 2881 4675
rect 2881 4641 2915 4675
rect 2915 4641 2924 4675
rect 2872 4632 2924 4641
rect 5632 4607 5684 4616
rect 5632 4573 5641 4607
rect 5641 4573 5675 4607
rect 5675 4573 5684 4607
rect 5632 4564 5684 4573
rect 5356 4496 5408 4548
rect 6552 4564 6604 4616
rect 6736 4564 6788 4616
rect 7288 4607 7340 4616
rect 7288 4573 7297 4607
rect 7297 4573 7331 4607
rect 7331 4573 7340 4607
rect 7288 4564 7340 4573
rect 6368 4496 6420 4548
rect 3608 4471 3660 4480
rect 3608 4437 3617 4471
rect 3617 4437 3651 4471
rect 3651 4437 3660 4471
rect 3608 4428 3660 4437
rect 5540 4428 5592 4480
rect 8392 4632 8444 4684
rect 9588 4632 9640 4684
rect 10600 4675 10652 4684
rect 10600 4641 10609 4675
rect 10609 4641 10643 4675
rect 10643 4641 10652 4675
rect 10600 4632 10652 4641
rect 13544 4675 13596 4684
rect 13544 4641 13553 4675
rect 13553 4641 13587 4675
rect 13587 4641 13596 4675
rect 13544 4632 13596 4641
rect 15384 4632 15436 4684
rect 16488 4675 16540 4684
rect 16488 4641 16497 4675
rect 16497 4641 16531 4675
rect 16531 4641 16540 4675
rect 16488 4632 16540 4641
rect 20628 4632 20680 4684
rect 11244 4564 11296 4616
rect 10508 4496 10560 4548
rect 17408 4564 17460 4616
rect 20168 4539 20220 4548
rect 12440 4471 12492 4480
rect 12440 4437 12449 4471
rect 12449 4437 12483 4471
rect 12483 4437 12492 4471
rect 12440 4428 12492 4437
rect 14004 4471 14056 4480
rect 14004 4437 14013 4471
rect 14013 4437 14047 4471
rect 14047 4437 14056 4471
rect 14004 4428 14056 4437
rect 16120 4471 16172 4480
rect 16120 4437 16129 4471
rect 16129 4437 16163 4471
rect 16163 4437 16172 4471
rect 20168 4505 20177 4539
rect 20177 4505 20211 4539
rect 20211 4505 20220 4539
rect 20168 4496 20220 4505
rect 16120 4428 16172 4437
rect 4982 4326 5034 4378
rect 5046 4326 5098 4378
rect 5110 4326 5162 4378
rect 5174 4326 5226 4378
rect 12982 4326 13034 4378
rect 13046 4326 13098 4378
rect 13110 4326 13162 4378
rect 13174 4326 13226 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 4804 4224 4856 4276
rect 5356 4267 5408 4276
rect 5356 4233 5365 4267
rect 5365 4233 5399 4267
rect 5399 4233 5408 4267
rect 5356 4224 5408 4233
rect 7748 4267 7800 4276
rect 7748 4233 7757 4267
rect 7757 4233 7791 4267
rect 7791 4233 7800 4267
rect 7748 4224 7800 4233
rect 8392 4267 8444 4276
rect 8392 4233 8401 4267
rect 8401 4233 8435 4267
rect 8435 4233 8444 4267
rect 8392 4224 8444 4233
rect 9312 4224 9364 4276
rect 9588 4224 9640 4276
rect 11704 4267 11756 4276
rect 11704 4233 11713 4267
rect 11713 4233 11747 4267
rect 11747 4233 11756 4267
rect 11704 4224 11756 4233
rect 2872 4156 2924 4208
rect 5816 4156 5868 4208
rect 8300 4156 8352 4208
rect 9680 4156 9732 4208
rect 11980 4156 12032 4208
rect 3424 4088 3476 4140
rect 3608 4063 3660 4072
rect 3608 4029 3617 4063
rect 3617 4029 3651 4063
rect 3651 4029 3660 4063
rect 3608 4020 3660 4029
rect 5632 4020 5684 4072
rect 3700 3952 3752 4004
rect 3148 3884 3200 3936
rect 6644 3952 6696 4004
rect 5540 3884 5592 3936
rect 8300 4020 8352 4072
rect 9496 4088 9548 4140
rect 9312 4020 9364 4072
rect 10600 4088 10652 4140
rect 15016 4156 15068 4208
rect 18788 4224 18840 4276
rect 20628 4224 20680 4276
rect 18236 4156 18288 4208
rect 18604 4156 18656 4208
rect 17316 4088 17368 4140
rect 20168 4131 20220 4140
rect 20168 4097 20177 4131
rect 20177 4097 20211 4131
rect 20211 4097 20220 4131
rect 20168 4088 20220 4097
rect 20352 4088 20404 4140
rect 7472 3952 7524 4004
rect 9404 3952 9456 4004
rect 9772 3952 9824 4004
rect 10876 3995 10928 4004
rect 10876 3961 10885 3995
rect 10885 3961 10919 3995
rect 10919 3961 10928 3995
rect 10876 3952 10928 3961
rect 11704 3952 11756 4004
rect 7380 3884 7432 3936
rect 11612 3884 11664 3936
rect 13636 4020 13688 4072
rect 13912 4020 13964 4072
rect 14096 4020 14148 4072
rect 14372 4063 14424 4072
rect 14372 4029 14381 4063
rect 14381 4029 14415 4063
rect 14415 4029 14424 4063
rect 14372 4020 14424 4029
rect 16212 4020 16264 4072
rect 16488 4020 16540 4072
rect 19340 4020 19392 4072
rect 13452 3927 13504 3936
rect 13452 3893 13461 3927
rect 13461 3893 13495 3927
rect 13495 3893 13504 3927
rect 17684 3952 17736 4004
rect 15384 3927 15436 3936
rect 13452 3884 13504 3893
rect 15384 3893 15393 3927
rect 15393 3893 15427 3927
rect 15427 3893 15436 3927
rect 15384 3884 15436 3893
rect 15752 3927 15804 3936
rect 15752 3893 15761 3927
rect 15761 3893 15795 3927
rect 15795 3893 15804 3927
rect 15752 3884 15804 3893
rect 16764 3884 16816 3936
rect 17408 3927 17460 3936
rect 17408 3893 17417 3927
rect 17417 3893 17451 3927
rect 17451 3893 17460 3927
rect 17408 3884 17460 3893
rect 8982 3782 9034 3834
rect 9046 3782 9098 3834
rect 9110 3782 9162 3834
rect 9174 3782 9226 3834
rect 16982 3782 17034 3834
rect 17046 3782 17098 3834
rect 17110 3782 17162 3834
rect 17174 3782 17226 3834
rect 3424 3723 3476 3732
rect 3424 3689 3433 3723
rect 3433 3689 3467 3723
rect 3467 3689 3476 3723
rect 3424 3680 3476 3689
rect 6276 3680 6328 3732
rect 7380 3723 7432 3732
rect 4436 3612 4488 3664
rect 5540 3612 5592 3664
rect 5632 3612 5684 3664
rect 7380 3689 7389 3723
rect 7389 3689 7423 3723
rect 7423 3689 7432 3723
rect 7380 3680 7432 3689
rect 7656 3680 7708 3732
rect 9496 3680 9548 3732
rect 9956 3723 10008 3732
rect 9956 3689 9965 3723
rect 9965 3689 9999 3723
rect 9999 3689 10008 3723
rect 9956 3680 10008 3689
rect 10600 3680 10652 3732
rect 10968 3680 11020 3732
rect 8116 3587 8168 3596
rect 8116 3553 8125 3587
rect 8125 3553 8159 3587
rect 8159 3553 8168 3587
rect 8116 3544 8168 3553
rect 8484 3544 8536 3596
rect 10232 3587 10284 3596
rect 4528 3519 4580 3528
rect 4528 3485 4537 3519
rect 4537 3485 4571 3519
rect 4571 3485 4580 3519
rect 4528 3476 4580 3485
rect 6368 3519 6420 3528
rect 6368 3485 6377 3519
rect 6377 3485 6411 3519
rect 6411 3485 6420 3519
rect 6368 3476 6420 3485
rect 5632 3408 5684 3460
rect 9588 3476 9640 3528
rect 10232 3553 10241 3587
rect 10241 3553 10275 3587
rect 10275 3553 10284 3587
rect 10232 3544 10284 3553
rect 12256 3680 12308 3732
rect 11520 3655 11572 3664
rect 11520 3621 11529 3655
rect 11529 3621 11563 3655
rect 11563 3621 11572 3655
rect 11520 3612 11572 3621
rect 13544 3680 13596 3732
rect 16028 3723 16080 3732
rect 16028 3689 16037 3723
rect 16037 3689 16071 3723
rect 16071 3689 16080 3723
rect 16028 3680 16080 3689
rect 17684 3723 17736 3732
rect 17684 3689 17693 3723
rect 17693 3689 17727 3723
rect 17727 3689 17736 3723
rect 17684 3680 17736 3689
rect 19340 3723 19392 3732
rect 19340 3689 19349 3723
rect 19349 3689 19383 3723
rect 19383 3689 19392 3723
rect 19340 3680 19392 3689
rect 19984 3680 20036 3732
rect 13912 3612 13964 3664
rect 13452 3544 13504 3596
rect 15660 3544 15712 3596
rect 15752 3544 15804 3596
rect 16212 3544 16264 3596
rect 16856 3544 16908 3596
rect 18236 3612 18288 3664
rect 19064 3612 19116 3664
rect 11704 3519 11756 3528
rect 11704 3485 11713 3519
rect 11713 3485 11747 3519
rect 11747 3485 11756 3519
rect 11704 3476 11756 3485
rect 15384 3476 15436 3528
rect 17776 3476 17828 3528
rect 20812 3476 20864 3528
rect 9680 3408 9732 3460
rect 8392 3340 8444 3392
rect 13268 3408 13320 3460
rect 13360 3408 13412 3460
rect 15476 3408 15528 3460
rect 16120 3408 16172 3460
rect 15936 3340 15988 3392
rect 16672 3383 16724 3392
rect 16672 3349 16681 3383
rect 16681 3349 16715 3383
rect 16715 3349 16724 3383
rect 16672 3340 16724 3349
rect 17316 3383 17368 3392
rect 17316 3349 17325 3383
rect 17325 3349 17359 3383
rect 17359 3349 17368 3383
rect 17316 3340 17368 3349
rect 18052 3383 18104 3392
rect 18052 3349 18061 3383
rect 18061 3349 18095 3383
rect 18095 3349 18104 3383
rect 18052 3340 18104 3349
rect 19892 3340 19944 3392
rect 4982 3238 5034 3290
rect 5046 3238 5098 3290
rect 5110 3238 5162 3290
rect 5174 3238 5226 3290
rect 12982 3238 13034 3290
rect 13046 3238 13098 3290
rect 13110 3238 13162 3290
rect 13174 3238 13226 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 4528 3136 4580 3188
rect 6276 3179 6328 3188
rect 6276 3145 6285 3179
rect 6285 3145 6319 3179
rect 6319 3145 6328 3179
rect 6276 3136 6328 3145
rect 8484 3136 8536 3188
rect 10232 3136 10284 3188
rect 10876 3179 10928 3188
rect 10876 3145 10885 3179
rect 10885 3145 10919 3179
rect 10919 3145 10928 3179
rect 10876 3136 10928 3145
rect 11520 3179 11572 3188
rect 11520 3145 11529 3179
rect 11529 3145 11563 3179
rect 11563 3145 11572 3179
rect 11520 3136 11572 3145
rect 12256 3179 12308 3188
rect 12256 3145 12265 3179
rect 12265 3145 12299 3179
rect 12299 3145 12308 3179
rect 12256 3136 12308 3145
rect 19064 3179 19116 3188
rect 19064 3145 19073 3179
rect 19073 3145 19107 3179
rect 19107 3145 19116 3179
rect 19064 3136 19116 3145
rect 20812 3136 20864 3188
rect 3424 3000 3476 3052
rect 9404 3068 9456 3120
rect 5632 3043 5684 3052
rect 5632 3009 5641 3043
rect 5641 3009 5675 3043
rect 5675 3009 5684 3043
rect 5632 3000 5684 3009
rect 9680 3000 9732 3052
rect 7104 2975 7156 2984
rect 7104 2941 7113 2975
rect 7113 2941 7147 2975
rect 7147 2941 7156 2975
rect 7104 2932 7156 2941
rect 8116 2932 8168 2984
rect 4620 2864 4672 2916
rect 4988 2907 5040 2916
rect 4988 2873 4997 2907
rect 4997 2873 5031 2907
rect 5031 2873 5040 2907
rect 4988 2864 5040 2873
rect 5080 2907 5132 2916
rect 5080 2873 5089 2907
rect 5089 2873 5123 2907
rect 5123 2873 5132 2907
rect 5080 2864 5132 2873
rect 8300 2907 8352 2916
rect 8300 2873 8309 2907
rect 8309 2873 8343 2907
rect 8343 2873 8352 2907
rect 8300 2864 8352 2873
rect 8392 2907 8444 2916
rect 8392 2873 8401 2907
rect 8401 2873 8435 2907
rect 8435 2873 8444 2907
rect 11060 3068 11112 3120
rect 16764 3068 16816 3120
rect 9956 3043 10008 3052
rect 9956 3009 9965 3043
rect 9965 3009 9999 3043
rect 9999 3009 10008 3043
rect 9956 3000 10008 3009
rect 15936 3043 15988 3052
rect 15936 3009 15945 3043
rect 15945 3009 15979 3043
rect 15979 3009 15988 3043
rect 15936 3000 15988 3009
rect 13084 2975 13136 2984
rect 13084 2941 13093 2975
rect 13093 2941 13127 2975
rect 13127 2941 13136 2975
rect 13084 2932 13136 2941
rect 13636 2975 13688 2984
rect 13636 2941 13645 2975
rect 13645 2941 13679 2975
rect 13679 2941 13688 2975
rect 13636 2932 13688 2941
rect 13912 2932 13964 2984
rect 14372 2932 14424 2984
rect 15384 2932 15436 2984
rect 16028 2932 16080 2984
rect 16672 2932 16724 2984
rect 18236 3068 18288 3120
rect 17408 3000 17460 3052
rect 18052 2975 18104 2984
rect 18052 2941 18061 2975
rect 18061 2941 18095 2975
rect 18095 2941 18104 2975
rect 18052 2932 18104 2941
rect 18236 2932 18288 2984
rect 19892 3043 19944 3052
rect 19892 3009 19901 3043
rect 19901 3009 19935 3043
rect 19935 3009 19944 3043
rect 19892 3000 19944 3009
rect 20352 3043 20404 3052
rect 20352 3009 20361 3043
rect 20361 3009 20395 3043
rect 20395 3009 20404 3043
rect 20352 3000 20404 3009
rect 8392 2864 8444 2873
rect 10600 2864 10652 2916
rect 15476 2864 15528 2916
rect 19984 2907 20036 2916
rect 4528 2839 4580 2848
rect 4528 2805 4537 2839
rect 4537 2805 4571 2839
rect 4571 2805 4580 2839
rect 4528 2796 4580 2805
rect 13452 2839 13504 2848
rect 13452 2805 13461 2839
rect 13461 2805 13495 2839
rect 13495 2805 13504 2839
rect 13452 2796 13504 2805
rect 15660 2839 15712 2848
rect 15660 2805 15669 2839
rect 15669 2805 15703 2839
rect 15703 2805 15712 2839
rect 15660 2796 15712 2805
rect 16028 2796 16080 2848
rect 18052 2796 18104 2848
rect 18144 2796 18196 2848
rect 19984 2873 19993 2907
rect 19993 2873 20027 2907
rect 20027 2873 20036 2907
rect 19984 2864 20036 2873
rect 8982 2694 9034 2746
rect 9046 2694 9098 2746
rect 9110 2694 9162 2746
rect 9174 2694 9226 2746
rect 16982 2694 17034 2746
rect 17046 2694 17098 2746
rect 17110 2694 17162 2746
rect 17174 2694 17226 2746
rect 1860 2592 1912 2644
rect 4988 2592 5040 2644
rect 6368 2635 6420 2644
rect 6368 2601 6377 2635
rect 6377 2601 6411 2635
rect 6411 2601 6420 2635
rect 6368 2592 6420 2601
rect 7472 2635 7524 2644
rect 7472 2601 7481 2635
rect 7481 2601 7515 2635
rect 7515 2601 7524 2635
rect 7472 2592 7524 2601
rect 8392 2592 8444 2644
rect 9588 2592 9640 2644
rect 10600 2635 10652 2644
rect 10600 2601 10609 2635
rect 10609 2601 10643 2635
rect 10643 2601 10652 2635
rect 10600 2592 10652 2601
rect 3424 2524 3476 2576
rect 4528 2524 4580 2576
rect 8300 2524 8352 2576
rect 11520 2592 11572 2644
rect 5080 2456 5132 2508
rect 7656 2499 7708 2508
rect 7656 2465 7665 2499
rect 7665 2465 7699 2499
rect 7699 2465 7708 2499
rect 7656 2456 7708 2465
rect 9680 2499 9732 2508
rect 9680 2465 9689 2499
rect 9689 2465 9723 2499
rect 9723 2465 9732 2499
rect 9680 2456 9732 2465
rect 13636 2635 13688 2644
rect 13636 2601 13645 2635
rect 13645 2601 13679 2635
rect 13679 2601 13688 2635
rect 13636 2592 13688 2601
rect 14372 2592 14424 2644
rect 16396 2635 16448 2644
rect 16396 2601 16405 2635
rect 16405 2601 16439 2635
rect 16439 2601 16448 2635
rect 16396 2592 16448 2601
rect 18052 2592 18104 2644
rect 15660 2524 15712 2576
rect 20812 2592 20864 2644
rect 13268 2456 13320 2508
rect 14188 2499 14240 2508
rect 14188 2465 14197 2499
rect 14197 2465 14231 2499
rect 14231 2465 14240 2499
rect 14188 2456 14240 2465
rect 16028 2456 16080 2508
rect 16212 2499 16264 2508
rect 16212 2465 16221 2499
rect 16221 2465 16255 2499
rect 16255 2465 16264 2499
rect 16212 2456 16264 2465
rect 16856 2456 16908 2508
rect 17132 2499 17184 2508
rect 17132 2465 17141 2499
rect 17141 2465 17175 2499
rect 17175 2465 17184 2499
rect 17132 2456 17184 2465
rect 18604 2499 18656 2508
rect 18604 2465 18613 2499
rect 18613 2465 18647 2499
rect 18647 2465 18656 2499
rect 18604 2456 18656 2465
rect 20444 2456 20496 2508
rect 13728 2388 13780 2440
rect 7104 2320 7156 2372
rect 9220 2320 9272 2372
rect 13268 2320 13320 2372
rect 3148 2252 3200 2304
rect 13728 2252 13780 2304
rect 17868 2388 17920 2440
rect 15936 2320 15988 2372
rect 20628 2320 20680 2372
rect 22652 2320 22704 2372
rect 16212 2252 16264 2304
rect 18604 2252 18656 2304
rect 4982 2150 5034 2202
rect 5046 2150 5098 2202
rect 5110 2150 5162 2202
rect 5174 2150 5226 2202
rect 12982 2150 13034 2202
rect 13046 2150 13098 2202
rect 13110 2150 13162 2202
rect 13174 2150 13226 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
rect 5172 1980 5224 2032
rect 11612 1980 11664 2032
<< metal2 >>
rect 1306 23610 1362 24000
rect 3974 23610 4030 24000
rect 6642 23610 6698 24000
rect 1306 23582 1532 23610
rect 1306 23520 1362 23582
rect 1122 21176 1178 21185
rect 1122 21111 1178 21120
rect 1136 14618 1164 21111
rect 1504 19825 1532 23582
rect 3974 23582 4200 23610
rect 3974 23520 4030 23582
rect 1582 22672 1638 22681
rect 1582 22607 1638 22616
rect 1596 20602 1624 22607
rect 1584 20596 1636 20602
rect 1584 20538 1636 20544
rect 4172 20534 4200 23582
rect 6380 23582 6698 23610
rect 4956 21788 5252 21808
rect 5012 21786 5036 21788
rect 5092 21786 5116 21788
rect 5172 21786 5196 21788
rect 5034 21734 5036 21786
rect 5098 21734 5110 21786
rect 5172 21734 5174 21786
rect 5012 21732 5036 21734
rect 5092 21732 5116 21734
rect 5172 21732 5196 21734
rect 4956 21712 5252 21732
rect 4956 20700 5252 20720
rect 5012 20698 5036 20700
rect 5092 20698 5116 20700
rect 5172 20698 5196 20700
rect 5034 20646 5036 20698
rect 5098 20646 5110 20698
rect 5172 20646 5174 20698
rect 5012 20644 5036 20646
rect 5092 20644 5116 20646
rect 5172 20644 5196 20646
rect 4956 20624 5252 20644
rect 6380 20602 6408 23582
rect 6642 23520 6698 23582
rect 9310 23610 9366 24000
rect 11978 23610 12034 24000
rect 9310 23582 9444 23610
rect 9310 23520 9366 23582
rect 8956 21244 9252 21264
rect 9012 21242 9036 21244
rect 9092 21242 9116 21244
rect 9172 21242 9196 21244
rect 9034 21190 9036 21242
rect 9098 21190 9110 21242
rect 9172 21190 9174 21242
rect 9012 21188 9036 21190
rect 9092 21188 9116 21190
rect 9172 21188 9196 21190
rect 8956 21168 9252 21188
rect 8208 20936 8260 20942
rect 8208 20878 8260 20884
rect 8220 20602 8248 20878
rect 6368 20596 6420 20602
rect 6368 20538 6420 20544
rect 8208 20596 8260 20602
rect 8208 20538 8260 20544
rect 8576 20596 8628 20602
rect 8576 20538 8628 20544
rect 4160 20528 4212 20534
rect 4160 20470 4212 20476
rect 8588 20466 8616 20538
rect 9416 20534 9444 23582
rect 11624 23582 12034 23610
rect 11624 20602 11652 23582
rect 11978 23520 12034 23582
rect 13820 23588 13872 23594
rect 13820 23530 13872 23536
rect 14646 23588 14702 24000
rect 14646 23536 14648 23588
rect 14700 23536 14702 23588
rect 12956 21788 13252 21808
rect 13012 21786 13036 21788
rect 13092 21786 13116 21788
rect 13172 21786 13196 21788
rect 13034 21734 13036 21786
rect 13098 21734 13110 21786
rect 13172 21734 13174 21786
rect 13012 21732 13036 21734
rect 13092 21732 13116 21734
rect 13172 21732 13196 21734
rect 12956 21712 13252 21732
rect 12956 20700 13252 20720
rect 13012 20698 13036 20700
rect 13092 20698 13116 20700
rect 13172 20698 13196 20700
rect 13034 20646 13036 20698
rect 13098 20646 13110 20698
rect 13172 20646 13174 20698
rect 13012 20644 13036 20646
rect 13092 20644 13116 20646
rect 13172 20644 13196 20646
rect 12956 20624 13252 20644
rect 11612 20596 11664 20602
rect 11612 20538 11664 20544
rect 9404 20528 9456 20534
rect 9404 20470 9456 20476
rect 8576 20460 8628 20466
rect 8576 20402 8628 20408
rect 5540 20392 5592 20398
rect 5540 20334 5592 20340
rect 5356 19984 5408 19990
rect 5356 19926 5408 19932
rect 4804 19848 4856 19854
rect 1490 19816 1546 19825
rect 4804 19790 4856 19796
rect 1490 19751 1546 19760
rect 1582 19680 1638 19689
rect 1582 19615 1638 19624
rect 1596 18970 1624 19615
rect 4816 19514 4844 19790
rect 4956 19612 5252 19632
rect 5012 19610 5036 19612
rect 5092 19610 5116 19612
rect 5172 19610 5196 19612
rect 5034 19558 5036 19610
rect 5098 19558 5110 19610
rect 5172 19558 5174 19610
rect 5012 19556 5036 19558
rect 5092 19556 5116 19558
rect 5172 19556 5196 19558
rect 4956 19536 5252 19556
rect 4804 19508 4856 19514
rect 4804 19450 4856 19456
rect 5368 19446 5396 19926
rect 5552 19854 5580 20334
rect 8760 20324 8812 20330
rect 8760 20266 8812 20272
rect 8772 20058 8800 20266
rect 8956 20156 9252 20176
rect 9012 20154 9036 20156
rect 9092 20154 9116 20156
rect 9172 20154 9196 20156
rect 9034 20102 9036 20154
rect 9098 20102 9110 20154
rect 9172 20102 9174 20154
rect 9012 20100 9036 20102
rect 9092 20100 9116 20102
rect 9172 20100 9196 20102
rect 8956 20080 9252 20100
rect 8760 20052 8812 20058
rect 8760 19994 8812 20000
rect 8668 19984 8720 19990
rect 8668 19926 8720 19932
rect 5540 19848 5592 19854
rect 5540 19790 5592 19796
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 5356 19440 5408 19446
rect 5356 19382 5408 19388
rect 3608 19168 3660 19174
rect 3608 19110 3660 19116
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 1584 18964 1636 18970
rect 1584 18906 1636 18912
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 1412 18426 1440 18770
rect 3516 18624 3568 18630
rect 3516 18566 3568 18572
rect 1400 18420 1452 18426
rect 1400 18362 1452 18368
rect 3528 18222 3556 18566
rect 3516 18216 3568 18222
rect 1398 18184 1454 18193
rect 3516 18158 3568 18164
rect 1398 18119 1454 18128
rect 1124 14612 1176 14618
rect 1124 14554 1176 14560
rect 110 14240 166 14249
rect 110 14175 166 14184
rect 124 14074 152 14175
rect 112 14068 164 14074
rect 112 14010 164 14016
rect 1412 13870 1440 18119
rect 3620 18086 3648 19110
rect 2872 18080 2924 18086
rect 2872 18022 2924 18028
rect 3608 18080 3660 18086
rect 3608 18022 3660 18028
rect 2884 17746 2912 18022
rect 4172 17814 4200 19110
rect 4712 18896 4764 18902
rect 4712 18838 4764 18844
rect 4724 18426 4752 18838
rect 5552 18766 5580 19790
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 6460 18964 6512 18970
rect 6460 18906 6512 18912
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 6092 18760 6144 18766
rect 6092 18702 6144 18708
rect 5448 18692 5500 18698
rect 5448 18634 5500 18640
rect 4956 18524 5252 18544
rect 5012 18522 5036 18524
rect 5092 18522 5116 18524
rect 5172 18522 5196 18524
rect 5034 18470 5036 18522
rect 5098 18470 5110 18522
rect 5172 18470 5174 18522
rect 5012 18468 5036 18470
rect 5092 18468 5116 18470
rect 5172 18468 5196 18470
rect 4956 18448 5252 18468
rect 4712 18420 4764 18426
rect 4712 18362 4764 18368
rect 4724 17882 4752 18362
rect 4988 18148 5040 18154
rect 4988 18090 5040 18096
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4712 17876 4764 17882
rect 4712 17818 4764 17824
rect 4160 17808 4212 17814
rect 4160 17750 4212 17756
rect 2596 17740 2648 17746
rect 2596 17682 2648 17688
rect 2872 17740 2924 17746
rect 2872 17682 2924 17688
rect 2608 17270 2636 17682
rect 2596 17264 2648 17270
rect 2596 17206 2648 17212
rect 2608 16998 2636 17206
rect 2884 17066 2912 17682
rect 3148 17672 3200 17678
rect 3148 17614 3200 17620
rect 3160 17338 3188 17614
rect 3148 17332 3200 17338
rect 3148 17274 3200 17280
rect 2872 17060 2924 17066
rect 2872 17002 2924 17008
rect 2596 16992 2648 16998
rect 2516 16952 2596 16980
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1412 13190 1440 13806
rect 2056 13734 2084 14418
rect 2044 13728 2096 13734
rect 2044 13670 2096 13676
rect 1400 13184 1452 13190
rect 1400 13126 1452 13132
rect 1676 13184 1728 13190
rect 1676 13126 1728 13132
rect 1688 12782 1716 13126
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 110 11248 166 11257
rect 110 11183 166 11192
rect 1676 11212 1728 11218
rect 124 11082 152 11183
rect 1676 11154 1728 11160
rect 112 11076 164 11082
rect 112 11018 164 11024
rect 756 11008 808 11014
rect 756 10950 808 10956
rect 110 8256 166 8265
rect 110 8191 166 8200
rect 124 7313 152 8191
rect 110 7304 166 7313
rect 110 7239 166 7248
rect 204 6656 256 6662
rect 204 6598 256 6604
rect 112 5296 164 5302
rect 18 5264 74 5273
rect 74 5244 112 5250
rect 74 5238 164 5244
rect 74 5222 152 5238
rect 18 5199 74 5208
rect 110 2272 166 2281
rect 216 2258 244 6598
rect 768 4185 796 10950
rect 1688 10742 1716 11154
rect 1952 11008 2004 11014
rect 1952 10950 2004 10956
rect 1676 10736 1728 10742
rect 1676 10678 1728 10684
rect 1688 10266 1716 10678
rect 1964 10538 1992 10950
rect 1952 10532 2004 10538
rect 1952 10474 2004 10480
rect 1964 10266 1992 10474
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 1860 10056 1912 10062
rect 2056 10033 2084 13670
rect 2516 12306 2544 16952
rect 2596 16934 2648 16940
rect 2884 16182 2912 17002
rect 4172 16998 4200 17750
rect 4712 17740 4764 17746
rect 4712 17682 4764 17688
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 2872 16176 2924 16182
rect 2872 16118 2924 16124
rect 2780 15632 2832 15638
rect 2780 15574 2832 15580
rect 2792 15162 2820 15574
rect 2884 15570 2912 16118
rect 3792 16040 3844 16046
rect 3792 15982 3844 15988
rect 3804 15910 3832 15982
rect 3792 15904 3844 15910
rect 3792 15846 3844 15852
rect 2872 15564 2924 15570
rect 2872 15506 2924 15512
rect 2780 15156 2832 15162
rect 2780 15098 2832 15104
rect 2884 15094 2912 15506
rect 3148 15496 3200 15502
rect 3148 15438 3200 15444
rect 3054 15192 3110 15201
rect 3160 15162 3188 15438
rect 3054 15127 3110 15136
rect 3148 15156 3200 15162
rect 2872 15088 2924 15094
rect 2872 15030 2924 15036
rect 3068 14958 3096 15127
rect 3148 15098 3200 15104
rect 3804 15065 3832 15846
rect 4172 15706 4200 16934
rect 4252 16652 4304 16658
rect 4252 16594 4304 16600
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 4264 15978 4292 16594
rect 4436 16448 4488 16454
rect 4436 16390 4488 16396
rect 4448 16114 4476 16390
rect 4632 16182 4660 16594
rect 4620 16176 4672 16182
rect 4620 16118 4672 16124
rect 4724 16114 4752 17682
rect 4816 17338 4844 18022
rect 5000 17746 5028 18090
rect 4988 17740 5040 17746
rect 4988 17682 5040 17688
rect 5460 17542 5488 18634
rect 5552 18358 5580 18702
rect 6104 18426 6132 18702
rect 6092 18420 6144 18426
rect 6092 18362 6144 18368
rect 5540 18352 5592 18358
rect 5540 18294 5592 18300
rect 6472 17746 6500 18906
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6748 18290 6776 18770
rect 7668 18630 7696 19246
rect 7852 19174 7880 19790
rect 8576 19304 8628 19310
rect 8576 19246 8628 19252
rect 7840 19168 7892 19174
rect 7840 19110 7892 19116
rect 8588 18834 8616 19246
rect 8680 19174 8708 19926
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 8576 18828 8628 18834
rect 8576 18770 8628 18776
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 7012 18284 7064 18290
rect 7012 18226 7064 18232
rect 6920 18148 6972 18154
rect 6920 18090 6972 18096
rect 6932 17882 6960 18090
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6736 17808 6788 17814
rect 6736 17750 6788 17756
rect 6460 17740 6512 17746
rect 6460 17682 6512 17688
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 4956 17436 5252 17456
rect 5012 17434 5036 17436
rect 5092 17434 5116 17436
rect 5172 17434 5196 17436
rect 5034 17382 5036 17434
rect 5098 17382 5110 17434
rect 5172 17382 5174 17434
rect 5012 17380 5036 17382
rect 5092 17380 5116 17382
rect 5172 17380 5196 17382
rect 4956 17360 5252 17380
rect 4804 17332 4856 17338
rect 4804 17274 4856 17280
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 5276 16726 5304 16934
rect 5264 16720 5316 16726
rect 5264 16662 5316 16668
rect 4956 16348 5252 16368
rect 5012 16346 5036 16348
rect 5092 16346 5116 16348
rect 5172 16346 5196 16348
rect 5034 16294 5036 16346
rect 5098 16294 5110 16346
rect 5172 16294 5174 16346
rect 5012 16292 5036 16294
rect 5092 16292 5116 16294
rect 5172 16292 5196 16294
rect 4956 16272 5252 16292
rect 5356 16176 5408 16182
rect 5356 16118 5408 16124
rect 4436 16108 4488 16114
rect 4436 16050 4488 16056
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 4252 15972 4304 15978
rect 4252 15914 4304 15920
rect 4528 15972 4580 15978
rect 4528 15914 4580 15920
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4172 15162 4200 15642
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 3790 15056 3846 15065
rect 3790 14991 3846 15000
rect 3056 14952 3108 14958
rect 3056 14894 3108 14900
rect 3516 14884 3568 14890
rect 3516 14826 3568 14832
rect 2780 13456 2832 13462
rect 2780 13398 2832 13404
rect 2596 13320 2648 13326
rect 2596 13262 2648 13268
rect 2608 12646 2636 13262
rect 2792 12986 2820 13398
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 3160 12986 3188 13262
rect 2780 12980 2832 12986
rect 2780 12922 2832 12928
rect 3148 12980 3200 12986
rect 3148 12922 3200 12928
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2608 12306 2636 12582
rect 2504 12300 2556 12306
rect 2504 12242 2556 12248
rect 2596 12300 2648 12306
rect 2596 12242 2648 12248
rect 2516 11694 2544 12242
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 2608 11558 2636 12242
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 3160 11762 3188 12174
rect 3148 11756 3200 11762
rect 3148 11698 3200 11704
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2688 11552 2740 11558
rect 2688 11494 2740 11500
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2424 10674 2452 11086
rect 2608 10674 2636 11494
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 2596 10192 2648 10198
rect 2700 10180 2728 11494
rect 3160 11354 3188 11698
rect 3148 11348 3200 11354
rect 3148 11290 3200 11296
rect 2648 10152 2728 10180
rect 2596 10134 2648 10140
rect 1860 9998 1912 10004
rect 2042 10024 2098 10033
rect 1872 9586 1900 9998
rect 2042 9959 2098 9968
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 2136 9512 2188 9518
rect 2136 9454 2188 9460
rect 2228 9512 2280 9518
rect 2228 9454 2280 9460
rect 2148 9042 2176 9454
rect 2240 9178 2268 9454
rect 2608 9382 2636 10134
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 1768 8560 1820 8566
rect 1768 8502 1820 8508
rect 1780 6866 1808 8502
rect 1872 8294 1900 8978
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 1860 8288 1912 8294
rect 1860 8230 1912 8236
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1780 6458 1808 6802
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 754 4176 810 4185
rect 754 4111 810 4120
rect 1872 2650 1900 8230
rect 2056 7410 2084 8434
rect 2424 7886 2452 9114
rect 2504 8356 2556 8362
rect 2504 8298 2556 8304
rect 2516 8090 2544 8298
rect 2608 8294 2636 9318
rect 3528 9081 3556 14826
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3514 9072 3570 9081
rect 2872 9036 2924 9042
rect 3514 9007 3570 9016
rect 2872 8978 2924 8984
rect 2884 8634 2912 8978
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2608 8022 2636 8230
rect 2596 8016 2648 8022
rect 2596 7958 2648 7964
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2424 7546 2452 7822
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 2608 7206 2636 7958
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 2688 6860 2740 6866
rect 2688 6802 2740 6808
rect 2700 6458 2728 6802
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 2976 6254 3004 6598
rect 2964 6248 3016 6254
rect 2870 6216 2926 6225
rect 2964 6190 3016 6196
rect 2870 6151 2926 6160
rect 1952 5160 2004 5166
rect 1950 5128 1952 5137
rect 2004 5128 2006 5137
rect 1950 5063 2006 5072
rect 1964 5030 1992 5063
rect 1952 5024 2004 5030
rect 1952 4966 2004 4972
rect 2884 4690 2912 6151
rect 2976 5030 3004 6190
rect 3160 6118 3188 7142
rect 3528 6866 3556 9007
rect 3620 7936 3648 11630
rect 3804 11082 3832 14991
rect 4172 14822 4200 15098
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 4068 14340 4120 14346
rect 4068 14282 4120 14288
rect 4080 14074 4108 14282
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 4172 13444 4200 14758
rect 4264 13977 4292 15914
rect 4540 15706 4568 15914
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 5000 15706 5028 15846
rect 4528 15700 4580 15706
rect 4528 15642 4580 15648
rect 4988 15700 5040 15706
rect 4988 15642 5040 15648
rect 4540 14890 4568 15642
rect 4956 15260 5252 15280
rect 5012 15258 5036 15260
rect 5092 15258 5116 15260
rect 5172 15258 5196 15260
rect 5034 15206 5036 15258
rect 5098 15206 5110 15258
rect 5172 15206 5174 15258
rect 5012 15204 5036 15206
rect 5092 15204 5116 15206
rect 5172 15204 5196 15206
rect 4956 15184 5252 15204
rect 4528 14884 4580 14890
rect 4528 14826 4580 14832
rect 4540 14618 4568 14826
rect 4528 14612 4580 14618
rect 4528 14554 4580 14560
rect 5368 14482 5396 16118
rect 5460 15094 5488 17478
rect 6472 17338 6500 17682
rect 6460 17332 6512 17338
rect 6460 17274 6512 17280
rect 6748 16998 6776 17750
rect 7024 17542 7052 18226
rect 7104 18148 7156 18154
rect 7104 18090 7156 18096
rect 7116 17542 7144 18090
rect 7194 17640 7250 17649
rect 7194 17575 7250 17584
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 7116 17066 7144 17478
rect 7104 17060 7156 17066
rect 7104 17002 7156 17008
rect 5816 16992 5868 16998
rect 5816 16934 5868 16940
rect 6736 16992 6788 16998
rect 6736 16934 6788 16940
rect 5828 15638 5856 16934
rect 7116 16794 7144 17002
rect 7104 16788 7156 16794
rect 7104 16730 7156 16736
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6184 16448 6236 16454
rect 6184 16390 6236 16396
rect 6196 16250 6224 16390
rect 6380 16250 6408 16526
rect 6184 16244 6236 16250
rect 6184 16186 6236 16192
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 5816 15632 5868 15638
rect 5816 15574 5868 15580
rect 5828 15162 5856 15574
rect 5908 15564 5960 15570
rect 5908 15506 5960 15512
rect 5816 15156 5868 15162
rect 5816 15098 5868 15104
rect 5448 15088 5500 15094
rect 5448 15030 5500 15036
rect 5356 14476 5408 14482
rect 5356 14418 5408 14424
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 4250 13968 4306 13977
rect 4356 13938 4384 14214
rect 4956 14172 5252 14192
rect 5012 14170 5036 14172
rect 5092 14170 5116 14172
rect 5172 14170 5196 14172
rect 5034 14118 5036 14170
rect 5098 14118 5110 14170
rect 5172 14118 5174 14170
rect 5012 14116 5036 14118
rect 5092 14116 5116 14118
rect 5172 14116 5196 14118
rect 4956 14096 5252 14116
rect 4436 14000 4488 14006
rect 4436 13942 4488 13948
rect 4250 13903 4306 13912
rect 4344 13932 4396 13938
rect 4264 13814 4292 13903
rect 4344 13874 4396 13880
rect 4264 13786 4384 13814
rect 4252 13456 4304 13462
rect 4172 13416 4252 13444
rect 4252 13398 4304 13404
rect 3976 12640 4028 12646
rect 3976 12582 4028 12588
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3896 11354 3924 12174
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3792 11076 3844 11082
rect 3792 11018 3844 11024
rect 3700 10600 3752 10606
rect 3700 10542 3752 10548
rect 3712 10470 3740 10542
rect 3700 10464 3752 10470
rect 3700 10406 3752 10412
rect 3712 10266 3740 10406
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3700 7948 3752 7954
rect 3620 7908 3700 7936
rect 3700 7890 3752 7896
rect 3712 7206 3740 7890
rect 3804 7342 3832 11018
rect 3988 9926 4016 12582
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4264 10674 4292 11086
rect 4252 10668 4304 10674
rect 4252 10610 4304 10616
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 3976 9920 4028 9926
rect 3976 9862 4028 9868
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3516 6860 3568 6866
rect 3516 6802 3568 6808
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3160 5574 3188 6054
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2872 4684 2924 4690
rect 2872 4626 2924 4632
rect 2884 4214 2912 4626
rect 2872 4208 2924 4214
rect 2872 4150 2924 4156
rect 3160 3942 3188 5510
rect 3424 5092 3476 5098
rect 3424 5034 3476 5040
rect 3436 4146 3464 5034
rect 3608 4480 3660 4486
rect 3608 4422 3660 4428
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 1860 2644 1912 2650
rect 1860 2586 1912 2592
rect 3160 2310 3188 3878
rect 3436 3738 3464 4082
rect 3620 4078 3648 4422
rect 3608 4072 3660 4078
rect 3608 4014 3660 4020
rect 3712 4010 3740 7142
rect 4080 5574 4108 9998
rect 4172 9518 4200 10542
rect 4264 10266 4292 10610
rect 4356 10470 4384 13786
rect 4448 12238 4476 13942
rect 5368 13802 5396 14418
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5552 13870 5580 14350
rect 5540 13864 5592 13870
rect 5540 13806 5592 13812
rect 4620 13796 4672 13802
rect 4620 13738 4672 13744
rect 5356 13796 5408 13802
rect 5356 13738 5408 13744
rect 4528 13252 4580 13258
rect 4528 13194 4580 13200
rect 4540 12850 4568 13194
rect 4632 13190 4660 13738
rect 5552 13530 5580 13806
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 4632 12714 4660 13126
rect 4956 13084 5252 13104
rect 5012 13082 5036 13084
rect 5092 13082 5116 13084
rect 5172 13082 5196 13084
rect 5034 13030 5036 13082
rect 5098 13030 5110 13082
rect 5172 13030 5174 13082
rect 5012 13028 5036 13030
rect 5092 13028 5116 13030
rect 5172 13028 5196 13030
rect 4956 13008 5252 13028
rect 5460 12986 5488 13126
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 4620 12708 4672 12714
rect 4620 12650 4672 12656
rect 5172 12708 5224 12714
rect 5172 12650 5224 12656
rect 4528 12640 4580 12646
rect 4580 12588 4660 12594
rect 4528 12582 4660 12588
rect 4540 12566 4660 12582
rect 4528 12368 4580 12374
rect 4528 12310 4580 12316
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 4540 11898 4568 12310
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4632 11286 4660 12566
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4724 11762 4752 12174
rect 5184 12170 5212 12650
rect 5920 12306 5948 15506
rect 6000 15496 6052 15502
rect 6000 15438 6052 15444
rect 6012 14822 6040 15438
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 6012 14550 6040 14758
rect 6000 14544 6052 14550
rect 6000 14486 6052 14492
rect 6564 13870 6592 13901
rect 6552 13864 6604 13870
rect 6550 13832 6552 13841
rect 6604 13832 6606 13841
rect 6748 13814 6776 16186
rect 7012 15972 7064 15978
rect 7012 15914 7064 15920
rect 7024 15706 7052 15914
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 7024 15162 7052 15642
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 7024 14890 7052 15098
rect 7012 14884 7064 14890
rect 7012 14826 7064 14832
rect 7208 14482 7236 17575
rect 7288 17060 7340 17066
rect 7288 17002 7340 17008
rect 7300 16182 7328 17002
rect 7668 16182 7696 18566
rect 8208 18352 8260 18358
rect 8208 18294 8260 18300
rect 8116 18080 8168 18086
rect 8116 18022 8168 18028
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 7760 16726 7788 17138
rect 7748 16720 7800 16726
rect 7748 16662 7800 16668
rect 7932 16652 7984 16658
rect 7932 16594 7984 16600
rect 7288 16176 7340 16182
rect 7288 16118 7340 16124
rect 7656 16176 7708 16182
rect 7656 16118 7708 16124
rect 7944 15910 7972 16594
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 7392 15026 7420 15302
rect 7944 15026 7972 15846
rect 8128 15502 8156 18022
rect 8220 17338 8248 18294
rect 8312 17542 8340 18770
rect 8588 18222 8616 18770
rect 8576 18216 8628 18222
rect 8576 18158 8628 18164
rect 8680 18086 8708 19110
rect 8956 19068 9252 19088
rect 9012 19066 9036 19068
rect 9092 19066 9116 19068
rect 9172 19066 9196 19068
rect 9034 19014 9036 19066
rect 9098 19014 9110 19066
rect 9172 19014 9174 19066
rect 9012 19012 9036 19014
rect 9092 19012 9116 19014
rect 9172 19012 9196 19014
rect 8956 18992 9252 19012
rect 8760 18760 8812 18766
rect 8760 18702 8812 18708
rect 8772 18290 8800 18702
rect 8760 18284 8812 18290
rect 8760 18226 8812 18232
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 8680 17814 8708 18022
rect 8772 17882 8800 18226
rect 8956 17980 9252 18000
rect 9012 17978 9036 17980
rect 9092 17978 9116 17980
rect 9172 17978 9196 17980
rect 9034 17926 9036 17978
rect 9098 17926 9110 17978
rect 9172 17926 9174 17978
rect 9012 17924 9036 17926
rect 9092 17924 9116 17926
rect 9172 17924 9196 17926
rect 8956 17904 9252 17924
rect 8760 17876 8812 17882
rect 8760 17818 8812 17824
rect 8668 17808 8720 17814
rect 8390 17776 8446 17785
rect 9416 17785 9444 20470
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 10784 19984 10836 19990
rect 10784 19926 10836 19932
rect 10600 19780 10652 19786
rect 10600 19722 10652 19728
rect 9956 19712 10008 19718
rect 9956 19654 10008 19660
rect 9968 19378 9996 19654
rect 9956 19372 10008 19378
rect 9956 19314 10008 19320
rect 9968 18970 9996 19314
rect 10612 19174 10640 19722
rect 10796 19514 10824 19926
rect 10784 19508 10836 19514
rect 10784 19450 10836 19456
rect 10600 19168 10652 19174
rect 10600 19110 10652 19116
rect 9956 18964 10008 18970
rect 9956 18906 10008 18912
rect 10140 18828 10192 18834
rect 10140 18770 10192 18776
rect 10048 18352 10100 18358
rect 10048 18294 10100 18300
rect 10060 17814 10088 18294
rect 10152 18222 10180 18770
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 10140 18216 10192 18222
rect 10140 18158 10192 18164
rect 10428 18086 10456 18702
rect 10416 18080 10468 18086
rect 10416 18022 10468 18028
rect 10048 17808 10100 17814
rect 8668 17750 8720 17756
rect 9402 17776 9458 17785
rect 8390 17711 8446 17720
rect 8484 17740 8536 17746
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 8312 16561 8340 17478
rect 8404 16658 8432 17711
rect 8484 17682 8536 17688
rect 8496 17338 8524 17682
rect 8484 17332 8536 17338
rect 8536 17292 8616 17320
rect 8484 17274 8536 17280
rect 8392 16652 8444 16658
rect 8392 16594 8444 16600
rect 8298 16552 8354 16561
rect 8298 16487 8354 16496
rect 8404 15910 8432 16594
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 7380 15020 7432 15026
rect 7380 14962 7432 14968
rect 7932 15020 7984 15026
rect 7932 14962 7984 14968
rect 7392 14618 7420 14962
rect 8128 14822 8156 15438
rect 8312 14822 8340 15506
rect 8116 14816 8168 14822
rect 8116 14758 8168 14764
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7012 14476 7064 14482
rect 7012 14418 7064 14424
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 6550 13767 6606 13776
rect 6656 13786 6776 13814
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 6196 12646 6224 13262
rect 6368 12912 6420 12918
rect 6368 12854 6420 12860
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 6196 12442 6224 12582
rect 6184 12436 6236 12442
rect 6184 12378 6236 12384
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 4804 12164 4856 12170
rect 4804 12106 4856 12112
rect 5172 12164 5224 12170
rect 5172 12106 5224 12112
rect 4816 11880 4844 12106
rect 4956 11996 5252 12016
rect 5012 11994 5036 11996
rect 5092 11994 5116 11996
rect 5172 11994 5196 11996
rect 5034 11942 5036 11994
rect 5098 11942 5110 11994
rect 5172 11942 5174 11994
rect 5012 11940 5036 11942
rect 5092 11940 5116 11942
rect 5172 11940 5196 11942
rect 4956 11920 5252 11940
rect 5920 11898 5948 12242
rect 5908 11892 5960 11898
rect 4816 11852 5028 11880
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4620 11280 4672 11286
rect 4620 11222 4672 11228
rect 4632 10588 4660 11222
rect 4724 10742 4752 11698
rect 5000 11626 5028 11852
rect 5908 11834 5960 11840
rect 4988 11620 5040 11626
rect 4988 11562 5040 11568
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4908 11354 4936 11494
rect 5920 11354 5948 11834
rect 6000 11620 6052 11626
rect 6000 11562 6052 11568
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5908 11348 5960 11354
rect 5908 11290 5960 11296
rect 4956 10908 5252 10928
rect 5012 10906 5036 10908
rect 5092 10906 5116 10908
rect 5172 10906 5196 10908
rect 5034 10854 5036 10906
rect 5098 10854 5110 10906
rect 5172 10854 5174 10906
rect 5012 10852 5036 10854
rect 5092 10852 5116 10854
rect 5172 10852 5196 10854
rect 4956 10832 5252 10852
rect 4712 10736 4764 10742
rect 4712 10678 4764 10684
rect 5460 10606 5488 11290
rect 6012 10674 6040 11562
rect 6276 11280 6328 11286
rect 6276 11222 6328 11228
rect 6288 10810 6316 11222
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 5448 10600 5500 10606
rect 4632 10560 4752 10588
rect 4724 10470 4752 10560
rect 5448 10542 5500 10548
rect 5724 10600 5776 10606
rect 5724 10542 5776 10548
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 4528 10464 4580 10470
rect 4712 10464 4764 10470
rect 4580 10424 4660 10452
rect 4528 10406 4580 10412
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4632 9926 4660 10424
rect 4712 10406 4764 10412
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 4724 10198 4752 10406
rect 4712 10192 4764 10198
rect 4712 10134 4764 10140
rect 5092 10130 5120 10406
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 4710 10024 4766 10033
rect 4710 9959 4766 9968
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4632 9518 4660 9862
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4528 9444 4580 9450
rect 4528 9386 4580 9392
rect 4540 9110 4568 9386
rect 4528 9104 4580 9110
rect 4528 9046 4580 9052
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 4264 8498 4292 8978
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4344 8424 4396 8430
rect 4344 8366 4396 8372
rect 4356 8090 4384 8366
rect 4344 8084 4396 8090
rect 4344 8026 4396 8032
rect 4540 7954 4568 9046
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 4540 7546 4568 7890
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4448 6798 4476 7142
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4528 6248 4580 6254
rect 4528 6190 4580 6196
rect 4540 5914 4568 6190
rect 4528 5908 4580 5914
rect 4528 5850 4580 5856
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4528 5772 4580 5778
rect 4528 5714 4580 5720
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4080 5234 4108 5510
rect 4172 5370 4200 5714
rect 4540 5370 4568 5714
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 4540 5166 4568 5306
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 3700 4004 3752 4010
rect 3700 3946 3752 3952
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3436 3058 3464 3674
rect 3712 3641 3740 3946
rect 4436 3664 4488 3670
rect 3698 3632 3754 3641
rect 4436 3606 4488 3612
rect 3698 3567 3754 3576
rect 3424 3052 3476 3058
rect 3424 2994 3476 3000
rect 3436 2582 3464 2994
rect 4448 2836 4476 3606
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4540 3194 4568 3470
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4632 2922 4660 9454
rect 4724 6390 4752 9959
rect 4816 9178 4844 10066
rect 5460 10062 5488 10542
rect 5632 10192 5684 10198
rect 5632 10134 5684 10140
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 4956 9820 5252 9840
rect 5012 9818 5036 9820
rect 5092 9818 5116 9820
rect 5172 9818 5196 9820
rect 5034 9766 5036 9818
rect 5098 9766 5110 9818
rect 5172 9766 5174 9818
rect 5012 9764 5036 9766
rect 5092 9764 5116 9766
rect 5172 9764 5196 9766
rect 4956 9744 5252 9764
rect 5356 9444 5408 9450
rect 5356 9386 5408 9392
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 5368 8974 5396 9386
rect 5644 9364 5672 10134
rect 5736 9586 5764 10542
rect 6276 10192 6328 10198
rect 6276 10134 6328 10140
rect 6288 9722 6316 10134
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5724 9376 5776 9382
rect 5644 9336 5724 9364
rect 5724 9318 5776 9324
rect 5736 9178 5764 9318
rect 5724 9172 5776 9178
rect 5724 9114 5776 9120
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 4956 8732 5252 8752
rect 5012 8730 5036 8732
rect 5092 8730 5116 8732
rect 5172 8730 5196 8732
rect 5034 8678 5036 8730
rect 5098 8678 5110 8730
rect 5172 8678 5174 8730
rect 5012 8676 5036 8678
rect 5092 8676 5116 8678
rect 5172 8676 5196 8678
rect 4956 8656 5252 8676
rect 5368 8634 5396 8910
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5736 8430 5764 9114
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5276 8022 5304 8230
rect 5264 8016 5316 8022
rect 5264 7958 5316 7964
rect 5908 8016 5960 8022
rect 5908 7958 5960 7964
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4816 7410 4844 7686
rect 4956 7644 5252 7664
rect 5012 7642 5036 7644
rect 5092 7642 5116 7644
rect 5172 7642 5196 7644
rect 5034 7590 5036 7642
rect 5098 7590 5110 7642
rect 5172 7590 5174 7642
rect 5012 7588 5036 7590
rect 5092 7588 5116 7590
rect 5172 7588 5196 7590
rect 4956 7568 5252 7588
rect 5920 7546 5948 7958
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6288 7546 6316 7822
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4816 7002 4844 7346
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 4804 6996 4856 7002
rect 4804 6938 4856 6944
rect 5000 6934 5028 7210
rect 4988 6928 5040 6934
rect 4988 6870 5040 6876
rect 5724 6928 5776 6934
rect 5724 6870 5776 6876
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 4712 6384 4764 6390
rect 4712 6326 4764 6332
rect 4816 5914 4844 6734
rect 4956 6556 5252 6576
rect 5012 6554 5036 6556
rect 5092 6554 5116 6556
rect 5172 6554 5196 6556
rect 5034 6502 5036 6554
rect 5098 6502 5110 6554
rect 5172 6502 5174 6554
rect 5012 6500 5036 6502
rect 5092 6500 5116 6502
rect 5172 6500 5196 6502
rect 4956 6480 5252 6500
rect 5736 6458 5764 6870
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 5920 5846 5948 6598
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 6012 5846 6040 6190
rect 5908 5840 5960 5846
rect 5908 5782 5960 5788
rect 6000 5840 6052 5846
rect 6000 5782 6052 5788
rect 4956 5468 5252 5488
rect 5012 5466 5036 5468
rect 5092 5466 5116 5468
rect 5172 5466 5196 5468
rect 5034 5414 5036 5466
rect 5098 5414 5110 5466
rect 5172 5414 5174 5466
rect 5012 5412 5036 5414
rect 5092 5412 5116 5414
rect 5172 5412 5196 5414
rect 4956 5392 5252 5412
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5540 5160 5592 5166
rect 5540 5102 5592 5108
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 4816 4282 4844 4694
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 4956 4380 5252 4400
rect 5012 4378 5036 4380
rect 5092 4378 5116 4380
rect 5172 4378 5196 4380
rect 5034 4326 5036 4378
rect 5098 4326 5110 4378
rect 5172 4326 5174 4378
rect 5012 4324 5036 4326
rect 5092 4324 5116 4326
rect 5172 4324 5196 4326
rect 4956 4304 5252 4324
rect 5368 4282 5396 4490
rect 5552 4486 5580 5102
rect 5644 4826 5672 5170
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5644 4078 5672 4558
rect 5828 4214 5856 5102
rect 5920 4826 5948 5782
rect 6012 5370 6040 5782
rect 6380 5370 6408 12854
rect 6460 12300 6512 12306
rect 6460 12242 6512 12248
rect 6472 11626 6500 12242
rect 6460 11620 6512 11626
rect 6460 11562 6512 11568
rect 6564 9518 6592 13767
rect 6656 10146 6684 13786
rect 7024 13734 7052 14418
rect 7208 14074 7236 14418
rect 7564 14272 7616 14278
rect 7564 14214 7616 14220
rect 7656 14272 7708 14278
rect 7656 14214 7708 14220
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6840 12646 6868 13466
rect 7024 13462 7052 13670
rect 7012 13456 7064 13462
rect 7012 13398 7064 13404
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6748 10674 6776 10950
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6932 10538 6960 10950
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6932 10198 6960 10474
rect 6920 10192 6972 10198
rect 6656 10118 6776 10146
rect 6920 10134 6972 10140
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6656 9110 6684 9998
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 6552 8560 6604 8566
rect 6552 8502 6604 8508
rect 6564 8022 6592 8502
rect 6748 8430 6776 10118
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6932 9110 6960 9454
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6472 6866 6500 7346
rect 6552 7268 6604 7274
rect 6552 7210 6604 7216
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6472 6390 6500 6802
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 6564 5778 6592 7210
rect 6840 7002 6868 8230
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6840 6390 6868 6938
rect 6932 6866 6960 9046
rect 7024 7313 7052 13398
rect 7208 11286 7236 14010
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7484 13530 7512 13874
rect 7576 13802 7604 14214
rect 7668 13938 7696 14214
rect 8128 13938 8156 14758
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 7564 13796 7616 13802
rect 7564 13738 7616 13744
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7576 13394 7604 13738
rect 7564 13388 7616 13394
rect 7564 13330 7616 13336
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7484 12850 7512 13126
rect 7576 12986 7604 13330
rect 8312 13297 8340 14758
rect 8404 14346 8432 15846
rect 8392 14340 8444 14346
rect 8392 14282 8444 14288
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 8298 13288 8354 13297
rect 8298 13223 8354 13232
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7576 12714 7604 12922
rect 7564 12708 7616 12714
rect 7564 12650 7616 12656
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7484 11558 7512 12582
rect 8220 12238 8248 12650
rect 8496 12646 8524 13330
rect 8588 12918 8616 17292
rect 8680 16266 8708 17750
rect 10048 17750 10100 17756
rect 9402 17711 9458 17720
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 9600 17338 9628 17478
rect 10060 17338 10088 17750
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 10048 17332 10100 17338
rect 10048 17274 10100 17280
rect 10428 17270 10456 18022
rect 10612 17610 10640 19110
rect 10784 18624 10836 18630
rect 10784 18566 10836 18572
rect 10796 18358 10824 18566
rect 10784 18352 10836 18358
rect 10784 18294 10836 18300
rect 10796 18154 10824 18294
rect 10692 18148 10744 18154
rect 10692 18090 10744 18096
rect 10784 18148 10836 18154
rect 10784 18090 10836 18096
rect 10600 17604 10652 17610
rect 10600 17546 10652 17552
rect 10416 17264 10468 17270
rect 10416 17206 10468 17212
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 9312 17128 9364 17134
rect 9310 17096 9312 17105
rect 9364 17096 9366 17105
rect 9310 17031 9366 17040
rect 9496 17060 9548 17066
rect 9324 16998 9352 17031
rect 9496 17002 9548 17008
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 8956 16892 9252 16912
rect 9012 16890 9036 16892
rect 9092 16890 9116 16892
rect 9172 16890 9196 16892
rect 9034 16838 9036 16890
rect 9098 16838 9110 16890
rect 9172 16838 9174 16890
rect 9012 16836 9036 16838
rect 9092 16836 9116 16838
rect 9172 16836 9196 16838
rect 8956 16816 9252 16836
rect 9036 16448 9088 16454
rect 9036 16390 9088 16396
rect 8680 16238 8800 16266
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 8680 15638 8708 16050
rect 8772 15978 8800 16238
rect 9048 16114 9076 16390
rect 9324 16250 9352 16934
rect 9508 16454 9536 17002
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 9310 16008 9366 16017
rect 8760 15972 8812 15978
rect 9310 15943 9366 15952
rect 8760 15914 8812 15920
rect 8772 15706 8800 15914
rect 8956 15804 9252 15824
rect 9012 15802 9036 15804
rect 9092 15802 9116 15804
rect 9172 15802 9196 15804
rect 9034 15750 9036 15802
rect 9098 15750 9110 15802
rect 9172 15750 9174 15802
rect 9012 15748 9036 15750
rect 9092 15748 9116 15750
rect 9172 15748 9196 15750
rect 8956 15728 9252 15748
rect 8760 15700 8812 15706
rect 8760 15642 8812 15648
rect 8668 15632 8720 15638
rect 8668 15574 8720 15580
rect 8758 15056 8814 15065
rect 8758 14991 8814 15000
rect 8772 14958 8800 14991
rect 9324 14958 9352 15943
rect 9508 15094 9536 16390
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9784 15162 9812 15438
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9496 15088 9548 15094
rect 9496 15030 9548 15036
rect 8760 14952 8812 14958
rect 8760 14894 8812 14900
rect 9312 14952 9364 14958
rect 9312 14894 9364 14900
rect 8956 14716 9252 14736
rect 9012 14714 9036 14716
rect 9092 14714 9116 14716
rect 9172 14714 9196 14716
rect 9034 14662 9036 14714
rect 9098 14662 9110 14714
rect 9172 14662 9174 14714
rect 9012 14660 9036 14662
rect 9092 14660 9116 14662
rect 9172 14660 9196 14662
rect 8956 14640 9252 14660
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 8760 14000 8812 14006
rect 8760 13942 8812 13948
rect 8576 12912 8628 12918
rect 8576 12854 8628 12860
rect 8772 12850 8800 13942
rect 9324 13870 9352 13901
rect 9312 13864 9364 13870
rect 9310 13832 9312 13841
rect 9364 13832 9366 13841
rect 9692 13802 9720 14350
rect 9310 13767 9366 13776
rect 9680 13796 9732 13802
rect 8956 13628 9252 13648
rect 9012 13626 9036 13628
rect 9092 13626 9116 13628
rect 9172 13626 9196 13628
rect 9034 13574 9036 13626
rect 9098 13574 9110 13626
rect 9172 13574 9174 13626
rect 9012 13572 9036 13574
rect 9092 13572 9116 13574
rect 9172 13572 9196 13574
rect 8956 13552 9252 13572
rect 9324 13530 9352 13767
rect 9680 13738 9732 13744
rect 9692 13530 9720 13738
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9968 13462 9996 17138
rect 10612 17066 10640 17546
rect 10704 17542 10732 18090
rect 10980 17649 11008 20334
rect 11336 20324 11388 20330
rect 11336 20266 11388 20272
rect 11348 19854 11376 20266
rect 11612 20256 11664 20262
rect 11612 20198 11664 20204
rect 13360 20256 13412 20262
rect 13360 20198 13412 20204
rect 11336 19848 11388 19854
rect 11624 19825 11652 20198
rect 11704 19848 11756 19854
rect 11336 19790 11388 19796
rect 11610 19816 11666 19825
rect 11704 19790 11756 19796
rect 11610 19751 11666 19760
rect 11520 18896 11572 18902
rect 11520 18838 11572 18844
rect 11428 18760 11480 18766
rect 11428 18702 11480 18708
rect 11440 18290 11468 18702
rect 11532 18358 11560 18838
rect 11716 18766 11744 19790
rect 12956 19612 13252 19632
rect 13012 19610 13036 19612
rect 13092 19610 13116 19612
rect 13172 19610 13196 19612
rect 13034 19558 13036 19610
rect 13098 19558 13110 19610
rect 13172 19558 13174 19610
rect 13012 19556 13036 19558
rect 13092 19556 13116 19558
rect 13172 19556 13196 19558
rect 12956 19536 13252 19556
rect 11704 18760 11756 18766
rect 11704 18702 11756 18708
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 11520 18352 11572 18358
rect 11520 18294 11572 18300
rect 11428 18284 11480 18290
rect 11428 18226 11480 18232
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 11440 17882 11468 18226
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11152 17672 11204 17678
rect 10966 17640 11022 17649
rect 11152 17614 11204 17620
rect 10966 17575 11022 17584
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10980 17270 11008 17575
rect 11164 17338 11192 17614
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 10876 17264 10928 17270
rect 10876 17206 10928 17212
rect 10968 17264 11020 17270
rect 10968 17206 11020 17212
rect 10600 17060 10652 17066
rect 10600 17002 10652 17008
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 10152 16726 10180 16934
rect 10140 16720 10192 16726
rect 10140 16662 10192 16668
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 10060 15706 10088 16526
rect 10152 16250 10180 16662
rect 10508 16448 10560 16454
rect 10508 16390 10560 16396
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 10060 14618 10088 15506
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 10060 13870 10088 14554
rect 10048 13864 10100 13870
rect 10048 13806 10100 13812
rect 9956 13456 10008 13462
rect 9956 13398 10008 13404
rect 10336 13394 10364 16186
rect 10520 15978 10548 16390
rect 10416 15972 10468 15978
rect 10416 15914 10468 15920
rect 10508 15972 10560 15978
rect 10508 15914 10560 15920
rect 10428 15366 10456 15914
rect 10520 15638 10548 15914
rect 10508 15632 10560 15638
rect 10508 15574 10560 15580
rect 10416 15360 10468 15366
rect 10416 15302 10468 15308
rect 10428 15162 10456 15302
rect 10520 15162 10548 15574
rect 10612 15502 10640 17002
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10508 15156 10560 15162
rect 10508 15098 10560 15104
rect 10414 15056 10470 15065
rect 10414 14991 10470 15000
rect 10428 14958 10456 14991
rect 10416 14952 10468 14958
rect 10416 14894 10468 14900
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8852 12708 8904 12714
rect 8852 12650 8904 12656
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7760 11694 7788 12038
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 7564 11620 7616 11626
rect 7564 11562 7616 11568
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7196 11280 7248 11286
rect 7196 11222 7248 11228
rect 7576 11218 7604 11562
rect 7760 11286 7788 11630
rect 8128 11558 8156 12174
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8128 11354 8156 11494
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7104 11076 7156 11082
rect 7104 11018 7156 11024
rect 7116 10810 7144 11018
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 7576 10742 7604 11154
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 7564 10736 7616 10742
rect 7564 10678 7616 10684
rect 7288 10532 7340 10538
rect 7288 10474 7340 10480
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 7196 9988 7248 9994
rect 7196 9930 7248 9936
rect 7116 9722 7144 9930
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7116 8090 7144 9114
rect 7208 9110 7236 9930
rect 7196 9104 7248 9110
rect 7196 9046 7248 9052
rect 7208 8634 7236 9046
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7300 7886 7328 10474
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7392 8265 7420 8298
rect 7378 8256 7434 8265
rect 7378 8191 7434 8200
rect 7484 8022 7512 8910
rect 7472 8016 7524 8022
rect 7472 7958 7524 7964
rect 7760 7954 7788 11086
rect 8496 10606 8524 12582
rect 8772 12374 8800 12582
rect 8864 12442 8892 12650
rect 10336 12646 10364 13330
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 8956 12540 9252 12560
rect 9012 12538 9036 12540
rect 9092 12538 9116 12540
rect 9172 12538 9196 12540
rect 9034 12486 9036 12538
rect 9098 12486 9110 12538
rect 9172 12486 9174 12538
rect 9012 12484 9036 12486
rect 9092 12484 9116 12486
rect 9172 12484 9196 12486
rect 8956 12464 9252 12484
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8760 12368 8812 12374
rect 8760 12310 8812 12316
rect 8772 11898 8800 12310
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8576 11620 8628 11626
rect 8576 11562 8628 11568
rect 8484 10600 8536 10606
rect 8484 10542 8536 10548
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 7944 10062 7972 10406
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 8022 9072 8078 9081
rect 8022 9007 8078 9016
rect 7840 8424 7892 8430
rect 7840 8366 7892 8372
rect 7852 8090 7880 8366
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7010 7304 7066 7313
rect 7010 7239 7066 7248
rect 7760 7002 7788 7890
rect 8036 7546 8064 9007
rect 8128 7954 8156 9522
rect 8588 9450 8616 11562
rect 9968 11558 9996 12242
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 8956 11452 9252 11472
rect 9012 11450 9036 11452
rect 9092 11450 9116 11452
rect 9172 11450 9196 11452
rect 9034 11398 9036 11450
rect 9098 11398 9110 11450
rect 9172 11398 9174 11450
rect 9012 11396 9036 11398
rect 9092 11396 9116 11398
rect 9172 11396 9196 11398
rect 8956 11376 9252 11396
rect 9312 11212 9364 11218
rect 9312 11154 9364 11160
rect 9324 10810 9352 11154
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 9312 10804 9364 10810
rect 9312 10746 9364 10752
rect 8956 10713 8984 10746
rect 8942 10704 8998 10713
rect 8852 10668 8904 10674
rect 8942 10639 8998 10648
rect 8852 10610 8904 10616
rect 8864 10130 8892 10610
rect 8956 10606 8984 10639
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 8956 10364 9252 10384
rect 9012 10362 9036 10364
rect 9092 10362 9116 10364
rect 9172 10362 9196 10364
rect 9034 10310 9036 10362
rect 9098 10310 9110 10362
rect 9172 10310 9174 10362
rect 9012 10308 9036 10310
rect 9092 10308 9116 10310
rect 9172 10308 9196 10310
rect 8956 10288 9252 10308
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8864 9722 8892 10066
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 8576 9444 8628 9450
rect 8576 9386 8628 9392
rect 8588 9178 8616 9386
rect 8956 9276 9252 9296
rect 9012 9274 9036 9276
rect 9092 9274 9116 9276
rect 9172 9274 9196 9276
rect 9034 9222 9036 9274
rect 9098 9222 9110 9274
rect 9172 9222 9174 9274
rect 9012 9220 9036 9222
rect 9092 9220 9116 9222
rect 9172 9220 9196 9222
rect 8956 9200 9252 9220
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8588 8566 8616 9114
rect 9600 8974 9628 10950
rect 9692 10538 9720 11018
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 9876 10538 9904 10950
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9864 10532 9916 10538
rect 9864 10474 9916 10480
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8588 8294 8616 8502
rect 8576 8288 8628 8294
rect 8576 8230 8628 8236
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 8036 7342 8064 7482
rect 8128 7478 8156 7890
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 8496 7342 8524 7686
rect 8588 7546 8616 8230
rect 8956 8188 9252 8208
rect 9012 8186 9036 8188
rect 9092 8186 9116 8188
rect 9172 8186 9196 8188
rect 9034 8134 9036 8186
rect 9098 8134 9110 8186
rect 9172 8134 9174 8186
rect 9012 8132 9036 8134
rect 9092 8132 9116 8134
rect 9172 8132 9196 8134
rect 8956 8112 9252 8132
rect 9600 8090 9628 8910
rect 9692 8906 9720 10474
rect 9876 10198 9904 10474
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9876 9722 9904 10134
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 9968 9518 9996 11494
rect 10336 11082 10364 12582
rect 10428 11898 10456 14894
rect 10520 14618 10548 15098
rect 10888 14618 10916 17206
rect 11440 16726 11468 17818
rect 11808 17134 11836 18226
rect 12544 18222 12572 18566
rect 12956 18524 13252 18544
rect 13012 18522 13036 18524
rect 13092 18522 13116 18524
rect 13172 18522 13196 18524
rect 13034 18470 13036 18522
rect 13098 18470 13110 18522
rect 13172 18470 13174 18522
rect 13012 18468 13036 18470
rect 13092 18468 13116 18470
rect 13172 18468 13196 18470
rect 12956 18448 13252 18468
rect 12532 18216 12584 18222
rect 12532 18158 12584 18164
rect 12544 17814 12572 18158
rect 12624 18080 12676 18086
rect 12808 18080 12860 18086
rect 12676 18040 12808 18068
rect 12624 18022 12676 18028
rect 12532 17808 12584 17814
rect 12532 17750 12584 17756
rect 11888 17740 11940 17746
rect 11888 17682 11940 17688
rect 12256 17740 12308 17746
rect 12256 17682 12308 17688
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 10968 16720 11020 16726
rect 10968 16662 11020 16668
rect 11428 16720 11480 16726
rect 11428 16662 11480 16668
rect 10980 16182 11008 16662
rect 11242 16552 11298 16561
rect 11242 16487 11298 16496
rect 10968 16176 11020 16182
rect 10968 16118 11020 16124
rect 10508 14612 10560 14618
rect 10508 14554 10560 14560
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10888 13870 10916 14554
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10876 13864 10928 13870
rect 10876 13806 10928 13812
rect 10796 13190 10824 13806
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10888 13530 10916 13670
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10508 12912 10560 12918
rect 10508 12854 10560 12860
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 10520 11830 10548 12854
rect 10796 12850 10824 13126
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 11060 12708 11112 12714
rect 11060 12650 11112 12656
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10704 12102 10732 12582
rect 11072 12442 11100 12650
rect 11060 12436 11112 12442
rect 11060 12378 11112 12384
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 10508 11824 10560 11830
rect 10508 11766 10560 11772
rect 10704 11626 10732 12038
rect 11164 11694 11192 12038
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 10692 11620 10744 11626
rect 10692 11562 10744 11568
rect 11164 11286 11192 11630
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 11256 11218 11284 16487
rect 11796 16448 11848 16454
rect 11900 16436 11928 17682
rect 12268 16998 12296 17682
rect 12530 17640 12586 17649
rect 12530 17575 12586 17584
rect 12440 17060 12492 17066
rect 12440 17002 12492 17008
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 11848 16408 11928 16436
rect 11796 16390 11848 16396
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11624 14550 11652 15846
rect 11612 14544 11664 14550
rect 11612 14486 11664 14492
rect 11624 14074 11652 14486
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11336 13932 11388 13938
rect 11336 13874 11388 13880
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 10324 11076 10376 11082
rect 10324 11018 10376 11024
rect 10336 10810 10364 11018
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10704 10742 10732 11154
rect 11256 10810 11284 11154
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 10232 10736 10284 10742
rect 10232 10678 10284 10684
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 10060 9722 10088 9998
rect 10048 9716 10100 9722
rect 10048 9658 10100 9664
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9876 8362 9904 9046
rect 10152 8498 10180 9318
rect 10244 8974 10272 10678
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10336 8566 10364 10474
rect 11256 10198 11284 10746
rect 11244 10192 11296 10198
rect 11244 10134 11296 10140
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10428 9110 10456 9998
rect 11152 9512 11204 9518
rect 11152 9454 11204 9460
rect 10416 9104 10468 9110
rect 10416 9046 10468 9052
rect 11164 8634 11192 9454
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 9864 8356 9916 8362
rect 9864 8298 9916 8304
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10428 8090 10456 8298
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8588 7342 8616 7482
rect 9968 7449 9996 7890
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10784 7744 10836 7750
rect 10784 7686 10836 7692
rect 9954 7440 10010 7449
rect 9954 7375 9956 7384
rect 10008 7375 10010 7384
rect 9956 7346 10008 7352
rect 8024 7336 8076 7342
rect 8024 7278 8076 7284
rect 8484 7336 8536 7342
rect 8484 7278 8536 7284
rect 8576 7336 8628 7342
rect 9968 7315 9996 7346
rect 8576 7278 8628 7284
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 6828 6384 6880 6390
rect 6828 6326 6880 6332
rect 7208 6322 7236 6734
rect 7196 6316 7248 6322
rect 7248 6276 7328 6304
rect 7196 6258 7248 6264
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6564 5370 6592 5714
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 6000 5364 6052 5370
rect 6000 5306 6052 5312
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6380 5166 6408 5306
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 6564 4622 6592 5306
rect 7208 5234 7236 5510
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 6736 5092 6788 5098
rect 6736 5034 6788 5040
rect 7012 5092 7064 5098
rect 7012 5034 7064 5040
rect 6748 4826 6776 5034
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6748 4622 6776 4762
rect 7024 4758 7052 5034
rect 7012 4752 7064 4758
rect 7012 4694 7064 4700
rect 7300 4622 7328 6276
rect 7576 5914 7604 6802
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7392 5234 7420 5306
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7760 5166 7788 6938
rect 8496 6934 8524 7278
rect 8484 6928 8536 6934
rect 8484 6870 8536 6876
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 7944 6118 7972 6802
rect 8588 6458 8616 7278
rect 8668 7268 8720 7274
rect 8668 7210 8720 7216
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7944 5778 7972 6054
rect 8496 5846 8524 6190
rect 8588 6186 8616 6394
rect 8576 6180 8628 6186
rect 8576 6122 8628 6128
rect 8484 5840 8536 5846
rect 8484 5782 8536 5788
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 8680 5710 8708 7210
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 8956 7100 9252 7120
rect 9012 7098 9036 7100
rect 9092 7098 9116 7100
rect 9172 7098 9196 7100
rect 9034 7046 9036 7098
rect 9098 7046 9110 7098
rect 9172 7046 9174 7098
rect 9012 7044 9036 7046
rect 9092 7044 9116 7046
rect 9172 7044 9196 7046
rect 8956 7024 9252 7044
rect 9692 7002 9720 7142
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9692 6458 9720 6938
rect 10336 6934 10364 7686
rect 10796 7410 10824 7686
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10324 6928 10376 6934
rect 10376 6888 10456 6916
rect 10324 6870 10376 6876
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 10336 6322 10364 6598
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 8956 6012 9252 6032
rect 9012 6010 9036 6012
rect 9092 6010 9116 6012
rect 9172 6010 9196 6012
rect 9034 5958 9036 6010
rect 9098 5958 9110 6010
rect 9172 5958 9174 6010
rect 9012 5956 9036 5958
rect 9092 5956 9116 5958
rect 9172 5956 9196 5958
rect 8956 5936 9252 5956
rect 10060 5846 10088 6190
rect 10428 5914 10456 6888
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 10612 5846 10640 6734
rect 10980 6322 11008 7346
rect 11164 6934 11192 8570
rect 11348 7954 11376 13874
rect 11624 13870 11652 14010
rect 11808 13977 11836 16390
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 11794 13968 11850 13977
rect 11794 13903 11850 13912
rect 11612 13864 11664 13870
rect 11612 13806 11664 13812
rect 11428 13728 11480 13734
rect 11428 13670 11480 13676
rect 11440 12782 11468 13670
rect 11624 13530 11652 13806
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11428 12776 11480 12782
rect 11428 12718 11480 12724
rect 11624 12646 11652 13466
rect 11808 12782 11836 13903
rect 11992 13734 12020 14350
rect 11980 13728 12032 13734
rect 11980 13670 12032 13676
rect 12176 13530 12204 14758
rect 12268 14006 12296 16934
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 12360 15910 12388 16526
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 12452 15706 12480 17002
rect 12544 16046 12572 17575
rect 12728 16794 12756 18040
rect 12808 18022 12860 18028
rect 13268 17604 13320 17610
rect 13268 17546 13320 17552
rect 12808 17536 12860 17542
rect 12808 17478 12860 17484
rect 12820 17066 12848 17478
rect 12956 17436 13252 17456
rect 13012 17434 13036 17436
rect 13092 17434 13116 17436
rect 13172 17434 13196 17436
rect 13034 17382 13036 17434
rect 13098 17382 13110 17434
rect 13172 17382 13174 17434
rect 13012 17380 13036 17382
rect 13092 17380 13116 17382
rect 13172 17380 13196 17382
rect 12956 17360 13252 17380
rect 13280 17066 13308 17546
rect 13372 17270 13400 20198
rect 13360 17264 13412 17270
rect 13360 17206 13412 17212
rect 12808 17060 12860 17066
rect 12808 17002 12860 17008
rect 13268 17060 13320 17066
rect 13268 17002 13320 17008
rect 13280 16794 13308 17002
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 12728 16114 12756 16730
rect 12956 16348 13252 16368
rect 13012 16346 13036 16348
rect 13092 16346 13116 16348
rect 13172 16346 13196 16348
rect 13034 16294 13036 16346
rect 13098 16294 13110 16346
rect 13172 16294 13174 16346
rect 13012 16292 13036 16294
rect 13092 16292 13116 16294
rect 13172 16292 13196 16294
rect 12956 16272 13252 16292
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12532 16040 12584 16046
rect 12532 15982 12584 15988
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 13280 15434 13308 15982
rect 13268 15428 13320 15434
rect 13268 15370 13320 15376
rect 12956 15260 13252 15280
rect 13012 15258 13036 15260
rect 13092 15258 13116 15260
rect 13172 15258 13196 15260
rect 13034 15206 13036 15258
rect 13098 15206 13110 15258
rect 13172 15206 13174 15258
rect 13012 15204 13036 15206
rect 13092 15204 13116 15206
rect 13172 15204 13196 15206
rect 12956 15184 13252 15204
rect 12532 14884 12584 14890
rect 12532 14826 12584 14832
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 12256 14000 12308 14006
rect 12256 13942 12308 13948
rect 12164 13524 12216 13530
rect 12164 13466 12216 13472
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11808 12374 11836 12582
rect 11796 12368 11848 12374
rect 11796 12310 11848 12316
rect 11808 11898 11836 12310
rect 12164 12232 12216 12238
rect 12164 12174 12216 12180
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 12176 11558 12204 12174
rect 12164 11552 12216 11558
rect 12164 11494 12216 11500
rect 12176 10810 12204 11494
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 11348 7546 11376 7890
rect 11336 7540 11388 7546
rect 11336 7482 11388 7488
rect 11152 6928 11204 6934
rect 11152 6870 11204 6876
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10048 5840 10100 5846
rect 10600 5840 10652 5846
rect 10048 5782 10100 5788
rect 10520 5800 10600 5828
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7852 4826 7880 5646
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8404 4826 8432 5102
rect 8496 5030 8524 5646
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 7840 4820 7892 4826
rect 8392 4820 8444 4826
rect 7840 4762 7892 4768
rect 8312 4780 8392 4808
rect 7748 4752 7800 4758
rect 7748 4694 7800 4700
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 6368 4548 6420 4554
rect 6368 4490 6420 4496
rect 5816 4208 5868 4214
rect 5816 4150 5868 4156
rect 5632 4072 5684 4078
rect 5632 4014 5684 4020
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5552 3670 5580 3878
rect 5644 3670 5672 4014
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 5632 3664 5684 3670
rect 5632 3606 5684 3612
rect 5644 3466 5672 3606
rect 5632 3460 5684 3466
rect 5632 3402 5684 3408
rect 4956 3292 5252 3312
rect 5012 3290 5036 3292
rect 5092 3290 5116 3292
rect 5172 3290 5196 3292
rect 5034 3238 5036 3290
rect 5098 3238 5110 3290
rect 5172 3238 5174 3290
rect 5012 3236 5036 3238
rect 5092 3236 5116 3238
rect 5172 3236 5196 3238
rect 4956 3216 5252 3236
rect 5644 3058 5672 3402
rect 6288 3194 6316 3674
rect 6380 3534 6408 4490
rect 7760 4282 7788 4694
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 8312 4214 8340 4780
rect 8392 4762 8444 4768
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 8404 4282 8432 4626
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8300 4208 8352 4214
rect 8300 4150 8352 4156
rect 8312 4078 8340 4150
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 7472 4004 7524 4010
rect 7472 3946 7524 3952
rect 6368 3528 6420 3534
rect 6368 3470 6420 3476
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 4620 2916 4672 2922
rect 4620 2858 4672 2864
rect 4988 2916 5040 2922
rect 4988 2858 5040 2864
rect 5080 2916 5132 2922
rect 5080 2858 5132 2864
rect 4528 2848 4580 2854
rect 4448 2808 4528 2836
rect 4528 2790 4580 2796
rect 4540 2582 4568 2790
rect 5000 2650 5028 2858
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 3424 2576 3476 2582
rect 3424 2518 3476 2524
rect 4528 2576 4580 2582
rect 4528 2518 4580 2524
rect 5092 2514 5120 2858
rect 6380 2650 6408 3470
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 5080 2508 5132 2514
rect 5080 2450 5132 2456
rect 166 2230 244 2258
rect 3148 2304 3200 2310
rect 3148 2246 3200 2252
rect 110 2207 166 2216
rect 1214 2000 1270 2009
rect 1214 1935 1270 1944
rect 938 82 994 480
rect 1228 82 1256 1935
rect 938 54 1256 82
rect 2870 82 2926 480
rect 3160 82 3188 2246
rect 4956 2204 5252 2224
rect 5012 2202 5036 2204
rect 5092 2202 5116 2204
rect 5172 2202 5196 2204
rect 5034 2150 5036 2202
rect 5098 2150 5110 2202
rect 5172 2150 5174 2202
rect 5012 2148 5036 2150
rect 5092 2148 5116 2150
rect 5172 2148 5196 2150
rect 4956 2128 5252 2148
rect 5172 2032 5224 2038
rect 5172 1974 5224 1980
rect 2870 54 3188 82
rect 4894 82 4950 480
rect 5184 82 5212 1974
rect 4894 54 5212 82
rect 6656 82 6684 3946
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7392 3738 7420 3878
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7116 2378 7144 2926
rect 7484 2650 7512 3946
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7668 2514 7696 3674
rect 8496 3602 8524 4966
rect 8956 4924 9252 4944
rect 9012 4922 9036 4924
rect 9092 4922 9116 4924
rect 9172 4922 9196 4924
rect 9034 4870 9036 4922
rect 9098 4870 9110 4922
rect 9172 4870 9174 4922
rect 9012 4868 9036 4870
rect 9092 4868 9116 4870
rect 9172 4868 9196 4870
rect 8956 4848 9252 4868
rect 9416 4758 9444 5646
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 9404 4752 9456 4758
rect 9404 4694 9456 4700
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9324 4078 9352 4218
rect 9508 4146 9536 5578
rect 10060 5370 10088 5782
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 9588 5092 9640 5098
rect 9588 5034 9640 5040
rect 10324 5092 10376 5098
rect 10324 5034 10376 5040
rect 9600 4690 9628 5034
rect 10336 4826 10364 5034
rect 10324 4820 10376 4826
rect 10324 4762 10376 4768
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9600 4282 9628 4626
rect 9678 4312 9734 4321
rect 9588 4276 9640 4282
rect 9678 4247 9734 4256
rect 9588 4218 9640 4224
rect 9692 4214 9720 4247
rect 9680 4208 9732 4214
rect 9680 4150 9732 4156
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 8956 3836 9252 3856
rect 9012 3834 9036 3836
rect 9092 3834 9116 3836
rect 9172 3834 9196 3836
rect 9034 3782 9036 3834
rect 9098 3782 9110 3834
rect 9172 3782 9174 3834
rect 9012 3780 9036 3782
rect 9092 3780 9116 3782
rect 9172 3780 9196 3782
rect 8956 3760 9252 3780
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8128 2990 8156 3538
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 7656 2508 7708 2514
rect 7656 2450 7708 2456
rect 8128 2417 8156 2926
rect 8404 2922 8432 3334
rect 8496 3194 8524 3538
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 9416 3126 9444 3946
rect 9508 3738 9536 4082
rect 9784 4010 9812 4694
rect 10520 4554 10548 5800
rect 10600 5782 10652 5788
rect 10980 5234 11008 6258
rect 11244 5296 11296 5302
rect 11244 5238 11296 5244
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10600 5024 10652 5030
rect 10600 4966 10652 4972
rect 10612 4690 10640 4966
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10508 4548 10560 4554
rect 10508 4490 10560 4496
rect 10520 4154 10548 4490
rect 10520 4146 10640 4154
rect 10520 4140 10652 4146
rect 10520 4126 10600 4140
rect 10600 4082 10652 4088
rect 9772 4004 9824 4010
rect 9772 3946 9824 3952
rect 10612 3738 10640 4082
rect 10876 4004 10928 4010
rect 10876 3946 10928 3952
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 9586 3632 9642 3641
rect 9586 3567 9642 3576
rect 9600 3534 9628 3567
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 8300 2916 8352 2922
rect 8300 2858 8352 2864
rect 8392 2916 8444 2922
rect 8392 2858 8444 2864
rect 8312 2582 8340 2858
rect 8404 2650 8432 2858
rect 8956 2748 9252 2768
rect 9012 2746 9036 2748
rect 9092 2746 9116 2748
rect 9172 2746 9196 2748
rect 9034 2694 9036 2746
rect 9098 2694 9110 2746
rect 9172 2694 9174 2746
rect 9012 2692 9036 2694
rect 9092 2692 9116 2694
rect 9172 2692 9196 2694
rect 8956 2672 9252 2692
rect 9600 2650 9628 3470
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9692 3058 9720 3402
rect 9968 3058 9996 3674
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10244 3194 10272 3538
rect 10888 3194 10916 3946
rect 10980 3738 11008 5170
rect 11256 4826 11284 5238
rect 11244 4820 11296 4826
rect 11244 4762 11296 4768
rect 11256 4622 11284 4762
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11440 4321 11468 10406
rect 11808 9586 11836 10406
rect 12268 10266 12296 13942
rect 12360 13462 12388 14214
rect 12348 13456 12400 13462
rect 12348 13398 12400 13404
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12452 12696 12480 13126
rect 12544 12918 12572 14826
rect 13280 14482 13308 15370
rect 13372 14890 13400 17206
rect 13832 16250 13860 23530
rect 14646 23520 14702 23536
rect 17314 23610 17370 24000
rect 19982 23610 20038 24000
rect 22650 23610 22706 24000
rect 17314 23582 17540 23610
rect 17314 23520 17370 23582
rect 14660 23499 14688 23520
rect 16956 21244 17252 21264
rect 17012 21242 17036 21244
rect 17092 21242 17116 21244
rect 17172 21242 17196 21244
rect 17034 21190 17036 21242
rect 17098 21190 17110 21242
rect 17172 21190 17174 21242
rect 17012 21188 17036 21190
rect 17092 21188 17116 21190
rect 17172 21188 17196 21190
rect 16956 21168 17252 21188
rect 16956 20156 17252 20176
rect 17012 20154 17036 20156
rect 17092 20154 17116 20156
rect 17172 20154 17196 20156
rect 17034 20102 17036 20154
rect 17098 20102 17110 20154
rect 17172 20102 17174 20154
rect 17012 20100 17036 20102
rect 17092 20100 17116 20102
rect 17172 20100 17196 20102
rect 16956 20080 17252 20100
rect 16672 19304 16724 19310
rect 16672 19246 16724 19252
rect 17316 19304 17368 19310
rect 17316 19246 17368 19252
rect 16212 19168 16264 19174
rect 16212 19110 16264 19116
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 14188 18352 14240 18358
rect 14188 18294 14240 18300
rect 13910 17776 13966 17785
rect 14200 17746 14228 18294
rect 15212 18290 15240 18770
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15200 18284 15252 18290
rect 15200 18226 15252 18232
rect 15016 18148 15068 18154
rect 15016 18090 15068 18096
rect 15028 17882 15056 18090
rect 15016 17876 15068 17882
rect 15016 17818 15068 17824
rect 13910 17711 13966 17720
rect 14004 17740 14056 17746
rect 13924 16658 13952 17711
rect 14188 17740 14240 17746
rect 14056 17700 14136 17728
rect 14004 17682 14056 17688
rect 14004 17060 14056 17066
rect 14004 17002 14056 17008
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13924 16250 13952 16594
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13912 16244 13964 16250
rect 13912 16186 13964 16192
rect 13820 15564 13872 15570
rect 14016 15552 14044 17002
rect 14108 16998 14136 17700
rect 14188 17682 14240 17688
rect 14200 17066 14228 17682
rect 15028 17338 15056 17818
rect 15292 17808 15344 17814
rect 15292 17750 15344 17756
rect 15016 17332 15068 17338
rect 15016 17274 15068 17280
rect 15108 17264 15160 17270
rect 15108 17206 15160 17212
rect 14188 17060 14240 17066
rect 14188 17002 14240 17008
rect 14096 16992 14148 16998
rect 14096 16934 14148 16940
rect 14108 16561 14136 16934
rect 14094 16552 14150 16561
rect 14094 16487 14150 16496
rect 14832 16040 14884 16046
rect 14832 15982 14884 15988
rect 14844 15638 14872 15982
rect 14832 15632 14884 15638
rect 14832 15574 14884 15580
rect 14096 15564 14148 15570
rect 14016 15524 14096 15552
rect 13820 15506 13872 15512
rect 14096 15506 14148 15512
rect 13360 14884 13412 14890
rect 13360 14826 13412 14832
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 12956 14172 13252 14192
rect 13012 14170 13036 14172
rect 13092 14170 13116 14172
rect 13172 14170 13196 14172
rect 13034 14118 13036 14170
rect 13098 14118 13110 14170
rect 13172 14118 13174 14170
rect 13012 14116 13036 14118
rect 13092 14116 13116 14118
rect 13172 14116 13196 14118
rect 12956 14096 13252 14116
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12532 12912 12584 12918
rect 12532 12854 12584 12860
rect 12532 12708 12584 12714
rect 12452 12668 12532 12696
rect 12532 12650 12584 12656
rect 12348 10532 12400 10538
rect 12348 10474 12400 10480
rect 12256 10260 12308 10266
rect 12256 10202 12308 10208
rect 12360 10130 12388 10474
rect 11980 10124 12032 10130
rect 11900 10084 11980 10112
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11900 9518 11928 10084
rect 11980 10066 12032 10072
rect 12348 10124 12400 10130
rect 12348 10066 12400 10072
rect 12072 9988 12124 9994
rect 12072 9930 12124 9936
rect 12084 9654 12112 9930
rect 12544 9722 12572 12650
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12072 9648 12124 9654
rect 12072 9590 12124 9596
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 11900 9042 11928 9454
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11520 8900 11572 8906
rect 11520 8842 11572 8848
rect 11532 8634 11560 8842
rect 11900 8838 11928 8978
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11532 6458 11560 8570
rect 11900 7732 11928 8774
rect 11992 8634 12020 8978
rect 12084 8634 12112 9590
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 11992 8090 12020 8570
rect 12636 8090 12664 13670
rect 13372 13326 13400 14826
rect 13832 14822 13860 15506
rect 14108 15162 14136 15506
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 15016 15156 15068 15162
rect 15016 15098 15068 15104
rect 14108 14890 14136 15098
rect 15028 15026 15056 15098
rect 15120 15094 15148 17206
rect 15304 16998 15332 17750
rect 15580 17202 15608 18566
rect 16224 18358 16252 19110
rect 16684 18630 16712 19246
rect 16956 19068 17252 19088
rect 17012 19066 17036 19068
rect 17092 19066 17116 19068
rect 17172 19066 17196 19068
rect 17034 19014 17036 19066
rect 17098 19014 17110 19066
rect 17172 19014 17174 19066
rect 17012 19012 17036 19014
rect 17092 19012 17116 19014
rect 17172 19012 17196 19014
rect 16956 18992 17252 19012
rect 17328 18902 17356 19246
rect 17408 19236 17460 19242
rect 17408 19178 17460 19184
rect 17316 18896 17368 18902
rect 17316 18838 17368 18844
rect 16856 18828 16908 18834
rect 16856 18770 16908 18776
rect 17040 18828 17092 18834
rect 17040 18770 17092 18776
rect 16672 18624 16724 18630
rect 16672 18566 16724 18572
rect 16212 18352 16264 18358
rect 16212 18294 16264 18300
rect 16028 18148 16080 18154
rect 16028 18090 16080 18096
rect 15752 18080 15804 18086
rect 15752 18022 15804 18028
rect 15568 17196 15620 17202
rect 15568 17138 15620 17144
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 15200 16448 15252 16454
rect 15200 16390 15252 16396
rect 15212 15502 15240 16390
rect 15304 15978 15332 16934
rect 15580 16794 15608 17138
rect 15764 17066 15792 18022
rect 15752 17060 15804 17066
rect 15752 17002 15804 17008
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 15764 16454 15792 17002
rect 15844 16720 15896 16726
rect 15844 16662 15896 16668
rect 15752 16448 15804 16454
rect 15752 16390 15804 16396
rect 15292 15972 15344 15978
rect 15292 15914 15344 15920
rect 15856 15910 15884 16662
rect 16040 16454 16068 18090
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 16224 17882 16252 18022
rect 16212 17876 16264 17882
rect 16212 17818 16264 17824
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 16500 17338 16528 17614
rect 16580 17536 16632 17542
rect 16580 17478 16632 17484
rect 16488 17332 16540 17338
rect 16488 17274 16540 17280
rect 16212 17060 16264 17066
rect 16212 17002 16264 17008
rect 16224 16522 16252 17002
rect 16592 16590 16620 17478
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16212 16516 16264 16522
rect 16212 16458 16264 16464
rect 16028 16448 16080 16454
rect 16028 16390 16080 16396
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15844 15904 15896 15910
rect 15844 15846 15896 15852
rect 15396 15638 15424 15846
rect 16040 15638 16068 16390
rect 16592 16250 16620 16526
rect 16580 16244 16632 16250
rect 16580 16186 16632 16192
rect 15384 15632 15436 15638
rect 15384 15574 15436 15580
rect 16028 15632 16080 15638
rect 16028 15574 16080 15580
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 15212 15094 15240 15438
rect 15396 15162 15424 15574
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 15108 15088 15160 15094
rect 15108 15030 15160 15036
rect 15200 15088 15252 15094
rect 15200 15030 15252 15036
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 14096 14884 14148 14890
rect 14372 14884 14424 14890
rect 14096 14826 14148 14832
rect 14292 14844 14372 14872
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13636 14476 13688 14482
rect 13636 14418 13688 14424
rect 13648 13841 13676 14418
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13740 13938 13768 14350
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 13634 13832 13690 13841
rect 13634 13767 13690 13776
rect 13648 13734 13676 13767
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13740 13530 13768 13874
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13452 13456 13504 13462
rect 13452 13398 13504 13404
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 12820 12374 12848 13262
rect 12956 13084 13252 13104
rect 13012 13082 13036 13084
rect 13092 13082 13116 13084
rect 13172 13082 13196 13084
rect 13034 13030 13036 13082
rect 13098 13030 13110 13082
rect 13172 13030 13174 13082
rect 13012 13028 13036 13030
rect 13092 13028 13116 13030
rect 13172 13028 13196 13030
rect 12956 13008 13252 13028
rect 13464 12986 13492 13398
rect 13832 13297 13860 14758
rect 14004 14340 14056 14346
rect 14004 14282 14056 14288
rect 13818 13288 13874 13297
rect 13818 13223 13874 13232
rect 13912 13252 13964 13258
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 12808 12368 12860 12374
rect 12714 12336 12770 12345
rect 12808 12310 12860 12316
rect 12714 12271 12770 12280
rect 12728 11694 12756 12271
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 12956 11996 13252 12016
rect 13012 11994 13036 11996
rect 13092 11994 13116 11996
rect 13172 11994 13196 11996
rect 13034 11942 13036 11994
rect 13098 11942 13110 11994
rect 13172 11942 13174 11994
rect 13012 11940 13036 11942
rect 13092 11940 13116 11942
rect 13172 11940 13196 11942
rect 12956 11920 13252 11940
rect 13464 11694 13492 12038
rect 13740 11762 13768 12174
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12624 7948 12676 7954
rect 12624 7890 12676 7896
rect 11980 7744 12032 7750
rect 11900 7704 11980 7732
rect 11980 7686 12032 7692
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11704 6180 11756 6186
rect 11704 6122 11756 6128
rect 11716 5778 11744 6122
rect 11704 5772 11756 5778
rect 11624 5732 11704 5760
rect 11624 5030 11652 5732
rect 11704 5714 11756 5720
rect 11808 5642 11836 6394
rect 11900 6390 11928 6802
rect 11888 6384 11940 6390
rect 11888 6326 11940 6332
rect 11796 5636 11848 5642
rect 11796 5578 11848 5584
rect 11808 5370 11836 5578
rect 11992 5574 12020 7686
rect 12636 7342 12664 7890
rect 12624 7336 12676 7342
rect 12624 7278 12676 7284
rect 12636 6662 12664 7278
rect 12728 7274 12756 11630
rect 13464 11286 13492 11630
rect 13740 11286 13768 11698
rect 13452 11280 13504 11286
rect 13452 11222 13504 11228
rect 13728 11280 13780 11286
rect 13728 11222 13780 11228
rect 13832 11200 13860 13223
rect 13912 13194 13964 13200
rect 13924 12850 13952 13194
rect 14016 13190 14044 14282
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 14016 12986 14044 13126
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13924 12374 13952 12582
rect 13912 12368 13964 12374
rect 13912 12310 13964 12316
rect 13912 11212 13964 11218
rect 13832 11172 13912 11200
rect 13912 11154 13964 11160
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12820 10742 12848 11086
rect 12956 10908 13252 10928
rect 13012 10906 13036 10908
rect 13092 10906 13116 10908
rect 13172 10906 13196 10908
rect 13034 10854 13036 10906
rect 13098 10854 13110 10906
rect 13172 10854 13174 10906
rect 13012 10852 13036 10854
rect 13092 10852 13116 10854
rect 13172 10852 13196 10854
rect 12956 10832 13252 10852
rect 12808 10736 12860 10742
rect 12808 10678 12860 10684
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 12820 9382 12848 10678
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13004 10130 13032 10542
rect 13280 10266 13308 10542
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 12956 9820 13252 9840
rect 13012 9818 13036 9820
rect 13092 9818 13116 9820
rect 13172 9818 13196 9820
rect 13034 9766 13036 9818
rect 13098 9766 13110 9818
rect 13172 9766 13174 9818
rect 13012 9764 13036 9766
rect 13092 9764 13116 9766
rect 13172 9764 13196 9766
rect 12956 9744 13252 9764
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12912 9178 12940 9522
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 13280 9110 13308 10202
rect 13268 9104 13320 9110
rect 13268 9046 13320 9052
rect 13372 8906 13400 10678
rect 13452 10192 13504 10198
rect 13452 10134 13504 10140
rect 13464 9654 13492 10134
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13452 9648 13504 9654
rect 13452 9590 13504 9596
rect 13556 9518 13584 9862
rect 13740 9586 13768 9930
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13556 9042 13584 9454
rect 13636 9444 13688 9450
rect 13636 9386 13688 9392
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13360 8900 13412 8906
rect 13360 8842 13412 8848
rect 12956 8732 13252 8752
rect 13012 8730 13036 8732
rect 13092 8730 13116 8732
rect 13172 8730 13196 8732
rect 13034 8678 13036 8730
rect 13098 8678 13110 8730
rect 13172 8678 13174 8730
rect 13012 8676 13036 8678
rect 13092 8676 13116 8678
rect 13172 8676 13196 8678
rect 12956 8656 13252 8676
rect 13372 8498 13400 8842
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 12808 8424 12860 8430
rect 12808 8366 12860 8372
rect 12820 7750 12848 8366
rect 13556 8276 13584 8978
rect 13648 8945 13676 9386
rect 13740 8974 13768 9522
rect 13728 8968 13780 8974
rect 13634 8936 13690 8945
rect 13728 8910 13780 8916
rect 13634 8871 13690 8880
rect 13636 8288 13688 8294
rect 13556 8248 13636 8276
rect 13636 8230 13688 8236
rect 13360 7812 13412 7818
rect 13360 7754 13412 7760
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12820 7546 12848 7686
rect 12956 7644 13252 7664
rect 13012 7642 13036 7644
rect 13092 7642 13116 7644
rect 13172 7642 13196 7644
rect 13034 7590 13036 7642
rect 13098 7590 13110 7642
rect 13172 7590 13174 7642
rect 13012 7588 13036 7590
rect 13092 7588 13116 7590
rect 13172 7588 13196 7590
rect 12956 7568 13252 7588
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 13372 7410 13400 7754
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 13360 7404 13412 7410
rect 13360 7346 13412 7352
rect 12716 7268 12768 7274
rect 12716 7210 12768 7216
rect 12728 7154 12756 7210
rect 12728 7126 12848 7154
rect 12820 6866 12848 7126
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12808 6656 12860 6662
rect 12912 6644 12940 7346
rect 13556 7342 13584 7686
rect 13648 7410 13676 8230
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13740 7449 13768 7482
rect 13726 7440 13782 7449
rect 13636 7404 13688 7410
rect 13726 7375 13782 7384
rect 13636 7346 13688 7352
rect 13544 7336 13596 7342
rect 13544 7278 13596 7284
rect 13648 6730 13676 7346
rect 13924 6866 13952 11154
rect 14016 11150 14044 12922
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 14108 10266 14136 14826
rect 14292 14278 14320 14844
rect 14372 14826 14424 14832
rect 14464 14816 14516 14822
rect 14464 14758 14516 14764
rect 14476 14278 14504 14758
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 14292 14006 14320 14214
rect 14476 14074 14504 14214
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 14372 12368 14424 12374
rect 14372 12310 14424 12316
rect 14384 11558 14412 12310
rect 14568 12238 14596 14962
rect 16408 14958 16436 15302
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 15580 14482 15608 14894
rect 16304 14816 16356 14822
rect 16304 14758 16356 14764
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 14832 13796 14884 13802
rect 14832 13738 14884 13744
rect 15108 13796 15160 13802
rect 15108 13738 15160 13744
rect 14844 12782 14872 13738
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 15120 12714 15148 13738
rect 15212 13734 15240 14418
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 15568 14000 15620 14006
rect 15568 13942 15620 13948
rect 15580 13802 15608 13942
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15200 13728 15252 13734
rect 15200 13670 15252 13676
rect 15384 13728 15436 13734
rect 15436 13688 15516 13716
rect 15384 13670 15436 13676
rect 15108 12708 15160 12714
rect 15108 12650 15160 12656
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14384 11354 14412 11494
rect 14372 11348 14424 11354
rect 14372 11290 14424 11296
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14188 11076 14240 11082
rect 14188 11018 14240 11024
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 14016 9518 14044 9998
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 13268 6724 13320 6730
rect 13268 6666 13320 6672
rect 13636 6724 13688 6730
rect 13636 6666 13688 6672
rect 12860 6616 12940 6644
rect 12808 6598 12860 6604
rect 12636 6254 12664 6598
rect 12716 6384 12768 6390
rect 12820 6372 12848 6598
rect 12956 6556 13252 6576
rect 13012 6554 13036 6556
rect 13092 6554 13116 6556
rect 13172 6554 13196 6556
rect 13034 6502 13036 6554
rect 13098 6502 13110 6554
rect 13172 6502 13174 6554
rect 13012 6500 13036 6502
rect 13092 6500 13116 6502
rect 13172 6500 13196 6502
rect 12956 6480 13252 6500
rect 12768 6344 12848 6372
rect 12716 6326 12768 6332
rect 12624 6248 12676 6254
rect 12624 6190 12676 6196
rect 12820 5846 12848 6344
rect 13280 6322 13308 6666
rect 13268 6316 13320 6322
rect 13268 6258 13320 6264
rect 13268 6180 13320 6186
rect 13268 6122 13320 6128
rect 13360 6180 13412 6186
rect 13360 6122 13412 6128
rect 12808 5840 12860 5846
rect 12808 5782 12860 5788
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 12544 5370 12572 5510
rect 12956 5468 13252 5488
rect 13012 5466 13036 5468
rect 13092 5466 13116 5468
rect 13172 5466 13196 5468
rect 13034 5414 13036 5466
rect 13098 5414 13110 5466
rect 13172 5414 13174 5466
rect 13012 5412 13036 5414
rect 13092 5412 13116 5414
rect 13172 5412 13196 5414
rect 12956 5392 13252 5412
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 12532 5364 12584 5370
rect 12532 5306 12584 5312
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11426 4312 11482 4321
rect 11426 4247 11482 4256
rect 11624 3942 11652 4966
rect 11704 4752 11756 4758
rect 11704 4694 11756 4700
rect 11716 4282 11744 4694
rect 11978 4312 12034 4321
rect 11704 4276 11756 4282
rect 11978 4247 12034 4256
rect 11704 4218 11756 4224
rect 11992 4214 12020 4247
rect 11980 4208 12032 4214
rect 11980 4150 12032 4156
rect 11704 4004 11756 4010
rect 11704 3946 11756 3952
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 11520 3664 11572 3670
rect 11520 3606 11572 3612
rect 11532 3194 11560 3606
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11060 3120 11112 3126
rect 11060 3062 11112 3068
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 9692 2514 9720 2994
rect 10600 2916 10652 2922
rect 10600 2858 10652 2864
rect 10612 2650 10640 2858
rect 10600 2644 10652 2650
rect 10600 2586 10652 2592
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 8114 2408 8170 2417
rect 7104 2372 7156 2378
rect 8114 2343 8170 2352
rect 9220 2372 9272 2378
rect 7104 2314 7156 2320
rect 9220 2314 9272 2320
rect 6918 82 6974 480
rect 6656 54 6974 82
rect 938 0 994 54
rect 2870 0 2926 54
rect 4894 0 4950 54
rect 6918 0 6974 54
rect 8942 82 8998 480
rect 9232 82 9260 2314
rect 8942 54 9260 82
rect 10874 82 10930 480
rect 11072 82 11100 3062
rect 11532 2650 11560 3130
rect 11520 2644 11572 2650
rect 11520 2586 11572 2592
rect 11624 2038 11652 3878
rect 11716 3534 11744 3946
rect 12268 3738 12296 5306
rect 12900 5160 12952 5166
rect 12900 5102 12952 5108
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12452 4486 12480 4966
rect 12912 4826 12940 5102
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 12268 3194 12296 3674
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 11612 2032 11664 2038
rect 12452 2009 12480 4422
rect 12956 4380 13252 4400
rect 13012 4378 13036 4380
rect 13092 4378 13116 4380
rect 13172 4378 13196 4380
rect 13034 4326 13036 4378
rect 13098 4326 13110 4378
rect 13172 4326 13174 4378
rect 13012 4324 13036 4326
rect 13092 4324 13116 4326
rect 13172 4324 13196 4326
rect 12956 4304 13252 4324
rect 13280 3466 13308 6122
rect 13372 5778 13400 6122
rect 13360 5772 13412 5778
rect 13360 5714 13412 5720
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 13372 5234 13400 5714
rect 13544 5636 13596 5642
rect 13544 5578 13596 5584
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13556 4690 13584 5578
rect 13648 5234 13676 5714
rect 14016 5710 14044 9454
rect 14200 7954 14228 11018
rect 14384 10810 14412 11086
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 14936 9654 14964 9862
rect 14924 9648 14976 9654
rect 14924 9590 14976 9596
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14292 9042 14320 9454
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14936 8430 14964 9590
rect 15120 9178 15148 12650
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 15212 11558 15240 12242
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 14096 7268 14148 7274
rect 14096 7210 14148 7216
rect 14108 6866 14136 7210
rect 14200 7206 14228 7890
rect 14936 7750 14964 8366
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 15212 7546 15240 11494
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15304 10266 15332 10406
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15396 9722 15424 10406
rect 15488 10198 15516 13688
rect 15580 13530 15608 13738
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 15764 12918 15792 13874
rect 15936 13728 15988 13734
rect 15936 13670 15988 13676
rect 15948 13530 15976 13670
rect 15936 13524 15988 13530
rect 15936 13466 15988 13472
rect 16132 13394 16160 14350
rect 16316 13462 16344 14758
rect 16684 14618 16712 18566
rect 16868 18086 16896 18770
rect 17052 18358 17080 18770
rect 17420 18426 17448 19178
rect 17408 18420 17460 18426
rect 17408 18362 17460 18368
rect 17040 18352 17092 18358
rect 17040 18294 17092 18300
rect 16856 18080 16908 18086
rect 16856 18022 16908 18028
rect 16868 17649 16896 18022
rect 16956 17980 17252 18000
rect 17012 17978 17036 17980
rect 17092 17978 17116 17980
rect 17172 17978 17196 17980
rect 17034 17926 17036 17978
rect 17098 17926 17110 17978
rect 17172 17926 17174 17978
rect 17012 17924 17036 17926
rect 17092 17924 17116 17926
rect 17172 17924 17196 17926
rect 16956 17904 17252 17924
rect 17132 17740 17184 17746
rect 17132 17682 17184 17688
rect 16854 17640 16910 17649
rect 16854 17575 16910 17584
rect 16672 14612 16724 14618
rect 16672 14554 16724 14560
rect 16868 14482 16896 17575
rect 17144 17270 17172 17682
rect 17132 17264 17184 17270
rect 17132 17206 17184 17212
rect 17512 17105 17540 23582
rect 19720 23582 20038 23610
rect 18420 20936 18472 20942
rect 18420 20878 18472 20884
rect 18432 19990 18460 20878
rect 19720 20602 19748 23582
rect 19982 23520 20038 23582
rect 22296 23582 22706 23610
rect 20350 22672 20406 22681
rect 20350 22607 20406 22616
rect 20364 20602 20392 22607
rect 20956 21788 21252 21808
rect 21012 21786 21036 21788
rect 21092 21786 21116 21788
rect 21172 21786 21196 21788
rect 21034 21734 21036 21786
rect 21098 21734 21110 21786
rect 21172 21734 21174 21786
rect 21012 21732 21036 21734
rect 21092 21732 21116 21734
rect 21172 21732 21196 21734
rect 20956 21712 21252 21732
rect 21362 21448 21418 21457
rect 21362 21383 21418 21392
rect 20956 20700 21252 20720
rect 21012 20698 21036 20700
rect 21092 20698 21116 20700
rect 21172 20698 21196 20700
rect 21034 20646 21036 20698
rect 21098 20646 21110 20698
rect 21172 20646 21174 20698
rect 21012 20644 21036 20646
rect 21092 20644 21116 20646
rect 21172 20644 21196 20646
rect 20956 20624 21252 20644
rect 19708 20596 19760 20602
rect 19708 20538 19760 20544
rect 20352 20596 20404 20602
rect 20352 20538 20404 20544
rect 18880 20392 18932 20398
rect 18880 20334 18932 20340
rect 19248 20392 19300 20398
rect 19248 20334 19300 20340
rect 18420 19984 18472 19990
rect 18420 19926 18472 19932
rect 18512 19984 18564 19990
rect 18512 19926 18564 19932
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 18064 19310 18092 19654
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 17776 19168 17828 19174
rect 17776 19110 17828 19116
rect 17788 18086 17816 19110
rect 18432 18970 18460 19926
rect 18524 19514 18552 19926
rect 18512 19508 18564 19514
rect 18512 19450 18564 19456
rect 18420 18964 18472 18970
rect 18420 18906 18472 18912
rect 18788 18896 18840 18902
rect 18788 18838 18840 18844
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 17776 18080 17828 18086
rect 17776 18022 17828 18028
rect 18512 18080 18564 18086
rect 18512 18022 18564 18028
rect 17788 17814 17816 18022
rect 18524 17814 18552 18022
rect 18708 17882 18736 18702
rect 18800 18426 18828 18838
rect 18788 18420 18840 18426
rect 18788 18362 18840 18368
rect 18696 17876 18748 17882
rect 18696 17818 18748 17824
rect 17776 17808 17828 17814
rect 17776 17750 17828 17756
rect 18512 17808 18564 17814
rect 18512 17750 18564 17756
rect 17788 17202 17816 17750
rect 17868 17740 17920 17746
rect 17868 17682 17920 17688
rect 17880 17338 17908 17682
rect 18052 17604 18104 17610
rect 18052 17546 18104 17552
rect 17868 17332 17920 17338
rect 17868 17274 17920 17280
rect 17776 17196 17828 17202
rect 17776 17138 17828 17144
rect 17498 17096 17554 17105
rect 17498 17031 17554 17040
rect 16956 16892 17252 16912
rect 17012 16890 17036 16892
rect 17092 16890 17116 16892
rect 17172 16890 17196 16892
rect 17034 16838 17036 16890
rect 17098 16838 17110 16890
rect 17172 16838 17174 16890
rect 17012 16836 17036 16838
rect 17092 16836 17116 16838
rect 17172 16836 17196 16838
rect 16956 16816 17252 16836
rect 16956 15804 17252 15824
rect 17012 15802 17036 15804
rect 17092 15802 17116 15804
rect 17172 15802 17196 15804
rect 17034 15750 17036 15802
rect 17098 15750 17110 15802
rect 17172 15750 17174 15802
rect 17012 15748 17036 15750
rect 17092 15748 17116 15750
rect 17172 15748 17196 15750
rect 16956 15728 17252 15748
rect 17408 15632 17460 15638
rect 17408 15574 17460 15580
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 17328 15026 17356 15438
rect 17316 15020 17368 15026
rect 17316 14962 17368 14968
rect 17420 14822 17448 15574
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 16956 14716 17252 14736
rect 17012 14714 17036 14716
rect 17092 14714 17116 14716
rect 17172 14714 17196 14716
rect 17034 14662 17036 14714
rect 17098 14662 17110 14714
rect 17172 14662 17174 14714
rect 17012 14660 17036 14662
rect 17092 14660 17116 14662
rect 17172 14660 17196 14662
rect 16956 14640 17252 14660
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 16408 13734 16436 14418
rect 16764 13864 16816 13870
rect 16764 13806 16816 13812
rect 16396 13728 16448 13734
rect 16396 13670 16448 13676
rect 16304 13456 16356 13462
rect 16304 13398 16356 13404
rect 16120 13388 16172 13394
rect 16120 13330 16172 13336
rect 16132 12986 16160 13330
rect 16316 12986 16344 13398
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 15752 12912 15804 12918
rect 15752 12854 15804 12860
rect 15936 12912 15988 12918
rect 15936 12854 15988 12860
rect 15568 10600 15620 10606
rect 15568 10542 15620 10548
rect 15476 10192 15528 10198
rect 15476 10134 15528 10140
rect 15580 9926 15608 10542
rect 15660 10056 15712 10062
rect 15660 9998 15712 10004
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15396 9586 15424 9658
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15672 9382 15700 9998
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 14648 7472 14700 7478
rect 14648 7414 14700 7420
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 14108 6458 14136 6802
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13544 4684 13596 4690
rect 13544 4626 13596 4632
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13358 3632 13414 3641
rect 13464 3602 13492 3878
rect 13556 3738 13584 4626
rect 14016 4486 14044 5646
rect 14096 5024 14148 5030
rect 14096 4966 14148 4972
rect 14108 4729 14136 4966
rect 14094 4720 14150 4729
rect 14094 4655 14150 4664
rect 14004 4480 14056 4486
rect 14004 4422 14056 4428
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13912 4072 13964 4078
rect 14016 4060 14044 4422
rect 14096 4072 14148 4078
rect 14016 4032 14096 4060
rect 13912 4014 13964 4020
rect 14096 4014 14148 4020
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13358 3567 13414 3576
rect 13452 3596 13504 3602
rect 13372 3466 13400 3567
rect 13452 3538 13504 3544
rect 13268 3460 13320 3466
rect 13268 3402 13320 3408
rect 13360 3460 13412 3466
rect 13360 3402 13412 3408
rect 12956 3292 13252 3312
rect 13012 3290 13036 3292
rect 13092 3290 13116 3292
rect 13172 3290 13196 3292
rect 13034 3238 13036 3290
rect 13098 3238 13110 3290
rect 13172 3238 13174 3290
rect 13012 3236 13036 3238
rect 13092 3236 13116 3238
rect 13172 3236 13196 3238
rect 12956 3216 13252 3236
rect 13082 3088 13138 3097
rect 13082 3023 13138 3032
rect 13096 2990 13124 3023
rect 13084 2984 13136 2990
rect 13084 2926 13136 2932
rect 13280 2514 13308 3402
rect 13464 2854 13492 3538
rect 13648 2990 13676 4014
rect 13924 3670 13952 4014
rect 13912 3664 13964 3670
rect 13912 3606 13964 3612
rect 13924 2990 13952 3606
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 13452 2848 13504 2854
rect 13452 2790 13504 2796
rect 13268 2508 13320 2514
rect 13268 2450 13320 2456
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 12956 2204 13252 2224
rect 13012 2202 13036 2204
rect 13092 2202 13116 2204
rect 13172 2202 13196 2204
rect 13034 2150 13036 2202
rect 13098 2150 13110 2202
rect 13172 2150 13174 2202
rect 13012 2148 13036 2150
rect 13092 2148 13116 2150
rect 13172 2148 13196 2150
rect 12956 2128 13252 2148
rect 11612 1974 11664 1980
rect 12438 2000 12494 2009
rect 12438 1935 12494 1944
rect 10874 54 11100 82
rect 12898 82 12954 480
rect 13280 82 13308 2314
rect 13464 1329 13492 2790
rect 13648 2650 13676 2926
rect 13636 2644 13688 2650
rect 13636 2586 13688 2592
rect 14200 2514 14228 7142
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14280 5636 14332 5642
rect 14280 5578 14332 5584
rect 14292 5302 14320 5578
rect 14384 5574 14412 6190
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 14280 5296 14332 5302
rect 14280 5238 14332 5244
rect 14384 4758 14412 5510
rect 14556 5160 14608 5166
rect 14556 5102 14608 5108
rect 14568 4826 14596 5102
rect 14556 4820 14608 4826
rect 14556 4762 14608 4768
rect 14372 4752 14424 4758
rect 14372 4694 14424 4700
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14384 2990 14412 4014
rect 14660 3505 14688 7414
rect 15396 6934 15424 8570
rect 15488 8362 15516 8910
rect 15672 8430 15700 9318
rect 15844 9036 15896 9042
rect 15844 8978 15896 8984
rect 15856 8634 15884 8978
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15476 8356 15528 8362
rect 15476 8298 15528 8304
rect 15488 8090 15516 8298
rect 15476 8084 15528 8090
rect 15476 8026 15528 8032
rect 15384 6928 15436 6934
rect 15384 6870 15436 6876
rect 15396 6458 15424 6870
rect 15476 6860 15528 6866
rect 15672 6848 15700 8366
rect 15844 8016 15896 8022
rect 15844 7958 15896 7964
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15528 6820 15700 6848
rect 15476 6802 15528 6808
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 14924 6112 14976 6118
rect 14924 6054 14976 6060
rect 14936 4729 14964 6054
rect 15396 5846 15424 6394
rect 15672 6186 15700 6820
rect 15660 6180 15712 6186
rect 15660 6122 15712 6128
rect 15672 5914 15700 6122
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15384 5840 15436 5846
rect 15384 5782 15436 5788
rect 15396 5370 15424 5782
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15660 5024 15712 5030
rect 15660 4966 15712 4972
rect 14922 4720 14978 4729
rect 14922 4655 14978 4664
rect 15384 4684 15436 4690
rect 15384 4626 15436 4632
rect 15016 4208 15068 4214
rect 15016 4150 15068 4156
rect 14646 3496 14702 3505
rect 14646 3431 14702 3440
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14384 2650 14412 2926
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 13740 2310 13768 2382
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 13450 1320 13506 1329
rect 13450 1255 13506 1264
rect 12898 54 13308 82
rect 14922 82 14978 480
rect 15028 82 15056 4150
rect 15396 3942 15424 4626
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 15396 3534 15424 3878
rect 15672 3602 15700 4966
rect 15764 4154 15792 7686
rect 15856 7274 15884 7958
rect 15844 7268 15896 7274
rect 15844 7210 15896 7216
rect 15948 6254 15976 12854
rect 16316 12782 16344 12922
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16316 11286 16344 12718
rect 16304 11280 16356 11286
rect 16304 11222 16356 11228
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 16132 10674 16160 11086
rect 16316 10810 16344 11222
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16132 9586 16160 10202
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 16212 9444 16264 9450
rect 16212 9386 16264 9392
rect 16224 9178 16252 9386
rect 16212 9172 16264 9178
rect 16212 9114 16264 9120
rect 16224 8634 16252 9114
rect 16316 9042 16344 10746
rect 16408 10606 16436 13670
rect 16580 13184 16632 13190
rect 16580 13126 16632 13132
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 16500 12442 16528 12786
rect 16592 12714 16620 13126
rect 16580 12708 16632 12714
rect 16580 12650 16632 12656
rect 16488 12436 16540 12442
rect 16488 12378 16540 12384
rect 16592 12374 16620 12650
rect 16580 12368 16632 12374
rect 16580 12310 16632 12316
rect 16776 12306 16804 13806
rect 16856 13728 16908 13734
rect 16856 13670 16908 13676
rect 16868 13530 16896 13670
rect 16956 13628 17252 13648
rect 17012 13626 17036 13628
rect 17092 13626 17116 13628
rect 17172 13626 17196 13628
rect 17034 13574 17036 13626
rect 17098 13574 17110 13626
rect 17172 13574 17174 13626
rect 17012 13572 17036 13574
rect 17092 13572 17116 13574
rect 17172 13572 17196 13574
rect 16956 13552 17252 13572
rect 17328 13530 17356 14418
rect 17604 13802 17632 14418
rect 18064 13870 18092 17546
rect 18328 16720 18380 16726
rect 18328 16662 18380 16668
rect 18236 16584 18288 16590
rect 18236 16526 18288 16532
rect 18248 16250 18276 16526
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18340 15978 18368 16662
rect 18708 16522 18736 17818
rect 18696 16516 18748 16522
rect 18696 16458 18748 16464
rect 18708 16182 18736 16458
rect 18696 16176 18748 16182
rect 18696 16118 18748 16124
rect 18328 15972 18380 15978
rect 18328 15914 18380 15920
rect 18144 15904 18196 15910
rect 18144 15846 18196 15852
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 18156 13814 18184 15846
rect 18340 15706 18368 15914
rect 18328 15700 18380 15706
rect 18328 15642 18380 15648
rect 18696 15564 18748 15570
rect 18696 15506 18748 15512
rect 18708 15162 18736 15506
rect 18696 15156 18748 15162
rect 18696 15098 18748 15104
rect 18708 15065 18736 15098
rect 18694 15056 18750 15065
rect 18694 14991 18750 15000
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 18340 14550 18368 14758
rect 18328 14544 18380 14550
rect 18328 14486 18380 14492
rect 18420 13864 18472 13870
rect 17592 13796 17644 13802
rect 18156 13786 18276 13814
rect 18472 13824 18644 13852
rect 18420 13806 18472 13812
rect 17592 13738 17644 13744
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 17684 13524 17736 13530
rect 17684 13466 17736 13472
rect 17328 12918 17356 13466
rect 17316 12912 17368 12918
rect 17316 12854 17368 12860
rect 17316 12708 17368 12714
rect 17316 12650 17368 12656
rect 16956 12540 17252 12560
rect 17012 12538 17036 12540
rect 17092 12538 17116 12540
rect 17172 12538 17196 12540
rect 17034 12486 17036 12538
rect 17098 12486 17110 12538
rect 17172 12486 17174 12538
rect 17012 12484 17036 12486
rect 17092 12484 17116 12486
rect 17172 12484 17196 12486
rect 16956 12464 17252 12484
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16764 12096 16816 12102
rect 16764 12038 16816 12044
rect 16776 11762 16804 12038
rect 17328 11830 17356 12650
rect 17408 12368 17460 12374
rect 17408 12310 17460 12316
rect 17420 11898 17448 12310
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 17316 11824 17368 11830
rect 17316 11766 17368 11772
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16580 11620 16632 11626
rect 16580 11562 16632 11568
rect 16592 11354 16620 11562
rect 16956 11452 17252 11472
rect 17012 11450 17036 11452
rect 17092 11450 17116 11452
rect 17172 11450 17196 11452
rect 17034 11398 17036 11450
rect 17098 11398 17110 11450
rect 17172 11398 17174 11450
rect 17012 11396 17036 11398
rect 17092 11396 17116 11398
rect 17172 11396 17196 11398
rect 16956 11376 17252 11396
rect 16580 11348 16632 11354
rect 16580 11290 16632 11296
rect 17316 11076 17368 11082
rect 17316 11018 17368 11024
rect 16396 10600 16448 10606
rect 16396 10542 16448 10548
rect 16956 10364 17252 10384
rect 17012 10362 17036 10364
rect 17092 10362 17116 10364
rect 17172 10362 17196 10364
rect 17034 10310 17036 10362
rect 17098 10310 17110 10362
rect 17172 10310 17174 10362
rect 17012 10308 17036 10310
rect 17092 10308 17116 10310
rect 17172 10308 17196 10310
rect 16956 10288 17252 10308
rect 16764 10192 16816 10198
rect 16764 10134 16816 10140
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16224 8294 16252 8570
rect 16684 8566 16712 9590
rect 16776 9382 16804 10134
rect 16856 10056 16908 10062
rect 16856 9998 16908 10004
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16776 8922 16804 9318
rect 16868 9042 16896 9998
rect 16956 9276 17252 9296
rect 17012 9274 17036 9276
rect 17092 9274 17116 9276
rect 17172 9274 17196 9276
rect 17034 9222 17036 9274
rect 17098 9222 17110 9274
rect 17172 9222 17174 9274
rect 17012 9220 17036 9222
rect 17092 9220 17116 9222
rect 17172 9220 17196 9222
rect 16956 9200 17252 9220
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 17328 8945 17356 11018
rect 17314 8936 17370 8945
rect 16776 8894 16896 8922
rect 16672 8560 16724 8566
rect 16672 8502 16724 8508
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 16212 8288 16264 8294
rect 16212 8230 16264 8236
rect 16592 8022 16620 8298
rect 16580 8016 16632 8022
rect 16580 7958 16632 7964
rect 16488 7880 16540 7886
rect 16488 7822 16540 7828
rect 16212 7268 16264 7274
rect 16212 7210 16264 7216
rect 16224 7002 16252 7210
rect 16500 7002 16528 7822
rect 16684 7478 16712 8502
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16776 7750 16804 8434
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 16672 7472 16724 7478
rect 16672 7414 16724 7420
rect 16776 7002 16804 7686
rect 16212 6996 16264 7002
rect 16212 6938 16264 6944
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 16764 6996 16816 7002
rect 16764 6938 16816 6944
rect 16580 6792 16632 6798
rect 16580 6734 16632 6740
rect 16592 6458 16620 6734
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16580 6452 16632 6458
rect 16580 6394 16632 6400
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 15936 6248 15988 6254
rect 15936 6190 15988 6196
rect 15948 5914 15976 6190
rect 15936 5908 15988 5914
rect 15936 5850 15988 5856
rect 16132 5778 16160 6258
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 16120 5772 16172 5778
rect 16040 5732 16120 5760
rect 16040 4826 16068 5732
rect 16120 5714 16172 5720
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 16132 4486 16160 5102
rect 16120 4480 16172 4486
rect 16120 4422 16172 4428
rect 15764 4126 16068 4154
rect 15752 3936 15804 3942
rect 15752 3878 15804 3884
rect 15764 3602 15792 3878
rect 16040 3738 16068 4126
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 15752 3596 15804 3602
rect 15752 3538 15804 3544
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15396 2990 15424 3470
rect 15476 3460 15528 3466
rect 15476 3402 15528 3408
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 15488 2922 15516 3402
rect 15476 2916 15528 2922
rect 15476 2858 15528 2864
rect 15672 2854 15700 3538
rect 16132 3466 16160 4422
rect 16316 4154 16344 5850
rect 16684 4826 16712 6598
rect 16868 5234 16896 8894
rect 17314 8871 17370 8880
rect 16956 8188 17252 8208
rect 17012 8186 17036 8188
rect 17092 8186 17116 8188
rect 17172 8186 17196 8188
rect 17034 8134 17036 8186
rect 17098 8134 17110 8186
rect 17172 8134 17174 8186
rect 17012 8132 17036 8134
rect 17092 8132 17116 8134
rect 17172 8132 17196 8134
rect 16956 8112 17252 8132
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 16960 7546 16988 7686
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 17328 7449 17356 8871
rect 17696 7954 17724 13466
rect 17868 12640 17920 12646
rect 17868 12582 17920 12588
rect 17880 12238 17908 12582
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17880 11898 17908 12174
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 18064 11354 18092 11494
rect 17776 11348 17828 11354
rect 17776 11290 17828 11296
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 17788 10810 17816 11290
rect 17776 10804 17828 10810
rect 17776 10746 17828 10752
rect 17788 10538 17816 10746
rect 18064 10742 18092 11290
rect 18248 11082 18276 13786
rect 18616 13530 18644 13824
rect 18788 13796 18840 13802
rect 18788 13738 18840 13744
rect 18604 13524 18656 13530
rect 18604 13466 18656 13472
rect 18800 12850 18828 13738
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 18800 12442 18828 12786
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18604 12368 18656 12374
rect 18604 12310 18656 12316
rect 18236 11076 18288 11082
rect 18236 11018 18288 11024
rect 18052 10736 18104 10742
rect 18052 10678 18104 10684
rect 18616 10674 18644 12310
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18604 10668 18656 10674
rect 18604 10610 18656 10616
rect 17776 10532 17828 10538
rect 17776 10474 17828 10480
rect 18708 10198 18736 11086
rect 18696 10192 18748 10198
rect 18696 10134 18748 10140
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 18156 9722 18184 10066
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 18144 9716 18196 9722
rect 18144 9658 18196 9664
rect 18248 9382 18276 9998
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 17776 9036 17828 9042
rect 17776 8978 17828 8984
rect 17788 8634 17816 8978
rect 18156 8974 18184 9114
rect 18144 8968 18196 8974
rect 18144 8910 18196 8916
rect 18156 8634 18184 8910
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17314 7440 17370 7449
rect 17314 7375 17370 7384
rect 17604 7206 17632 7822
rect 17696 7546 17724 7890
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17774 7304 17830 7313
rect 17774 7239 17830 7248
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 16956 7100 17252 7120
rect 17012 7098 17036 7100
rect 17092 7098 17116 7100
rect 17172 7098 17196 7100
rect 17034 7046 17036 7098
rect 17098 7046 17110 7098
rect 17172 7046 17174 7098
rect 17012 7044 17036 7046
rect 17092 7044 17116 7046
rect 17172 7044 17196 7046
rect 16956 7024 17252 7044
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 17144 6458 17172 6802
rect 17132 6452 17184 6458
rect 17132 6394 17184 6400
rect 17604 6254 17632 7142
rect 17592 6248 17644 6254
rect 17592 6190 17644 6196
rect 16956 6012 17252 6032
rect 17012 6010 17036 6012
rect 17092 6010 17116 6012
rect 17172 6010 17196 6012
rect 17034 5958 17036 6010
rect 17098 5958 17110 6010
rect 17172 5958 17174 6010
rect 17012 5956 17036 5958
rect 17092 5956 17116 5958
rect 17172 5956 17196 5958
rect 16956 5936 17252 5956
rect 17500 5704 17552 5710
rect 17500 5646 17552 5652
rect 17512 5370 17540 5646
rect 17500 5364 17552 5370
rect 17500 5306 17552 5312
rect 17604 5234 17632 6190
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 17592 5228 17644 5234
rect 17592 5170 17644 5176
rect 17316 5024 17368 5030
rect 17316 4966 17368 4972
rect 16956 4924 17252 4944
rect 17012 4922 17036 4924
rect 17092 4922 17116 4924
rect 17172 4922 17196 4924
rect 17034 4870 17036 4922
rect 17098 4870 17110 4922
rect 17172 4870 17174 4922
rect 17012 4868 17036 4870
rect 17092 4868 17116 4870
rect 17172 4868 17196 4870
rect 16956 4848 17252 4868
rect 16672 4820 16724 4826
rect 16672 4762 16724 4768
rect 16488 4684 16540 4690
rect 16488 4626 16540 4632
rect 16316 4126 16436 4154
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16224 3602 16252 4014
rect 16212 3596 16264 3602
rect 16212 3538 16264 3544
rect 16120 3460 16172 3466
rect 16120 3402 16172 3408
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 15948 3058 15976 3334
rect 15936 3052 15988 3058
rect 15936 2994 15988 3000
rect 15660 2848 15712 2854
rect 15660 2790 15712 2796
rect 15672 2582 15700 2790
rect 15660 2576 15712 2582
rect 15660 2518 15712 2524
rect 15948 2378 15976 2994
rect 16028 2984 16080 2990
rect 16028 2926 16080 2932
rect 16040 2854 16068 2926
rect 16028 2848 16080 2854
rect 16028 2790 16080 2796
rect 16040 2514 16068 2790
rect 16224 2514 16252 3538
rect 16408 2650 16436 4126
rect 16500 4078 16528 4626
rect 17328 4146 17356 4966
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 16488 4072 16540 4078
rect 16488 4014 16540 4020
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16672 3392 16724 3398
rect 16672 3334 16724 3340
rect 16684 2990 16712 3334
rect 16776 3126 16804 3878
rect 16956 3836 17252 3856
rect 17012 3834 17036 3836
rect 17092 3834 17116 3836
rect 17172 3834 17196 3836
rect 17034 3782 17036 3834
rect 17098 3782 17110 3834
rect 17172 3782 17174 3834
rect 17012 3780 17036 3782
rect 17092 3780 17116 3782
rect 17172 3780 17196 3782
rect 16956 3760 17252 3780
rect 16856 3596 16908 3602
rect 16856 3538 16908 3544
rect 16764 3120 16816 3126
rect 16764 3062 16816 3068
rect 16672 2984 16724 2990
rect 16672 2926 16724 2932
rect 16396 2644 16448 2650
rect 16396 2586 16448 2592
rect 16028 2508 16080 2514
rect 16028 2450 16080 2456
rect 16212 2508 16264 2514
rect 16212 2450 16264 2456
rect 15936 2372 15988 2378
rect 15936 2314 15988 2320
rect 16224 2310 16252 2450
rect 16408 2417 16436 2586
rect 16868 2514 16896 3538
rect 17328 3482 17356 4082
rect 17420 3942 17448 4558
rect 17684 4004 17736 4010
rect 17684 3946 17736 3952
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17696 3738 17724 3946
rect 17684 3732 17736 3738
rect 17684 3674 17736 3680
rect 17788 3534 17816 7239
rect 17776 3528 17828 3534
rect 17328 3454 17448 3482
rect 17776 3470 17828 3476
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 16956 2748 17252 2768
rect 17012 2746 17036 2748
rect 17092 2746 17116 2748
rect 17172 2746 17196 2748
rect 17034 2694 17036 2746
rect 17098 2694 17110 2746
rect 17172 2694 17174 2746
rect 17012 2692 17036 2694
rect 17092 2692 17116 2694
rect 17172 2692 17196 2694
rect 16956 2672 17252 2692
rect 16856 2508 16908 2514
rect 16856 2450 16908 2456
rect 17132 2508 17184 2514
rect 17132 2450 17184 2456
rect 17144 2417 17172 2450
rect 16394 2408 16450 2417
rect 16394 2343 16450 2352
rect 17130 2408 17186 2417
rect 17130 2343 17186 2352
rect 16212 2304 16264 2310
rect 16212 2246 16264 2252
rect 14922 54 15056 82
rect 16946 82 17002 480
rect 17328 82 17356 3334
rect 17420 3058 17448 3454
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17880 2446 17908 7482
rect 18156 6934 18184 8570
rect 18144 6928 18196 6934
rect 18064 6888 18144 6916
rect 18064 6458 18092 6888
rect 18144 6870 18196 6876
rect 18144 6792 18196 6798
rect 18144 6734 18196 6740
rect 18052 6452 18104 6458
rect 18052 6394 18104 6400
rect 18156 6186 18184 6734
rect 18248 6662 18276 9318
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18236 6656 18288 6662
rect 18236 6598 18288 6604
rect 18432 6322 18460 7822
rect 18512 7472 18564 7478
rect 18512 7414 18564 7420
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 18144 6180 18196 6186
rect 18144 6122 18196 6128
rect 18052 5840 18104 5846
rect 18052 5782 18104 5788
rect 18064 5370 18092 5782
rect 18052 5364 18104 5370
rect 18052 5306 18104 5312
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 18064 4826 18092 5102
rect 18156 5030 18184 6122
rect 18432 5914 18460 6258
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 18524 5642 18552 7414
rect 18604 6180 18656 6186
rect 18604 6122 18656 6128
rect 18512 5636 18564 5642
rect 18512 5578 18564 5584
rect 18524 5137 18552 5578
rect 18510 5128 18566 5137
rect 18510 5063 18566 5072
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 18616 4826 18644 6122
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 18604 4820 18656 4826
rect 18604 4762 18656 4768
rect 18064 4154 18092 4762
rect 18616 4214 18644 4762
rect 18800 4282 18828 11494
rect 18892 7993 18920 20334
rect 19260 19854 19288 20334
rect 21270 20224 21326 20233
rect 21270 20159 21326 20168
rect 19248 19848 19300 19854
rect 19248 19790 19300 19796
rect 19260 18698 19288 19790
rect 20956 19612 21252 19632
rect 21012 19610 21036 19612
rect 21092 19610 21116 19612
rect 21172 19610 21196 19612
rect 21034 19558 21036 19610
rect 21098 19558 21110 19610
rect 21172 19558 21174 19610
rect 21012 19556 21036 19558
rect 21092 19556 21116 19558
rect 21172 19556 21196 19558
rect 20956 19536 21252 19556
rect 21284 19514 21312 20159
rect 21272 19508 21324 19514
rect 21272 19450 21324 19456
rect 21270 18864 21326 18873
rect 21270 18799 21326 18808
rect 19248 18692 19300 18698
rect 19248 18634 19300 18640
rect 19064 17536 19116 17542
rect 19064 17478 19116 17484
rect 18972 17196 19024 17202
rect 18972 17138 19024 17144
rect 18984 16522 19012 17138
rect 19076 17066 19104 17478
rect 19260 17202 19288 18634
rect 20956 18524 21252 18544
rect 21012 18522 21036 18524
rect 21092 18522 21116 18524
rect 21172 18522 21196 18524
rect 21034 18470 21036 18522
rect 21098 18470 21110 18522
rect 21172 18470 21174 18522
rect 21012 18468 21036 18470
rect 21092 18468 21116 18470
rect 21172 18468 21196 18470
rect 20956 18448 21252 18468
rect 19800 18216 19852 18222
rect 19800 18158 19852 18164
rect 19812 17610 19840 18158
rect 19892 18080 19944 18086
rect 19892 18022 19944 18028
rect 19904 17746 19932 18022
rect 21284 17882 21312 18799
rect 21272 17876 21324 17882
rect 21272 17818 21324 17824
rect 19892 17740 19944 17746
rect 19892 17682 19944 17688
rect 20720 17740 20772 17746
rect 20720 17682 20772 17688
rect 19800 17604 19852 17610
rect 19800 17546 19852 17552
rect 20536 17264 20588 17270
rect 20536 17206 20588 17212
rect 19248 17196 19300 17202
rect 19248 17138 19300 17144
rect 19524 17128 19576 17134
rect 19524 17070 19576 17076
rect 19064 17060 19116 17066
rect 19064 17002 19116 17008
rect 18972 16516 19024 16522
rect 18972 16458 19024 16464
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19260 15638 19288 16186
rect 19536 15910 19564 17070
rect 19524 15904 19576 15910
rect 19524 15846 19576 15852
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 18972 15632 19024 15638
rect 18972 15574 19024 15580
rect 19248 15632 19300 15638
rect 19248 15574 19300 15580
rect 18984 14890 19012 15574
rect 19996 15162 20024 15846
rect 19984 15156 20036 15162
rect 19984 15098 20036 15104
rect 18972 14884 19024 14890
rect 18972 14826 19024 14832
rect 18972 14476 19024 14482
rect 18972 14418 19024 14424
rect 19064 14476 19116 14482
rect 19064 14418 19116 14424
rect 18984 14006 19012 14418
rect 19076 14074 19104 14418
rect 19248 14408 19300 14414
rect 19248 14350 19300 14356
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 18972 14000 19024 14006
rect 18972 13942 19024 13948
rect 19076 13870 19104 14010
rect 19064 13864 19116 13870
rect 19064 13806 19116 13812
rect 19064 13456 19116 13462
rect 19064 13398 19116 13404
rect 19076 12986 19104 13398
rect 19260 13326 19288 14350
rect 20168 14272 20220 14278
rect 20168 14214 20220 14220
rect 19800 13932 19852 13938
rect 19800 13874 19852 13880
rect 19248 13320 19300 13326
rect 19248 13262 19300 13268
rect 19064 12980 19116 12986
rect 19064 12922 19116 12928
rect 19076 12714 19104 12922
rect 19064 12708 19116 12714
rect 19064 12650 19116 12656
rect 19076 12306 19104 12650
rect 19064 12300 19116 12306
rect 19064 12242 19116 12248
rect 19340 12300 19392 12306
rect 19340 12242 19392 12248
rect 19076 11354 19104 12242
rect 19352 11558 19380 12242
rect 19708 12096 19760 12102
rect 19708 12038 19760 12044
rect 19616 11620 19668 11626
rect 19616 11562 19668 11568
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 19524 11552 19576 11558
rect 19524 11494 19576 11500
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 19076 10810 19104 11290
rect 19064 10804 19116 10810
rect 19064 10746 19116 10752
rect 19064 9920 19116 9926
rect 19064 9862 19116 9868
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19076 9450 19104 9862
rect 19260 9586 19288 9862
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 19064 9444 19116 9450
rect 19064 9386 19116 9392
rect 19076 9178 19104 9386
rect 19260 9178 19288 9522
rect 19064 9172 19116 9178
rect 19064 9114 19116 9120
rect 19248 9172 19300 9178
rect 19248 9114 19300 9120
rect 18972 8832 19024 8838
rect 18972 8774 19024 8780
rect 18984 8498 19012 8774
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 19076 8362 19104 9114
rect 19352 9081 19380 11494
rect 19536 11218 19564 11494
rect 19628 11354 19656 11562
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19524 11212 19576 11218
rect 19524 11154 19576 11160
rect 19536 10810 19564 11154
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 19536 10538 19564 10746
rect 19720 10674 19748 12038
rect 19812 10713 19840 13874
rect 20180 13802 20208 14214
rect 20548 13954 20576 17206
rect 20732 16998 20760 17682
rect 21270 17640 21326 17649
rect 21270 17575 21326 17584
rect 20956 17436 21252 17456
rect 21012 17434 21036 17436
rect 21092 17434 21116 17436
rect 21172 17434 21196 17436
rect 21034 17382 21036 17434
rect 21098 17382 21110 17434
rect 21172 17382 21174 17434
rect 21012 17380 21036 17382
rect 21092 17380 21116 17382
rect 21172 17380 21196 17382
rect 20956 17360 21252 17380
rect 21284 17338 21312 17575
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 20732 16017 20760 16934
rect 20956 16348 21252 16368
rect 21012 16346 21036 16348
rect 21092 16346 21116 16348
rect 21172 16346 21196 16348
rect 21034 16294 21036 16346
rect 21098 16294 21110 16346
rect 21172 16294 21174 16346
rect 21012 16292 21036 16294
rect 21092 16292 21116 16294
rect 21172 16292 21196 16294
rect 20956 16272 21252 16292
rect 20718 16008 20774 16017
rect 20718 15943 20774 15952
rect 20956 15260 21252 15280
rect 21012 15258 21036 15260
rect 21092 15258 21116 15260
rect 21172 15258 21196 15260
rect 21034 15206 21036 15258
rect 21098 15206 21110 15258
rect 21172 15206 21174 15258
rect 21012 15204 21036 15206
rect 21092 15204 21116 15206
rect 21172 15204 21196 15206
rect 20956 15184 21252 15204
rect 21272 15088 21324 15094
rect 21272 15030 21324 15036
rect 20628 14816 20680 14822
rect 20628 14758 20680 14764
rect 20640 14618 20668 14758
rect 20628 14612 20680 14618
rect 20628 14554 20680 14560
rect 20812 14476 20864 14482
rect 20812 14418 20864 14424
rect 20824 14006 20852 14418
rect 20956 14172 21252 14192
rect 21012 14170 21036 14172
rect 21092 14170 21116 14172
rect 21172 14170 21196 14172
rect 21034 14118 21036 14170
rect 21098 14118 21110 14170
rect 21172 14118 21174 14170
rect 21012 14116 21036 14118
rect 21092 14116 21116 14118
rect 21172 14116 21196 14118
rect 20956 14096 21252 14116
rect 21284 14056 21312 15030
rect 21192 14028 21312 14056
rect 20812 14000 20864 14006
rect 20626 13968 20682 13977
rect 20548 13926 20626 13954
rect 20812 13942 20864 13948
rect 20626 13903 20682 13912
rect 20168 13796 20220 13802
rect 20168 13738 20220 13744
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19996 13530 20024 13670
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 20180 11830 20208 13738
rect 20260 13320 20312 13326
rect 20260 13262 20312 13268
rect 20272 12918 20300 13262
rect 20260 12912 20312 12918
rect 20260 12854 20312 12860
rect 20168 11824 20220 11830
rect 20168 11766 20220 11772
rect 19798 10704 19854 10713
rect 19708 10668 19760 10674
rect 20180 10674 20208 11766
rect 19798 10639 19854 10648
rect 20168 10668 20220 10674
rect 19708 10610 19760 10616
rect 19524 10532 19576 10538
rect 19524 10474 19576 10480
rect 19720 10266 19748 10610
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 19812 10130 19840 10639
rect 20168 10610 20220 10616
rect 20444 10464 20496 10470
rect 20444 10406 20496 10412
rect 19800 10124 19852 10130
rect 19800 10066 19852 10072
rect 19812 9450 19840 10066
rect 19524 9444 19576 9450
rect 19524 9386 19576 9392
rect 19800 9444 19852 9450
rect 19800 9386 19852 9392
rect 19338 9072 19394 9081
rect 19338 9007 19394 9016
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19064 8356 19116 8362
rect 19064 8298 19116 8304
rect 19076 8090 19104 8298
rect 19064 8084 19116 8090
rect 19064 8026 19116 8032
rect 19156 8016 19208 8022
rect 18878 7984 18934 7993
rect 19156 7958 19208 7964
rect 18878 7919 18934 7928
rect 18892 6866 18920 7919
rect 19168 7546 19196 7958
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 19168 7002 19196 7482
rect 19260 7410 19288 8434
rect 19536 8294 19564 9386
rect 19812 9353 19840 9386
rect 19798 9344 19854 9353
rect 19798 9279 19854 9288
rect 19708 9036 19760 9042
rect 19708 8978 19760 8984
rect 19720 8634 19748 8978
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19524 8288 19576 8294
rect 19524 8230 19576 8236
rect 19536 7886 19564 8230
rect 19524 7880 19576 7886
rect 19524 7822 19576 7828
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 19156 6996 19208 7002
rect 19156 6938 19208 6944
rect 18880 6860 18932 6866
rect 18880 6802 18932 6808
rect 19352 6458 19380 7142
rect 19536 7002 19564 7822
rect 19616 7812 19668 7818
rect 19616 7754 19668 7760
rect 19628 7478 19656 7754
rect 20456 7750 20484 10406
rect 20444 7744 20496 7750
rect 20444 7686 20496 7692
rect 19616 7472 19668 7478
rect 19616 7414 19668 7420
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 20352 5568 20404 5574
rect 20352 5510 20404 5516
rect 20364 5098 20392 5510
rect 20352 5092 20404 5098
rect 20352 5034 20404 5040
rect 20168 4548 20220 4554
rect 20168 4490 20220 4496
rect 18788 4276 18840 4282
rect 18788 4218 18840 4224
rect 18236 4208 18288 4214
rect 18064 4126 18184 4154
rect 18236 4150 18288 4156
rect 18604 4208 18656 4214
rect 18604 4150 18656 4156
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 18064 2990 18092 3334
rect 18052 2984 18104 2990
rect 18052 2926 18104 2932
rect 18064 2854 18092 2926
rect 18156 2854 18184 4126
rect 18248 3670 18276 4150
rect 18236 3664 18288 3670
rect 18236 3606 18288 3612
rect 18236 3120 18288 3126
rect 18236 3062 18288 3068
rect 18248 2990 18276 3062
rect 18236 2984 18288 2990
rect 18236 2926 18288 2932
rect 18052 2848 18104 2854
rect 18052 2790 18104 2796
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 18064 2650 18092 2790
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 17868 2440 17920 2446
rect 18248 2417 18276 2926
rect 18604 2508 18656 2514
rect 18604 2450 18656 2456
rect 17868 2382 17920 2388
rect 18234 2408 18290 2417
rect 18234 2343 18290 2352
rect 18616 2310 18644 2450
rect 18604 2304 18656 2310
rect 18604 2246 18656 2252
rect 18616 1193 18644 2246
rect 18602 1184 18658 1193
rect 18602 1119 18658 1128
rect 16946 54 17356 82
rect 18800 82 18828 4218
rect 20180 4146 20208 4490
rect 20364 4146 20392 5034
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 19352 3738 19380 4014
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 19984 3732 20036 3738
rect 19984 3674 20036 3680
rect 19064 3664 19116 3670
rect 19064 3606 19116 3612
rect 19076 3194 19104 3606
rect 19892 3392 19944 3398
rect 19892 3334 19944 3340
rect 19064 3188 19116 3194
rect 19064 3130 19116 3136
rect 19904 3058 19932 3334
rect 19892 3052 19944 3058
rect 19892 2994 19944 3000
rect 19996 2922 20024 3674
rect 20364 3058 20392 4082
rect 20352 3052 20404 3058
rect 20352 2994 20404 3000
rect 19984 2916 20036 2922
rect 19984 2858 20036 2864
rect 20456 2514 20484 7686
rect 20640 4690 20668 13903
rect 21192 13870 21220 14028
rect 21180 13864 21232 13870
rect 21376 13814 21404 21383
rect 21456 19304 21508 19310
rect 21456 19246 21508 19252
rect 21468 15026 21496 19246
rect 21546 16416 21602 16425
rect 21546 16351 21602 16360
rect 21456 15020 21508 15026
rect 21456 14962 21508 14968
rect 21180 13806 21232 13812
rect 20812 13456 20864 13462
rect 20812 13398 20864 13404
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20732 12442 20760 13262
rect 20824 12986 20852 13398
rect 21192 13326 21220 13806
rect 21284 13786 21404 13814
rect 21180 13320 21232 13326
rect 21180 13262 21232 13268
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 20812 12980 20864 12986
rect 20812 12922 20864 12928
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20732 11762 20760 12378
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20812 11212 20864 11218
rect 20812 11154 20864 11160
rect 20824 10470 20852 11154
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 21086 10160 21142 10169
rect 20812 10124 20864 10130
rect 21086 10095 21142 10104
rect 20812 10066 20864 10072
rect 20824 9364 20852 10066
rect 21100 9994 21128 10095
rect 21088 9988 21140 9994
rect 21088 9930 21140 9936
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 20904 9376 20956 9382
rect 20824 9336 20904 9364
rect 20904 9318 20956 9324
rect 20916 9081 20944 9318
rect 20902 9072 20958 9081
rect 20902 9007 20958 9016
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20732 5098 20760 6054
rect 20824 5846 20852 7142
rect 21284 7002 21312 13786
rect 21362 13152 21418 13161
rect 21362 13087 21418 13096
rect 21376 12986 21404 13087
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 21560 12782 21588 16351
rect 21640 15564 21692 15570
rect 21640 15506 21692 15512
rect 21548 12776 21600 12782
rect 21548 12718 21600 12724
rect 21362 11928 21418 11937
rect 21652 11898 21680 15506
rect 22296 14618 22324 23582
rect 22650 23520 22706 23582
rect 23570 15736 23626 15745
rect 23570 15671 23626 15680
rect 23584 15570 23612 15671
rect 23572 15564 23624 15570
rect 23572 15506 23624 15512
rect 22284 14612 22336 14618
rect 22284 14554 22336 14560
rect 21362 11863 21418 11872
rect 21640 11892 21692 11898
rect 21376 11830 21404 11863
rect 21640 11834 21692 11840
rect 21364 11824 21416 11830
rect 21364 11766 21416 11772
rect 21652 11694 21680 11834
rect 21640 11688 21692 11694
rect 21640 11630 21692 11636
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 21456 6860 21508 6866
rect 21456 6802 21508 6808
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 21468 6458 21496 6802
rect 21456 6452 21508 6458
rect 21456 6394 21508 6400
rect 21180 6180 21232 6186
rect 21180 6122 21232 6128
rect 21192 5846 21220 6122
rect 20812 5840 20864 5846
rect 20812 5782 20864 5788
rect 21180 5840 21232 5846
rect 21232 5800 21312 5828
rect 21180 5782 21232 5788
rect 20824 5370 20852 5782
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 21284 5370 21312 5800
rect 21468 5710 21496 6394
rect 21456 5704 21508 5710
rect 21456 5646 21508 5652
rect 21362 5400 21418 5409
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 21272 5364 21324 5370
rect 21362 5335 21418 5344
rect 21272 5306 21324 5312
rect 21376 5302 21404 5335
rect 21364 5296 21416 5302
rect 21364 5238 21416 5244
rect 21468 5234 21496 5646
rect 21456 5228 21508 5234
rect 21456 5170 21508 5176
rect 20720 5092 20772 5098
rect 20720 5034 20772 5040
rect 20732 4826 20760 5034
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 20628 4684 20680 4690
rect 20628 4626 20680 4632
rect 20640 4282 20668 4626
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 20628 4276 20680 4282
rect 20628 4218 20680 4224
rect 20640 3097 20668 4218
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 20824 3194 20852 3470
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 20626 3088 20682 3097
rect 20626 3023 20682 3032
rect 20824 2650 20852 3130
rect 20812 2644 20864 2650
rect 20812 2586 20864 2592
rect 20444 2508 20496 2514
rect 20444 2450 20496 2456
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 22652 2372 22704 2378
rect 22652 2314 22704 2320
rect 18878 82 18934 480
rect 18800 54 18934 82
rect 20640 82 20668 2314
rect 20956 2204 21252 2224
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 20902 82 20958 480
rect 20640 54 20958 82
rect 22664 82 22692 2314
rect 22926 82 22982 480
rect 22664 54 22982 82
rect 8942 0 8998 54
rect 10874 0 10930 54
rect 12898 0 12954 54
rect 14922 0 14978 54
rect 16946 0 17002 54
rect 18878 0 18934 54
rect 20902 0 20958 54
rect 22926 0 22982 54
<< via2 >>
rect 1122 21120 1178 21176
rect 1582 22616 1638 22672
rect 4956 21786 5012 21788
rect 5036 21786 5092 21788
rect 5116 21786 5172 21788
rect 5196 21786 5252 21788
rect 4956 21734 4982 21786
rect 4982 21734 5012 21786
rect 5036 21734 5046 21786
rect 5046 21734 5092 21786
rect 5116 21734 5162 21786
rect 5162 21734 5172 21786
rect 5196 21734 5226 21786
rect 5226 21734 5252 21786
rect 4956 21732 5012 21734
rect 5036 21732 5092 21734
rect 5116 21732 5172 21734
rect 5196 21732 5252 21734
rect 4956 20698 5012 20700
rect 5036 20698 5092 20700
rect 5116 20698 5172 20700
rect 5196 20698 5252 20700
rect 4956 20646 4982 20698
rect 4982 20646 5012 20698
rect 5036 20646 5046 20698
rect 5046 20646 5092 20698
rect 5116 20646 5162 20698
rect 5162 20646 5172 20698
rect 5196 20646 5226 20698
rect 5226 20646 5252 20698
rect 4956 20644 5012 20646
rect 5036 20644 5092 20646
rect 5116 20644 5172 20646
rect 5196 20644 5252 20646
rect 8956 21242 9012 21244
rect 9036 21242 9092 21244
rect 9116 21242 9172 21244
rect 9196 21242 9252 21244
rect 8956 21190 8982 21242
rect 8982 21190 9012 21242
rect 9036 21190 9046 21242
rect 9046 21190 9092 21242
rect 9116 21190 9162 21242
rect 9162 21190 9172 21242
rect 9196 21190 9226 21242
rect 9226 21190 9252 21242
rect 8956 21188 9012 21190
rect 9036 21188 9092 21190
rect 9116 21188 9172 21190
rect 9196 21188 9252 21190
rect 12956 21786 13012 21788
rect 13036 21786 13092 21788
rect 13116 21786 13172 21788
rect 13196 21786 13252 21788
rect 12956 21734 12982 21786
rect 12982 21734 13012 21786
rect 13036 21734 13046 21786
rect 13046 21734 13092 21786
rect 13116 21734 13162 21786
rect 13162 21734 13172 21786
rect 13196 21734 13226 21786
rect 13226 21734 13252 21786
rect 12956 21732 13012 21734
rect 13036 21732 13092 21734
rect 13116 21732 13172 21734
rect 13196 21732 13252 21734
rect 12956 20698 13012 20700
rect 13036 20698 13092 20700
rect 13116 20698 13172 20700
rect 13196 20698 13252 20700
rect 12956 20646 12982 20698
rect 12982 20646 13012 20698
rect 13036 20646 13046 20698
rect 13046 20646 13092 20698
rect 13116 20646 13162 20698
rect 13162 20646 13172 20698
rect 13196 20646 13226 20698
rect 13226 20646 13252 20698
rect 12956 20644 13012 20646
rect 13036 20644 13092 20646
rect 13116 20644 13172 20646
rect 13196 20644 13252 20646
rect 1490 19760 1546 19816
rect 1582 19624 1638 19680
rect 4956 19610 5012 19612
rect 5036 19610 5092 19612
rect 5116 19610 5172 19612
rect 5196 19610 5252 19612
rect 4956 19558 4982 19610
rect 4982 19558 5012 19610
rect 5036 19558 5046 19610
rect 5046 19558 5092 19610
rect 5116 19558 5162 19610
rect 5162 19558 5172 19610
rect 5196 19558 5226 19610
rect 5226 19558 5252 19610
rect 4956 19556 5012 19558
rect 5036 19556 5092 19558
rect 5116 19556 5172 19558
rect 5196 19556 5252 19558
rect 8956 20154 9012 20156
rect 9036 20154 9092 20156
rect 9116 20154 9172 20156
rect 9196 20154 9252 20156
rect 8956 20102 8982 20154
rect 8982 20102 9012 20154
rect 9036 20102 9046 20154
rect 9046 20102 9092 20154
rect 9116 20102 9162 20154
rect 9162 20102 9172 20154
rect 9196 20102 9226 20154
rect 9226 20102 9252 20154
rect 8956 20100 9012 20102
rect 9036 20100 9092 20102
rect 9116 20100 9172 20102
rect 9196 20100 9252 20102
rect 1398 18128 1454 18184
rect 110 14184 166 14240
rect 4956 18522 5012 18524
rect 5036 18522 5092 18524
rect 5116 18522 5172 18524
rect 5196 18522 5252 18524
rect 4956 18470 4982 18522
rect 4982 18470 5012 18522
rect 5036 18470 5046 18522
rect 5046 18470 5092 18522
rect 5116 18470 5162 18522
rect 5162 18470 5172 18522
rect 5196 18470 5226 18522
rect 5226 18470 5252 18522
rect 4956 18468 5012 18470
rect 5036 18468 5092 18470
rect 5116 18468 5172 18470
rect 5196 18468 5252 18470
rect 110 11192 166 11248
rect 110 8200 166 8256
rect 110 7248 166 7304
rect 18 5208 74 5264
rect 110 2216 166 2272
rect 3054 15136 3110 15192
rect 4956 17434 5012 17436
rect 5036 17434 5092 17436
rect 5116 17434 5172 17436
rect 5196 17434 5252 17436
rect 4956 17382 4982 17434
rect 4982 17382 5012 17434
rect 5036 17382 5046 17434
rect 5046 17382 5092 17434
rect 5116 17382 5162 17434
rect 5162 17382 5172 17434
rect 5196 17382 5226 17434
rect 5226 17382 5252 17434
rect 4956 17380 5012 17382
rect 5036 17380 5092 17382
rect 5116 17380 5172 17382
rect 5196 17380 5252 17382
rect 4956 16346 5012 16348
rect 5036 16346 5092 16348
rect 5116 16346 5172 16348
rect 5196 16346 5252 16348
rect 4956 16294 4982 16346
rect 4982 16294 5012 16346
rect 5036 16294 5046 16346
rect 5046 16294 5092 16346
rect 5116 16294 5162 16346
rect 5162 16294 5172 16346
rect 5196 16294 5226 16346
rect 5226 16294 5252 16346
rect 4956 16292 5012 16294
rect 5036 16292 5092 16294
rect 5116 16292 5172 16294
rect 5196 16292 5252 16294
rect 3790 15000 3846 15056
rect 2042 9968 2098 10024
rect 754 4120 810 4176
rect 3514 9016 3570 9072
rect 2870 6160 2926 6216
rect 1950 5108 1952 5128
rect 1952 5108 2004 5128
rect 2004 5108 2006 5128
rect 1950 5072 2006 5108
rect 4956 15258 5012 15260
rect 5036 15258 5092 15260
rect 5116 15258 5172 15260
rect 5196 15258 5252 15260
rect 4956 15206 4982 15258
rect 4982 15206 5012 15258
rect 5036 15206 5046 15258
rect 5046 15206 5092 15258
rect 5116 15206 5162 15258
rect 5162 15206 5172 15258
rect 5196 15206 5226 15258
rect 5226 15206 5252 15258
rect 4956 15204 5012 15206
rect 5036 15204 5092 15206
rect 5116 15204 5172 15206
rect 5196 15204 5252 15206
rect 7194 17584 7250 17640
rect 4250 13912 4306 13968
rect 4956 14170 5012 14172
rect 5036 14170 5092 14172
rect 5116 14170 5172 14172
rect 5196 14170 5252 14172
rect 4956 14118 4982 14170
rect 4982 14118 5012 14170
rect 5036 14118 5046 14170
rect 5046 14118 5092 14170
rect 5116 14118 5162 14170
rect 5162 14118 5172 14170
rect 5196 14118 5226 14170
rect 5226 14118 5252 14170
rect 4956 14116 5012 14118
rect 5036 14116 5092 14118
rect 5116 14116 5172 14118
rect 5196 14116 5252 14118
rect 4956 13082 5012 13084
rect 5036 13082 5092 13084
rect 5116 13082 5172 13084
rect 5196 13082 5252 13084
rect 4956 13030 4982 13082
rect 4982 13030 5012 13082
rect 5036 13030 5046 13082
rect 5046 13030 5092 13082
rect 5116 13030 5162 13082
rect 5162 13030 5172 13082
rect 5196 13030 5226 13082
rect 5226 13030 5252 13082
rect 4956 13028 5012 13030
rect 5036 13028 5092 13030
rect 5116 13028 5172 13030
rect 5196 13028 5252 13030
rect 6550 13812 6552 13832
rect 6552 13812 6604 13832
rect 6604 13812 6606 13832
rect 8956 19066 9012 19068
rect 9036 19066 9092 19068
rect 9116 19066 9172 19068
rect 9196 19066 9252 19068
rect 8956 19014 8982 19066
rect 8982 19014 9012 19066
rect 9036 19014 9046 19066
rect 9046 19014 9092 19066
rect 9116 19014 9162 19066
rect 9162 19014 9172 19066
rect 9196 19014 9226 19066
rect 9226 19014 9252 19066
rect 8956 19012 9012 19014
rect 9036 19012 9092 19014
rect 9116 19012 9172 19014
rect 9196 19012 9252 19014
rect 8956 17978 9012 17980
rect 9036 17978 9092 17980
rect 9116 17978 9172 17980
rect 9196 17978 9252 17980
rect 8956 17926 8982 17978
rect 8982 17926 9012 17978
rect 9036 17926 9046 17978
rect 9046 17926 9092 17978
rect 9116 17926 9162 17978
rect 9162 17926 9172 17978
rect 9196 17926 9226 17978
rect 9226 17926 9252 17978
rect 8956 17924 9012 17926
rect 9036 17924 9092 17926
rect 9116 17924 9172 17926
rect 9196 17924 9252 17926
rect 8390 17720 8446 17776
rect 8298 16496 8354 16552
rect 6550 13776 6606 13812
rect 4956 11994 5012 11996
rect 5036 11994 5092 11996
rect 5116 11994 5172 11996
rect 5196 11994 5252 11996
rect 4956 11942 4982 11994
rect 4982 11942 5012 11994
rect 5036 11942 5046 11994
rect 5046 11942 5092 11994
rect 5116 11942 5162 11994
rect 5162 11942 5172 11994
rect 5196 11942 5226 11994
rect 5226 11942 5252 11994
rect 4956 11940 5012 11942
rect 5036 11940 5092 11942
rect 5116 11940 5172 11942
rect 5196 11940 5252 11942
rect 4956 10906 5012 10908
rect 5036 10906 5092 10908
rect 5116 10906 5172 10908
rect 5196 10906 5252 10908
rect 4956 10854 4982 10906
rect 4982 10854 5012 10906
rect 5036 10854 5046 10906
rect 5046 10854 5092 10906
rect 5116 10854 5162 10906
rect 5162 10854 5172 10906
rect 5196 10854 5226 10906
rect 5226 10854 5252 10906
rect 4956 10852 5012 10854
rect 5036 10852 5092 10854
rect 5116 10852 5172 10854
rect 5196 10852 5252 10854
rect 4710 9968 4766 10024
rect 3698 3576 3754 3632
rect 4956 9818 5012 9820
rect 5036 9818 5092 9820
rect 5116 9818 5172 9820
rect 5196 9818 5252 9820
rect 4956 9766 4982 9818
rect 4982 9766 5012 9818
rect 5036 9766 5046 9818
rect 5046 9766 5092 9818
rect 5116 9766 5162 9818
rect 5162 9766 5172 9818
rect 5196 9766 5226 9818
rect 5226 9766 5252 9818
rect 4956 9764 5012 9766
rect 5036 9764 5092 9766
rect 5116 9764 5172 9766
rect 5196 9764 5252 9766
rect 4956 8730 5012 8732
rect 5036 8730 5092 8732
rect 5116 8730 5172 8732
rect 5196 8730 5252 8732
rect 4956 8678 4982 8730
rect 4982 8678 5012 8730
rect 5036 8678 5046 8730
rect 5046 8678 5092 8730
rect 5116 8678 5162 8730
rect 5162 8678 5172 8730
rect 5196 8678 5226 8730
rect 5226 8678 5252 8730
rect 4956 8676 5012 8678
rect 5036 8676 5092 8678
rect 5116 8676 5172 8678
rect 5196 8676 5252 8678
rect 4956 7642 5012 7644
rect 5036 7642 5092 7644
rect 5116 7642 5172 7644
rect 5196 7642 5252 7644
rect 4956 7590 4982 7642
rect 4982 7590 5012 7642
rect 5036 7590 5046 7642
rect 5046 7590 5092 7642
rect 5116 7590 5162 7642
rect 5162 7590 5172 7642
rect 5196 7590 5226 7642
rect 5226 7590 5252 7642
rect 4956 7588 5012 7590
rect 5036 7588 5092 7590
rect 5116 7588 5172 7590
rect 5196 7588 5252 7590
rect 4956 6554 5012 6556
rect 5036 6554 5092 6556
rect 5116 6554 5172 6556
rect 5196 6554 5252 6556
rect 4956 6502 4982 6554
rect 4982 6502 5012 6554
rect 5036 6502 5046 6554
rect 5046 6502 5092 6554
rect 5116 6502 5162 6554
rect 5162 6502 5172 6554
rect 5196 6502 5226 6554
rect 5226 6502 5252 6554
rect 4956 6500 5012 6502
rect 5036 6500 5092 6502
rect 5116 6500 5172 6502
rect 5196 6500 5252 6502
rect 4956 5466 5012 5468
rect 5036 5466 5092 5468
rect 5116 5466 5172 5468
rect 5196 5466 5252 5468
rect 4956 5414 4982 5466
rect 4982 5414 5012 5466
rect 5036 5414 5046 5466
rect 5046 5414 5092 5466
rect 5116 5414 5162 5466
rect 5162 5414 5172 5466
rect 5196 5414 5226 5466
rect 5226 5414 5252 5466
rect 4956 5412 5012 5414
rect 5036 5412 5092 5414
rect 5116 5412 5172 5414
rect 5196 5412 5252 5414
rect 4956 4378 5012 4380
rect 5036 4378 5092 4380
rect 5116 4378 5172 4380
rect 5196 4378 5252 4380
rect 4956 4326 4982 4378
rect 4982 4326 5012 4378
rect 5036 4326 5046 4378
rect 5046 4326 5092 4378
rect 5116 4326 5162 4378
rect 5162 4326 5172 4378
rect 5196 4326 5226 4378
rect 5226 4326 5252 4378
rect 4956 4324 5012 4326
rect 5036 4324 5092 4326
rect 5116 4324 5172 4326
rect 5196 4324 5252 4326
rect 8298 13232 8354 13288
rect 9402 17720 9458 17776
rect 9310 17076 9312 17096
rect 9312 17076 9364 17096
rect 9364 17076 9366 17096
rect 9310 17040 9366 17076
rect 8956 16890 9012 16892
rect 9036 16890 9092 16892
rect 9116 16890 9172 16892
rect 9196 16890 9252 16892
rect 8956 16838 8982 16890
rect 8982 16838 9012 16890
rect 9036 16838 9046 16890
rect 9046 16838 9092 16890
rect 9116 16838 9162 16890
rect 9162 16838 9172 16890
rect 9196 16838 9226 16890
rect 9226 16838 9252 16890
rect 8956 16836 9012 16838
rect 9036 16836 9092 16838
rect 9116 16836 9172 16838
rect 9196 16836 9252 16838
rect 9310 15952 9366 16008
rect 8956 15802 9012 15804
rect 9036 15802 9092 15804
rect 9116 15802 9172 15804
rect 9196 15802 9252 15804
rect 8956 15750 8982 15802
rect 8982 15750 9012 15802
rect 9036 15750 9046 15802
rect 9046 15750 9092 15802
rect 9116 15750 9162 15802
rect 9162 15750 9172 15802
rect 9196 15750 9226 15802
rect 9226 15750 9252 15802
rect 8956 15748 9012 15750
rect 9036 15748 9092 15750
rect 9116 15748 9172 15750
rect 9196 15748 9252 15750
rect 8758 15000 8814 15056
rect 8956 14714 9012 14716
rect 9036 14714 9092 14716
rect 9116 14714 9172 14716
rect 9196 14714 9252 14716
rect 8956 14662 8982 14714
rect 8982 14662 9012 14714
rect 9036 14662 9046 14714
rect 9046 14662 9092 14714
rect 9116 14662 9162 14714
rect 9162 14662 9172 14714
rect 9196 14662 9226 14714
rect 9226 14662 9252 14714
rect 8956 14660 9012 14662
rect 9036 14660 9092 14662
rect 9116 14660 9172 14662
rect 9196 14660 9252 14662
rect 9310 13812 9312 13832
rect 9312 13812 9364 13832
rect 9364 13812 9366 13832
rect 9310 13776 9366 13812
rect 8956 13626 9012 13628
rect 9036 13626 9092 13628
rect 9116 13626 9172 13628
rect 9196 13626 9252 13628
rect 8956 13574 8982 13626
rect 8982 13574 9012 13626
rect 9036 13574 9046 13626
rect 9046 13574 9092 13626
rect 9116 13574 9162 13626
rect 9162 13574 9172 13626
rect 9196 13574 9226 13626
rect 9226 13574 9252 13626
rect 8956 13572 9012 13574
rect 9036 13572 9092 13574
rect 9116 13572 9172 13574
rect 9196 13572 9252 13574
rect 11610 19760 11666 19816
rect 12956 19610 13012 19612
rect 13036 19610 13092 19612
rect 13116 19610 13172 19612
rect 13196 19610 13252 19612
rect 12956 19558 12982 19610
rect 12982 19558 13012 19610
rect 13036 19558 13046 19610
rect 13046 19558 13092 19610
rect 13116 19558 13162 19610
rect 13162 19558 13172 19610
rect 13196 19558 13226 19610
rect 13226 19558 13252 19610
rect 12956 19556 13012 19558
rect 13036 19556 13092 19558
rect 13116 19556 13172 19558
rect 13196 19556 13252 19558
rect 10966 17584 11022 17640
rect 10414 15000 10470 15056
rect 7378 8200 7434 8256
rect 8956 12538 9012 12540
rect 9036 12538 9092 12540
rect 9116 12538 9172 12540
rect 9196 12538 9252 12540
rect 8956 12486 8982 12538
rect 8982 12486 9012 12538
rect 9036 12486 9046 12538
rect 9046 12486 9092 12538
rect 9116 12486 9162 12538
rect 9162 12486 9172 12538
rect 9196 12486 9226 12538
rect 9226 12486 9252 12538
rect 8956 12484 9012 12486
rect 9036 12484 9092 12486
rect 9116 12484 9172 12486
rect 9196 12484 9252 12486
rect 8022 9016 8078 9072
rect 7010 7248 7066 7304
rect 8956 11450 9012 11452
rect 9036 11450 9092 11452
rect 9116 11450 9172 11452
rect 9196 11450 9252 11452
rect 8956 11398 8982 11450
rect 8982 11398 9012 11450
rect 9036 11398 9046 11450
rect 9046 11398 9092 11450
rect 9116 11398 9162 11450
rect 9162 11398 9172 11450
rect 9196 11398 9226 11450
rect 9226 11398 9252 11450
rect 8956 11396 9012 11398
rect 9036 11396 9092 11398
rect 9116 11396 9172 11398
rect 9196 11396 9252 11398
rect 8942 10648 8998 10704
rect 8956 10362 9012 10364
rect 9036 10362 9092 10364
rect 9116 10362 9172 10364
rect 9196 10362 9252 10364
rect 8956 10310 8982 10362
rect 8982 10310 9012 10362
rect 9036 10310 9046 10362
rect 9046 10310 9092 10362
rect 9116 10310 9162 10362
rect 9162 10310 9172 10362
rect 9196 10310 9226 10362
rect 9226 10310 9252 10362
rect 8956 10308 9012 10310
rect 9036 10308 9092 10310
rect 9116 10308 9172 10310
rect 9196 10308 9252 10310
rect 8956 9274 9012 9276
rect 9036 9274 9092 9276
rect 9116 9274 9172 9276
rect 9196 9274 9252 9276
rect 8956 9222 8982 9274
rect 8982 9222 9012 9274
rect 9036 9222 9046 9274
rect 9046 9222 9092 9274
rect 9116 9222 9162 9274
rect 9162 9222 9172 9274
rect 9196 9222 9226 9274
rect 9226 9222 9252 9274
rect 8956 9220 9012 9222
rect 9036 9220 9092 9222
rect 9116 9220 9172 9222
rect 9196 9220 9252 9222
rect 8956 8186 9012 8188
rect 9036 8186 9092 8188
rect 9116 8186 9172 8188
rect 9196 8186 9252 8188
rect 8956 8134 8982 8186
rect 8982 8134 9012 8186
rect 9036 8134 9046 8186
rect 9046 8134 9092 8186
rect 9116 8134 9162 8186
rect 9162 8134 9172 8186
rect 9196 8134 9226 8186
rect 9226 8134 9252 8186
rect 8956 8132 9012 8134
rect 9036 8132 9092 8134
rect 9116 8132 9172 8134
rect 9196 8132 9252 8134
rect 12956 18522 13012 18524
rect 13036 18522 13092 18524
rect 13116 18522 13172 18524
rect 13196 18522 13252 18524
rect 12956 18470 12982 18522
rect 12982 18470 13012 18522
rect 13036 18470 13046 18522
rect 13046 18470 13092 18522
rect 13116 18470 13162 18522
rect 13162 18470 13172 18522
rect 13196 18470 13226 18522
rect 13226 18470 13252 18522
rect 12956 18468 13012 18470
rect 13036 18468 13092 18470
rect 13116 18468 13172 18470
rect 13196 18468 13252 18470
rect 11242 16496 11298 16552
rect 12530 17584 12586 17640
rect 9954 7404 10010 7440
rect 9954 7384 9956 7404
rect 9956 7384 10008 7404
rect 10008 7384 10010 7404
rect 8956 7098 9012 7100
rect 9036 7098 9092 7100
rect 9116 7098 9172 7100
rect 9196 7098 9252 7100
rect 8956 7046 8982 7098
rect 8982 7046 9012 7098
rect 9036 7046 9046 7098
rect 9046 7046 9092 7098
rect 9116 7046 9162 7098
rect 9162 7046 9172 7098
rect 9196 7046 9226 7098
rect 9226 7046 9252 7098
rect 8956 7044 9012 7046
rect 9036 7044 9092 7046
rect 9116 7044 9172 7046
rect 9196 7044 9252 7046
rect 8956 6010 9012 6012
rect 9036 6010 9092 6012
rect 9116 6010 9172 6012
rect 9196 6010 9252 6012
rect 8956 5958 8982 6010
rect 8982 5958 9012 6010
rect 9036 5958 9046 6010
rect 9046 5958 9092 6010
rect 9116 5958 9162 6010
rect 9162 5958 9172 6010
rect 9196 5958 9226 6010
rect 9226 5958 9252 6010
rect 8956 5956 9012 5958
rect 9036 5956 9092 5958
rect 9116 5956 9172 5958
rect 9196 5956 9252 5958
rect 11794 13912 11850 13968
rect 12956 17434 13012 17436
rect 13036 17434 13092 17436
rect 13116 17434 13172 17436
rect 13196 17434 13252 17436
rect 12956 17382 12982 17434
rect 12982 17382 13012 17434
rect 13036 17382 13046 17434
rect 13046 17382 13092 17434
rect 13116 17382 13162 17434
rect 13162 17382 13172 17434
rect 13196 17382 13226 17434
rect 13226 17382 13252 17434
rect 12956 17380 13012 17382
rect 13036 17380 13092 17382
rect 13116 17380 13172 17382
rect 13196 17380 13252 17382
rect 12956 16346 13012 16348
rect 13036 16346 13092 16348
rect 13116 16346 13172 16348
rect 13196 16346 13252 16348
rect 12956 16294 12982 16346
rect 12982 16294 13012 16346
rect 13036 16294 13046 16346
rect 13046 16294 13092 16346
rect 13116 16294 13162 16346
rect 13162 16294 13172 16346
rect 13196 16294 13226 16346
rect 13226 16294 13252 16346
rect 12956 16292 13012 16294
rect 13036 16292 13092 16294
rect 13116 16292 13172 16294
rect 13196 16292 13252 16294
rect 12956 15258 13012 15260
rect 13036 15258 13092 15260
rect 13116 15258 13172 15260
rect 13196 15258 13252 15260
rect 12956 15206 12982 15258
rect 12982 15206 13012 15258
rect 13036 15206 13046 15258
rect 13046 15206 13092 15258
rect 13116 15206 13162 15258
rect 13162 15206 13172 15258
rect 13196 15206 13226 15258
rect 13226 15206 13252 15258
rect 12956 15204 13012 15206
rect 13036 15204 13092 15206
rect 13116 15204 13172 15206
rect 13196 15204 13252 15206
rect 4956 3290 5012 3292
rect 5036 3290 5092 3292
rect 5116 3290 5172 3292
rect 5196 3290 5252 3292
rect 4956 3238 4982 3290
rect 4982 3238 5012 3290
rect 5036 3238 5046 3290
rect 5046 3238 5092 3290
rect 5116 3238 5162 3290
rect 5162 3238 5172 3290
rect 5196 3238 5226 3290
rect 5226 3238 5252 3290
rect 4956 3236 5012 3238
rect 5036 3236 5092 3238
rect 5116 3236 5172 3238
rect 5196 3236 5252 3238
rect 1214 1944 1270 2000
rect 4956 2202 5012 2204
rect 5036 2202 5092 2204
rect 5116 2202 5172 2204
rect 5196 2202 5252 2204
rect 4956 2150 4982 2202
rect 4982 2150 5012 2202
rect 5036 2150 5046 2202
rect 5046 2150 5092 2202
rect 5116 2150 5162 2202
rect 5162 2150 5172 2202
rect 5196 2150 5226 2202
rect 5226 2150 5252 2202
rect 4956 2148 5012 2150
rect 5036 2148 5092 2150
rect 5116 2148 5172 2150
rect 5196 2148 5252 2150
rect 8956 4922 9012 4924
rect 9036 4922 9092 4924
rect 9116 4922 9172 4924
rect 9196 4922 9252 4924
rect 8956 4870 8982 4922
rect 8982 4870 9012 4922
rect 9036 4870 9046 4922
rect 9046 4870 9092 4922
rect 9116 4870 9162 4922
rect 9162 4870 9172 4922
rect 9196 4870 9226 4922
rect 9226 4870 9252 4922
rect 8956 4868 9012 4870
rect 9036 4868 9092 4870
rect 9116 4868 9172 4870
rect 9196 4868 9252 4870
rect 9678 4256 9734 4312
rect 8956 3834 9012 3836
rect 9036 3834 9092 3836
rect 9116 3834 9172 3836
rect 9196 3834 9252 3836
rect 8956 3782 8982 3834
rect 8982 3782 9012 3834
rect 9036 3782 9046 3834
rect 9046 3782 9092 3834
rect 9116 3782 9162 3834
rect 9162 3782 9172 3834
rect 9196 3782 9226 3834
rect 9226 3782 9252 3834
rect 8956 3780 9012 3782
rect 9036 3780 9092 3782
rect 9116 3780 9172 3782
rect 9196 3780 9252 3782
rect 9586 3576 9642 3632
rect 8956 2746 9012 2748
rect 9036 2746 9092 2748
rect 9116 2746 9172 2748
rect 9196 2746 9252 2748
rect 8956 2694 8982 2746
rect 8982 2694 9012 2746
rect 9036 2694 9046 2746
rect 9046 2694 9092 2746
rect 9116 2694 9162 2746
rect 9162 2694 9172 2746
rect 9196 2694 9226 2746
rect 9226 2694 9252 2746
rect 8956 2692 9012 2694
rect 9036 2692 9092 2694
rect 9116 2692 9172 2694
rect 9196 2692 9252 2694
rect 16956 21242 17012 21244
rect 17036 21242 17092 21244
rect 17116 21242 17172 21244
rect 17196 21242 17252 21244
rect 16956 21190 16982 21242
rect 16982 21190 17012 21242
rect 17036 21190 17046 21242
rect 17046 21190 17092 21242
rect 17116 21190 17162 21242
rect 17162 21190 17172 21242
rect 17196 21190 17226 21242
rect 17226 21190 17252 21242
rect 16956 21188 17012 21190
rect 17036 21188 17092 21190
rect 17116 21188 17172 21190
rect 17196 21188 17252 21190
rect 16956 20154 17012 20156
rect 17036 20154 17092 20156
rect 17116 20154 17172 20156
rect 17196 20154 17252 20156
rect 16956 20102 16982 20154
rect 16982 20102 17012 20154
rect 17036 20102 17046 20154
rect 17046 20102 17092 20154
rect 17116 20102 17162 20154
rect 17162 20102 17172 20154
rect 17196 20102 17226 20154
rect 17226 20102 17252 20154
rect 16956 20100 17012 20102
rect 17036 20100 17092 20102
rect 17116 20100 17172 20102
rect 17196 20100 17252 20102
rect 13910 17720 13966 17776
rect 14094 16496 14150 16552
rect 12956 14170 13012 14172
rect 13036 14170 13092 14172
rect 13116 14170 13172 14172
rect 13196 14170 13252 14172
rect 12956 14118 12982 14170
rect 12982 14118 13012 14170
rect 13036 14118 13046 14170
rect 13046 14118 13092 14170
rect 13116 14118 13162 14170
rect 13162 14118 13172 14170
rect 13196 14118 13226 14170
rect 13226 14118 13252 14170
rect 12956 14116 13012 14118
rect 13036 14116 13092 14118
rect 13116 14116 13172 14118
rect 13196 14116 13252 14118
rect 16956 19066 17012 19068
rect 17036 19066 17092 19068
rect 17116 19066 17172 19068
rect 17196 19066 17252 19068
rect 16956 19014 16982 19066
rect 16982 19014 17012 19066
rect 17036 19014 17046 19066
rect 17046 19014 17092 19066
rect 17116 19014 17162 19066
rect 17162 19014 17172 19066
rect 17196 19014 17226 19066
rect 17226 19014 17252 19066
rect 16956 19012 17012 19014
rect 17036 19012 17092 19014
rect 17116 19012 17172 19014
rect 17196 19012 17252 19014
rect 13634 13776 13690 13832
rect 12956 13082 13012 13084
rect 13036 13082 13092 13084
rect 13116 13082 13172 13084
rect 13196 13082 13252 13084
rect 12956 13030 12982 13082
rect 12982 13030 13012 13082
rect 13036 13030 13046 13082
rect 13046 13030 13092 13082
rect 13116 13030 13162 13082
rect 13162 13030 13172 13082
rect 13196 13030 13226 13082
rect 13226 13030 13252 13082
rect 12956 13028 13012 13030
rect 13036 13028 13092 13030
rect 13116 13028 13172 13030
rect 13196 13028 13252 13030
rect 13818 13232 13874 13288
rect 12714 12280 12770 12336
rect 12956 11994 13012 11996
rect 13036 11994 13092 11996
rect 13116 11994 13172 11996
rect 13196 11994 13252 11996
rect 12956 11942 12982 11994
rect 12982 11942 13012 11994
rect 13036 11942 13046 11994
rect 13046 11942 13092 11994
rect 13116 11942 13162 11994
rect 13162 11942 13172 11994
rect 13196 11942 13226 11994
rect 13226 11942 13252 11994
rect 12956 11940 13012 11942
rect 13036 11940 13092 11942
rect 13116 11940 13172 11942
rect 13196 11940 13252 11942
rect 12956 10906 13012 10908
rect 13036 10906 13092 10908
rect 13116 10906 13172 10908
rect 13196 10906 13252 10908
rect 12956 10854 12982 10906
rect 12982 10854 13012 10906
rect 13036 10854 13046 10906
rect 13046 10854 13092 10906
rect 13116 10854 13162 10906
rect 13162 10854 13172 10906
rect 13196 10854 13226 10906
rect 13226 10854 13252 10906
rect 12956 10852 13012 10854
rect 13036 10852 13092 10854
rect 13116 10852 13172 10854
rect 13196 10852 13252 10854
rect 12956 9818 13012 9820
rect 13036 9818 13092 9820
rect 13116 9818 13172 9820
rect 13196 9818 13252 9820
rect 12956 9766 12982 9818
rect 12982 9766 13012 9818
rect 13036 9766 13046 9818
rect 13046 9766 13092 9818
rect 13116 9766 13162 9818
rect 13162 9766 13172 9818
rect 13196 9766 13226 9818
rect 13226 9766 13252 9818
rect 12956 9764 13012 9766
rect 13036 9764 13092 9766
rect 13116 9764 13172 9766
rect 13196 9764 13252 9766
rect 12956 8730 13012 8732
rect 13036 8730 13092 8732
rect 13116 8730 13172 8732
rect 13196 8730 13252 8732
rect 12956 8678 12982 8730
rect 12982 8678 13012 8730
rect 13036 8678 13046 8730
rect 13046 8678 13092 8730
rect 13116 8678 13162 8730
rect 13162 8678 13172 8730
rect 13196 8678 13226 8730
rect 13226 8678 13252 8730
rect 12956 8676 13012 8678
rect 13036 8676 13092 8678
rect 13116 8676 13172 8678
rect 13196 8676 13252 8678
rect 13634 8880 13690 8936
rect 12956 7642 13012 7644
rect 13036 7642 13092 7644
rect 13116 7642 13172 7644
rect 13196 7642 13252 7644
rect 12956 7590 12982 7642
rect 12982 7590 13012 7642
rect 13036 7590 13046 7642
rect 13046 7590 13092 7642
rect 13116 7590 13162 7642
rect 13162 7590 13172 7642
rect 13196 7590 13226 7642
rect 13226 7590 13252 7642
rect 12956 7588 13012 7590
rect 13036 7588 13092 7590
rect 13116 7588 13172 7590
rect 13196 7588 13252 7590
rect 13726 7384 13782 7440
rect 12956 6554 13012 6556
rect 13036 6554 13092 6556
rect 13116 6554 13172 6556
rect 13196 6554 13252 6556
rect 12956 6502 12982 6554
rect 12982 6502 13012 6554
rect 13036 6502 13046 6554
rect 13046 6502 13092 6554
rect 13116 6502 13162 6554
rect 13162 6502 13172 6554
rect 13196 6502 13226 6554
rect 13226 6502 13252 6554
rect 12956 6500 13012 6502
rect 13036 6500 13092 6502
rect 13116 6500 13172 6502
rect 13196 6500 13252 6502
rect 12956 5466 13012 5468
rect 13036 5466 13092 5468
rect 13116 5466 13172 5468
rect 13196 5466 13252 5468
rect 12956 5414 12982 5466
rect 12982 5414 13012 5466
rect 13036 5414 13046 5466
rect 13046 5414 13092 5466
rect 13116 5414 13162 5466
rect 13162 5414 13172 5466
rect 13196 5414 13226 5466
rect 13226 5414 13252 5466
rect 12956 5412 13012 5414
rect 13036 5412 13092 5414
rect 13116 5412 13172 5414
rect 13196 5412 13252 5414
rect 11426 4256 11482 4312
rect 11978 4256 12034 4312
rect 8114 2352 8170 2408
rect 12956 4378 13012 4380
rect 13036 4378 13092 4380
rect 13116 4378 13172 4380
rect 13196 4378 13252 4380
rect 12956 4326 12982 4378
rect 12982 4326 13012 4378
rect 13036 4326 13046 4378
rect 13046 4326 13092 4378
rect 13116 4326 13162 4378
rect 13162 4326 13172 4378
rect 13196 4326 13226 4378
rect 13226 4326 13252 4378
rect 12956 4324 13012 4326
rect 13036 4324 13092 4326
rect 13116 4324 13172 4326
rect 13196 4324 13252 4326
rect 16956 17978 17012 17980
rect 17036 17978 17092 17980
rect 17116 17978 17172 17980
rect 17196 17978 17252 17980
rect 16956 17926 16982 17978
rect 16982 17926 17012 17978
rect 17036 17926 17046 17978
rect 17046 17926 17092 17978
rect 17116 17926 17162 17978
rect 17162 17926 17172 17978
rect 17196 17926 17226 17978
rect 17226 17926 17252 17978
rect 16956 17924 17012 17926
rect 17036 17924 17092 17926
rect 17116 17924 17172 17926
rect 17196 17924 17252 17926
rect 16854 17584 16910 17640
rect 20350 22616 20406 22672
rect 20956 21786 21012 21788
rect 21036 21786 21092 21788
rect 21116 21786 21172 21788
rect 21196 21786 21252 21788
rect 20956 21734 20982 21786
rect 20982 21734 21012 21786
rect 21036 21734 21046 21786
rect 21046 21734 21092 21786
rect 21116 21734 21162 21786
rect 21162 21734 21172 21786
rect 21196 21734 21226 21786
rect 21226 21734 21252 21786
rect 20956 21732 21012 21734
rect 21036 21732 21092 21734
rect 21116 21732 21172 21734
rect 21196 21732 21252 21734
rect 21362 21392 21418 21448
rect 20956 20698 21012 20700
rect 21036 20698 21092 20700
rect 21116 20698 21172 20700
rect 21196 20698 21252 20700
rect 20956 20646 20982 20698
rect 20982 20646 21012 20698
rect 21036 20646 21046 20698
rect 21046 20646 21092 20698
rect 21116 20646 21162 20698
rect 21162 20646 21172 20698
rect 21196 20646 21226 20698
rect 21226 20646 21252 20698
rect 20956 20644 21012 20646
rect 21036 20644 21092 20646
rect 21116 20644 21172 20646
rect 21196 20644 21252 20646
rect 17498 17040 17554 17096
rect 16956 16890 17012 16892
rect 17036 16890 17092 16892
rect 17116 16890 17172 16892
rect 17196 16890 17252 16892
rect 16956 16838 16982 16890
rect 16982 16838 17012 16890
rect 17036 16838 17046 16890
rect 17046 16838 17092 16890
rect 17116 16838 17162 16890
rect 17162 16838 17172 16890
rect 17196 16838 17226 16890
rect 17226 16838 17252 16890
rect 16956 16836 17012 16838
rect 17036 16836 17092 16838
rect 17116 16836 17172 16838
rect 17196 16836 17252 16838
rect 16956 15802 17012 15804
rect 17036 15802 17092 15804
rect 17116 15802 17172 15804
rect 17196 15802 17252 15804
rect 16956 15750 16982 15802
rect 16982 15750 17012 15802
rect 17036 15750 17046 15802
rect 17046 15750 17092 15802
rect 17116 15750 17162 15802
rect 17162 15750 17172 15802
rect 17196 15750 17226 15802
rect 17226 15750 17252 15802
rect 16956 15748 17012 15750
rect 17036 15748 17092 15750
rect 17116 15748 17172 15750
rect 17196 15748 17252 15750
rect 16956 14714 17012 14716
rect 17036 14714 17092 14716
rect 17116 14714 17172 14716
rect 17196 14714 17252 14716
rect 16956 14662 16982 14714
rect 16982 14662 17012 14714
rect 17036 14662 17046 14714
rect 17046 14662 17092 14714
rect 17116 14662 17162 14714
rect 17162 14662 17172 14714
rect 17196 14662 17226 14714
rect 17226 14662 17252 14714
rect 16956 14660 17012 14662
rect 17036 14660 17092 14662
rect 17116 14660 17172 14662
rect 17196 14660 17252 14662
rect 13358 3576 13414 3632
rect 14094 4664 14150 4720
rect 12956 3290 13012 3292
rect 13036 3290 13092 3292
rect 13116 3290 13172 3292
rect 13196 3290 13252 3292
rect 12956 3238 12982 3290
rect 12982 3238 13012 3290
rect 13036 3238 13046 3290
rect 13046 3238 13092 3290
rect 13116 3238 13162 3290
rect 13162 3238 13172 3290
rect 13196 3238 13226 3290
rect 13226 3238 13252 3290
rect 12956 3236 13012 3238
rect 13036 3236 13092 3238
rect 13116 3236 13172 3238
rect 13196 3236 13252 3238
rect 13082 3032 13138 3088
rect 12956 2202 13012 2204
rect 13036 2202 13092 2204
rect 13116 2202 13172 2204
rect 13196 2202 13252 2204
rect 12956 2150 12982 2202
rect 12982 2150 13012 2202
rect 13036 2150 13046 2202
rect 13046 2150 13092 2202
rect 13116 2150 13162 2202
rect 13162 2150 13172 2202
rect 13196 2150 13226 2202
rect 13226 2150 13252 2202
rect 12956 2148 13012 2150
rect 13036 2148 13092 2150
rect 13116 2148 13172 2150
rect 13196 2148 13252 2150
rect 12438 1944 12494 2000
rect 14922 4664 14978 4720
rect 14646 3440 14702 3496
rect 13450 1264 13506 1320
rect 16956 13626 17012 13628
rect 17036 13626 17092 13628
rect 17116 13626 17172 13628
rect 17196 13626 17252 13628
rect 16956 13574 16982 13626
rect 16982 13574 17012 13626
rect 17036 13574 17046 13626
rect 17046 13574 17092 13626
rect 17116 13574 17162 13626
rect 17162 13574 17172 13626
rect 17196 13574 17226 13626
rect 17226 13574 17252 13626
rect 16956 13572 17012 13574
rect 17036 13572 17092 13574
rect 17116 13572 17172 13574
rect 17196 13572 17252 13574
rect 18694 15000 18750 15056
rect 16956 12538 17012 12540
rect 17036 12538 17092 12540
rect 17116 12538 17172 12540
rect 17196 12538 17252 12540
rect 16956 12486 16982 12538
rect 16982 12486 17012 12538
rect 17036 12486 17046 12538
rect 17046 12486 17092 12538
rect 17116 12486 17162 12538
rect 17162 12486 17172 12538
rect 17196 12486 17226 12538
rect 17226 12486 17252 12538
rect 16956 12484 17012 12486
rect 17036 12484 17092 12486
rect 17116 12484 17172 12486
rect 17196 12484 17252 12486
rect 16956 11450 17012 11452
rect 17036 11450 17092 11452
rect 17116 11450 17172 11452
rect 17196 11450 17252 11452
rect 16956 11398 16982 11450
rect 16982 11398 17012 11450
rect 17036 11398 17046 11450
rect 17046 11398 17092 11450
rect 17116 11398 17162 11450
rect 17162 11398 17172 11450
rect 17196 11398 17226 11450
rect 17226 11398 17252 11450
rect 16956 11396 17012 11398
rect 17036 11396 17092 11398
rect 17116 11396 17172 11398
rect 17196 11396 17252 11398
rect 16956 10362 17012 10364
rect 17036 10362 17092 10364
rect 17116 10362 17172 10364
rect 17196 10362 17252 10364
rect 16956 10310 16982 10362
rect 16982 10310 17012 10362
rect 17036 10310 17046 10362
rect 17046 10310 17092 10362
rect 17116 10310 17162 10362
rect 17162 10310 17172 10362
rect 17196 10310 17226 10362
rect 17226 10310 17252 10362
rect 16956 10308 17012 10310
rect 17036 10308 17092 10310
rect 17116 10308 17172 10310
rect 17196 10308 17252 10310
rect 16956 9274 17012 9276
rect 17036 9274 17092 9276
rect 17116 9274 17172 9276
rect 17196 9274 17252 9276
rect 16956 9222 16982 9274
rect 16982 9222 17012 9274
rect 17036 9222 17046 9274
rect 17046 9222 17092 9274
rect 17116 9222 17162 9274
rect 17162 9222 17172 9274
rect 17196 9222 17226 9274
rect 17226 9222 17252 9274
rect 16956 9220 17012 9222
rect 17036 9220 17092 9222
rect 17116 9220 17172 9222
rect 17196 9220 17252 9222
rect 17314 8880 17370 8936
rect 16956 8186 17012 8188
rect 17036 8186 17092 8188
rect 17116 8186 17172 8188
rect 17196 8186 17252 8188
rect 16956 8134 16982 8186
rect 16982 8134 17012 8186
rect 17036 8134 17046 8186
rect 17046 8134 17092 8186
rect 17116 8134 17162 8186
rect 17162 8134 17172 8186
rect 17196 8134 17226 8186
rect 17226 8134 17252 8186
rect 16956 8132 17012 8134
rect 17036 8132 17092 8134
rect 17116 8132 17172 8134
rect 17196 8132 17252 8134
rect 17314 7384 17370 7440
rect 17774 7248 17830 7304
rect 16956 7098 17012 7100
rect 17036 7098 17092 7100
rect 17116 7098 17172 7100
rect 17196 7098 17252 7100
rect 16956 7046 16982 7098
rect 16982 7046 17012 7098
rect 17036 7046 17046 7098
rect 17046 7046 17092 7098
rect 17116 7046 17162 7098
rect 17162 7046 17172 7098
rect 17196 7046 17226 7098
rect 17226 7046 17252 7098
rect 16956 7044 17012 7046
rect 17036 7044 17092 7046
rect 17116 7044 17172 7046
rect 17196 7044 17252 7046
rect 16956 6010 17012 6012
rect 17036 6010 17092 6012
rect 17116 6010 17172 6012
rect 17196 6010 17252 6012
rect 16956 5958 16982 6010
rect 16982 5958 17012 6010
rect 17036 5958 17046 6010
rect 17046 5958 17092 6010
rect 17116 5958 17162 6010
rect 17162 5958 17172 6010
rect 17196 5958 17226 6010
rect 17226 5958 17252 6010
rect 16956 5956 17012 5958
rect 17036 5956 17092 5958
rect 17116 5956 17172 5958
rect 17196 5956 17252 5958
rect 16956 4922 17012 4924
rect 17036 4922 17092 4924
rect 17116 4922 17172 4924
rect 17196 4922 17252 4924
rect 16956 4870 16982 4922
rect 16982 4870 17012 4922
rect 17036 4870 17046 4922
rect 17046 4870 17092 4922
rect 17116 4870 17162 4922
rect 17162 4870 17172 4922
rect 17196 4870 17226 4922
rect 17226 4870 17252 4922
rect 16956 4868 17012 4870
rect 17036 4868 17092 4870
rect 17116 4868 17172 4870
rect 17196 4868 17252 4870
rect 16956 3834 17012 3836
rect 17036 3834 17092 3836
rect 17116 3834 17172 3836
rect 17196 3834 17252 3836
rect 16956 3782 16982 3834
rect 16982 3782 17012 3834
rect 17036 3782 17046 3834
rect 17046 3782 17092 3834
rect 17116 3782 17162 3834
rect 17162 3782 17172 3834
rect 17196 3782 17226 3834
rect 17226 3782 17252 3834
rect 16956 3780 17012 3782
rect 17036 3780 17092 3782
rect 17116 3780 17172 3782
rect 17196 3780 17252 3782
rect 16956 2746 17012 2748
rect 17036 2746 17092 2748
rect 17116 2746 17172 2748
rect 17196 2746 17252 2748
rect 16956 2694 16982 2746
rect 16982 2694 17012 2746
rect 17036 2694 17046 2746
rect 17046 2694 17092 2746
rect 17116 2694 17162 2746
rect 17162 2694 17172 2746
rect 17196 2694 17226 2746
rect 17226 2694 17252 2746
rect 16956 2692 17012 2694
rect 17036 2692 17092 2694
rect 17116 2692 17172 2694
rect 17196 2692 17252 2694
rect 16394 2352 16450 2408
rect 17130 2352 17186 2408
rect 18510 5072 18566 5128
rect 21270 20168 21326 20224
rect 20956 19610 21012 19612
rect 21036 19610 21092 19612
rect 21116 19610 21172 19612
rect 21196 19610 21252 19612
rect 20956 19558 20982 19610
rect 20982 19558 21012 19610
rect 21036 19558 21046 19610
rect 21046 19558 21092 19610
rect 21116 19558 21162 19610
rect 21162 19558 21172 19610
rect 21196 19558 21226 19610
rect 21226 19558 21252 19610
rect 20956 19556 21012 19558
rect 21036 19556 21092 19558
rect 21116 19556 21172 19558
rect 21196 19556 21252 19558
rect 21270 18808 21326 18864
rect 20956 18522 21012 18524
rect 21036 18522 21092 18524
rect 21116 18522 21172 18524
rect 21196 18522 21252 18524
rect 20956 18470 20982 18522
rect 20982 18470 21012 18522
rect 21036 18470 21046 18522
rect 21046 18470 21092 18522
rect 21116 18470 21162 18522
rect 21162 18470 21172 18522
rect 21196 18470 21226 18522
rect 21226 18470 21252 18522
rect 20956 18468 21012 18470
rect 21036 18468 21092 18470
rect 21116 18468 21172 18470
rect 21196 18468 21252 18470
rect 21270 17584 21326 17640
rect 20956 17434 21012 17436
rect 21036 17434 21092 17436
rect 21116 17434 21172 17436
rect 21196 17434 21252 17436
rect 20956 17382 20982 17434
rect 20982 17382 21012 17434
rect 21036 17382 21046 17434
rect 21046 17382 21092 17434
rect 21116 17382 21162 17434
rect 21162 17382 21172 17434
rect 21196 17382 21226 17434
rect 21226 17382 21252 17434
rect 20956 17380 21012 17382
rect 21036 17380 21092 17382
rect 21116 17380 21172 17382
rect 21196 17380 21252 17382
rect 20956 16346 21012 16348
rect 21036 16346 21092 16348
rect 21116 16346 21172 16348
rect 21196 16346 21252 16348
rect 20956 16294 20982 16346
rect 20982 16294 21012 16346
rect 21036 16294 21046 16346
rect 21046 16294 21092 16346
rect 21116 16294 21162 16346
rect 21162 16294 21172 16346
rect 21196 16294 21226 16346
rect 21226 16294 21252 16346
rect 20956 16292 21012 16294
rect 21036 16292 21092 16294
rect 21116 16292 21172 16294
rect 21196 16292 21252 16294
rect 20718 15952 20774 16008
rect 20956 15258 21012 15260
rect 21036 15258 21092 15260
rect 21116 15258 21172 15260
rect 21196 15258 21252 15260
rect 20956 15206 20982 15258
rect 20982 15206 21012 15258
rect 21036 15206 21046 15258
rect 21046 15206 21092 15258
rect 21116 15206 21162 15258
rect 21162 15206 21172 15258
rect 21196 15206 21226 15258
rect 21226 15206 21252 15258
rect 20956 15204 21012 15206
rect 21036 15204 21092 15206
rect 21116 15204 21172 15206
rect 21196 15204 21252 15206
rect 20956 14170 21012 14172
rect 21036 14170 21092 14172
rect 21116 14170 21172 14172
rect 21196 14170 21252 14172
rect 20956 14118 20982 14170
rect 20982 14118 21012 14170
rect 21036 14118 21046 14170
rect 21046 14118 21092 14170
rect 21116 14118 21162 14170
rect 21162 14118 21172 14170
rect 21196 14118 21226 14170
rect 21226 14118 21252 14170
rect 20956 14116 21012 14118
rect 21036 14116 21092 14118
rect 21116 14116 21172 14118
rect 21196 14116 21252 14118
rect 20626 13912 20682 13968
rect 19798 10648 19854 10704
rect 19338 9016 19394 9072
rect 18878 7928 18934 7984
rect 19798 9288 19854 9344
rect 18234 2352 18290 2408
rect 18602 1128 18658 1184
rect 21546 16360 21602 16416
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 21086 10104 21142 10160
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 20902 9016 20958 9072
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 21362 13096 21418 13152
rect 21362 11872 21418 11928
rect 23570 15680 23626 15736
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 21362 5344 21418 5400
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 20626 3032 20682 3088
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
<< metal3 >>
rect 0 23128 480 23248
rect 23520 23128 24000 23248
rect 62 22674 122 23128
rect 1577 22674 1643 22677
rect 62 22672 1643 22674
rect 62 22616 1582 22672
rect 1638 22616 1643 22672
rect 62 22614 1643 22616
rect 1577 22611 1643 22614
rect 20345 22674 20411 22677
rect 23614 22674 23674 23128
rect 20345 22672 23674 22674
rect 20345 22616 20350 22672
rect 20406 22616 23674 22672
rect 20345 22614 23674 22616
rect 20345 22611 20411 22614
rect 23520 21904 24000 22024
rect 4944 21792 5264 21793
rect 0 21632 480 21752
rect 4944 21728 4952 21792
rect 5016 21728 5032 21792
rect 5096 21728 5112 21792
rect 5176 21728 5192 21792
rect 5256 21728 5264 21792
rect 4944 21727 5264 21728
rect 12944 21792 13264 21793
rect 12944 21728 12952 21792
rect 13016 21728 13032 21792
rect 13096 21728 13112 21792
rect 13176 21728 13192 21792
rect 13256 21728 13264 21792
rect 12944 21727 13264 21728
rect 20944 21792 21264 21793
rect 20944 21728 20952 21792
rect 21016 21728 21032 21792
rect 21096 21728 21112 21792
rect 21176 21728 21192 21792
rect 21256 21728 21264 21792
rect 20944 21727 21264 21728
rect 62 21178 122 21632
rect 21357 21450 21423 21453
rect 23614 21450 23674 21904
rect 21357 21448 23674 21450
rect 21357 21392 21362 21448
rect 21418 21392 23674 21448
rect 21357 21390 23674 21392
rect 21357 21387 21423 21390
rect 8944 21248 9264 21249
rect 8944 21184 8952 21248
rect 9016 21184 9032 21248
rect 9096 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9264 21248
rect 8944 21183 9264 21184
rect 16944 21248 17264 21249
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 21183 17264 21184
rect 1117 21178 1183 21181
rect 62 21176 1183 21178
rect 62 21120 1122 21176
rect 1178 21120 1183 21176
rect 62 21118 1183 21120
rect 1117 21115 1183 21118
rect 4944 20704 5264 20705
rect 4944 20640 4952 20704
rect 5016 20640 5032 20704
rect 5096 20640 5112 20704
rect 5176 20640 5192 20704
rect 5256 20640 5264 20704
rect 4944 20639 5264 20640
rect 12944 20704 13264 20705
rect 12944 20640 12952 20704
rect 13016 20640 13032 20704
rect 13096 20640 13112 20704
rect 13176 20640 13192 20704
rect 13256 20640 13264 20704
rect 12944 20639 13264 20640
rect 20944 20704 21264 20705
rect 20944 20640 20952 20704
rect 21016 20640 21032 20704
rect 21096 20640 21112 20704
rect 21176 20640 21192 20704
rect 21256 20640 21264 20704
rect 23520 20680 24000 20800
rect 20944 20639 21264 20640
rect 0 20136 480 20256
rect 21265 20226 21331 20229
rect 23614 20226 23674 20680
rect 21265 20224 23674 20226
rect 21265 20168 21270 20224
rect 21326 20168 23674 20224
rect 21265 20166 23674 20168
rect 21265 20163 21331 20166
rect 8944 20160 9264 20161
rect 62 19682 122 20136
rect 8944 20096 8952 20160
rect 9016 20096 9032 20160
rect 9096 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9264 20160
rect 8944 20095 9264 20096
rect 16944 20160 17264 20161
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 16944 20095 17264 20096
rect 1485 19818 1551 19821
rect 11605 19818 11671 19821
rect 1485 19816 11671 19818
rect 1485 19760 1490 19816
rect 1546 19760 11610 19816
rect 11666 19760 11671 19816
rect 1485 19758 11671 19760
rect 1485 19755 1551 19758
rect 11605 19755 11671 19758
rect 1577 19682 1643 19685
rect 62 19680 1643 19682
rect 62 19624 1582 19680
rect 1638 19624 1643 19680
rect 62 19622 1643 19624
rect 1577 19619 1643 19622
rect 4944 19616 5264 19617
rect 4944 19552 4952 19616
rect 5016 19552 5032 19616
rect 5096 19552 5112 19616
rect 5176 19552 5192 19616
rect 5256 19552 5264 19616
rect 4944 19551 5264 19552
rect 12944 19616 13264 19617
rect 12944 19552 12952 19616
rect 13016 19552 13032 19616
rect 13096 19552 13112 19616
rect 13176 19552 13192 19616
rect 13256 19552 13264 19616
rect 12944 19551 13264 19552
rect 20944 19616 21264 19617
rect 20944 19552 20952 19616
rect 21016 19552 21032 19616
rect 21096 19552 21112 19616
rect 21176 19552 21192 19616
rect 21256 19552 21264 19616
rect 20944 19551 21264 19552
rect 23520 19320 24000 19440
rect 8944 19072 9264 19073
rect 8944 19008 8952 19072
rect 9016 19008 9032 19072
rect 9096 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9264 19072
rect 8944 19007 9264 19008
rect 16944 19072 17264 19073
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 19007 17264 19008
rect 21265 18866 21331 18869
rect 23614 18866 23674 19320
rect 21265 18864 23674 18866
rect 21265 18808 21270 18864
rect 21326 18808 23674 18864
rect 21265 18806 23674 18808
rect 21265 18803 21331 18806
rect 0 18640 480 18760
rect 62 18186 122 18640
rect 4944 18528 5264 18529
rect 4944 18464 4952 18528
rect 5016 18464 5032 18528
rect 5096 18464 5112 18528
rect 5176 18464 5192 18528
rect 5256 18464 5264 18528
rect 4944 18463 5264 18464
rect 12944 18528 13264 18529
rect 12944 18464 12952 18528
rect 13016 18464 13032 18528
rect 13096 18464 13112 18528
rect 13176 18464 13192 18528
rect 13256 18464 13264 18528
rect 12944 18463 13264 18464
rect 20944 18528 21264 18529
rect 20944 18464 20952 18528
rect 21016 18464 21032 18528
rect 21096 18464 21112 18528
rect 21176 18464 21192 18528
rect 21256 18464 21264 18528
rect 20944 18463 21264 18464
rect 1393 18186 1459 18189
rect 62 18184 1459 18186
rect 62 18128 1398 18184
rect 1454 18128 1459 18184
rect 62 18126 1459 18128
rect 1393 18123 1459 18126
rect 23520 18096 24000 18216
rect 8944 17984 9264 17985
rect 8944 17920 8952 17984
rect 9016 17920 9032 17984
rect 9096 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9264 17984
rect 8944 17919 9264 17920
rect 16944 17984 17264 17985
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 17919 17264 17920
rect 8385 17778 8451 17781
rect 9397 17778 9463 17781
rect 13905 17778 13971 17781
rect 8385 17776 13971 17778
rect 8385 17720 8390 17776
rect 8446 17720 9402 17776
rect 9458 17720 13910 17776
rect 13966 17720 13971 17776
rect 8385 17718 13971 17720
rect 8385 17715 8451 17718
rect 9397 17715 9463 17718
rect 13905 17715 13971 17718
rect 7189 17642 7255 17645
rect 10961 17642 11027 17645
rect 62 17640 11027 17642
rect 62 17584 7194 17640
rect 7250 17584 10966 17640
rect 11022 17584 11027 17640
rect 62 17582 11027 17584
rect 62 17264 122 17582
rect 7189 17579 7255 17582
rect 10961 17579 11027 17582
rect 12525 17642 12591 17645
rect 16849 17642 16915 17645
rect 12525 17640 16915 17642
rect 12525 17584 12530 17640
rect 12586 17584 16854 17640
rect 16910 17584 16915 17640
rect 12525 17582 16915 17584
rect 12525 17579 12591 17582
rect 16849 17579 16915 17582
rect 21265 17642 21331 17645
rect 23614 17642 23674 18096
rect 21265 17640 23674 17642
rect 21265 17584 21270 17640
rect 21326 17584 23674 17640
rect 21265 17582 23674 17584
rect 21265 17579 21331 17582
rect 4944 17440 5264 17441
rect 4944 17376 4952 17440
rect 5016 17376 5032 17440
rect 5096 17376 5112 17440
rect 5176 17376 5192 17440
rect 5256 17376 5264 17440
rect 4944 17375 5264 17376
rect 12944 17440 13264 17441
rect 12944 17376 12952 17440
rect 13016 17376 13032 17440
rect 13096 17376 13112 17440
rect 13176 17376 13192 17440
rect 13256 17376 13264 17440
rect 12944 17375 13264 17376
rect 20944 17440 21264 17441
rect 20944 17376 20952 17440
rect 21016 17376 21032 17440
rect 21096 17376 21112 17440
rect 21176 17376 21192 17440
rect 21256 17376 21264 17440
rect 20944 17375 21264 17376
rect 0 17144 480 17264
rect 9305 17098 9371 17101
rect 17493 17098 17559 17101
rect 9305 17096 17559 17098
rect 9305 17040 9310 17096
rect 9366 17040 17498 17096
rect 17554 17040 17559 17096
rect 9305 17038 17559 17040
rect 9305 17035 9371 17038
rect 17493 17035 17559 17038
rect 8944 16896 9264 16897
rect 8944 16832 8952 16896
rect 9016 16832 9032 16896
rect 9096 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9264 16896
rect 8944 16831 9264 16832
rect 16944 16896 17264 16897
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 23520 16872 24000 16992
rect 16944 16831 17264 16832
rect 8293 16554 8359 16557
rect 11237 16554 11303 16557
rect 14089 16554 14155 16557
rect 8293 16552 14155 16554
rect 8293 16496 8298 16552
rect 8354 16496 11242 16552
rect 11298 16496 14094 16552
rect 14150 16496 14155 16552
rect 8293 16494 14155 16496
rect 8293 16491 8359 16494
rect 11237 16491 11303 16494
rect 14089 16491 14155 16494
rect 21541 16418 21607 16421
rect 23614 16418 23674 16872
rect 21541 16416 23674 16418
rect 21541 16360 21546 16416
rect 21602 16360 23674 16416
rect 21541 16358 23674 16360
rect 21541 16355 21607 16358
rect 4944 16352 5264 16353
rect 4944 16288 4952 16352
rect 5016 16288 5032 16352
rect 5096 16288 5112 16352
rect 5176 16288 5192 16352
rect 5256 16288 5264 16352
rect 4944 16287 5264 16288
rect 12944 16352 13264 16353
rect 12944 16288 12952 16352
rect 13016 16288 13032 16352
rect 13096 16288 13112 16352
rect 13176 16288 13192 16352
rect 13256 16288 13264 16352
rect 12944 16287 13264 16288
rect 20944 16352 21264 16353
rect 20944 16288 20952 16352
rect 21016 16288 21032 16352
rect 21096 16288 21112 16352
rect 21176 16288 21192 16352
rect 21256 16288 21264 16352
rect 20944 16287 21264 16288
rect 9305 16010 9371 16013
rect 20713 16010 20779 16013
rect 9305 16008 20779 16010
rect 9305 15952 9310 16008
rect 9366 15952 20718 16008
rect 20774 15952 20779 16008
rect 9305 15950 20779 15952
rect 9305 15947 9371 15950
rect 20713 15947 20779 15950
rect 8944 15808 9264 15809
rect 0 15648 480 15768
rect 8944 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9264 15808
rect 8944 15743 9264 15744
rect 16944 15808 17264 15809
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 15743 17264 15744
rect 23520 15738 24000 15768
rect 23484 15736 24000 15738
rect 23484 15680 23570 15736
rect 23626 15680 24000 15736
rect 23484 15678 24000 15680
rect 23520 15648 24000 15678
rect 62 15194 122 15648
rect 4944 15264 5264 15265
rect 4944 15200 4952 15264
rect 5016 15200 5032 15264
rect 5096 15200 5112 15264
rect 5176 15200 5192 15264
rect 5256 15200 5264 15264
rect 4944 15199 5264 15200
rect 12944 15264 13264 15265
rect 12944 15200 12952 15264
rect 13016 15200 13032 15264
rect 13096 15200 13112 15264
rect 13176 15200 13192 15264
rect 13256 15200 13264 15264
rect 12944 15199 13264 15200
rect 20944 15264 21264 15265
rect 20944 15200 20952 15264
rect 21016 15200 21032 15264
rect 21096 15200 21112 15264
rect 21176 15200 21192 15264
rect 21256 15200 21264 15264
rect 20944 15199 21264 15200
rect 3049 15194 3115 15197
rect 62 15192 3115 15194
rect 62 15136 3054 15192
rect 3110 15136 3115 15192
rect 62 15134 3115 15136
rect 3049 15131 3115 15134
rect 3785 15058 3851 15061
rect 8753 15058 8819 15061
rect 3785 15056 8819 15058
rect 3785 15000 3790 15056
rect 3846 15000 8758 15056
rect 8814 15000 8819 15056
rect 3785 14998 8819 15000
rect 3785 14995 3851 14998
rect 8753 14995 8819 14998
rect 10409 15058 10475 15061
rect 18689 15058 18755 15061
rect 10409 15056 18755 15058
rect 10409 15000 10414 15056
rect 10470 15000 18694 15056
rect 18750 15000 18755 15056
rect 10409 14998 18755 15000
rect 10409 14995 10475 14998
rect 18689 14995 18755 14998
rect 8944 14720 9264 14721
rect 8944 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9264 14720
rect 8944 14655 9264 14656
rect 16944 14720 17264 14721
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 14655 17264 14656
rect 23520 14288 24000 14408
rect 0 14240 480 14272
rect 0 14184 110 14240
rect 166 14184 480 14240
rect 0 14152 480 14184
rect 4944 14176 5264 14177
rect 4944 14112 4952 14176
rect 5016 14112 5032 14176
rect 5096 14112 5112 14176
rect 5176 14112 5192 14176
rect 5256 14112 5264 14176
rect 4944 14111 5264 14112
rect 12944 14176 13264 14177
rect 12944 14112 12952 14176
rect 13016 14112 13032 14176
rect 13096 14112 13112 14176
rect 13176 14112 13192 14176
rect 13256 14112 13264 14176
rect 12944 14111 13264 14112
rect 20944 14176 21264 14177
rect 20944 14112 20952 14176
rect 21016 14112 21032 14176
rect 21096 14112 21112 14176
rect 21176 14112 21192 14176
rect 21256 14112 21264 14176
rect 20944 14111 21264 14112
rect 4245 13970 4311 13973
rect 11789 13970 11855 13973
rect 4245 13968 11855 13970
rect 4245 13912 4250 13968
rect 4306 13912 11794 13968
rect 11850 13912 11855 13968
rect 4245 13910 11855 13912
rect 4245 13907 4311 13910
rect 11789 13907 11855 13910
rect 20621 13970 20687 13973
rect 23614 13970 23674 14288
rect 20621 13968 23674 13970
rect 20621 13912 20626 13968
rect 20682 13912 23674 13968
rect 20621 13910 23674 13912
rect 20621 13907 20687 13910
rect 6545 13834 6611 13837
rect 9305 13834 9371 13837
rect 13629 13834 13695 13837
rect 6545 13832 13695 13834
rect 6545 13776 6550 13832
rect 6606 13776 9310 13832
rect 9366 13776 13634 13832
rect 13690 13776 13695 13832
rect 6545 13774 13695 13776
rect 6545 13771 6611 13774
rect 9305 13771 9371 13774
rect 13629 13771 13695 13774
rect 8944 13632 9264 13633
rect 8944 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9264 13632
rect 8944 13567 9264 13568
rect 16944 13632 17264 13633
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 13567 17264 13568
rect 8293 13290 8359 13293
rect 13813 13290 13879 13293
rect 8293 13288 13879 13290
rect 8293 13232 8298 13288
rect 8354 13232 13818 13288
rect 13874 13232 13879 13288
rect 8293 13230 13879 13232
rect 8293 13227 8359 13230
rect 13813 13227 13879 13230
rect 21357 13154 21423 13157
rect 23520 13154 24000 13184
rect 21357 13152 24000 13154
rect 21357 13096 21362 13152
rect 21418 13096 24000 13152
rect 21357 13094 24000 13096
rect 21357 13091 21423 13094
rect 4944 13088 5264 13089
rect 4944 13024 4952 13088
rect 5016 13024 5032 13088
rect 5096 13024 5112 13088
rect 5176 13024 5192 13088
rect 5256 13024 5264 13088
rect 4944 13023 5264 13024
rect 12944 13088 13264 13089
rect 12944 13024 12952 13088
rect 13016 13024 13032 13088
rect 13096 13024 13112 13088
rect 13176 13024 13192 13088
rect 13256 13024 13264 13088
rect 12944 13023 13264 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 23520 13064 24000 13094
rect 20944 13023 21264 13024
rect 0 12748 480 12776
rect 0 12684 60 12748
rect 124 12684 480 12748
rect 0 12656 480 12684
rect 8944 12544 9264 12545
rect 8944 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9264 12544
rect 8944 12479 9264 12480
rect 16944 12544 17264 12545
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 12479 17264 12480
rect 54 12276 60 12340
rect 124 12338 130 12340
rect 12709 12338 12775 12341
rect 124 12336 12775 12338
rect 124 12280 12714 12336
rect 12770 12280 12775 12336
rect 124 12278 12775 12280
rect 124 12276 130 12278
rect 12709 12275 12775 12278
rect 4944 12000 5264 12001
rect 4944 11936 4952 12000
rect 5016 11936 5032 12000
rect 5096 11936 5112 12000
rect 5176 11936 5192 12000
rect 5256 11936 5264 12000
rect 4944 11935 5264 11936
rect 12944 12000 13264 12001
rect 12944 11936 12952 12000
rect 13016 11936 13032 12000
rect 13096 11936 13112 12000
rect 13176 11936 13192 12000
rect 13256 11936 13264 12000
rect 12944 11935 13264 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 21357 11930 21423 11933
rect 23520 11930 24000 11960
rect 21357 11928 24000 11930
rect 21357 11872 21362 11928
rect 21418 11872 24000 11928
rect 21357 11870 24000 11872
rect 21357 11867 21423 11870
rect 23520 11840 24000 11870
rect 8944 11456 9264 11457
rect 8944 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9264 11456
rect 8944 11391 9264 11392
rect 16944 11456 17264 11457
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 11391 17264 11392
rect 0 11248 480 11280
rect 0 11192 110 11248
rect 166 11192 480 11248
rect 0 11160 480 11192
rect 4944 10912 5264 10913
rect 4944 10848 4952 10912
rect 5016 10848 5032 10912
rect 5096 10848 5112 10912
rect 5176 10848 5192 10912
rect 5256 10848 5264 10912
rect 4944 10847 5264 10848
rect 12944 10912 13264 10913
rect 12944 10848 12952 10912
rect 13016 10848 13032 10912
rect 13096 10848 13112 10912
rect 13176 10848 13192 10912
rect 13256 10848 13264 10912
rect 12944 10847 13264 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 8937 10706 9003 10709
rect 19793 10706 19859 10709
rect 8937 10704 19859 10706
rect 8937 10648 8942 10704
rect 8998 10648 19798 10704
rect 19854 10648 19859 10704
rect 8937 10646 19859 10648
rect 8937 10643 9003 10646
rect 19793 10643 19859 10646
rect 23520 10616 24000 10736
rect 8944 10368 9264 10369
rect 8944 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9264 10368
rect 8944 10303 9264 10304
rect 16944 10368 17264 10369
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 10303 17264 10304
rect 21081 10162 21147 10165
rect 23614 10162 23674 10616
rect 21081 10160 23674 10162
rect 21081 10104 21086 10160
rect 21142 10104 23674 10160
rect 21081 10102 23674 10104
rect 21081 10099 21147 10102
rect 54 9964 60 10028
rect 124 10026 130 10028
rect 2037 10026 2103 10029
rect 4705 10026 4771 10029
rect 124 10024 4771 10026
rect 124 9968 2042 10024
rect 2098 9968 4710 10024
rect 4766 9968 4771 10024
rect 124 9966 4771 9968
rect 124 9964 130 9966
rect 2037 9963 2103 9966
rect 4705 9963 4771 9966
rect 4944 9824 5264 9825
rect 0 9756 480 9784
rect 4944 9760 4952 9824
rect 5016 9760 5032 9824
rect 5096 9760 5112 9824
rect 5176 9760 5192 9824
rect 5256 9760 5264 9824
rect 4944 9759 5264 9760
rect 12944 9824 13264 9825
rect 12944 9760 12952 9824
rect 13016 9760 13032 9824
rect 13096 9760 13112 9824
rect 13176 9760 13192 9824
rect 13256 9760 13264 9824
rect 12944 9759 13264 9760
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 0 9692 60 9756
rect 124 9692 480 9756
rect 0 9664 480 9692
rect 19793 9346 19859 9349
rect 23520 9346 24000 9376
rect 19793 9344 24000 9346
rect 19793 9288 19798 9344
rect 19854 9288 24000 9344
rect 19793 9286 24000 9288
rect 19793 9283 19859 9286
rect 8944 9280 9264 9281
rect 8944 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9264 9280
rect 8944 9215 9264 9216
rect 16944 9280 17264 9281
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 23520 9256 24000 9286
rect 16944 9215 17264 9216
rect 3509 9074 3575 9077
rect 8017 9074 8083 9077
rect 19333 9074 19399 9077
rect 20897 9074 20963 9077
rect 3509 9072 20963 9074
rect 3509 9016 3514 9072
rect 3570 9016 8022 9072
rect 8078 9016 19338 9072
rect 19394 9016 20902 9072
rect 20958 9016 20963 9072
rect 3509 9014 20963 9016
rect 3509 9011 3575 9014
rect 8017 9011 8083 9014
rect 19333 9011 19399 9014
rect 20897 9011 20963 9014
rect 13629 8938 13695 8941
rect 17309 8938 17375 8941
rect 13629 8936 17375 8938
rect 13629 8880 13634 8936
rect 13690 8880 17314 8936
rect 17370 8880 17375 8936
rect 13629 8878 17375 8880
rect 13629 8875 13695 8878
rect 17309 8875 17375 8878
rect 4944 8736 5264 8737
rect 4944 8672 4952 8736
rect 5016 8672 5032 8736
rect 5096 8672 5112 8736
rect 5176 8672 5192 8736
rect 5256 8672 5264 8736
rect 4944 8671 5264 8672
rect 12944 8736 13264 8737
rect 12944 8672 12952 8736
rect 13016 8672 13032 8736
rect 13096 8672 13112 8736
rect 13176 8672 13192 8736
rect 13256 8672 13264 8736
rect 12944 8671 13264 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 0 8256 480 8288
rect 0 8200 110 8256
rect 166 8200 480 8256
rect 0 8168 480 8200
rect 7373 8258 7439 8261
rect 7598 8258 7604 8260
rect 7373 8256 7604 8258
rect 7373 8200 7378 8256
rect 7434 8200 7604 8256
rect 7373 8198 7604 8200
rect 7373 8195 7439 8198
rect 7598 8196 7604 8198
rect 7668 8196 7674 8260
rect 8944 8192 9264 8193
rect 8944 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9264 8192
rect 8944 8127 9264 8128
rect 16944 8192 17264 8193
rect 16944 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17264 8192
rect 16944 8127 17264 8128
rect 23520 8124 24000 8152
rect 23520 8122 23612 8124
rect 23484 8062 23612 8122
rect 23520 8060 23612 8062
rect 23676 8060 24000 8124
rect 23520 8032 24000 8060
rect 18873 7986 18939 7989
rect 18873 7984 19350 7986
rect 18873 7928 18878 7984
rect 18934 7928 19350 7984
rect 18873 7926 19350 7928
rect 18873 7923 18939 7926
rect 19290 7850 19350 7926
rect 23606 7850 23612 7852
rect 19290 7790 23612 7850
rect 23606 7788 23612 7790
rect 23676 7788 23682 7852
rect 4944 7648 5264 7649
rect 4944 7584 4952 7648
rect 5016 7584 5032 7648
rect 5096 7584 5112 7648
rect 5176 7584 5192 7648
rect 5256 7584 5264 7648
rect 4944 7583 5264 7584
rect 12944 7648 13264 7649
rect 12944 7584 12952 7648
rect 13016 7584 13032 7648
rect 13096 7584 13112 7648
rect 13176 7584 13192 7648
rect 13256 7584 13264 7648
rect 12944 7583 13264 7584
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 9949 7442 10015 7445
rect 13721 7442 13787 7445
rect 9949 7440 13787 7442
rect 9949 7384 9954 7440
rect 10010 7384 13726 7440
rect 13782 7384 13787 7440
rect 9949 7382 13787 7384
rect 9949 7379 10015 7382
rect 13721 7379 13787 7382
rect 17309 7442 17375 7445
rect 17309 7440 23674 7442
rect 17309 7384 17314 7440
rect 17370 7384 23674 7440
rect 17309 7382 23674 7384
rect 17309 7379 17375 7382
rect 105 7306 171 7309
rect 7005 7306 7071 7309
rect 17769 7306 17835 7309
rect 105 7304 17835 7306
rect 105 7248 110 7304
rect 166 7248 7010 7304
rect 7066 7248 17774 7304
rect 17830 7248 17835 7304
rect 105 7246 17835 7248
rect 105 7243 171 7246
rect 7005 7243 7071 7246
rect 17769 7243 17835 7246
rect 8944 7104 9264 7105
rect 8944 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9264 7104
rect 8944 7039 9264 7040
rect 16944 7104 17264 7105
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 7039 17264 7040
rect 23614 6928 23674 7382
rect 23520 6808 24000 6928
rect 0 6672 480 6792
rect 62 6218 122 6672
rect 4944 6560 5264 6561
rect 4944 6496 4952 6560
rect 5016 6496 5032 6560
rect 5096 6496 5112 6560
rect 5176 6496 5192 6560
rect 5256 6496 5264 6560
rect 4944 6495 5264 6496
rect 12944 6560 13264 6561
rect 12944 6496 12952 6560
rect 13016 6496 13032 6560
rect 13096 6496 13112 6560
rect 13176 6496 13192 6560
rect 13256 6496 13264 6560
rect 12944 6495 13264 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 2865 6218 2931 6221
rect 62 6216 2931 6218
rect 62 6160 2870 6216
rect 2926 6160 2931 6216
rect 62 6158 2931 6160
rect 2865 6155 2931 6158
rect 8944 6016 9264 6017
rect 8944 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9264 6016
rect 8944 5951 9264 5952
rect 16944 6016 17264 6017
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 5951 17264 5952
rect 23520 5584 24000 5704
rect 4944 5472 5264 5473
rect 4944 5408 4952 5472
rect 5016 5408 5032 5472
rect 5096 5408 5112 5472
rect 5176 5408 5192 5472
rect 5256 5408 5264 5472
rect 4944 5407 5264 5408
rect 12944 5472 13264 5473
rect 12944 5408 12952 5472
rect 13016 5408 13032 5472
rect 13096 5408 13112 5472
rect 13176 5408 13192 5472
rect 13256 5408 13264 5472
rect 12944 5407 13264 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 21357 5402 21423 5405
rect 23614 5402 23674 5584
rect 21357 5400 23674 5402
rect 21357 5344 21362 5400
rect 21418 5344 23674 5400
rect 21357 5342 23674 5344
rect 21357 5339 21423 5342
rect 0 5264 480 5296
rect 0 5208 18 5264
rect 74 5208 480 5264
rect 0 5176 480 5208
rect 1945 5130 2011 5133
rect 18505 5130 18571 5133
rect 1945 5128 18571 5130
rect 1945 5072 1950 5128
rect 2006 5072 18510 5128
rect 18566 5072 18571 5128
rect 1945 5070 18571 5072
rect 1945 5067 2011 5070
rect 18505 5067 18571 5070
rect 8944 4928 9264 4929
rect 8944 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9264 4928
rect 8944 4863 9264 4864
rect 16944 4928 17264 4929
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 4863 17264 4864
rect 14089 4722 14155 4725
rect 14917 4722 14983 4725
rect 14089 4720 23674 4722
rect 14089 4664 14094 4720
rect 14150 4664 14922 4720
rect 14978 4664 23674 4720
rect 14089 4662 23674 4664
rect 14089 4659 14155 4662
rect 14917 4659 14983 4662
rect 4944 4384 5264 4385
rect 4944 4320 4952 4384
rect 5016 4320 5032 4384
rect 5096 4320 5112 4384
rect 5176 4320 5192 4384
rect 5256 4320 5264 4384
rect 4944 4319 5264 4320
rect 12944 4384 13264 4385
rect 12944 4320 12952 4384
rect 13016 4320 13032 4384
rect 13096 4320 13112 4384
rect 13176 4320 13192 4384
rect 13256 4320 13264 4384
rect 12944 4319 13264 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 23614 4344 23674 4662
rect 20944 4319 21264 4320
rect 9673 4314 9739 4317
rect 11421 4314 11487 4317
rect 11973 4314 12039 4317
rect 9673 4312 12039 4314
rect 9673 4256 9678 4312
rect 9734 4256 11426 4312
rect 11482 4256 11978 4312
rect 12034 4256 12039 4312
rect 9673 4254 12039 4256
rect 9673 4251 9739 4254
rect 11421 4251 11487 4254
rect 11973 4251 12039 4254
rect 23520 4224 24000 4344
rect 749 4178 815 4181
rect 62 4176 815 4178
rect 62 4120 754 4176
rect 810 4120 815 4176
rect 62 4118 815 4120
rect 62 3800 122 4118
rect 749 4115 815 4118
rect 8944 3840 9264 3841
rect 0 3680 480 3800
rect 8944 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9264 3840
rect 8944 3775 9264 3776
rect 16944 3840 17264 3841
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 3775 17264 3776
rect 3693 3634 3759 3637
rect 9581 3634 9647 3637
rect 13353 3634 13419 3637
rect 3693 3632 13419 3634
rect 3693 3576 3698 3632
rect 3754 3576 9586 3632
rect 9642 3576 13358 3632
rect 13414 3576 13419 3632
rect 3693 3574 13419 3576
rect 3693 3571 3759 3574
rect 9581 3571 9647 3574
rect 13353 3571 13419 3574
rect 14641 3498 14707 3501
rect 14641 3496 23674 3498
rect 14641 3440 14646 3496
rect 14702 3440 23674 3496
rect 14641 3438 23674 3440
rect 14641 3435 14707 3438
rect 4944 3296 5264 3297
rect 4944 3232 4952 3296
rect 5016 3232 5032 3296
rect 5096 3232 5112 3296
rect 5176 3232 5192 3296
rect 5256 3232 5264 3296
rect 4944 3231 5264 3232
rect 12944 3296 13264 3297
rect 12944 3232 12952 3296
rect 13016 3232 13032 3296
rect 13096 3232 13112 3296
rect 13176 3232 13192 3296
rect 13256 3232 13264 3296
rect 12944 3231 13264 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 23614 3120 23674 3438
rect 13077 3090 13143 3093
rect 20621 3090 20687 3093
rect 13077 3088 20687 3090
rect 13077 3032 13082 3088
rect 13138 3032 20626 3088
rect 20682 3032 20687 3088
rect 13077 3030 20687 3032
rect 13077 3027 13143 3030
rect 20621 3027 20687 3030
rect 23520 3000 24000 3120
rect 8944 2752 9264 2753
rect 8944 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9264 2752
rect 8944 2687 9264 2688
rect 16944 2752 17264 2753
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 16944 2687 17264 2688
rect 8109 2410 8175 2413
rect 16389 2410 16455 2413
rect 8109 2408 16455 2410
rect 8109 2352 8114 2408
rect 8170 2352 16394 2408
rect 16450 2352 16455 2408
rect 8109 2350 16455 2352
rect 8109 2347 8175 2350
rect 16389 2347 16455 2350
rect 16614 2348 16620 2412
rect 16684 2410 16690 2412
rect 17125 2410 17191 2413
rect 16684 2408 17191 2410
rect 16684 2352 17130 2408
rect 17186 2352 17191 2408
rect 16684 2350 17191 2352
rect 16684 2348 16690 2350
rect 17125 2347 17191 2350
rect 18229 2410 18295 2413
rect 18229 2408 23674 2410
rect 18229 2352 18234 2408
rect 18290 2352 23674 2408
rect 18229 2350 23674 2352
rect 18229 2347 18295 2350
rect 0 2272 480 2304
rect 0 2216 110 2272
rect 166 2216 480 2272
rect 0 2184 480 2216
rect 4944 2208 5264 2209
rect 4944 2144 4952 2208
rect 5016 2144 5032 2208
rect 5096 2144 5112 2208
rect 5176 2144 5192 2208
rect 5256 2144 5264 2208
rect 4944 2143 5264 2144
rect 12944 2208 13264 2209
rect 12944 2144 12952 2208
rect 13016 2144 13032 2208
rect 13096 2144 13112 2208
rect 13176 2144 13192 2208
rect 13256 2144 13264 2208
rect 12944 2143 13264 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 1209 2002 1275 2005
rect 12433 2002 12499 2005
rect 1209 2000 12499 2002
rect 1209 1944 1214 2000
rect 1270 1944 12438 2000
rect 12494 1944 12499 2000
rect 1209 1942 12499 1944
rect 1209 1939 1275 1942
rect 12433 1939 12499 1942
rect 23614 1896 23674 2350
rect 23520 1776 24000 1896
rect 13445 1322 13511 1325
rect 62 1320 13511 1322
rect 62 1264 13450 1320
rect 13506 1264 13511 1320
rect 62 1262 13511 1264
rect 62 808 122 1262
rect 13445 1259 13511 1262
rect 18597 1186 18663 1189
rect 18597 1184 23674 1186
rect 18597 1128 18602 1184
rect 18658 1128 23674 1184
rect 18597 1126 23674 1128
rect 18597 1123 18663 1126
rect 0 688 480 808
rect 23614 672 23674 1126
rect 23520 552 24000 672
<< via3 >>
rect 4952 21788 5016 21792
rect 4952 21732 4956 21788
rect 4956 21732 5012 21788
rect 5012 21732 5016 21788
rect 4952 21728 5016 21732
rect 5032 21788 5096 21792
rect 5032 21732 5036 21788
rect 5036 21732 5092 21788
rect 5092 21732 5096 21788
rect 5032 21728 5096 21732
rect 5112 21788 5176 21792
rect 5112 21732 5116 21788
rect 5116 21732 5172 21788
rect 5172 21732 5176 21788
rect 5112 21728 5176 21732
rect 5192 21788 5256 21792
rect 5192 21732 5196 21788
rect 5196 21732 5252 21788
rect 5252 21732 5256 21788
rect 5192 21728 5256 21732
rect 12952 21788 13016 21792
rect 12952 21732 12956 21788
rect 12956 21732 13012 21788
rect 13012 21732 13016 21788
rect 12952 21728 13016 21732
rect 13032 21788 13096 21792
rect 13032 21732 13036 21788
rect 13036 21732 13092 21788
rect 13092 21732 13096 21788
rect 13032 21728 13096 21732
rect 13112 21788 13176 21792
rect 13112 21732 13116 21788
rect 13116 21732 13172 21788
rect 13172 21732 13176 21788
rect 13112 21728 13176 21732
rect 13192 21788 13256 21792
rect 13192 21732 13196 21788
rect 13196 21732 13252 21788
rect 13252 21732 13256 21788
rect 13192 21728 13256 21732
rect 20952 21788 21016 21792
rect 20952 21732 20956 21788
rect 20956 21732 21012 21788
rect 21012 21732 21016 21788
rect 20952 21728 21016 21732
rect 21032 21788 21096 21792
rect 21032 21732 21036 21788
rect 21036 21732 21092 21788
rect 21092 21732 21096 21788
rect 21032 21728 21096 21732
rect 21112 21788 21176 21792
rect 21112 21732 21116 21788
rect 21116 21732 21172 21788
rect 21172 21732 21176 21788
rect 21112 21728 21176 21732
rect 21192 21788 21256 21792
rect 21192 21732 21196 21788
rect 21196 21732 21252 21788
rect 21252 21732 21256 21788
rect 21192 21728 21256 21732
rect 8952 21244 9016 21248
rect 8952 21188 8956 21244
rect 8956 21188 9012 21244
rect 9012 21188 9016 21244
rect 8952 21184 9016 21188
rect 9032 21244 9096 21248
rect 9032 21188 9036 21244
rect 9036 21188 9092 21244
rect 9092 21188 9096 21244
rect 9032 21184 9096 21188
rect 9112 21244 9176 21248
rect 9112 21188 9116 21244
rect 9116 21188 9172 21244
rect 9172 21188 9176 21244
rect 9112 21184 9176 21188
rect 9192 21244 9256 21248
rect 9192 21188 9196 21244
rect 9196 21188 9252 21244
rect 9252 21188 9256 21244
rect 9192 21184 9256 21188
rect 16952 21244 17016 21248
rect 16952 21188 16956 21244
rect 16956 21188 17012 21244
rect 17012 21188 17016 21244
rect 16952 21184 17016 21188
rect 17032 21244 17096 21248
rect 17032 21188 17036 21244
rect 17036 21188 17092 21244
rect 17092 21188 17096 21244
rect 17032 21184 17096 21188
rect 17112 21244 17176 21248
rect 17112 21188 17116 21244
rect 17116 21188 17172 21244
rect 17172 21188 17176 21244
rect 17112 21184 17176 21188
rect 17192 21244 17256 21248
rect 17192 21188 17196 21244
rect 17196 21188 17252 21244
rect 17252 21188 17256 21244
rect 17192 21184 17256 21188
rect 4952 20700 5016 20704
rect 4952 20644 4956 20700
rect 4956 20644 5012 20700
rect 5012 20644 5016 20700
rect 4952 20640 5016 20644
rect 5032 20700 5096 20704
rect 5032 20644 5036 20700
rect 5036 20644 5092 20700
rect 5092 20644 5096 20700
rect 5032 20640 5096 20644
rect 5112 20700 5176 20704
rect 5112 20644 5116 20700
rect 5116 20644 5172 20700
rect 5172 20644 5176 20700
rect 5112 20640 5176 20644
rect 5192 20700 5256 20704
rect 5192 20644 5196 20700
rect 5196 20644 5252 20700
rect 5252 20644 5256 20700
rect 5192 20640 5256 20644
rect 12952 20700 13016 20704
rect 12952 20644 12956 20700
rect 12956 20644 13012 20700
rect 13012 20644 13016 20700
rect 12952 20640 13016 20644
rect 13032 20700 13096 20704
rect 13032 20644 13036 20700
rect 13036 20644 13092 20700
rect 13092 20644 13096 20700
rect 13032 20640 13096 20644
rect 13112 20700 13176 20704
rect 13112 20644 13116 20700
rect 13116 20644 13172 20700
rect 13172 20644 13176 20700
rect 13112 20640 13176 20644
rect 13192 20700 13256 20704
rect 13192 20644 13196 20700
rect 13196 20644 13252 20700
rect 13252 20644 13256 20700
rect 13192 20640 13256 20644
rect 20952 20700 21016 20704
rect 20952 20644 20956 20700
rect 20956 20644 21012 20700
rect 21012 20644 21016 20700
rect 20952 20640 21016 20644
rect 21032 20700 21096 20704
rect 21032 20644 21036 20700
rect 21036 20644 21092 20700
rect 21092 20644 21096 20700
rect 21032 20640 21096 20644
rect 21112 20700 21176 20704
rect 21112 20644 21116 20700
rect 21116 20644 21172 20700
rect 21172 20644 21176 20700
rect 21112 20640 21176 20644
rect 21192 20700 21256 20704
rect 21192 20644 21196 20700
rect 21196 20644 21252 20700
rect 21252 20644 21256 20700
rect 21192 20640 21256 20644
rect 8952 20156 9016 20160
rect 8952 20100 8956 20156
rect 8956 20100 9012 20156
rect 9012 20100 9016 20156
rect 8952 20096 9016 20100
rect 9032 20156 9096 20160
rect 9032 20100 9036 20156
rect 9036 20100 9092 20156
rect 9092 20100 9096 20156
rect 9032 20096 9096 20100
rect 9112 20156 9176 20160
rect 9112 20100 9116 20156
rect 9116 20100 9172 20156
rect 9172 20100 9176 20156
rect 9112 20096 9176 20100
rect 9192 20156 9256 20160
rect 9192 20100 9196 20156
rect 9196 20100 9252 20156
rect 9252 20100 9256 20156
rect 9192 20096 9256 20100
rect 16952 20156 17016 20160
rect 16952 20100 16956 20156
rect 16956 20100 17012 20156
rect 17012 20100 17016 20156
rect 16952 20096 17016 20100
rect 17032 20156 17096 20160
rect 17032 20100 17036 20156
rect 17036 20100 17092 20156
rect 17092 20100 17096 20156
rect 17032 20096 17096 20100
rect 17112 20156 17176 20160
rect 17112 20100 17116 20156
rect 17116 20100 17172 20156
rect 17172 20100 17176 20156
rect 17112 20096 17176 20100
rect 17192 20156 17256 20160
rect 17192 20100 17196 20156
rect 17196 20100 17252 20156
rect 17252 20100 17256 20156
rect 17192 20096 17256 20100
rect 4952 19612 5016 19616
rect 4952 19556 4956 19612
rect 4956 19556 5012 19612
rect 5012 19556 5016 19612
rect 4952 19552 5016 19556
rect 5032 19612 5096 19616
rect 5032 19556 5036 19612
rect 5036 19556 5092 19612
rect 5092 19556 5096 19612
rect 5032 19552 5096 19556
rect 5112 19612 5176 19616
rect 5112 19556 5116 19612
rect 5116 19556 5172 19612
rect 5172 19556 5176 19612
rect 5112 19552 5176 19556
rect 5192 19612 5256 19616
rect 5192 19556 5196 19612
rect 5196 19556 5252 19612
rect 5252 19556 5256 19612
rect 5192 19552 5256 19556
rect 12952 19612 13016 19616
rect 12952 19556 12956 19612
rect 12956 19556 13012 19612
rect 13012 19556 13016 19612
rect 12952 19552 13016 19556
rect 13032 19612 13096 19616
rect 13032 19556 13036 19612
rect 13036 19556 13092 19612
rect 13092 19556 13096 19612
rect 13032 19552 13096 19556
rect 13112 19612 13176 19616
rect 13112 19556 13116 19612
rect 13116 19556 13172 19612
rect 13172 19556 13176 19612
rect 13112 19552 13176 19556
rect 13192 19612 13256 19616
rect 13192 19556 13196 19612
rect 13196 19556 13252 19612
rect 13252 19556 13256 19612
rect 13192 19552 13256 19556
rect 20952 19612 21016 19616
rect 20952 19556 20956 19612
rect 20956 19556 21012 19612
rect 21012 19556 21016 19612
rect 20952 19552 21016 19556
rect 21032 19612 21096 19616
rect 21032 19556 21036 19612
rect 21036 19556 21092 19612
rect 21092 19556 21096 19612
rect 21032 19552 21096 19556
rect 21112 19612 21176 19616
rect 21112 19556 21116 19612
rect 21116 19556 21172 19612
rect 21172 19556 21176 19612
rect 21112 19552 21176 19556
rect 21192 19612 21256 19616
rect 21192 19556 21196 19612
rect 21196 19556 21252 19612
rect 21252 19556 21256 19612
rect 21192 19552 21256 19556
rect 8952 19068 9016 19072
rect 8952 19012 8956 19068
rect 8956 19012 9012 19068
rect 9012 19012 9016 19068
rect 8952 19008 9016 19012
rect 9032 19068 9096 19072
rect 9032 19012 9036 19068
rect 9036 19012 9092 19068
rect 9092 19012 9096 19068
rect 9032 19008 9096 19012
rect 9112 19068 9176 19072
rect 9112 19012 9116 19068
rect 9116 19012 9172 19068
rect 9172 19012 9176 19068
rect 9112 19008 9176 19012
rect 9192 19068 9256 19072
rect 9192 19012 9196 19068
rect 9196 19012 9252 19068
rect 9252 19012 9256 19068
rect 9192 19008 9256 19012
rect 16952 19068 17016 19072
rect 16952 19012 16956 19068
rect 16956 19012 17012 19068
rect 17012 19012 17016 19068
rect 16952 19008 17016 19012
rect 17032 19068 17096 19072
rect 17032 19012 17036 19068
rect 17036 19012 17092 19068
rect 17092 19012 17096 19068
rect 17032 19008 17096 19012
rect 17112 19068 17176 19072
rect 17112 19012 17116 19068
rect 17116 19012 17172 19068
rect 17172 19012 17176 19068
rect 17112 19008 17176 19012
rect 17192 19068 17256 19072
rect 17192 19012 17196 19068
rect 17196 19012 17252 19068
rect 17252 19012 17256 19068
rect 17192 19008 17256 19012
rect 4952 18524 5016 18528
rect 4952 18468 4956 18524
rect 4956 18468 5012 18524
rect 5012 18468 5016 18524
rect 4952 18464 5016 18468
rect 5032 18524 5096 18528
rect 5032 18468 5036 18524
rect 5036 18468 5092 18524
rect 5092 18468 5096 18524
rect 5032 18464 5096 18468
rect 5112 18524 5176 18528
rect 5112 18468 5116 18524
rect 5116 18468 5172 18524
rect 5172 18468 5176 18524
rect 5112 18464 5176 18468
rect 5192 18524 5256 18528
rect 5192 18468 5196 18524
rect 5196 18468 5252 18524
rect 5252 18468 5256 18524
rect 5192 18464 5256 18468
rect 12952 18524 13016 18528
rect 12952 18468 12956 18524
rect 12956 18468 13012 18524
rect 13012 18468 13016 18524
rect 12952 18464 13016 18468
rect 13032 18524 13096 18528
rect 13032 18468 13036 18524
rect 13036 18468 13092 18524
rect 13092 18468 13096 18524
rect 13032 18464 13096 18468
rect 13112 18524 13176 18528
rect 13112 18468 13116 18524
rect 13116 18468 13172 18524
rect 13172 18468 13176 18524
rect 13112 18464 13176 18468
rect 13192 18524 13256 18528
rect 13192 18468 13196 18524
rect 13196 18468 13252 18524
rect 13252 18468 13256 18524
rect 13192 18464 13256 18468
rect 20952 18524 21016 18528
rect 20952 18468 20956 18524
rect 20956 18468 21012 18524
rect 21012 18468 21016 18524
rect 20952 18464 21016 18468
rect 21032 18524 21096 18528
rect 21032 18468 21036 18524
rect 21036 18468 21092 18524
rect 21092 18468 21096 18524
rect 21032 18464 21096 18468
rect 21112 18524 21176 18528
rect 21112 18468 21116 18524
rect 21116 18468 21172 18524
rect 21172 18468 21176 18524
rect 21112 18464 21176 18468
rect 21192 18524 21256 18528
rect 21192 18468 21196 18524
rect 21196 18468 21252 18524
rect 21252 18468 21256 18524
rect 21192 18464 21256 18468
rect 8952 17980 9016 17984
rect 8952 17924 8956 17980
rect 8956 17924 9012 17980
rect 9012 17924 9016 17980
rect 8952 17920 9016 17924
rect 9032 17980 9096 17984
rect 9032 17924 9036 17980
rect 9036 17924 9092 17980
rect 9092 17924 9096 17980
rect 9032 17920 9096 17924
rect 9112 17980 9176 17984
rect 9112 17924 9116 17980
rect 9116 17924 9172 17980
rect 9172 17924 9176 17980
rect 9112 17920 9176 17924
rect 9192 17980 9256 17984
rect 9192 17924 9196 17980
rect 9196 17924 9252 17980
rect 9252 17924 9256 17980
rect 9192 17920 9256 17924
rect 16952 17980 17016 17984
rect 16952 17924 16956 17980
rect 16956 17924 17012 17980
rect 17012 17924 17016 17980
rect 16952 17920 17016 17924
rect 17032 17980 17096 17984
rect 17032 17924 17036 17980
rect 17036 17924 17092 17980
rect 17092 17924 17096 17980
rect 17032 17920 17096 17924
rect 17112 17980 17176 17984
rect 17112 17924 17116 17980
rect 17116 17924 17172 17980
rect 17172 17924 17176 17980
rect 17112 17920 17176 17924
rect 17192 17980 17256 17984
rect 17192 17924 17196 17980
rect 17196 17924 17252 17980
rect 17252 17924 17256 17980
rect 17192 17920 17256 17924
rect 4952 17436 5016 17440
rect 4952 17380 4956 17436
rect 4956 17380 5012 17436
rect 5012 17380 5016 17436
rect 4952 17376 5016 17380
rect 5032 17436 5096 17440
rect 5032 17380 5036 17436
rect 5036 17380 5092 17436
rect 5092 17380 5096 17436
rect 5032 17376 5096 17380
rect 5112 17436 5176 17440
rect 5112 17380 5116 17436
rect 5116 17380 5172 17436
rect 5172 17380 5176 17436
rect 5112 17376 5176 17380
rect 5192 17436 5256 17440
rect 5192 17380 5196 17436
rect 5196 17380 5252 17436
rect 5252 17380 5256 17436
rect 5192 17376 5256 17380
rect 12952 17436 13016 17440
rect 12952 17380 12956 17436
rect 12956 17380 13012 17436
rect 13012 17380 13016 17436
rect 12952 17376 13016 17380
rect 13032 17436 13096 17440
rect 13032 17380 13036 17436
rect 13036 17380 13092 17436
rect 13092 17380 13096 17436
rect 13032 17376 13096 17380
rect 13112 17436 13176 17440
rect 13112 17380 13116 17436
rect 13116 17380 13172 17436
rect 13172 17380 13176 17436
rect 13112 17376 13176 17380
rect 13192 17436 13256 17440
rect 13192 17380 13196 17436
rect 13196 17380 13252 17436
rect 13252 17380 13256 17436
rect 13192 17376 13256 17380
rect 20952 17436 21016 17440
rect 20952 17380 20956 17436
rect 20956 17380 21012 17436
rect 21012 17380 21016 17436
rect 20952 17376 21016 17380
rect 21032 17436 21096 17440
rect 21032 17380 21036 17436
rect 21036 17380 21092 17436
rect 21092 17380 21096 17436
rect 21032 17376 21096 17380
rect 21112 17436 21176 17440
rect 21112 17380 21116 17436
rect 21116 17380 21172 17436
rect 21172 17380 21176 17436
rect 21112 17376 21176 17380
rect 21192 17436 21256 17440
rect 21192 17380 21196 17436
rect 21196 17380 21252 17436
rect 21252 17380 21256 17436
rect 21192 17376 21256 17380
rect 8952 16892 9016 16896
rect 8952 16836 8956 16892
rect 8956 16836 9012 16892
rect 9012 16836 9016 16892
rect 8952 16832 9016 16836
rect 9032 16892 9096 16896
rect 9032 16836 9036 16892
rect 9036 16836 9092 16892
rect 9092 16836 9096 16892
rect 9032 16832 9096 16836
rect 9112 16892 9176 16896
rect 9112 16836 9116 16892
rect 9116 16836 9172 16892
rect 9172 16836 9176 16892
rect 9112 16832 9176 16836
rect 9192 16892 9256 16896
rect 9192 16836 9196 16892
rect 9196 16836 9252 16892
rect 9252 16836 9256 16892
rect 9192 16832 9256 16836
rect 16952 16892 17016 16896
rect 16952 16836 16956 16892
rect 16956 16836 17012 16892
rect 17012 16836 17016 16892
rect 16952 16832 17016 16836
rect 17032 16892 17096 16896
rect 17032 16836 17036 16892
rect 17036 16836 17092 16892
rect 17092 16836 17096 16892
rect 17032 16832 17096 16836
rect 17112 16892 17176 16896
rect 17112 16836 17116 16892
rect 17116 16836 17172 16892
rect 17172 16836 17176 16892
rect 17112 16832 17176 16836
rect 17192 16892 17256 16896
rect 17192 16836 17196 16892
rect 17196 16836 17252 16892
rect 17252 16836 17256 16892
rect 17192 16832 17256 16836
rect 4952 16348 5016 16352
rect 4952 16292 4956 16348
rect 4956 16292 5012 16348
rect 5012 16292 5016 16348
rect 4952 16288 5016 16292
rect 5032 16348 5096 16352
rect 5032 16292 5036 16348
rect 5036 16292 5092 16348
rect 5092 16292 5096 16348
rect 5032 16288 5096 16292
rect 5112 16348 5176 16352
rect 5112 16292 5116 16348
rect 5116 16292 5172 16348
rect 5172 16292 5176 16348
rect 5112 16288 5176 16292
rect 5192 16348 5256 16352
rect 5192 16292 5196 16348
rect 5196 16292 5252 16348
rect 5252 16292 5256 16348
rect 5192 16288 5256 16292
rect 12952 16348 13016 16352
rect 12952 16292 12956 16348
rect 12956 16292 13012 16348
rect 13012 16292 13016 16348
rect 12952 16288 13016 16292
rect 13032 16348 13096 16352
rect 13032 16292 13036 16348
rect 13036 16292 13092 16348
rect 13092 16292 13096 16348
rect 13032 16288 13096 16292
rect 13112 16348 13176 16352
rect 13112 16292 13116 16348
rect 13116 16292 13172 16348
rect 13172 16292 13176 16348
rect 13112 16288 13176 16292
rect 13192 16348 13256 16352
rect 13192 16292 13196 16348
rect 13196 16292 13252 16348
rect 13252 16292 13256 16348
rect 13192 16288 13256 16292
rect 20952 16348 21016 16352
rect 20952 16292 20956 16348
rect 20956 16292 21012 16348
rect 21012 16292 21016 16348
rect 20952 16288 21016 16292
rect 21032 16348 21096 16352
rect 21032 16292 21036 16348
rect 21036 16292 21092 16348
rect 21092 16292 21096 16348
rect 21032 16288 21096 16292
rect 21112 16348 21176 16352
rect 21112 16292 21116 16348
rect 21116 16292 21172 16348
rect 21172 16292 21176 16348
rect 21112 16288 21176 16292
rect 21192 16348 21256 16352
rect 21192 16292 21196 16348
rect 21196 16292 21252 16348
rect 21252 16292 21256 16348
rect 21192 16288 21256 16292
rect 8952 15804 9016 15808
rect 8952 15748 8956 15804
rect 8956 15748 9012 15804
rect 9012 15748 9016 15804
rect 8952 15744 9016 15748
rect 9032 15804 9096 15808
rect 9032 15748 9036 15804
rect 9036 15748 9092 15804
rect 9092 15748 9096 15804
rect 9032 15744 9096 15748
rect 9112 15804 9176 15808
rect 9112 15748 9116 15804
rect 9116 15748 9172 15804
rect 9172 15748 9176 15804
rect 9112 15744 9176 15748
rect 9192 15804 9256 15808
rect 9192 15748 9196 15804
rect 9196 15748 9252 15804
rect 9252 15748 9256 15804
rect 9192 15744 9256 15748
rect 16952 15804 17016 15808
rect 16952 15748 16956 15804
rect 16956 15748 17012 15804
rect 17012 15748 17016 15804
rect 16952 15744 17016 15748
rect 17032 15804 17096 15808
rect 17032 15748 17036 15804
rect 17036 15748 17092 15804
rect 17092 15748 17096 15804
rect 17032 15744 17096 15748
rect 17112 15804 17176 15808
rect 17112 15748 17116 15804
rect 17116 15748 17172 15804
rect 17172 15748 17176 15804
rect 17112 15744 17176 15748
rect 17192 15804 17256 15808
rect 17192 15748 17196 15804
rect 17196 15748 17252 15804
rect 17252 15748 17256 15804
rect 17192 15744 17256 15748
rect 4952 15260 5016 15264
rect 4952 15204 4956 15260
rect 4956 15204 5012 15260
rect 5012 15204 5016 15260
rect 4952 15200 5016 15204
rect 5032 15260 5096 15264
rect 5032 15204 5036 15260
rect 5036 15204 5092 15260
rect 5092 15204 5096 15260
rect 5032 15200 5096 15204
rect 5112 15260 5176 15264
rect 5112 15204 5116 15260
rect 5116 15204 5172 15260
rect 5172 15204 5176 15260
rect 5112 15200 5176 15204
rect 5192 15260 5256 15264
rect 5192 15204 5196 15260
rect 5196 15204 5252 15260
rect 5252 15204 5256 15260
rect 5192 15200 5256 15204
rect 12952 15260 13016 15264
rect 12952 15204 12956 15260
rect 12956 15204 13012 15260
rect 13012 15204 13016 15260
rect 12952 15200 13016 15204
rect 13032 15260 13096 15264
rect 13032 15204 13036 15260
rect 13036 15204 13092 15260
rect 13092 15204 13096 15260
rect 13032 15200 13096 15204
rect 13112 15260 13176 15264
rect 13112 15204 13116 15260
rect 13116 15204 13172 15260
rect 13172 15204 13176 15260
rect 13112 15200 13176 15204
rect 13192 15260 13256 15264
rect 13192 15204 13196 15260
rect 13196 15204 13252 15260
rect 13252 15204 13256 15260
rect 13192 15200 13256 15204
rect 20952 15260 21016 15264
rect 20952 15204 20956 15260
rect 20956 15204 21012 15260
rect 21012 15204 21016 15260
rect 20952 15200 21016 15204
rect 21032 15260 21096 15264
rect 21032 15204 21036 15260
rect 21036 15204 21092 15260
rect 21092 15204 21096 15260
rect 21032 15200 21096 15204
rect 21112 15260 21176 15264
rect 21112 15204 21116 15260
rect 21116 15204 21172 15260
rect 21172 15204 21176 15260
rect 21112 15200 21176 15204
rect 21192 15260 21256 15264
rect 21192 15204 21196 15260
rect 21196 15204 21252 15260
rect 21252 15204 21256 15260
rect 21192 15200 21256 15204
rect 8952 14716 9016 14720
rect 8952 14660 8956 14716
rect 8956 14660 9012 14716
rect 9012 14660 9016 14716
rect 8952 14656 9016 14660
rect 9032 14716 9096 14720
rect 9032 14660 9036 14716
rect 9036 14660 9092 14716
rect 9092 14660 9096 14716
rect 9032 14656 9096 14660
rect 9112 14716 9176 14720
rect 9112 14660 9116 14716
rect 9116 14660 9172 14716
rect 9172 14660 9176 14716
rect 9112 14656 9176 14660
rect 9192 14716 9256 14720
rect 9192 14660 9196 14716
rect 9196 14660 9252 14716
rect 9252 14660 9256 14716
rect 9192 14656 9256 14660
rect 16952 14716 17016 14720
rect 16952 14660 16956 14716
rect 16956 14660 17012 14716
rect 17012 14660 17016 14716
rect 16952 14656 17016 14660
rect 17032 14716 17096 14720
rect 17032 14660 17036 14716
rect 17036 14660 17092 14716
rect 17092 14660 17096 14716
rect 17032 14656 17096 14660
rect 17112 14716 17176 14720
rect 17112 14660 17116 14716
rect 17116 14660 17172 14716
rect 17172 14660 17176 14716
rect 17112 14656 17176 14660
rect 17192 14716 17256 14720
rect 17192 14660 17196 14716
rect 17196 14660 17252 14716
rect 17252 14660 17256 14716
rect 17192 14656 17256 14660
rect 4952 14172 5016 14176
rect 4952 14116 4956 14172
rect 4956 14116 5012 14172
rect 5012 14116 5016 14172
rect 4952 14112 5016 14116
rect 5032 14172 5096 14176
rect 5032 14116 5036 14172
rect 5036 14116 5092 14172
rect 5092 14116 5096 14172
rect 5032 14112 5096 14116
rect 5112 14172 5176 14176
rect 5112 14116 5116 14172
rect 5116 14116 5172 14172
rect 5172 14116 5176 14172
rect 5112 14112 5176 14116
rect 5192 14172 5256 14176
rect 5192 14116 5196 14172
rect 5196 14116 5252 14172
rect 5252 14116 5256 14172
rect 5192 14112 5256 14116
rect 12952 14172 13016 14176
rect 12952 14116 12956 14172
rect 12956 14116 13012 14172
rect 13012 14116 13016 14172
rect 12952 14112 13016 14116
rect 13032 14172 13096 14176
rect 13032 14116 13036 14172
rect 13036 14116 13092 14172
rect 13092 14116 13096 14172
rect 13032 14112 13096 14116
rect 13112 14172 13176 14176
rect 13112 14116 13116 14172
rect 13116 14116 13172 14172
rect 13172 14116 13176 14172
rect 13112 14112 13176 14116
rect 13192 14172 13256 14176
rect 13192 14116 13196 14172
rect 13196 14116 13252 14172
rect 13252 14116 13256 14172
rect 13192 14112 13256 14116
rect 20952 14172 21016 14176
rect 20952 14116 20956 14172
rect 20956 14116 21012 14172
rect 21012 14116 21016 14172
rect 20952 14112 21016 14116
rect 21032 14172 21096 14176
rect 21032 14116 21036 14172
rect 21036 14116 21092 14172
rect 21092 14116 21096 14172
rect 21032 14112 21096 14116
rect 21112 14172 21176 14176
rect 21112 14116 21116 14172
rect 21116 14116 21172 14172
rect 21172 14116 21176 14172
rect 21112 14112 21176 14116
rect 21192 14172 21256 14176
rect 21192 14116 21196 14172
rect 21196 14116 21252 14172
rect 21252 14116 21256 14172
rect 21192 14112 21256 14116
rect 8952 13628 9016 13632
rect 8952 13572 8956 13628
rect 8956 13572 9012 13628
rect 9012 13572 9016 13628
rect 8952 13568 9016 13572
rect 9032 13628 9096 13632
rect 9032 13572 9036 13628
rect 9036 13572 9092 13628
rect 9092 13572 9096 13628
rect 9032 13568 9096 13572
rect 9112 13628 9176 13632
rect 9112 13572 9116 13628
rect 9116 13572 9172 13628
rect 9172 13572 9176 13628
rect 9112 13568 9176 13572
rect 9192 13628 9256 13632
rect 9192 13572 9196 13628
rect 9196 13572 9252 13628
rect 9252 13572 9256 13628
rect 9192 13568 9256 13572
rect 16952 13628 17016 13632
rect 16952 13572 16956 13628
rect 16956 13572 17012 13628
rect 17012 13572 17016 13628
rect 16952 13568 17016 13572
rect 17032 13628 17096 13632
rect 17032 13572 17036 13628
rect 17036 13572 17092 13628
rect 17092 13572 17096 13628
rect 17032 13568 17096 13572
rect 17112 13628 17176 13632
rect 17112 13572 17116 13628
rect 17116 13572 17172 13628
rect 17172 13572 17176 13628
rect 17112 13568 17176 13572
rect 17192 13628 17256 13632
rect 17192 13572 17196 13628
rect 17196 13572 17252 13628
rect 17252 13572 17256 13628
rect 17192 13568 17256 13572
rect 4952 13084 5016 13088
rect 4952 13028 4956 13084
rect 4956 13028 5012 13084
rect 5012 13028 5016 13084
rect 4952 13024 5016 13028
rect 5032 13084 5096 13088
rect 5032 13028 5036 13084
rect 5036 13028 5092 13084
rect 5092 13028 5096 13084
rect 5032 13024 5096 13028
rect 5112 13084 5176 13088
rect 5112 13028 5116 13084
rect 5116 13028 5172 13084
rect 5172 13028 5176 13084
rect 5112 13024 5176 13028
rect 5192 13084 5256 13088
rect 5192 13028 5196 13084
rect 5196 13028 5252 13084
rect 5252 13028 5256 13084
rect 5192 13024 5256 13028
rect 12952 13084 13016 13088
rect 12952 13028 12956 13084
rect 12956 13028 13012 13084
rect 13012 13028 13016 13084
rect 12952 13024 13016 13028
rect 13032 13084 13096 13088
rect 13032 13028 13036 13084
rect 13036 13028 13092 13084
rect 13092 13028 13096 13084
rect 13032 13024 13096 13028
rect 13112 13084 13176 13088
rect 13112 13028 13116 13084
rect 13116 13028 13172 13084
rect 13172 13028 13176 13084
rect 13112 13024 13176 13028
rect 13192 13084 13256 13088
rect 13192 13028 13196 13084
rect 13196 13028 13252 13084
rect 13252 13028 13256 13084
rect 13192 13024 13256 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 60 12684 124 12748
rect 8952 12540 9016 12544
rect 8952 12484 8956 12540
rect 8956 12484 9012 12540
rect 9012 12484 9016 12540
rect 8952 12480 9016 12484
rect 9032 12540 9096 12544
rect 9032 12484 9036 12540
rect 9036 12484 9092 12540
rect 9092 12484 9096 12540
rect 9032 12480 9096 12484
rect 9112 12540 9176 12544
rect 9112 12484 9116 12540
rect 9116 12484 9172 12540
rect 9172 12484 9176 12540
rect 9112 12480 9176 12484
rect 9192 12540 9256 12544
rect 9192 12484 9196 12540
rect 9196 12484 9252 12540
rect 9252 12484 9256 12540
rect 9192 12480 9256 12484
rect 16952 12540 17016 12544
rect 16952 12484 16956 12540
rect 16956 12484 17012 12540
rect 17012 12484 17016 12540
rect 16952 12480 17016 12484
rect 17032 12540 17096 12544
rect 17032 12484 17036 12540
rect 17036 12484 17092 12540
rect 17092 12484 17096 12540
rect 17032 12480 17096 12484
rect 17112 12540 17176 12544
rect 17112 12484 17116 12540
rect 17116 12484 17172 12540
rect 17172 12484 17176 12540
rect 17112 12480 17176 12484
rect 17192 12540 17256 12544
rect 17192 12484 17196 12540
rect 17196 12484 17252 12540
rect 17252 12484 17256 12540
rect 17192 12480 17256 12484
rect 60 12276 124 12340
rect 4952 11996 5016 12000
rect 4952 11940 4956 11996
rect 4956 11940 5012 11996
rect 5012 11940 5016 11996
rect 4952 11936 5016 11940
rect 5032 11996 5096 12000
rect 5032 11940 5036 11996
rect 5036 11940 5092 11996
rect 5092 11940 5096 11996
rect 5032 11936 5096 11940
rect 5112 11996 5176 12000
rect 5112 11940 5116 11996
rect 5116 11940 5172 11996
rect 5172 11940 5176 11996
rect 5112 11936 5176 11940
rect 5192 11996 5256 12000
rect 5192 11940 5196 11996
rect 5196 11940 5252 11996
rect 5252 11940 5256 11996
rect 5192 11936 5256 11940
rect 12952 11996 13016 12000
rect 12952 11940 12956 11996
rect 12956 11940 13012 11996
rect 13012 11940 13016 11996
rect 12952 11936 13016 11940
rect 13032 11996 13096 12000
rect 13032 11940 13036 11996
rect 13036 11940 13092 11996
rect 13092 11940 13096 11996
rect 13032 11936 13096 11940
rect 13112 11996 13176 12000
rect 13112 11940 13116 11996
rect 13116 11940 13172 11996
rect 13172 11940 13176 11996
rect 13112 11936 13176 11940
rect 13192 11996 13256 12000
rect 13192 11940 13196 11996
rect 13196 11940 13252 11996
rect 13252 11940 13256 11996
rect 13192 11936 13256 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 8952 11452 9016 11456
rect 8952 11396 8956 11452
rect 8956 11396 9012 11452
rect 9012 11396 9016 11452
rect 8952 11392 9016 11396
rect 9032 11452 9096 11456
rect 9032 11396 9036 11452
rect 9036 11396 9092 11452
rect 9092 11396 9096 11452
rect 9032 11392 9096 11396
rect 9112 11452 9176 11456
rect 9112 11396 9116 11452
rect 9116 11396 9172 11452
rect 9172 11396 9176 11452
rect 9112 11392 9176 11396
rect 9192 11452 9256 11456
rect 9192 11396 9196 11452
rect 9196 11396 9252 11452
rect 9252 11396 9256 11452
rect 9192 11392 9256 11396
rect 16952 11452 17016 11456
rect 16952 11396 16956 11452
rect 16956 11396 17012 11452
rect 17012 11396 17016 11452
rect 16952 11392 17016 11396
rect 17032 11452 17096 11456
rect 17032 11396 17036 11452
rect 17036 11396 17092 11452
rect 17092 11396 17096 11452
rect 17032 11392 17096 11396
rect 17112 11452 17176 11456
rect 17112 11396 17116 11452
rect 17116 11396 17172 11452
rect 17172 11396 17176 11452
rect 17112 11392 17176 11396
rect 17192 11452 17256 11456
rect 17192 11396 17196 11452
rect 17196 11396 17252 11452
rect 17252 11396 17256 11452
rect 17192 11392 17256 11396
rect 4952 10908 5016 10912
rect 4952 10852 4956 10908
rect 4956 10852 5012 10908
rect 5012 10852 5016 10908
rect 4952 10848 5016 10852
rect 5032 10908 5096 10912
rect 5032 10852 5036 10908
rect 5036 10852 5092 10908
rect 5092 10852 5096 10908
rect 5032 10848 5096 10852
rect 5112 10908 5176 10912
rect 5112 10852 5116 10908
rect 5116 10852 5172 10908
rect 5172 10852 5176 10908
rect 5112 10848 5176 10852
rect 5192 10908 5256 10912
rect 5192 10852 5196 10908
rect 5196 10852 5252 10908
rect 5252 10852 5256 10908
rect 5192 10848 5256 10852
rect 12952 10908 13016 10912
rect 12952 10852 12956 10908
rect 12956 10852 13012 10908
rect 13012 10852 13016 10908
rect 12952 10848 13016 10852
rect 13032 10908 13096 10912
rect 13032 10852 13036 10908
rect 13036 10852 13092 10908
rect 13092 10852 13096 10908
rect 13032 10848 13096 10852
rect 13112 10908 13176 10912
rect 13112 10852 13116 10908
rect 13116 10852 13172 10908
rect 13172 10852 13176 10908
rect 13112 10848 13176 10852
rect 13192 10908 13256 10912
rect 13192 10852 13196 10908
rect 13196 10852 13252 10908
rect 13252 10852 13256 10908
rect 13192 10848 13256 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 8952 10364 9016 10368
rect 8952 10308 8956 10364
rect 8956 10308 9012 10364
rect 9012 10308 9016 10364
rect 8952 10304 9016 10308
rect 9032 10364 9096 10368
rect 9032 10308 9036 10364
rect 9036 10308 9092 10364
rect 9092 10308 9096 10364
rect 9032 10304 9096 10308
rect 9112 10364 9176 10368
rect 9112 10308 9116 10364
rect 9116 10308 9172 10364
rect 9172 10308 9176 10364
rect 9112 10304 9176 10308
rect 9192 10364 9256 10368
rect 9192 10308 9196 10364
rect 9196 10308 9252 10364
rect 9252 10308 9256 10364
rect 9192 10304 9256 10308
rect 16952 10364 17016 10368
rect 16952 10308 16956 10364
rect 16956 10308 17012 10364
rect 17012 10308 17016 10364
rect 16952 10304 17016 10308
rect 17032 10364 17096 10368
rect 17032 10308 17036 10364
rect 17036 10308 17092 10364
rect 17092 10308 17096 10364
rect 17032 10304 17096 10308
rect 17112 10364 17176 10368
rect 17112 10308 17116 10364
rect 17116 10308 17172 10364
rect 17172 10308 17176 10364
rect 17112 10304 17176 10308
rect 17192 10364 17256 10368
rect 17192 10308 17196 10364
rect 17196 10308 17252 10364
rect 17252 10308 17256 10364
rect 17192 10304 17256 10308
rect 60 9964 124 10028
rect 4952 9820 5016 9824
rect 4952 9764 4956 9820
rect 4956 9764 5012 9820
rect 5012 9764 5016 9820
rect 4952 9760 5016 9764
rect 5032 9820 5096 9824
rect 5032 9764 5036 9820
rect 5036 9764 5092 9820
rect 5092 9764 5096 9820
rect 5032 9760 5096 9764
rect 5112 9820 5176 9824
rect 5112 9764 5116 9820
rect 5116 9764 5172 9820
rect 5172 9764 5176 9820
rect 5112 9760 5176 9764
rect 5192 9820 5256 9824
rect 5192 9764 5196 9820
rect 5196 9764 5252 9820
rect 5252 9764 5256 9820
rect 5192 9760 5256 9764
rect 12952 9820 13016 9824
rect 12952 9764 12956 9820
rect 12956 9764 13012 9820
rect 13012 9764 13016 9820
rect 12952 9760 13016 9764
rect 13032 9820 13096 9824
rect 13032 9764 13036 9820
rect 13036 9764 13092 9820
rect 13092 9764 13096 9820
rect 13032 9760 13096 9764
rect 13112 9820 13176 9824
rect 13112 9764 13116 9820
rect 13116 9764 13172 9820
rect 13172 9764 13176 9820
rect 13112 9760 13176 9764
rect 13192 9820 13256 9824
rect 13192 9764 13196 9820
rect 13196 9764 13252 9820
rect 13252 9764 13256 9820
rect 13192 9760 13256 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 60 9692 124 9756
rect 8952 9276 9016 9280
rect 8952 9220 8956 9276
rect 8956 9220 9012 9276
rect 9012 9220 9016 9276
rect 8952 9216 9016 9220
rect 9032 9276 9096 9280
rect 9032 9220 9036 9276
rect 9036 9220 9092 9276
rect 9092 9220 9096 9276
rect 9032 9216 9096 9220
rect 9112 9276 9176 9280
rect 9112 9220 9116 9276
rect 9116 9220 9172 9276
rect 9172 9220 9176 9276
rect 9112 9216 9176 9220
rect 9192 9276 9256 9280
rect 9192 9220 9196 9276
rect 9196 9220 9252 9276
rect 9252 9220 9256 9276
rect 9192 9216 9256 9220
rect 16952 9276 17016 9280
rect 16952 9220 16956 9276
rect 16956 9220 17012 9276
rect 17012 9220 17016 9276
rect 16952 9216 17016 9220
rect 17032 9276 17096 9280
rect 17032 9220 17036 9276
rect 17036 9220 17092 9276
rect 17092 9220 17096 9276
rect 17032 9216 17096 9220
rect 17112 9276 17176 9280
rect 17112 9220 17116 9276
rect 17116 9220 17172 9276
rect 17172 9220 17176 9276
rect 17112 9216 17176 9220
rect 17192 9276 17256 9280
rect 17192 9220 17196 9276
rect 17196 9220 17252 9276
rect 17252 9220 17256 9276
rect 17192 9216 17256 9220
rect 4952 8732 5016 8736
rect 4952 8676 4956 8732
rect 4956 8676 5012 8732
rect 5012 8676 5016 8732
rect 4952 8672 5016 8676
rect 5032 8732 5096 8736
rect 5032 8676 5036 8732
rect 5036 8676 5092 8732
rect 5092 8676 5096 8732
rect 5032 8672 5096 8676
rect 5112 8732 5176 8736
rect 5112 8676 5116 8732
rect 5116 8676 5172 8732
rect 5172 8676 5176 8732
rect 5112 8672 5176 8676
rect 5192 8732 5256 8736
rect 5192 8676 5196 8732
rect 5196 8676 5252 8732
rect 5252 8676 5256 8732
rect 5192 8672 5256 8676
rect 12952 8732 13016 8736
rect 12952 8676 12956 8732
rect 12956 8676 13012 8732
rect 13012 8676 13016 8732
rect 12952 8672 13016 8676
rect 13032 8732 13096 8736
rect 13032 8676 13036 8732
rect 13036 8676 13092 8732
rect 13092 8676 13096 8732
rect 13032 8672 13096 8676
rect 13112 8732 13176 8736
rect 13112 8676 13116 8732
rect 13116 8676 13172 8732
rect 13172 8676 13176 8732
rect 13112 8672 13176 8676
rect 13192 8732 13256 8736
rect 13192 8676 13196 8732
rect 13196 8676 13252 8732
rect 13252 8676 13256 8732
rect 13192 8672 13256 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 7604 8196 7668 8260
rect 8952 8188 9016 8192
rect 8952 8132 8956 8188
rect 8956 8132 9012 8188
rect 9012 8132 9016 8188
rect 8952 8128 9016 8132
rect 9032 8188 9096 8192
rect 9032 8132 9036 8188
rect 9036 8132 9092 8188
rect 9092 8132 9096 8188
rect 9032 8128 9096 8132
rect 9112 8188 9176 8192
rect 9112 8132 9116 8188
rect 9116 8132 9172 8188
rect 9172 8132 9176 8188
rect 9112 8128 9176 8132
rect 9192 8188 9256 8192
rect 9192 8132 9196 8188
rect 9196 8132 9252 8188
rect 9252 8132 9256 8188
rect 9192 8128 9256 8132
rect 16952 8188 17016 8192
rect 16952 8132 16956 8188
rect 16956 8132 17012 8188
rect 17012 8132 17016 8188
rect 16952 8128 17016 8132
rect 17032 8188 17096 8192
rect 17032 8132 17036 8188
rect 17036 8132 17092 8188
rect 17092 8132 17096 8188
rect 17032 8128 17096 8132
rect 17112 8188 17176 8192
rect 17112 8132 17116 8188
rect 17116 8132 17172 8188
rect 17172 8132 17176 8188
rect 17112 8128 17176 8132
rect 17192 8188 17256 8192
rect 17192 8132 17196 8188
rect 17196 8132 17252 8188
rect 17252 8132 17256 8188
rect 17192 8128 17256 8132
rect 23612 8060 23676 8124
rect 23612 7788 23676 7852
rect 4952 7644 5016 7648
rect 4952 7588 4956 7644
rect 4956 7588 5012 7644
rect 5012 7588 5016 7644
rect 4952 7584 5016 7588
rect 5032 7644 5096 7648
rect 5032 7588 5036 7644
rect 5036 7588 5092 7644
rect 5092 7588 5096 7644
rect 5032 7584 5096 7588
rect 5112 7644 5176 7648
rect 5112 7588 5116 7644
rect 5116 7588 5172 7644
rect 5172 7588 5176 7644
rect 5112 7584 5176 7588
rect 5192 7644 5256 7648
rect 5192 7588 5196 7644
rect 5196 7588 5252 7644
rect 5252 7588 5256 7644
rect 5192 7584 5256 7588
rect 12952 7644 13016 7648
rect 12952 7588 12956 7644
rect 12956 7588 13012 7644
rect 13012 7588 13016 7644
rect 12952 7584 13016 7588
rect 13032 7644 13096 7648
rect 13032 7588 13036 7644
rect 13036 7588 13092 7644
rect 13092 7588 13096 7644
rect 13032 7584 13096 7588
rect 13112 7644 13176 7648
rect 13112 7588 13116 7644
rect 13116 7588 13172 7644
rect 13172 7588 13176 7644
rect 13112 7584 13176 7588
rect 13192 7644 13256 7648
rect 13192 7588 13196 7644
rect 13196 7588 13252 7644
rect 13252 7588 13256 7644
rect 13192 7584 13256 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 8952 7100 9016 7104
rect 8952 7044 8956 7100
rect 8956 7044 9012 7100
rect 9012 7044 9016 7100
rect 8952 7040 9016 7044
rect 9032 7100 9096 7104
rect 9032 7044 9036 7100
rect 9036 7044 9092 7100
rect 9092 7044 9096 7100
rect 9032 7040 9096 7044
rect 9112 7100 9176 7104
rect 9112 7044 9116 7100
rect 9116 7044 9172 7100
rect 9172 7044 9176 7100
rect 9112 7040 9176 7044
rect 9192 7100 9256 7104
rect 9192 7044 9196 7100
rect 9196 7044 9252 7100
rect 9252 7044 9256 7100
rect 9192 7040 9256 7044
rect 16952 7100 17016 7104
rect 16952 7044 16956 7100
rect 16956 7044 17012 7100
rect 17012 7044 17016 7100
rect 16952 7040 17016 7044
rect 17032 7100 17096 7104
rect 17032 7044 17036 7100
rect 17036 7044 17092 7100
rect 17092 7044 17096 7100
rect 17032 7040 17096 7044
rect 17112 7100 17176 7104
rect 17112 7044 17116 7100
rect 17116 7044 17172 7100
rect 17172 7044 17176 7100
rect 17112 7040 17176 7044
rect 17192 7100 17256 7104
rect 17192 7044 17196 7100
rect 17196 7044 17252 7100
rect 17252 7044 17256 7100
rect 17192 7040 17256 7044
rect 4952 6556 5016 6560
rect 4952 6500 4956 6556
rect 4956 6500 5012 6556
rect 5012 6500 5016 6556
rect 4952 6496 5016 6500
rect 5032 6556 5096 6560
rect 5032 6500 5036 6556
rect 5036 6500 5092 6556
rect 5092 6500 5096 6556
rect 5032 6496 5096 6500
rect 5112 6556 5176 6560
rect 5112 6500 5116 6556
rect 5116 6500 5172 6556
rect 5172 6500 5176 6556
rect 5112 6496 5176 6500
rect 5192 6556 5256 6560
rect 5192 6500 5196 6556
rect 5196 6500 5252 6556
rect 5252 6500 5256 6556
rect 5192 6496 5256 6500
rect 12952 6556 13016 6560
rect 12952 6500 12956 6556
rect 12956 6500 13012 6556
rect 13012 6500 13016 6556
rect 12952 6496 13016 6500
rect 13032 6556 13096 6560
rect 13032 6500 13036 6556
rect 13036 6500 13092 6556
rect 13092 6500 13096 6556
rect 13032 6496 13096 6500
rect 13112 6556 13176 6560
rect 13112 6500 13116 6556
rect 13116 6500 13172 6556
rect 13172 6500 13176 6556
rect 13112 6496 13176 6500
rect 13192 6556 13256 6560
rect 13192 6500 13196 6556
rect 13196 6500 13252 6556
rect 13252 6500 13256 6556
rect 13192 6496 13256 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 8952 6012 9016 6016
rect 8952 5956 8956 6012
rect 8956 5956 9012 6012
rect 9012 5956 9016 6012
rect 8952 5952 9016 5956
rect 9032 6012 9096 6016
rect 9032 5956 9036 6012
rect 9036 5956 9092 6012
rect 9092 5956 9096 6012
rect 9032 5952 9096 5956
rect 9112 6012 9176 6016
rect 9112 5956 9116 6012
rect 9116 5956 9172 6012
rect 9172 5956 9176 6012
rect 9112 5952 9176 5956
rect 9192 6012 9256 6016
rect 9192 5956 9196 6012
rect 9196 5956 9252 6012
rect 9252 5956 9256 6012
rect 9192 5952 9256 5956
rect 16952 6012 17016 6016
rect 16952 5956 16956 6012
rect 16956 5956 17012 6012
rect 17012 5956 17016 6012
rect 16952 5952 17016 5956
rect 17032 6012 17096 6016
rect 17032 5956 17036 6012
rect 17036 5956 17092 6012
rect 17092 5956 17096 6012
rect 17032 5952 17096 5956
rect 17112 6012 17176 6016
rect 17112 5956 17116 6012
rect 17116 5956 17172 6012
rect 17172 5956 17176 6012
rect 17112 5952 17176 5956
rect 17192 6012 17256 6016
rect 17192 5956 17196 6012
rect 17196 5956 17252 6012
rect 17252 5956 17256 6012
rect 17192 5952 17256 5956
rect 4952 5468 5016 5472
rect 4952 5412 4956 5468
rect 4956 5412 5012 5468
rect 5012 5412 5016 5468
rect 4952 5408 5016 5412
rect 5032 5468 5096 5472
rect 5032 5412 5036 5468
rect 5036 5412 5092 5468
rect 5092 5412 5096 5468
rect 5032 5408 5096 5412
rect 5112 5468 5176 5472
rect 5112 5412 5116 5468
rect 5116 5412 5172 5468
rect 5172 5412 5176 5468
rect 5112 5408 5176 5412
rect 5192 5468 5256 5472
rect 5192 5412 5196 5468
rect 5196 5412 5252 5468
rect 5252 5412 5256 5468
rect 5192 5408 5256 5412
rect 12952 5468 13016 5472
rect 12952 5412 12956 5468
rect 12956 5412 13012 5468
rect 13012 5412 13016 5468
rect 12952 5408 13016 5412
rect 13032 5468 13096 5472
rect 13032 5412 13036 5468
rect 13036 5412 13092 5468
rect 13092 5412 13096 5468
rect 13032 5408 13096 5412
rect 13112 5468 13176 5472
rect 13112 5412 13116 5468
rect 13116 5412 13172 5468
rect 13172 5412 13176 5468
rect 13112 5408 13176 5412
rect 13192 5468 13256 5472
rect 13192 5412 13196 5468
rect 13196 5412 13252 5468
rect 13252 5412 13256 5468
rect 13192 5408 13256 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 8952 4924 9016 4928
rect 8952 4868 8956 4924
rect 8956 4868 9012 4924
rect 9012 4868 9016 4924
rect 8952 4864 9016 4868
rect 9032 4924 9096 4928
rect 9032 4868 9036 4924
rect 9036 4868 9092 4924
rect 9092 4868 9096 4924
rect 9032 4864 9096 4868
rect 9112 4924 9176 4928
rect 9112 4868 9116 4924
rect 9116 4868 9172 4924
rect 9172 4868 9176 4924
rect 9112 4864 9176 4868
rect 9192 4924 9256 4928
rect 9192 4868 9196 4924
rect 9196 4868 9252 4924
rect 9252 4868 9256 4924
rect 9192 4864 9256 4868
rect 16952 4924 17016 4928
rect 16952 4868 16956 4924
rect 16956 4868 17012 4924
rect 17012 4868 17016 4924
rect 16952 4864 17016 4868
rect 17032 4924 17096 4928
rect 17032 4868 17036 4924
rect 17036 4868 17092 4924
rect 17092 4868 17096 4924
rect 17032 4864 17096 4868
rect 17112 4924 17176 4928
rect 17112 4868 17116 4924
rect 17116 4868 17172 4924
rect 17172 4868 17176 4924
rect 17112 4864 17176 4868
rect 17192 4924 17256 4928
rect 17192 4868 17196 4924
rect 17196 4868 17252 4924
rect 17252 4868 17256 4924
rect 17192 4864 17256 4868
rect 4952 4380 5016 4384
rect 4952 4324 4956 4380
rect 4956 4324 5012 4380
rect 5012 4324 5016 4380
rect 4952 4320 5016 4324
rect 5032 4380 5096 4384
rect 5032 4324 5036 4380
rect 5036 4324 5092 4380
rect 5092 4324 5096 4380
rect 5032 4320 5096 4324
rect 5112 4380 5176 4384
rect 5112 4324 5116 4380
rect 5116 4324 5172 4380
rect 5172 4324 5176 4380
rect 5112 4320 5176 4324
rect 5192 4380 5256 4384
rect 5192 4324 5196 4380
rect 5196 4324 5252 4380
rect 5252 4324 5256 4380
rect 5192 4320 5256 4324
rect 12952 4380 13016 4384
rect 12952 4324 12956 4380
rect 12956 4324 13012 4380
rect 13012 4324 13016 4380
rect 12952 4320 13016 4324
rect 13032 4380 13096 4384
rect 13032 4324 13036 4380
rect 13036 4324 13092 4380
rect 13092 4324 13096 4380
rect 13032 4320 13096 4324
rect 13112 4380 13176 4384
rect 13112 4324 13116 4380
rect 13116 4324 13172 4380
rect 13172 4324 13176 4380
rect 13112 4320 13176 4324
rect 13192 4380 13256 4384
rect 13192 4324 13196 4380
rect 13196 4324 13252 4380
rect 13252 4324 13256 4380
rect 13192 4320 13256 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 8952 3836 9016 3840
rect 8952 3780 8956 3836
rect 8956 3780 9012 3836
rect 9012 3780 9016 3836
rect 8952 3776 9016 3780
rect 9032 3836 9096 3840
rect 9032 3780 9036 3836
rect 9036 3780 9092 3836
rect 9092 3780 9096 3836
rect 9032 3776 9096 3780
rect 9112 3836 9176 3840
rect 9112 3780 9116 3836
rect 9116 3780 9172 3836
rect 9172 3780 9176 3836
rect 9112 3776 9176 3780
rect 9192 3836 9256 3840
rect 9192 3780 9196 3836
rect 9196 3780 9252 3836
rect 9252 3780 9256 3836
rect 9192 3776 9256 3780
rect 16952 3836 17016 3840
rect 16952 3780 16956 3836
rect 16956 3780 17012 3836
rect 17012 3780 17016 3836
rect 16952 3776 17016 3780
rect 17032 3836 17096 3840
rect 17032 3780 17036 3836
rect 17036 3780 17092 3836
rect 17092 3780 17096 3836
rect 17032 3776 17096 3780
rect 17112 3836 17176 3840
rect 17112 3780 17116 3836
rect 17116 3780 17172 3836
rect 17172 3780 17176 3836
rect 17112 3776 17176 3780
rect 17192 3836 17256 3840
rect 17192 3780 17196 3836
rect 17196 3780 17252 3836
rect 17252 3780 17256 3836
rect 17192 3776 17256 3780
rect 4952 3292 5016 3296
rect 4952 3236 4956 3292
rect 4956 3236 5012 3292
rect 5012 3236 5016 3292
rect 4952 3232 5016 3236
rect 5032 3292 5096 3296
rect 5032 3236 5036 3292
rect 5036 3236 5092 3292
rect 5092 3236 5096 3292
rect 5032 3232 5096 3236
rect 5112 3292 5176 3296
rect 5112 3236 5116 3292
rect 5116 3236 5172 3292
rect 5172 3236 5176 3292
rect 5112 3232 5176 3236
rect 5192 3292 5256 3296
rect 5192 3236 5196 3292
rect 5196 3236 5252 3292
rect 5252 3236 5256 3292
rect 5192 3232 5256 3236
rect 12952 3292 13016 3296
rect 12952 3236 12956 3292
rect 12956 3236 13012 3292
rect 13012 3236 13016 3292
rect 12952 3232 13016 3236
rect 13032 3292 13096 3296
rect 13032 3236 13036 3292
rect 13036 3236 13092 3292
rect 13092 3236 13096 3292
rect 13032 3232 13096 3236
rect 13112 3292 13176 3296
rect 13112 3236 13116 3292
rect 13116 3236 13172 3292
rect 13172 3236 13176 3292
rect 13112 3232 13176 3236
rect 13192 3292 13256 3296
rect 13192 3236 13196 3292
rect 13196 3236 13252 3292
rect 13252 3236 13256 3292
rect 13192 3232 13256 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 8952 2748 9016 2752
rect 8952 2692 8956 2748
rect 8956 2692 9012 2748
rect 9012 2692 9016 2748
rect 8952 2688 9016 2692
rect 9032 2748 9096 2752
rect 9032 2692 9036 2748
rect 9036 2692 9092 2748
rect 9092 2692 9096 2748
rect 9032 2688 9096 2692
rect 9112 2748 9176 2752
rect 9112 2692 9116 2748
rect 9116 2692 9172 2748
rect 9172 2692 9176 2748
rect 9112 2688 9176 2692
rect 9192 2748 9256 2752
rect 9192 2692 9196 2748
rect 9196 2692 9252 2748
rect 9252 2692 9256 2748
rect 9192 2688 9256 2692
rect 16952 2748 17016 2752
rect 16952 2692 16956 2748
rect 16956 2692 17012 2748
rect 17012 2692 17016 2748
rect 16952 2688 17016 2692
rect 17032 2748 17096 2752
rect 17032 2692 17036 2748
rect 17036 2692 17092 2748
rect 17092 2692 17096 2748
rect 17032 2688 17096 2692
rect 17112 2748 17176 2752
rect 17112 2692 17116 2748
rect 17116 2692 17172 2748
rect 17172 2692 17176 2748
rect 17112 2688 17176 2692
rect 17192 2748 17256 2752
rect 17192 2692 17196 2748
rect 17196 2692 17252 2748
rect 17252 2692 17256 2748
rect 17192 2688 17256 2692
rect 16620 2348 16684 2412
rect 4952 2204 5016 2208
rect 4952 2148 4956 2204
rect 4956 2148 5012 2204
rect 5012 2148 5016 2204
rect 4952 2144 5016 2148
rect 5032 2204 5096 2208
rect 5032 2148 5036 2204
rect 5036 2148 5092 2204
rect 5092 2148 5096 2204
rect 5032 2144 5096 2148
rect 5112 2204 5176 2208
rect 5112 2148 5116 2204
rect 5116 2148 5172 2204
rect 5172 2148 5176 2204
rect 5112 2144 5176 2148
rect 5192 2204 5256 2208
rect 5192 2148 5196 2204
rect 5196 2148 5252 2204
rect 5252 2148 5256 2204
rect 5192 2144 5256 2148
rect 12952 2204 13016 2208
rect 12952 2148 12956 2204
rect 12956 2148 13012 2204
rect 13012 2148 13016 2204
rect 12952 2144 13016 2148
rect 13032 2204 13096 2208
rect 13032 2148 13036 2204
rect 13036 2148 13092 2204
rect 13092 2148 13096 2204
rect 13032 2144 13096 2148
rect 13112 2204 13176 2208
rect 13112 2148 13116 2204
rect 13116 2148 13172 2204
rect 13172 2148 13176 2204
rect 13112 2144 13176 2148
rect 13192 2204 13256 2208
rect 13192 2148 13196 2204
rect 13196 2148 13252 2204
rect 13252 2148 13256 2204
rect 13192 2144 13256 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
<< metal4 >>
rect 4944 21792 5264 21808
rect 4944 21728 4952 21792
rect 5016 21728 5032 21792
rect 5096 21728 5112 21792
rect 5176 21728 5192 21792
rect 5256 21728 5264 21792
rect 4944 20704 5264 21728
rect 4944 20640 4952 20704
rect 5016 20640 5032 20704
rect 5096 20640 5112 20704
rect 5176 20640 5192 20704
rect 5256 20640 5264 20704
rect 4944 19616 5264 20640
rect 4944 19552 4952 19616
rect 5016 19552 5032 19616
rect 5096 19552 5112 19616
rect 5176 19552 5192 19616
rect 5256 19552 5264 19616
rect 4944 18528 5264 19552
rect 4944 18464 4952 18528
rect 5016 18464 5032 18528
rect 5096 18464 5112 18528
rect 5176 18464 5192 18528
rect 5256 18464 5264 18528
rect 4944 17440 5264 18464
rect 4944 17376 4952 17440
rect 5016 17376 5032 17440
rect 5096 17376 5112 17440
rect 5176 17376 5192 17440
rect 5256 17376 5264 17440
rect 4944 16352 5264 17376
rect 4944 16288 4952 16352
rect 5016 16288 5032 16352
rect 5096 16288 5112 16352
rect 5176 16288 5192 16352
rect 5256 16288 5264 16352
rect 4944 15264 5264 16288
rect 4944 15200 4952 15264
rect 5016 15200 5032 15264
rect 5096 15200 5112 15264
rect 5176 15200 5192 15264
rect 5256 15200 5264 15264
rect 4944 14176 5264 15200
rect 4944 14112 4952 14176
rect 5016 14112 5032 14176
rect 5096 14112 5112 14176
rect 5176 14112 5192 14176
rect 5256 14112 5264 14176
rect 4944 13088 5264 14112
rect 4944 13024 4952 13088
rect 5016 13024 5032 13088
rect 5096 13024 5112 13088
rect 5176 13024 5192 13088
rect 5256 13024 5264 13088
rect 59 12748 125 12749
rect 59 12684 60 12748
rect 124 12684 125 12748
rect 59 12683 125 12684
rect 62 12341 122 12683
rect 59 12340 125 12341
rect 59 12276 60 12340
rect 124 12276 125 12340
rect 59 12275 125 12276
rect 4944 12000 5264 13024
rect 4944 11936 4952 12000
rect 5016 11936 5032 12000
rect 5096 11936 5112 12000
rect 5176 11936 5192 12000
rect 5256 11936 5264 12000
rect 4944 10912 5264 11936
rect 4944 10848 4952 10912
rect 5016 10848 5032 10912
rect 5096 10848 5112 10912
rect 5176 10848 5192 10912
rect 5256 10848 5264 10912
rect 59 10028 125 10029
rect 59 9964 60 10028
rect 124 9964 125 10028
rect 59 9963 125 9964
rect 62 9757 122 9963
rect 4944 9824 5264 10848
rect 4944 9760 4952 9824
rect 5016 9760 5032 9824
rect 5096 9760 5112 9824
rect 5176 9760 5192 9824
rect 5256 9760 5264 9824
rect 59 9756 125 9757
rect 59 9692 60 9756
rect 124 9692 125 9756
rect 59 9691 125 9692
rect 4944 8736 5264 9760
rect 4944 8672 4952 8736
rect 5016 8672 5032 8736
rect 5096 8672 5112 8736
rect 5176 8672 5192 8736
rect 5256 8672 5264 8736
rect 4944 7648 5264 8672
rect 8944 21248 9264 21808
rect 8944 21184 8952 21248
rect 9016 21184 9032 21248
rect 9096 21184 9112 21248
rect 9176 21184 9192 21248
rect 9256 21184 9264 21248
rect 8944 20160 9264 21184
rect 8944 20096 8952 20160
rect 9016 20096 9032 20160
rect 9096 20096 9112 20160
rect 9176 20096 9192 20160
rect 9256 20096 9264 20160
rect 8944 19072 9264 20096
rect 8944 19008 8952 19072
rect 9016 19008 9032 19072
rect 9096 19008 9112 19072
rect 9176 19008 9192 19072
rect 9256 19008 9264 19072
rect 8944 17984 9264 19008
rect 8944 17920 8952 17984
rect 9016 17920 9032 17984
rect 9096 17920 9112 17984
rect 9176 17920 9192 17984
rect 9256 17920 9264 17984
rect 8944 16896 9264 17920
rect 8944 16832 8952 16896
rect 9016 16832 9032 16896
rect 9096 16832 9112 16896
rect 9176 16832 9192 16896
rect 9256 16832 9264 16896
rect 8944 15808 9264 16832
rect 8944 15744 8952 15808
rect 9016 15744 9032 15808
rect 9096 15744 9112 15808
rect 9176 15744 9192 15808
rect 9256 15744 9264 15808
rect 8944 14720 9264 15744
rect 8944 14656 8952 14720
rect 9016 14656 9032 14720
rect 9096 14656 9112 14720
rect 9176 14656 9192 14720
rect 9256 14656 9264 14720
rect 8944 13632 9264 14656
rect 8944 13568 8952 13632
rect 9016 13568 9032 13632
rect 9096 13568 9112 13632
rect 9176 13568 9192 13632
rect 9256 13568 9264 13632
rect 8944 12544 9264 13568
rect 8944 12480 8952 12544
rect 9016 12480 9032 12544
rect 9096 12480 9112 12544
rect 9176 12480 9192 12544
rect 9256 12480 9264 12544
rect 8944 11456 9264 12480
rect 8944 11392 8952 11456
rect 9016 11392 9032 11456
rect 9096 11392 9112 11456
rect 9176 11392 9192 11456
rect 9256 11392 9264 11456
rect 8944 10368 9264 11392
rect 8944 10304 8952 10368
rect 9016 10304 9032 10368
rect 9096 10304 9112 10368
rect 9176 10304 9192 10368
rect 9256 10304 9264 10368
rect 8944 9280 9264 10304
rect 8944 9216 8952 9280
rect 9016 9216 9032 9280
rect 9096 9216 9112 9280
rect 9176 9216 9192 9280
rect 9256 9216 9264 9280
rect 7603 8260 7669 8261
rect 7603 8196 7604 8260
rect 7668 8196 7669 8260
rect 7603 8195 7669 8196
rect 4944 7584 4952 7648
rect 5016 7584 5032 7648
rect 5096 7584 5112 7648
rect 5176 7584 5192 7648
rect 5256 7584 5264 7648
rect 4944 6560 5264 7584
rect 4944 6496 4952 6560
rect 5016 6496 5032 6560
rect 5096 6496 5112 6560
rect 5176 6496 5192 6560
rect 5256 6496 5264 6560
rect 4944 5472 5264 6496
rect 4944 5408 4952 5472
rect 5016 5408 5032 5472
rect 5096 5408 5112 5472
rect 5176 5408 5192 5472
rect 5256 5408 5264 5472
rect 4944 4384 5264 5408
rect 4944 4320 4952 4384
rect 5016 4320 5032 4384
rect 5096 4320 5112 4384
rect 5176 4320 5192 4384
rect 5256 4320 5264 4384
rect 4944 3296 5264 4320
rect 4944 3232 4952 3296
rect 5016 3232 5032 3296
rect 5096 3232 5112 3296
rect 5176 3232 5192 3296
rect 5256 3232 5264 3296
rect 4944 2208 5264 3232
rect 7606 2498 7666 8195
rect 8944 8192 9264 9216
rect 8944 8128 8952 8192
rect 9016 8128 9032 8192
rect 9096 8128 9112 8192
rect 9176 8128 9192 8192
rect 9256 8128 9264 8192
rect 8944 7104 9264 8128
rect 8944 7040 8952 7104
rect 9016 7040 9032 7104
rect 9096 7040 9112 7104
rect 9176 7040 9192 7104
rect 9256 7040 9264 7104
rect 8944 6016 9264 7040
rect 8944 5952 8952 6016
rect 9016 5952 9032 6016
rect 9096 5952 9112 6016
rect 9176 5952 9192 6016
rect 9256 5952 9264 6016
rect 8944 4928 9264 5952
rect 8944 4864 8952 4928
rect 9016 4864 9032 4928
rect 9096 4864 9112 4928
rect 9176 4864 9192 4928
rect 9256 4864 9264 4928
rect 8944 3840 9264 4864
rect 8944 3776 8952 3840
rect 9016 3776 9032 3840
rect 9096 3776 9112 3840
rect 9176 3776 9192 3840
rect 9256 3776 9264 3840
rect 8944 2752 9264 3776
rect 8944 2688 8952 2752
rect 9016 2688 9032 2752
rect 9096 2688 9112 2752
rect 9176 2688 9192 2752
rect 9256 2688 9264 2752
rect 4944 2144 4952 2208
rect 5016 2144 5032 2208
rect 5096 2144 5112 2208
rect 5176 2144 5192 2208
rect 5256 2144 5264 2208
rect 4944 2128 5264 2144
rect 8944 2128 9264 2688
rect 12944 21792 13264 21808
rect 12944 21728 12952 21792
rect 13016 21728 13032 21792
rect 13096 21728 13112 21792
rect 13176 21728 13192 21792
rect 13256 21728 13264 21792
rect 12944 20704 13264 21728
rect 12944 20640 12952 20704
rect 13016 20640 13032 20704
rect 13096 20640 13112 20704
rect 13176 20640 13192 20704
rect 13256 20640 13264 20704
rect 12944 19616 13264 20640
rect 12944 19552 12952 19616
rect 13016 19552 13032 19616
rect 13096 19552 13112 19616
rect 13176 19552 13192 19616
rect 13256 19552 13264 19616
rect 12944 18528 13264 19552
rect 12944 18464 12952 18528
rect 13016 18464 13032 18528
rect 13096 18464 13112 18528
rect 13176 18464 13192 18528
rect 13256 18464 13264 18528
rect 12944 17440 13264 18464
rect 12944 17376 12952 17440
rect 13016 17376 13032 17440
rect 13096 17376 13112 17440
rect 13176 17376 13192 17440
rect 13256 17376 13264 17440
rect 12944 16352 13264 17376
rect 12944 16288 12952 16352
rect 13016 16288 13032 16352
rect 13096 16288 13112 16352
rect 13176 16288 13192 16352
rect 13256 16288 13264 16352
rect 12944 15264 13264 16288
rect 12944 15200 12952 15264
rect 13016 15200 13032 15264
rect 13096 15200 13112 15264
rect 13176 15200 13192 15264
rect 13256 15200 13264 15264
rect 12944 14176 13264 15200
rect 12944 14112 12952 14176
rect 13016 14112 13032 14176
rect 13096 14112 13112 14176
rect 13176 14112 13192 14176
rect 13256 14112 13264 14176
rect 12944 13088 13264 14112
rect 12944 13024 12952 13088
rect 13016 13024 13032 13088
rect 13096 13024 13112 13088
rect 13176 13024 13192 13088
rect 13256 13024 13264 13088
rect 12944 12000 13264 13024
rect 12944 11936 12952 12000
rect 13016 11936 13032 12000
rect 13096 11936 13112 12000
rect 13176 11936 13192 12000
rect 13256 11936 13264 12000
rect 12944 10912 13264 11936
rect 12944 10848 12952 10912
rect 13016 10848 13032 10912
rect 13096 10848 13112 10912
rect 13176 10848 13192 10912
rect 13256 10848 13264 10912
rect 12944 9824 13264 10848
rect 12944 9760 12952 9824
rect 13016 9760 13032 9824
rect 13096 9760 13112 9824
rect 13176 9760 13192 9824
rect 13256 9760 13264 9824
rect 12944 8736 13264 9760
rect 12944 8672 12952 8736
rect 13016 8672 13032 8736
rect 13096 8672 13112 8736
rect 13176 8672 13192 8736
rect 13256 8672 13264 8736
rect 12944 7648 13264 8672
rect 12944 7584 12952 7648
rect 13016 7584 13032 7648
rect 13096 7584 13112 7648
rect 13176 7584 13192 7648
rect 13256 7584 13264 7648
rect 12944 6560 13264 7584
rect 12944 6496 12952 6560
rect 13016 6496 13032 6560
rect 13096 6496 13112 6560
rect 13176 6496 13192 6560
rect 13256 6496 13264 6560
rect 12944 5472 13264 6496
rect 12944 5408 12952 5472
rect 13016 5408 13032 5472
rect 13096 5408 13112 5472
rect 13176 5408 13192 5472
rect 13256 5408 13264 5472
rect 12944 4384 13264 5408
rect 12944 4320 12952 4384
rect 13016 4320 13032 4384
rect 13096 4320 13112 4384
rect 13176 4320 13192 4384
rect 13256 4320 13264 4384
rect 12944 3296 13264 4320
rect 12944 3232 12952 3296
rect 13016 3232 13032 3296
rect 13096 3232 13112 3296
rect 13176 3232 13192 3296
rect 13256 3232 13264 3296
rect 12944 2208 13264 3232
rect 16944 21248 17264 21808
rect 16944 21184 16952 21248
rect 17016 21184 17032 21248
rect 17096 21184 17112 21248
rect 17176 21184 17192 21248
rect 17256 21184 17264 21248
rect 16944 20160 17264 21184
rect 16944 20096 16952 20160
rect 17016 20096 17032 20160
rect 17096 20096 17112 20160
rect 17176 20096 17192 20160
rect 17256 20096 17264 20160
rect 16944 19072 17264 20096
rect 16944 19008 16952 19072
rect 17016 19008 17032 19072
rect 17096 19008 17112 19072
rect 17176 19008 17192 19072
rect 17256 19008 17264 19072
rect 16944 17984 17264 19008
rect 16944 17920 16952 17984
rect 17016 17920 17032 17984
rect 17096 17920 17112 17984
rect 17176 17920 17192 17984
rect 17256 17920 17264 17984
rect 16944 16896 17264 17920
rect 16944 16832 16952 16896
rect 17016 16832 17032 16896
rect 17096 16832 17112 16896
rect 17176 16832 17192 16896
rect 17256 16832 17264 16896
rect 16944 15808 17264 16832
rect 16944 15744 16952 15808
rect 17016 15744 17032 15808
rect 17096 15744 17112 15808
rect 17176 15744 17192 15808
rect 17256 15744 17264 15808
rect 16944 14720 17264 15744
rect 16944 14656 16952 14720
rect 17016 14656 17032 14720
rect 17096 14656 17112 14720
rect 17176 14656 17192 14720
rect 17256 14656 17264 14720
rect 16944 13632 17264 14656
rect 16944 13568 16952 13632
rect 17016 13568 17032 13632
rect 17096 13568 17112 13632
rect 17176 13568 17192 13632
rect 17256 13568 17264 13632
rect 16944 12544 17264 13568
rect 16944 12480 16952 12544
rect 17016 12480 17032 12544
rect 17096 12480 17112 12544
rect 17176 12480 17192 12544
rect 17256 12480 17264 12544
rect 16944 11456 17264 12480
rect 16944 11392 16952 11456
rect 17016 11392 17032 11456
rect 17096 11392 17112 11456
rect 17176 11392 17192 11456
rect 17256 11392 17264 11456
rect 16944 10368 17264 11392
rect 16944 10304 16952 10368
rect 17016 10304 17032 10368
rect 17096 10304 17112 10368
rect 17176 10304 17192 10368
rect 17256 10304 17264 10368
rect 16944 9280 17264 10304
rect 16944 9216 16952 9280
rect 17016 9216 17032 9280
rect 17096 9216 17112 9280
rect 17176 9216 17192 9280
rect 17256 9216 17264 9280
rect 16944 8192 17264 9216
rect 16944 8128 16952 8192
rect 17016 8128 17032 8192
rect 17096 8128 17112 8192
rect 17176 8128 17192 8192
rect 17256 8128 17264 8192
rect 16944 7104 17264 8128
rect 16944 7040 16952 7104
rect 17016 7040 17032 7104
rect 17096 7040 17112 7104
rect 17176 7040 17192 7104
rect 17256 7040 17264 7104
rect 16944 6016 17264 7040
rect 16944 5952 16952 6016
rect 17016 5952 17032 6016
rect 17096 5952 17112 6016
rect 17176 5952 17192 6016
rect 17256 5952 17264 6016
rect 16944 4928 17264 5952
rect 16944 4864 16952 4928
rect 17016 4864 17032 4928
rect 17096 4864 17112 4928
rect 17176 4864 17192 4928
rect 17256 4864 17264 4928
rect 16944 3840 17264 4864
rect 16944 3776 16952 3840
rect 17016 3776 17032 3840
rect 17096 3776 17112 3840
rect 17176 3776 17192 3840
rect 17256 3776 17264 3840
rect 16944 2752 17264 3776
rect 16944 2688 16952 2752
rect 17016 2688 17032 2752
rect 17096 2688 17112 2752
rect 17176 2688 17192 2752
rect 17256 2688 17264 2752
rect 12944 2144 12952 2208
rect 13016 2144 13032 2208
rect 13096 2144 13112 2208
rect 13176 2144 13192 2208
rect 13256 2144 13264 2208
rect 12944 2128 13264 2144
rect 16944 2128 17264 2688
rect 20944 21792 21264 21808
rect 20944 21728 20952 21792
rect 21016 21728 21032 21792
rect 21096 21728 21112 21792
rect 21176 21728 21192 21792
rect 21256 21728 21264 21792
rect 20944 20704 21264 21728
rect 20944 20640 20952 20704
rect 21016 20640 21032 20704
rect 21096 20640 21112 20704
rect 21176 20640 21192 20704
rect 21256 20640 21264 20704
rect 20944 19616 21264 20640
rect 20944 19552 20952 19616
rect 21016 19552 21032 19616
rect 21096 19552 21112 19616
rect 21176 19552 21192 19616
rect 21256 19552 21264 19616
rect 20944 18528 21264 19552
rect 20944 18464 20952 18528
rect 21016 18464 21032 18528
rect 21096 18464 21112 18528
rect 21176 18464 21192 18528
rect 21256 18464 21264 18528
rect 20944 17440 21264 18464
rect 20944 17376 20952 17440
rect 21016 17376 21032 17440
rect 21096 17376 21112 17440
rect 21176 17376 21192 17440
rect 21256 17376 21264 17440
rect 20944 16352 21264 17376
rect 20944 16288 20952 16352
rect 21016 16288 21032 16352
rect 21096 16288 21112 16352
rect 21176 16288 21192 16352
rect 21256 16288 21264 16352
rect 20944 15264 21264 16288
rect 20944 15200 20952 15264
rect 21016 15200 21032 15264
rect 21096 15200 21112 15264
rect 21176 15200 21192 15264
rect 21256 15200 21264 15264
rect 20944 14176 21264 15200
rect 20944 14112 20952 14176
rect 21016 14112 21032 14176
rect 21096 14112 21112 14176
rect 21176 14112 21192 14176
rect 21256 14112 21264 14176
rect 20944 13088 21264 14112
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 23611 8124 23677 8125
rect 23611 8060 23612 8124
rect 23676 8060 23677 8124
rect 23611 8059 23677 8060
rect 23614 7853 23674 8059
rect 23611 7852 23677 7853
rect 23611 7788 23612 7852
rect 23676 7788 23677 7852
rect 23611 7787 23677 7788
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 2208 21264 3232
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
<< via4 >>
rect 7518 2262 7754 2498
rect 16534 2412 16770 2498
rect 16534 2348 16620 2412
rect 16620 2348 16684 2412
rect 16684 2348 16770 2412
rect 16534 2262 16770 2348
<< metal5 >>
rect 7476 2498 16812 2540
rect 7476 2262 7518 2498
rect 7754 2262 16534 2498
rect 16770 2262 16812 2498
rect 7476 2220 16812 2262
use scs8hd_fill_1  FILLER_0_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_0_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__063__B tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_6  FILLER_1_15 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_10 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use scs8hd_nor2_4  _063_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_1  FILLER_1_21
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 3128 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_33
timestamp 1586364061
transform 1 0 4140 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_72 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_5_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1050 592
use scs8hd_nor2_4  _064_
timestamp 1586364061
transform 1 0 3312 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_39
timestamp 1586364061
transform 1 0 4692 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_43
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_50
timestamp 1586364061
transform 1 0 5704 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_47
timestamp 1586364061
transform 1 0 5428 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5612 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5888 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 222 592
use scs8hd_conb_1  _134_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4876 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_58
timestamp 1586364061
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_54
timestamp 1586364061
transform 1 0 6072 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6256 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_69
timestamp 1586364061
transform 1 0 7452 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_67
timestamp 1586364061
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 6992 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use scs8hd_conb_1  _138_
timestamp 1586364061
transform 1 0 7176 0 1 2720
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7636 0 -1 2720
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__092__B
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8832 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_82
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_86
timestamp 1586364061
transform 1 0 9016 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_75
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_86
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_92
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_97
timestamp 1586364061
transform 1 0 10028 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_90
timestamp 1586364061
transform 1 0 9384 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__B
timestamp 1586364061
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9752 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_107
timestamp 1586364061
transform 1 0 10948 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_101
timestamp 1586364061
transform 1 0 10396 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 10212 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_4_.latch
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9936 0 1 2720
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_1_111
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11132 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_115
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_119
timestamp 1586364061
transform 1 0 12052 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _147_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_131
timestamp 1586364061
transform 1 0 13156 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_127
timestamp 1586364061
transform 1 0 12788 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__C
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__039__A
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _145_
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use scs8hd_nor4_4  _106_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 13616 0 1 2720
box -38 -48 1602 592
use scs8hd_nor2_4  _093_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_0_146
timestamp 1586364061
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_150
timestamp 1586364061
transform 1 0 14904 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 14720 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_1_153
timestamp 1586364061
transform 1 0 15180 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_156
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__048__A
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__060__C
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_160
timestamp 1586364061
transform 1 0 15824 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 15640 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_178
timestamp 1586364061
transform 1 0 17480 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_174
timestamp 1586364061
transform 1 0 17112 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_170
timestamp 1586364061
transform 1 0 16744 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_176
timestamp 1586364061
transform 1 0 17296 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_170
timestamp 1586364061
transform 1 0 16744 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 17112 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__043__A
timestamp 1586364061
transform 1 0 17296 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__060__B
timestamp 1586364061
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use scs8hd_or3_4  _048_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15916 0 -1 2720
box -38 -48 866 592
use scs8hd_inv_8  _043_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15916 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__B
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__A
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__C
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_193
timestamp 1586364061
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use scs8hd_or3_4  _054_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use scs8hd_or3_4  _052_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_201
timestamp 1586364061
transform 1 0 19596 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_197
timestamp 1586364061
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_200
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__B
timestamp 1586364061
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__A
timestamp 1586364061
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__048__C
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _156_
timestamp 1586364061
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_212
timestamp 1586364061
transform 1 0 20608 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_212
timestamp 1586364061
transform 1 0 20608 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_208
timestamp 1586364061
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 20424 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19780 0 1 2720
box -38 -48 866 592
use scs8hd_buf_2  _149_
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 21712 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_216
timestamp 1586364061
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_222
timestamp 1586364061
transform 1 0 21528 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_226
timestamp 1586364061
transform 1 0 21896 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_217
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_229
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 22816 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 22816 0 1 2720
box -38 -48 314 592
use scs8hd_fill_1  FILLER_0_232
timestamp 1586364061
transform 1 0 22448 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__065__B
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_9
timestamp 1586364061
transform 1 0 1932 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_12
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__064__B
timestamp 1586364061
transform 1 0 3312 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_26
timestamp 1586364061
transform 1 0 3496 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_30
timestamp 1586364061
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4508 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5704 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_36
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_48
timestamp 1586364061
transform 1 0 5520 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_52
timestamp 1586364061
transform 1 0 5888 0 -1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6256 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_65
timestamp 1586364061
transform 1 0 7084 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_69
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _092_
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__068__B
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_82
timestamp 1586364061
transform 1 0 8648 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_86
timestamp 1586364061
transform 1 0 9016 0 -1 3808
box -38 -48 406 592
use scs8hd_nor2_4  _094_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_102
timestamp 1586364061
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_106
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11316 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_120
timestamp 1586364061
transform 1 0 12144 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_124
timestamp 1586364061
transform 1 0 12512 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_8  _039_
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__045__A
timestamp 1586364061
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__D
timestamp 1586364061
transform 1 0 13432 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_127
timestamp 1586364061
transform 1 0 12788 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_131
timestamp 1586364061
transform 1 0 13156 0 -1 3808
box -38 -48 314 592
use scs8hd_or3_4  _060_
timestamp 1586364061
transform 1 0 15548 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__048__B
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_3  FILLER_2_154
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use scs8hd_buf_2  _143_
timestamp 1586364061
transform 1 0 17112 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__058__B
timestamp 1586364061
transform 1 0 16560 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_166
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_170
timestamp 1586364061
transform 1 0 16744 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_178
timestamp 1586364061
transform 1 0 17480 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18400 0 -1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__054__C
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17664 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_182
timestamp 1586364061
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_186
timestamp 1586364061
transform 1 0 18216 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20148 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_199
timestamp 1586364061
transform 1 0 19412 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_205
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_209
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_213
timestamp 1586364061
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_218
timestamp 1586364061
transform 1 0 21160 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_2_230
timestamp 1586364061
transform 1 0 22264 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 22816 0 -1 3808
box -38 -48 314 592
use scs8hd_nor2_4  _065_
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_23
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4876 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_38
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_43
timestamp 1586364061
transform 1 0 5060 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_47
timestamp 1586364061
transform 1 0 5428 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_52
timestamp 1586364061
transform 1 0 5888 0 1 3808
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_nor2_4  _068_
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_73
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_77
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_90
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_99
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 314 592
use scs8hd_buf_2  _144_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11684 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_113
timestamp 1586364061
transform 1 0 11500 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_117
timestamp 1586364061
transform 1 0 11868 0 1 3808
box -38 -48 314 592
use scs8hd_nor4_4  _107_
timestamp 1586364061
transform 1 0 13524 0 1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__107__D
timestamp 1586364061
transform 1 0 13340 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 12972 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_127
timestamp 1586364061
transform 1 0 12788 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_131
timestamp 1586364061
transform 1 0 13156 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__042__A
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__C
timestamp 1586364061
transform 1 0 15272 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_152
timestamp 1586364061
transform 1 0 15088 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_160
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use scs8hd_inv_8  _042_
timestamp 1586364061
transform 1 0 16192 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_173
timestamp 1586364061
transform 1 0 17020 0 1 3808
box -38 -48 406 592
use scs8hd_inv_8  _041_
timestamp 1586364061
transform 1 0 18492 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 18216 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__041__A
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_179
timestamp 1586364061
transform 1 0 17572 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_188
timestamp 1586364061
transform 1 0 18400 0 1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20056 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19872 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_198
timestamp 1586364061
transform 1 0 19320 0 1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_215
timestamp 1586364061
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_219
timestamp 1586364061
transform 1 0 21252 0 1 3808
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_3_231
timestamp 1586364061
transform 1 0 22356 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 22816 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_19
timestamp 1586364061
transform 1 0 2852 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_29
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_32 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_40
timestamp 1586364061
transform 1 0 4784 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_50
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6716 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_54
timestamp 1586364061
transform 1 0 6072 0 -1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_4_60
timestamp 1586364061
transform 1 0 6624 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 7912 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_72
timestamp 1586364061
transform 1 0 7728 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_76
timestamp 1586364061
transform 1 0 8096 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_6  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_104
timestamp 1586364061
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11408 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__049__A
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_108
timestamp 1586364061
transform 1 0 11040 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_121
timestamp 1586364061
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_8  _045_
timestamp 1586364061
transform 1 0 12972 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__107__C
timestamp 1586364061
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__B
timestamp 1586364061
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_125
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_138
timestamp 1586364061
transform 1 0 13800 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_142
timestamp 1586364061
transform 1 0 14168 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__044__A
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_147
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_4  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_160
timestamp 1586364061
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use scs8hd_or3_4  _058_
timestamp 1586364061
transform 1 0 16192 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__056__B
timestamp 1586364061
transform 1 0 16008 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_173
timestamp 1586364061
transform 1 0 17020 0 -1 4896
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_181
timestamp 1586364061
transform 1 0 17756 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20516 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_197
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_205
timestamp 1586364061
transform 1 0 19964 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_4_208
timestamp 1586364061
transform 1 0 20240 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_4_213
timestamp 1586364061
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_12  FILLER_4_218
timestamp 1586364061
transform 1 0 21160 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_4_230
timestamp 1586364061
transform 1 0 22264 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 22816 0 -1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__067__B
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_6
timestamp 1586364061
transform 1 0 1656 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_10
timestamp 1586364061
transform 1 0 2024 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_14
timestamp 1586364061
transform 1 0 2392 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_17
timestamp 1586364061
transform 1 0 2668 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _067_
timestamp 1586364061
transform 1 0 3036 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_30
timestamp 1586364061
transform 1 0 3864 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_34
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4692 0 1 4896
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__B
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5520 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_38
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_42
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_46
timestamp 1586364061
transform 1 0 5336 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_71
timestamp 1586364061
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _097_
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__B
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_75
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_88
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_92
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_95
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use scs8hd_nand3_4  _049_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1326 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__C
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__B
timestamp 1586364061
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_108
timestamp 1586364061
transform 1 0 11040 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_112
timestamp 1586364061
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_116
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__105__C
timestamp 1586364061
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_137
timestamp 1586364061
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_141
timestamp 1586364061
transform 1 0 14076 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _044_
timestamp 1586364061
transform 1 0 14444 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__056__C
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__B
timestamp 1586364061
transform 1 0 14260 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_154
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_158
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_or3_4  _056_
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__056__A
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_171
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_175
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _087_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20516 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20332 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_197
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21528 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_220
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_5_224
timestamp 1586364061
transform 1 0 21712 0 1 4896
box -38 -48 774 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 22816 0 1 4896
box -38 -48 314 592
use scs8hd_fill_1  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2576 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_6_15
timestamp 1586364061
transform 1 0 2484 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_20
timestamp 1586364061
transform 1 0 2944 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2760 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_33
timestamp 1586364061
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_29
timestamp 1586364061
transform 1 0 3772 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_28
timestamp 1586364061
transform 1 0 3680 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2760 0 1 5984
box -38 -48 1050 592
use scs8hd_nor2_4  _066_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4508 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_45
timestamp 1586364061
transform 1 0 5244 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_48
timestamp 1586364061
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_52
timestamp 1586364061
transform 1 0 5888 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_60
timestamp 1586364061
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_60
timestamp 1586364061
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6440 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_71
timestamp 1586364061
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_68
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_64
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 7544 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use scs8hd_nor2_4  _096_
timestamp 1586364061
transform 1 0 7728 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8464 0 1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8280 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_81
timestamp 1586364061
transform 1 0 8556 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_85
timestamp 1586364061
transform 1 0 8924 0 -1 5984
box -38 -48 590 592
use scs8hd_decap_3  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_95
timestamp 1586364061
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_91
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_91
timestamp 1586364061
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_104
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_108
timestamp 1586364061
transform 1 0 11040 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_6_108
timestamp 1586364061
transform 1 0 11040 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__062__C
timestamp 1586364061
transform 1 0 11408 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_123
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_or4_4  _091_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12512 0 1 5984
box -38 -48 866 592
use scs8hd_or3_4  _062_
timestamp 1586364061
transform 1 0 11592 0 -1 5984
box -38 -48 866 592
use scs8hd_or2_4  _083_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14076 0 1 5984
box -38 -48 682 592
use scs8hd_or3_4  _105_
timestamp 1586364061
transform 1 0 13340 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 13156 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__C
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_127
timestamp 1586364061
transform 1 0 12788 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_142
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_133
timestamp 1586364061
transform 1 0 13340 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_148
timestamp 1586364061
transform 1 0 14720 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_146
timestamp 1586364061
transform 1 0 14536 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_156
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_152
timestamp 1586364061
transform 1 0 15088 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_159
timestamp 1586364061
transform 1 0 15732 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_152
timestamp 1586364061
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 15548 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_nor2_4  _085_
timestamp 1586364061
transform 1 0 15548 0 1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_5_.latch
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 15916 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_174
timestamp 1586364061
transform 1 0 17112 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_166
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_170
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_184
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 18216 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_6_195
timestamp 1586364061
transform 1 0 19044 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_191
timestamp 1586364061
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18860 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17848 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_4_.latch
timestamp 1586364061
transform 1 0 18400 0 1 5984
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_7_199
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 774 592
use scs8hd_decap_8  FILLER_6_202
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 774 592
use scs8hd_conb_1  _137_
timestamp 1586364061
transform 1 0 19412 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_7_207
timestamp 1586364061
transform 1 0 20148 0 1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_213
timestamp 1586364061
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_210
timestamp 1586364061
transform 1 0 20424 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__040__A
timestamp 1586364061
transform 1 0 20240 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_inv_8  _040_
timestamp 1586364061
transform 1 0 20424 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_224
timestamp 1586364061
transform 1 0 21712 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_219
timestamp 1586364061
transform 1 0 21252 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_7_223
timestamp 1586364061
transform 1 0 21620 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_231
timestamp 1586364061
transform 1 0 22356 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 22816 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 22816 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_232
timestamp 1586364061
transform 1 0 22448 0 -1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 2944 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2760 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_6  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4692 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_38
timestamp 1586364061
transform 1 0 4600 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_50
timestamp 1586364061
transform 1 0 5704 0 -1 7072
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_61
timestamp 1586364061
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_65
timestamp 1586364061
transform 1 0 7084 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_69
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 7728 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_8  FILLER_8_81
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_89
timestamp 1586364061
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10212 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10028 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_93
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11776 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__091__D
timestamp 1586364061
transform 1 0 12512 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_108
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_4  FILLER_8_119
timestamp 1586364061
transform 1 0 12052 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_123
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 130 592
use scs8hd_nor2_4  _089_
timestamp 1586364061
transform 1 0 13616 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 13248 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__C
timestamp 1586364061
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_126
timestamp 1586364061
transform 1 0 12696 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_130
timestamp 1586364061
transform 1 0 13064 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_134
timestamp 1586364061
transform 1 0 13432 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_149
timestamp 1586364061
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17020 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16468 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_165
timestamp 1586364061
transform 1 0 16284 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_169
timestamp 1586364061
transform 1 0 16652 0 -1 7072
box -38 -48 406 592
use scs8hd_decap_8  FILLER_8_176
timestamp 1586364061
transform 1 0 17296 0 -1 7072
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18308 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_8_184
timestamp 1586364061
transform 1 0 18032 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19504 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_198
timestamp 1586364061
transform 1 0 19320 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_218
timestamp 1586364061
transform 1 0 21160 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_8_230
timestamp 1586364061
transform 1 0 22264 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 22816 0 -1 7072
box -38 -48 314 592
use scs8hd_conb_1  _132_
timestamp 1586364061
transform 1 0 2024 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 2484 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_3
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 590 592
use scs8hd_fill_1  FILLER_9_9
timestamp 1586364061
transform 1 0 1932 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_13
timestamp 1586364061
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_17
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3680 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 3496 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_21
timestamp 1586364061
transform 1 0 3036 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_25
timestamp 1586364061
transform 1 0 3404 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_31
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5796 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_48
timestamp 1586364061
transform 1 0 5520 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 406 592
use scs8hd_decap_4  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_66
timestamp 1586364061
transform 1 0 7176 0 1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_6.LATCH_2_.latch
timestamp 1586364061
transform 1 0 8464 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7912 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_72
timestamp 1586364061
transform 1 0 7728 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_76
timestamp 1586364061
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10672 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_91
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_95
timestamp 1586364061
transform 1 0 9844 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_98
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__D
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_113
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_117
timestamp 1586364061
transform 1 0 11868 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_123
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use scs8hd_or4_4  _084_
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__098__B
timestamp 1586364061
transform 1 0 12604 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 13064 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_127
timestamp 1586364061
transform 1 0 12788 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_141
timestamp 1586364061
transform 1 0 14076 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14996 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14260 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_145
timestamp 1586364061
transform 1 0 14444 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_154
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_158
timestamp 1586364061
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__086__B
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_171
timestamp 1586364061
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18492 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_184
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_188
timestamp 1586364061
transform 1 0 18400 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_191
timestamp 1586364061
transform 1 0 18676 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _130_
timestamp 1586364061
transform 1 0 20792 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_204
timestamp 1586364061
transform 1 0 19872 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_217
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_9_229
timestamp 1586364061
transform 1 0 22172 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 22816 0 1 7072
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 1050 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_3
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _125_
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_21
timestamp 1586364061
transform 1 0 3036 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_29
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5796 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_45
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_49
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 7544 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7084 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_60
timestamp 1586364061
transform 1 0 6624 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_64
timestamp 1586364061
transform 1 0 6992 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_67
timestamp 1586364061
transform 1 0 7268 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_6.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8556 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_79
timestamp 1586364061
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_83
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_89
timestamp 1586364061
transform 1 0 9292 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9936 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10396 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_99
timestamp 1586364061
transform 1 0 10212 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_103
timestamp 1586364061
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_107
timestamp 1586364061
transform 1 0 10948 0 -1 8160
box -38 -48 130 592
use scs8hd_or4_4  _098_
timestamp 1586364061
transform 1 0 12512 0 -1 8160
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_6.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11040 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 12328 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__C
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_111
timestamp 1586364061
transform 1 0 11316 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_3  FILLER_10_119
timestamp 1586364061
transform 1 0 12052 0 -1 8160
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__084__D
timestamp 1586364061
transform 1 0 13524 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__C
timestamp 1586364061
transform 1 0 13892 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_133
timestamp 1586364061
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_137
timestamp 1586364061
transform 1 0 13708 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_141
timestamp 1586364061
transform 1 0 14076 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 14720 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15456 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  FILLER_10_150
timestamp 1586364061
transform 1 0 14904 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _086_
timestamp 1586364061
transform 1 0 17388 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16652 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_167
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_171
timestamp 1586364061
transform 1 0 16836 0 -1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18952 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18676 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_186
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_190
timestamp 1586364061
transform 1 0 18584 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_193
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_203
timestamp 1586364061
transform 1 0 19780 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  FILLER_10_211
timestamp 1586364061
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 22816 0 -1 8160
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_fill_2  FILLER_11_9
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4324 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 3772 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_22
timestamp 1586364061
transform 1 0 3128 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_26
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_31
timestamp 1586364061
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5888 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_46
timestamp 1586364061
transform 1 0 5336 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_50
timestamp 1586364061
transform 1 0 5704 0 1 8160
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_54
timestamp 1586364061
transform 1 0 6072 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_58
timestamp 1586364061
transform 1 0 6440 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_65
timestamp 1586364061
transform 1 0 7084 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_69
timestamp 1586364061
transform 1 0 7452 0 1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8280 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7728 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_74
timestamp 1586364061
transform 1 0 7912 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_89
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10028 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_95
timestamp 1586364061
transform 1 0 9844 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_106
timestamp 1586364061
transform 1 0 10856 0 1 8160
box -38 -48 222 592
use scs8hd_inv_8  _047_
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__047__A
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_110
timestamp 1586364061
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__046__A
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_11_136
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 774 592
use scs8hd_nor2_4  _090_
timestamp 1586364061
transform 1 0 14720 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__B
timestamp 1586364061
transform 1 0 14536 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_144
timestamp 1586364061
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_157
timestamp 1586364061
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16284 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_161
timestamp 1586364061
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_11_174
timestamp 1586364061
transform 1 0 17112 0 1 8160
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 18216 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_5.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_180
timestamp 1586364061
transform 1 0 17664 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_188
timestamp 1586364061
transform 1 0 18400 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19688 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_200
timestamp 1586364061
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_204
timestamp 1586364061
transform 1 0 19872 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_216
timestamp 1586364061
transform 1 0 20976 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_11_228
timestamp 1586364061
transform 1 0 22080 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 22816 0 1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 2300 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__077__B
timestamp 1586364061
transform 1 0 2116 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4324 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_22
timestamp 1586364061
transform 1 0 3128 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_30
timestamp 1586364061
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 5336 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4968 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_38
timestamp 1586364061
transform 1 0 4600 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7084 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 6900 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_57
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_61
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 8464 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_74
timestamp 1586364061
transform 1 0 7912 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_8  FILLER_12_82
timestamp 1586364061
transform 1 0 8648 0 -1 9248
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_90
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 1142 592
use scs8hd_or3_4  _076_
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__069__C
timestamp 1586364061
transform 1 0 11684 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_114
timestamp 1586364061
transform 1 0 11592 0 -1 9248
box -38 -48 130 592
use scs8hd_inv_8  _046_
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__050__B
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__050__C
timestamp 1586364061
transform 1 0 13248 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_126
timestamp 1586364061
transform 1 0 12696 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_130
timestamp 1586364061
transform 1 0 13064 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15364 0 -1 9248
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__108__B
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_143
timestamp 1586364061
transform 1 0 14260 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_147
timestamp 1586364061
transform 1 0 14628 0 -1 9248
box -38 -48 590 592
use scs8hd_fill_1  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16560 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_170
timestamp 1586364061
transform 1 0 16744 0 -1 9248
box -38 -48 1142 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_5.LATCH_2_.latch
timestamp 1586364061
transform 1 0 17940 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19136 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_182
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_12_194
timestamp 1586364061
transform 1 0 18952 0 -1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19504 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_198
timestamp 1586364061
transform 1 0 19320 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_205
timestamp 1586364061
transform 1 0 19964 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_213
timestamp 1586364061
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 590 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 22816 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_7
timestamp 1586364061
transform 1 0 1748 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 1840 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_13_10
timestamp 1586364061
transform 1 0 2024 0 1 9248
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_5_.latch
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 1050 592
use scs8hd_nor2_4  _077_
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_19
timestamp 1586364061
transform 1 0 2852 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_24
timestamp 1586364061
transform 1 0 3312 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_20
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_29
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_28
timestamp 1586364061
transform 1 0 3680 0 1 9248
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_40
timestamp 1586364061
transform 1 0 4784 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_36
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 4600 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__B
timestamp 1586364061
transform 1 0 4416 0 1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_14_53
timestamp 1586364061
transform 1 0 5980 0 -1 10336
box -38 -48 774 592
use scs8hd_decap_4  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_47
timestamp 1586364061
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4968 0 -1 10336
box -38 -48 1050 592
use scs8hd_nor2_4  _124_
timestamp 1586364061
transform 1 0 4600 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _126_
timestamp 1586364061
transform 1 0 6900 0 1 9248
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6716 0 -1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_14_70
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 8464 0 1 9248
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8280 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_72
timestamp 1586364061
transform 1 0 7728 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_76
timestamp 1586364061
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_78
timestamp 1586364061
transform 1 0 8280 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_95
timestamp 1586364061
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_91
timestamp 1586364061
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_106
timestamp 1586364061
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_102
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10672 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_114
timestamp 1586364061
transform 1 0 11592 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_113
timestamp 1586364061
transform 1 0 11500 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_120
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_117
timestamp 1586364061
transform 1 0 11868 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 11776 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__069__B
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_or3_4  _069_
timestamp 1586364061
transform 1 0 11960 0 -1 10336
box -38 -48 866 592
use scs8hd_or3_4  _050_
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_or3_4  _108_
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 866 592
use scs8hd_or3_4  _115_
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__115__B
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__050__A
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_138
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_127
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_131
timestamp 1586364061
transform 1 0 13156 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_145
timestamp 1586364061
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__C
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_149
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_149
timestamp 1586364061
transform 1 0 14812 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 14996 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_13_157
timestamp 1586364061
transform 1 0 15548 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_153
timestamp 1586364061
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 15548 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__C
timestamp 1586364061
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_159
timestamp 1586364061
transform 1 0 15732 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__B
timestamp 1586364061
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _088_
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16008 0 1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 17020 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15916 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_175
timestamp 1586364061
transform 1 0 17204 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_172
timestamp 1586364061
transform 1 0 16928 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_182
timestamp 1586364061
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_179
timestamp 1586364061
transform 1 0 17572 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 18216 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__113__B
timestamp 1586364061
transform 1 0 17664 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_193
timestamp 1586364061
transform 1 0 18860 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_189
timestamp 1586364061
transform 1 0 18492 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_188
timestamp 1586364061
transform 1 0 18400 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18676 0 -1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_5.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 1 9248
box -38 -48 866 592
use scs8hd_nor2_4  _113_
timestamp 1586364061
transform 1 0 17664 0 -1 10336
box -38 -48 866 592
use scs8hd_decap_8  FILLER_14_204
timestamp 1586364061
transform 1 0 19872 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_2  FILLER_14_200
timestamp 1586364061
transform 1 0 19504 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_8  FILLER_13_204
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_13_200
timestamp 1586364061
transform 1 0 19504 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19688 0 1 9248
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19228 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_212
timestamp 1586364061
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_212
timestamp 1586364061
transform 1 0 20608 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_buf_2  _148_
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_217
timestamp 1586364061
transform 1 0 21068 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_13_229
timestamp 1586364061
transform 1 0 22172 0 1 9248
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_219
timestamp 1586364061
transform 1 0 21252 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_231
timestamp 1586364061
transform 1 0 22356 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 22816 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 22816 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1840 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1656 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_17
timestamp 1586364061
transform 1 0 2668 0 1 10336
box -38 -48 774 592
use scs8hd_nor2_4  _078_
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _127_
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__B
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_36
timestamp 1586364061
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_40
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8372 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_75
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_82
timestamp 1586364061
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9568 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__B
timestamp 1586364061
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_90
timestamp 1586364061
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_101
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_105
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_109
timestamp 1586364061
transform 1 0 11132 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_113
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_117
timestamp 1586364061
transform 1 0 11868 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use scs8hd_or3_4  _122_
timestamp 1586364061
transform 1 0 12972 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__122__C
timestamp 1586364061
transform 1 0 12788 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_138
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_142
timestamp 1586364061
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _114_
timestamp 1586364061
transform 1 0 15548 0 1 10336
box -38 -48 866 592
use scs8hd_inv_1  mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14536 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_5.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_149
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_153
timestamp 1586364061
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16560 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16928 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_166
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_170
timestamp 1586364061
transform 1 0 16744 0 1 10336
box -38 -48 222 592
use scs8hd_decap_6  FILLER_15_174
timestamp 1586364061
transform 1 0 17112 0 1 10336
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_180
timestamp 1586364061
transform 1 0 17664 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_193
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19596 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_197
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_210
timestamp 1586364061
transform 1 0 20424 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_214
timestamp 1586364061
transform 1 0 20792 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_217
timestamp 1586364061
transform 1 0 21068 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_15_229
timestamp 1586364061
transform 1 0 22172 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 22816 0 1 10336
box -38 -48 314 592
use scs8hd_conb_1  _136_
timestamp 1586364061
transform 1 0 2392 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_4.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_6
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_10
timestamp 1586364061
transform 1 0 2024 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_4  FILLER_16_17
timestamp 1586364061
transform 1 0 2668 0 -1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3128 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_21
timestamp 1586364061
transform 1 0 3036 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_24
timestamp 1586364061
transform 1 0 3312 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_28
timestamp 1586364061
transform 1 0 3680 0 -1 11424
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5796 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_43
timestamp 1586364061
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_47
timestamp 1586364061
transform 1 0 5428 0 -1 11424
box -38 -48 406 592
use scs8hd_nor2_4  _082_
timestamp 1586364061
transform 1 0 6992 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_54
timestamp 1586364061
transform 1 0 6072 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_73
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_77
timestamp 1586364061
transform 1 0 8188 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_8  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 774 592
use scs8hd_nor2_4  _061_
timestamp 1586364061
transform 1 0 10396 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_97
timestamp 1586364061
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__B
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_110
timestamp 1586364061
transform 1 0 11224 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_16_122
timestamp 1586364061
transform 1 0 12328 0 -1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _059_
timestamp 1586364061
transform 1 0 12696 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_135
timestamp 1586364061
transform 1 0 13524 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_139
timestamp 1586364061
transform 1 0 13892 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_143
timestamp 1586364061
transform 1 0 14260 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_16_151
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_16_162
timestamp 1586364061
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_174
timestamp 1586364061
transform 1 0 17112 0 -1 11424
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18676 0 -1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_182
timestamp 1586364061
transform 1 0 17848 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19872 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_218
timestamp 1586364061
transform 1 0 21160 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_16_230
timestamp 1586364061
transform 1 0 22264 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 22816 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 2024 0 1 11424
box -38 -48 222 592
use scs8hd_decap_6  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_9
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_12
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_16
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_3_.latch
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4324 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_33
timestamp 1586364061
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_37
timestamp 1586364061
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_50
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7636 0 1 11424
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 6256 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_54
timestamp 1586364061
transform 1 0 6072 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_58
timestamp 1586364061
transform 1 0 6440 0 1 11424
box -38 -48 314 592
use scs8hd_decap_6  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 590 592
use scs8hd_fill_1  FILLER_17_68
timestamp 1586364061
transform 1 0 7360 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8832 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_82
timestamp 1586364061
transform 1 0 8648 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10580 0 1 11424
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9384 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_93
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_97
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_101
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_118
timestamp 1586364061
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_126
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_130
timestamp 1586364061
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15364 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15180 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_145
timestamp 1586364061
transform 1 0 14444 0 1 11424
box -38 -48 774 592
use scs8hd_fill_2  FILLER_17_158
timestamp 1586364061
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_162
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_175
timestamp 1586364061
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18952 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_179
timestamp 1586364061
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_187
timestamp 1586364061
transform 1 0 18308 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_191
timestamp 1586364061
transform 1 0 18676 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19504 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19320 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_209
timestamp 1586364061
transform 1 0 20332 0 1 11424
box -38 -48 774 592
use scs8hd_buf_2  _142_
timestamp 1586364061
transform 1 0 21068 0 1 11424
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 21620 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_221
timestamp 1586364061
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use scs8hd_decap_8  FILLER_17_225
timestamp 1586364061
transform 1 0 21804 0 1 11424
box -38 -48 774 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 22816 0 1 11424
box -38 -48 314 592
use scs8hd_nor2_4  _079_
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_11
timestamp 1586364061
transform 1 0 2116 0 -1 12512
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4324 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_3  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 314 592
use scs8hd_nor2_4  _081_
timestamp 1586364061
transform 1 0 5888 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_48
timestamp 1586364061
transform 1 0 5520 0 -1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_61
timestamp 1586364061
transform 1 0 6716 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_18_69
timestamp 1586364061
transform 1 0 7452 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_73
timestamp 1586364061
transform 1 0 7820 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_84
timestamp 1586364061
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_88
timestamp 1586364061
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10580 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__053__B
timestamp 1586364061
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_96
timestamp 1586364061
transform 1 0 9936 0 -1 12512
box -38 -48 590 592
use scs8hd_fill_1  FILLER_18_102
timestamp 1586364061
transform 1 0 10488 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11592 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11316 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_109
timestamp 1586364061
transform 1 0 11132 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_113
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_6  FILLER_18_123
timestamp 1586364061
transform 1 0 12420 0 -1 12512
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13432 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_131
timestamp 1586364061
transform 1 0 13156 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 774 592
use scs8hd_decap_8  FILLER_18_157
timestamp 1586364061
transform 1 0 15548 0 -1 12512
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_165
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_168
timestamp 1586364061
transform 1 0 16560 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_172
timestamp 1586364061
transform 1 0 16928 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 19044 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_182
timestamp 1586364061
transform 1 0 17848 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_194
timestamp 1586364061
transform 1 0 18952 0 -1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19320 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19780 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_197
timestamp 1586364061
transform 1 0 19228 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_201
timestamp 1586364061
transform 1 0 19596 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_18_205
timestamp 1586364061
transform 1 0 19964 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_213
timestamp 1586364061
transform 1 0 20700 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21068 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_18_219
timestamp 1586364061
transform 1 0 21252 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_18_231
timestamp 1586364061
transform 1 0 22356 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 22816 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_6  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_13
timestamp 1586364061
transform 1 0 2300 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_16
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_11
timestamp 1586364061
transform 1 0 2116 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__080__B
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use scs8hd_nor2_4  _080_
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use scs8hd_decap_8  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_19_20
timestamp 1586364061
transform 1 0 2944 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3404 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_32
timestamp 1586364061
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_28
timestamp 1586364061
transform 1 0 3680 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 4232 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3864 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_2_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4416 0 1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5428 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_45
timestamp 1586364061
transform 1 0 5244 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_49
timestamp 1586364061
transform 1 0 5612 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_43
timestamp 1586364061
transform 1 0 5060 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_47
timestamp 1586364061
transform 1 0 5428 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  FILLER_20_55
timestamp 1586364061
transform 1 0 6164 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_19_60
timestamp 1586364061
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_56
timestamp 1586364061
transform 1 0 6256 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_4.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6440 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_69
timestamp 1586364061
transform 1 0 7452 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_4.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6440 0 -1 13600
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_20_80
timestamp 1586364061
transform 1 0 8464 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_73
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_77
timestamp 1586364061
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8188 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_81
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 8924 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_97
timestamp 1586364061
transform 1 0 10028 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_91
timestamp 1586364061
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_94
timestamp 1586364061
transform 1 0 9752 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9844 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_101
timestamp 1586364061
transform 1 0 10396 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__053__A
timestamp 1586364061
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10212 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10212 0 -1 13600
box -38 -48 314 592
use scs8hd_nor2_4  _053_
timestamp 1586364061
transform 1 0 10672 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_113
timestamp 1586364061
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_121
timestamp 1586364061
transform 1 0 12236 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_117
timestamp 1586364061
transform 1 0 11868 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 11224 0 -1 13600
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_142
timestamp 1586364061
transform 1 0 14168 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_138
timestamp 1586364061
transform 1 0 13800 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_136
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 13984 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 866 592
use scs8hd_decap_6  FILLER_20_146
timestamp 1586364061
transform 1 0 14536 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_149
timestamp 1586364061
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_152
timestamp 1586364061
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_6  FILLER_19_153
timestamp 1586364061
transform 1 0 15180 0 1 12512
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_158
timestamp 1586364061
transform 1 0 15640 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15824 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_20_162
timestamp 1586364061
transform 1 0 16008 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_165
timestamp 1586364061
transform 1 0 16284 0 1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_161
timestamp 1586364061
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 16100 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_178
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_20_174
timestamp 1586364061
transform 1 0 17112 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 17296 0 -1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 12512
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_20_186
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_187
timestamp 1586364061
transform 1 0 18308 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_194
timestamp 1586364061
transform 1 0 18952 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_191
timestamp 1586364061
transform 1 0 18676 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 12512
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 19044 0 -1 13600
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20700 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_206
timestamp 1586364061
transform 1 0 20056 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_210
timestamp 1586364061
transform 1 0 20424 0 1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 774 592
use scs8hd_buf_2  _140_
timestamp 1586364061
transform 1 0 20884 0 1 12512
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 21436 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_219
timestamp 1586364061
transform 1 0 21252 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_19_223
timestamp 1586364061
transform 1 0 21620 0 1 12512
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_231
timestamp 1586364061
transform 1 0 22356 0 1 12512
box -38 -48 222 592
use scs8hd_decap_8  FILLER_20_224
timestamp 1586364061
transform 1 0 21712 0 -1 13600
box -38 -48 774 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 22816 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 22816 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_232
timestamp 1586364061
transform 1 0 22448 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_2  _141_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_11
timestamp 1586364061
transform 1 0 2116 0 1 13600
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4140 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3220 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_25
timestamp 1586364061
transform 1 0 3404 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_29
timestamp 1586364061
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__B
timestamp 1586364061
transform 1 0 5244 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 5612 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_42
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_47
timestamp 1586364061
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use scs8hd_decap_8  FILLER_21_51
timestamp 1586364061
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6992 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_66
timestamp 1586364061
transform 1 0 7176 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _073_
timestamp 1586364061
transform 1 0 8924 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__B
timestamp 1586364061
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_77
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_81
timestamp 1586364061
transform 1 0 8556 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _055_
timestamp 1586364061
transform 1 0 10580 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 9936 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__A
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_94
timestamp 1586364061
transform 1 0 9752 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_98
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_112
timestamp 1586364061
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_116
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_120
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12604 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13064 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_128
timestamp 1586364061
transform 1 0 12880 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_132
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 15180 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__B
timestamp 1586364061
transform 1 0 14812 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_147
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_151
timestamp 1586364061
transform 1 0 14996 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 16376 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_164
timestamp 1586364061
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_168
timestamp 1586364061
transform 1 0 16560 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _110_
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__111__B
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_193
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20056 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19872 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_197
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_201
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 21068 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_215
timestamp 1586364061
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_219
timestamp 1586364061
transform 1 0 21252 0 1 13600
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_21_231
timestamp 1586364061
transform 1 0 22356 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 22816 0 1 13600
box -38 -48 314 592
use scs8hd_buf_2  _153_
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_19
timestamp 1586364061
transform 1 0 2852 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_22_35
timestamp 1586364061
transform 1 0 4324 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _102_
timestamp 1586364061
transform 1 0 5244 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_39
timestamp 1586364061
transform 1 0 4692 0 -1 14688
box -38 -48 590 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_22_54
timestamp 1586364061
transform 1 0 6072 0 -1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_22_65
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  FILLER_22_70
timestamp 1586364061
transform 1 0 7544 0 -1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_4.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_22_76
timestamp 1586364061
transform 1 0 8096 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_2_.latch
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__055__B
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_104
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 1050 592
use scs8hd_decap_4  FILLER_22_108
timestamp 1586364061
transform 1 0 11040 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_8  FILLER_22_123
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _057_
timestamp 1586364061
transform 1 0 13156 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_140
timestamp 1586364061
transform 1 0 13984 0 -1 14688
box -38 -48 222 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 15548 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_144
timestamp 1586364061
transform 1 0 14352 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_148
timestamp 1586364061
transform 1 0 14720 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_152
timestamp 1586364061
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 17112 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 774 592
use scs8hd_nor2_4  _111_
timestamp 1586364061
transform 1 0 18676 0 -1 14688
box -38 -48 866 592
use scs8hd_decap_8  FILLER_22_183
timestamp 1586364061
transform 1 0 17940 0 -1 14688
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_200
timestamp 1586364061
transform 1 0 19504 0 -1 14688
box -38 -48 590 592
use scs8hd_decap_4  FILLER_22_208
timestamp 1586364061
transform 1 0 20240 0 -1 14688
box -38 -48 406 592
use scs8hd_buf_2  _150_
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_22_219
timestamp 1586364061
transform 1 0 21252 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_22_231
timestamp 1586364061
transform 1 0 22356 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 22816 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use scs8hd_decap_8  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  FILLER_23_11
timestamp 1586364061
transform 1 0 2116 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_16
timestamp 1586364061
transform 1 0 2576 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3312 0 1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4324 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 4140 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 2760 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3128 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_20
timestamp 1586364061
transform 1 0 2944 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_31
timestamp 1586364061
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5336 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_44
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_48
timestamp 1586364061
transform 1 0 5520 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_71
timestamp 1586364061
transform 1 0 7636 0 1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8832 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9292 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_76
timestamp 1586364061
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_80
timestamp 1586364061
transform 1 0 8464 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_87
timestamp 1586364061
transform 1 0 9108 0 1 14688
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10856 0 1 14688
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9844 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10304 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_91
timestamp 1586364061
transform 1 0 9476 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_98
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_102
timestamp 1586364061
transform 1 0 10488 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_109
timestamp 1586364061
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_113
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_118
timestamp 1586364061
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 13616 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 13984 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_132
timestamp 1586364061
transform 1 0 13248 0 1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_23_138
timestamp 1586364061
transform 1 0 13800 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_151
timestamp 1586364061
transform 1 0 14996 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_156
timestamp 1586364061
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_160
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 406 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 16376 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 16192 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18676 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18308 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_189
timestamp 1586364061
transform 1 0 18492 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 20608 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20424 0 1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_23_204
timestamp 1586364061
transform 1 0 19872 0 1 14688
box -38 -48 590 592
use scs8hd_decap_12  FILLER_23_221
timestamp 1586364061
transform 1 0 21436 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 22816 0 1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_3  FILLER_24_11
timestamp 1586364061
transform 1 0 2116 0 -1 15776
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_2_.latch
timestamp 1586364061
transform 1 0 5796 0 -1 15776
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_24_43
timestamp 1586364061
transform 1 0 5060 0 -1 15776
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_62
timestamp 1586364061
transform 1 0 6808 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_66
timestamp 1586364061
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_70
timestamp 1586364061
transform 1 0 7544 0 -1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _074_
timestamp 1586364061
transform 1 0 7912 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8924 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_83
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_87
timestamp 1586364061
transform 1 0 9108 0 -1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9936 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_91
timestamp 1586364061
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_24_107
timestamp 1586364061
transform 1 0 10948 0 -1 15776
box -38 -48 222 592
use scs8hd_conb_1  _133_
timestamp 1586364061
transform 1 0 12420 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_111
timestamp 1586364061
transform 1 0 11316 0 -1 15776
box -38 -48 1142 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__051__B
timestamp 1586364061
transform 1 0 12880 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_126
timestamp 1586364061
transform 1 0 12696 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_24_130
timestamp 1586364061
transform 1 0 13064 0 -1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_151
timestamp 1586364061
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 17296 0 -1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_24_163
timestamp 1586364061
transform 1 0 16100 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_168
timestamp 1586364061
transform 1 0 16560 0 -1 15776
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 18860 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18492 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_187
timestamp 1586364061
transform 1 0 18308 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_191
timestamp 1586364061
transform 1 0 18676 0 -1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_198
timestamp 1586364061
transform 1 0 19320 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_24_210
timestamp 1586364061
transform 1 0 20424 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 590 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 22816 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 590 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3312 0 1 15776
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3772 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__B
timestamp 1586364061
transform 1 0 4140 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 3128 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_21
timestamp 1586364061
transform 1 0 3036 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_31
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5336 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_44
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_48
timestamp 1586364061
transform 1 0 5520 0 1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6440 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6072 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_56
timestamp 1586364061
transform 1 0 6256 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_60
timestamp 1586364061
transform 1 0 6624 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_71
timestamp 1586364061
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8372 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_75
timestamp 1586364061
transform 1 0 8004 0 1 15776
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_92
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _051_
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__051__A
timestamp 1586364061
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use scs8hd_decap_3  FILLER_25_109
timestamp 1586364061
transform 1 0 11132 0 1 15776
box -38 -48 314 592
use scs8hd_fill_2  FILLER_25_114
timestamp 1586364061
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_118
timestamp 1586364061
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14076 0 1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_25_132
timestamp 1586364061
transform 1 0 13248 0 1 15776
box -38 -48 774 592
use scs8hd_fill_1  FILLER_25_140
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 14812 0 1 15776
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_143
timestamp 1586364061
transform 1 0 14260 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_160
timestamp 1586364061
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16928 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_164
timestamp 1586364061
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_168
timestamp 1586364061
transform 1 0 16560 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_175
timestamp 1586364061
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_179
timestamp 1586364061
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_193
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use scs8hd_conb_1  _129_
timestamp 1586364061
transform 1 0 19964 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_197
timestamp 1586364061
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_201
timestamp 1586364061
transform 1 0 19596 0 1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_220
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 22816 0 1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  FILLER_27_11
timestamp 1586364061
transform 1 0 2116 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_16
timestamp 1586364061
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_24
timestamp 1586364061
transform 1 0 3312 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_20
timestamp 1586364061
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3128 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_28
timestamp 1586364061
transform 1 0 3680 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_4_.latch
timestamp 1586364061
transform 1 0 4048 0 1 16864
box -38 -48 1050 592
use scs8hd_nor2_4  _100_
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5244 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_45
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_43
timestamp 1586364061
transform 1 0 5060 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_47
timestamp 1586364061
transform 1 0 5428 0 1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_60
timestamp 1586364061
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_56
timestamp 1586364061
transform 1 0 6256 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_61
timestamp 1586364061
transform 1 0 6716 0 -1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_57
timestamp 1586364061
transform 1 0 6348 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6072 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6440 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6440 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_26_66
timestamp 1586364061
transform 1 0 7176 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6992 0 -1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7452 0 -1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6992 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_79
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_73
timestamp 1586364061
transform 1 0 7820 0 1 16864
box -38 -48 406 592
use scs8hd_fill_1  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_26_72
timestamp 1586364061
transform 1 0 7728 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_88
timestamp 1586364061
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_84
timestamp 1586364061
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9200 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 16864
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_90
timestamp 1586364061
transform 1 0 9384 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_107
timestamp 1586364061
transform 1 0 10948 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_103
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10948 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9936 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9752 0 1 16864
box -38 -48 866 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_115
timestamp 1586364061
transform 1 0 11684 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_26_109
timestamp 1586364061
transform 1 0 11132 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11132 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_118
timestamp 1586364061
transform 1 0 11960 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 11776 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__B
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 12328 0 -1 16864
box -38 -48 1050 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 13708 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 14076 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_133
timestamp 1586364061
transform 1 0 13340 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_139
timestamp 1586364061
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_150
timestamp 1586364061
transform 1 0 14904 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_146
timestamp 1586364061
transform 1 0 14536 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_150
timestamp 1586364061
transform 1 0 14904 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_26_144
timestamp 1586364061
transform 1 0 14352 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14720 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14260 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15456 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16468 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_167
timestamp 1586364061
transform 1 0 16468 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_165
timestamp 1586364061
transform 1 0 16284 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_169
timestamp 1586364061
transform 1 0 16652 0 1 16864
box -38 -48 406 592
use scs8hd_decap_6  FILLER_27_175
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_179
timestamp 1586364061
transform 1 0 17572 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 18216 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_188
timestamp 1586364061
transform 1 0 18400 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_194
timestamp 1586364061
transform 1 0 18952 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19136 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18584 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18768 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18124 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 20700 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_198
timestamp 1586364061
transform 1 0 19320 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_26_210
timestamp 1586364061
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_27_201
timestamp 1586364061
transform 1 0 19596 0 1 16864
box -38 -48 1142 592
use scs8hd_buf_2  _155_
timestamp 1586364061
transform 1 0 20884 0 1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_27_219
timestamp 1586364061
transform 1 0 21252 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_27_223
timestamp 1586364061
transform 1 0 21620 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_231
timestamp 1586364061
transform 1 0 22356 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 22816 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 22816 0 1 16864
box -38 -48 314 592
use scs8hd_nor2_4  _101_
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_3  FILLER_28_11
timestamp 1586364061
transform 1 0 2116 0 -1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_3_.latch
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5612 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_43
timestamp 1586364061
transform 1 0 5060 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_47
timestamp 1586364061
transform 1 0 5428 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_51
timestamp 1586364061
transform 1 0 5796 0 -1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6440 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_55
timestamp 1586364061
transform 1 0 6164 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_69
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8188 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 8004 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_73
timestamp 1586364061
transform 1 0 7820 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_6  FILLER_28_86
timestamp 1586364061
transform 1 0 9016 0 -1 17952
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9844 0 -1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10856 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_104
timestamp 1586364061
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _071_
timestamp 1586364061
transform 1 0 11776 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11316 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_108
timestamp 1586364061
transform 1 0 11040 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_113
timestamp 1586364061
transform 1 0 11500 0 -1 17952
box -38 -48 314 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 13616 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13156 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_125
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_133
timestamp 1586364061
transform 1 0 13340 0 -1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14904 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_28_149
timestamp 1586364061
transform 1 0 14812 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_152
timestamp 1586364061
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17020 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_165
timestamp 1586364061
transform 1 0 16284 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_8  FILLER_28_176
timestamp 1586364061
transform 1 0 17296 0 -1 17952
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 18124 0 -1 17952
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_28_184
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_28_196
timestamp 1586364061
transform 1 0 19136 0 -1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 19780 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19320 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_200
timestamp 1586364061
transform 1 0 19504 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_205
timestamp 1586364061
transform 1 0 19964 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_1  FILLER_28_213
timestamp 1586364061
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use scs8hd_buf_2  _152_
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_219
timestamp 1586364061
transform 1 0 21252 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_28_231
timestamp 1586364061
transform 1 0 22356 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 22816 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 1564 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_7
timestamp 1586364061
transform 1 0 1748 0 1 17952
box -38 -48 1142 592
use scs8hd_nor2_4  _099_
timestamp 1586364061
transform 1 0 3312 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4324 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_19
timestamp 1586364061
transform 1 0 2852 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_33
timestamp 1586364061
transform 1 0 4140 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4876 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_37
timestamp 1586364061
transform 1 0 4508 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_50
timestamp 1586364061
transform 1 0 5704 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_55
timestamp 1586364061
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_71
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8832 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8648 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__075__B
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_77
timestamp 1586364061
transform 1 0 8188 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_81
timestamp 1586364061
transform 1 0 8556 0 1 17952
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_95
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_99
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_112
timestamp 1586364061
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_116
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_29_134
timestamp 1586364061
transform 1 0 13432 0 1 17952
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14904 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14720 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_146
timestamp 1586364061
transform 1 0 14536 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15916 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 16560 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_29_163
timestamp 1586364061
transform 1 0 16100 0 1 17952
box -38 -48 406 592
use scs8hd_fill_1  FILLER_29_167
timestamp 1586364061
transform 1 0 16468 0 1 17952
box -38 -48 130 592
use scs8hd_fill_2  FILLER_29_170
timestamp 1586364061
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_174
timestamp 1586364061
transform 1 0 17112 0 1 17952
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_179
timestamp 1586364061
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_195
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _117_
timestamp 1586364061
transform 1 0 19780 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__117__B
timestamp 1586364061
transform 1 0 19596 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_199
timestamp 1586364061
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_212
timestamp 1586364061
transform 1 0 20608 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_224
timestamp 1586364061
transform 1 0 21712 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 22816 0 1 17952
box -38 -48 314 592
use scs8hd_fill_1  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 130 592
use scs8hd_buf_2  _157_
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_7
timestamp 1586364061
transform 1 0 1748 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 3312 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_19
timestamp 1586364061
transform 1 0 2852 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_23
timestamp 1586364061
transform 1 0 3220 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_26
timestamp 1586364061
transform 1 0 3496 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_30
timestamp 1586364061
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4784 0 -1 19040
box -38 -48 866 592
use scs8hd_decap_8  FILLER_30_49
timestamp 1586364061
transform 1 0 5612 0 -1 19040
box -38 -48 774 592
use scs8hd_nor2_4  _104_
timestamp 1586364061
transform 1 0 6348 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_66
timestamp 1586364061
transform 1 0 7176 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_70
timestamp 1586364061
transform 1 0 7544 0 -1 19040
box -38 -48 130 592
use scs8hd_nor2_4  _075_
timestamp 1586364061
transform 1 0 8004 0 -1 19040
box -38 -48 866 592
use scs8hd_fill_2  FILLER_30_73
timestamp 1586364061
transform 1 0 7820 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 774 592
use scs8hd_nor2_4  _072_
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_102
timestamp 1586364061
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_106
timestamp 1586364061
transform 1 0 10856 0 -1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11316 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_110
timestamp 1586364061
transform 1 0 11224 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_30_120
timestamp 1586364061
transform 1 0 12144 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_125
timestamp 1586364061
transform 1 0 12604 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_137
timestamp 1586364061
transform 1 0 13708 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_149
timestamp 1586364061
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_8  FILLER_30_157
timestamp 1586364061
transform 1 0 15548 0 -1 19040
box -38 -48 774 592
use scs8hd_nor2_4  _116_
timestamp 1586364061
transform 1 0 16560 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_165
timestamp 1586364061
transform 1 0 16284 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_8  FILLER_30_177
timestamp 1586364061
transform 1 0 17388 0 -1 19040
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18308 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_185
timestamp 1586364061
transform 1 0 18124 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_30_189
timestamp 1586364061
transform 1 0 18492 0 -1 19040
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_199
timestamp 1586364061
transform 1 0 19412 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_30_211
timestamp 1586364061
transform 1 0 20516 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 590 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 22816 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_7.LATCH_5_.latch
timestamp 1586364061
transform 1 0 4048 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 3864 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_7.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3496 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_23
timestamp 1586364061
transform 1 0 3220 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_28
timestamp 1586364061
transform 1 0 3680 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5612 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_43
timestamp 1586364061
transform 1 0 5060 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_47
timestamp 1586364061
transform 1 0 5428 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_nor2_4  _070_
timestamp 1586364061
transform 1 0 7636 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__070__B
timestamp 1586364061
transform 1 0 7452 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7084 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_67
timestamp 1586364061
transform 1 0 7268 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 8648 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_80
timestamp 1586364061
transform 1 0 8464 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_84
timestamp 1586364061
transform 1 0 8832 0 1 19040
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_3_.latch
timestamp 1586364061
transform 1 0 9936 0 1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_92
timestamp 1586364061
transform 1 0 9568 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_107
timestamp 1586364061
transform 1 0 10948 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_111
timestamp 1586364061
transform 1 0 11316 0 1 19040
box -38 -48 222 592
use scs8hd_decap_6  FILLER_31_115
timestamp 1586364061
transform 1 0 11684 0 1 19040
box -38 -48 590 592
use scs8hd_fill_1  FILLER_31_121
timestamp 1586364061
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 16376 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 16192 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_163
timestamp 1586364061
transform 1 0 16100 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_175
timestamp 1586364061
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_31_195
timestamp 1586364061
transform 1 0 19044 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_207
timestamp 1586364061
transform 1 0 20148 0 1 19040
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_218
timestamp 1586364061
transform 1 0 21160 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_222
timestamp 1586364061
transform 1 0 21528 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_31_230
timestamp 1586364061
transform 1 0 22264 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 22816 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_conb_1  _139_
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_8  FILLER_32_35
timestamp 1586364061
transform 1 0 4324 0 -1 20128
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_ipin_7.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5060 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_12  FILLER_32_52
timestamp 1586364061
transform 1 0 5888 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_32_64
timestamp 1586364061
transform 1 0 6992 0 -1 20128
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_3.LATCH_5_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 20128
box -38 -48 1050 592
use scs8hd_fill_1  FILLER_32_72
timestamp 1586364061
transform 1 0 7728 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_3.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9936 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_32_98
timestamp 1586364061
transform 1 0 10120 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_102
timestamp 1586364061
transform 1 0 10488 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_112
timestamp 1586364061
transform 1 0 11408 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_124
timestamp 1586364061
transform 1 0 12512 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_136
timestamp 1586364061
transform 1 0 13616 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_148
timestamp 1586364061
transform 1 0 14720 0 -1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_32_152
timestamp 1586364061
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_32_186
timestamp 1586364061
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_196
timestamp 1586364061
transform 1 0 19136 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_6  FILLER_32_208
timestamp 1586364061
transform 1 0 20240 0 -1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 590 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 22816 0 -1 20128
box -38 -48 314 592
use scs8hd_buf_2  _151_
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 1932 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_7
timestamp 1586364061
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_11
timestamp 1586364061
transform 1 0 2116 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_23
timestamp 1586364061
transform 1 0 3220 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_35
timestamp 1586364061
transform 1 0 4324 0 1 20128
box -38 -48 774 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5336 0 1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_33_43
timestamp 1586364061
transform 1 0 5060 0 1 20128
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_49
timestamp 1586364061
transform 1 0 5612 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_33_53
timestamp 1586364061
transform 1 0 5980 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7452 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_66
timestamp 1586364061
transform 1 0 7176 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 774 592
use scs8hd_conb_1  _135_
timestamp 1586364061
transform 1 0 8188 0 -1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8464 0 1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_72
timestamp 1586364061
transform 1 0 7728 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_76
timestamp 1586364061
transform 1 0 8096 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_89
timestamp 1586364061
transform 1 0 9292 0 1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_76
timestamp 1586364061
transform 1 0 8096 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_buf_2  _146_
timestamp 1586364061
transform 1 0 10948 0 1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_33_101
timestamp 1586364061
transform 1 0 10396 0 1 20128
box -38 -48 590 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 11500 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_111
timestamp 1586364061
transform 1 0 11316 0 1 20128
box -38 -48 222 592
use scs8hd_decap_6  FILLER_33_115
timestamp 1586364061
transform 1 0 11684 0 1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_33_121
timestamp 1586364061
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_126
timestamp 1586364061
transform 1 0 12696 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_130
timestamp 1586364061
transform 1 0 13064 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_142
timestamp 1586364061
transform 1 0 14168 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_154
timestamp 1586364061
transform 1 0 15272 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_166
timestamp 1586364061
transform 1 0 16376 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_33_178
timestamp 1586364061
transform 1 0 17480 0 1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 774 592
use scs8hd_conb_1  _131_
timestamp 1586364061
transform 1 0 18308 0 -1 21216
box -38 -48 314 592
use scs8hd_buf_2  _154_
timestamp 1586364061
transform 1 0 18952 0 1 20128
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_33_182
timestamp 1586364061
transform 1 0 17848 0 1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_192
timestamp 1586364061
transform 1 0 18768 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_186
timestamp 1586364061
transform 1 0 18216 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20056 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 19504 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20516 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_198
timestamp 1586364061
transform 1 0 19320 0 1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_202
timestamp 1586364061
transform 1 0 19688 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_209
timestamp 1586364061
transform 1 0 20332 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_213
timestamp 1586364061
transform 1 0 20700 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_225
timestamp 1586364061
transform 1 0 21804 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 590 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 22816 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 22816 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use scs8hd_decap_4  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_35_32
timestamp 1586364061
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_44
timestamp 1586364061
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_56
timestamp 1586364061
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_63
timestamp 1586364061
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_75
timestamp 1586364061
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_87
timestamp 1586364061
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_94
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_106
timestamp 1586364061
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_118
timestamp 1586364061
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_125
timestamp 1586364061
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_137
timestamp 1586364061
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_149
timestamp 1586364061
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_156
timestamp 1586364061
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_168
timestamp 1586364061
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_35_180
timestamp 1586364061
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use scs8hd_decap_12  FILLER_35_187
timestamp 1586364061
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_199
timestamp 1586364061
transform 1 0 19412 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_35_211
timestamp 1586364061
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_218
timestamp 1586364061
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_35_230
timestamp 1586364061
transform 1 0 22264 0 1 21216
box -38 -48 314 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 22816 0 1 21216
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 688 480 808 6 address[0]
port 0 nsew default input
rlabel metal3 s 23520 552 24000 672 6 address[1]
port 1 nsew default input
rlabel metal3 s 23520 1776 24000 1896 6 address[2]
port 2 nsew default input
rlabel metal3 s 23520 3000 24000 3120 6 address[3]
port 3 nsew default input
rlabel metal2 s 4894 0 4950 480 6 address[4]
port 4 nsew default input
rlabel metal3 s 23520 4224 24000 4344 6 address[5]
port 5 nsew default input
rlabel metal3 s 23520 5584 24000 5704 6 address[6]
port 6 nsew default input
rlabel metal3 s 0 2184 480 2304 6 bottom_grid_pin_0_
port 7 nsew default tristate
rlabel metal3 s 0 5176 480 5296 6 bottom_grid_pin_10_
port 8 nsew default tristate
rlabel metal2 s 8942 0 8998 480 6 bottom_grid_pin_12_
port 9 nsew default tristate
rlabel metal2 s 6642 23520 6698 24000 6 bottom_grid_pin_14_
port 10 nsew default tristate
rlabel metal2 s 1306 23520 1362 24000 6 bottom_grid_pin_2_
port 11 nsew default tristate
rlabel metal2 s 6918 0 6974 480 6 bottom_grid_pin_4_
port 12 nsew default tristate
rlabel metal2 s 3974 23520 4030 24000 6 bottom_grid_pin_6_
port 13 nsew default tristate
rlabel metal3 s 0 3680 480 3800 6 bottom_grid_pin_8_
port 14 nsew default tristate
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[0]
port 15 nsew default input
rlabel metal3 s 0 8168 480 8288 6 chanx_left_in[1]
port 16 nsew default input
rlabel metal3 s 23520 6808 24000 6928 6 chanx_left_in[2]
port 17 nsew default input
rlabel metal3 s 23520 8032 24000 8152 6 chanx_left_in[3]
port 18 nsew default input
rlabel metal3 s 0 9664 480 9784 6 chanx_left_in[4]
port 19 nsew default input
rlabel metal3 s 0 11160 480 11280 6 chanx_left_in[5]
port 20 nsew default input
rlabel metal2 s 9310 23520 9366 24000 6 chanx_left_in[6]
port 21 nsew default input
rlabel metal3 s 23520 9256 24000 9376 6 chanx_left_in[7]
port 22 nsew default input
rlabel metal3 s 0 12656 480 12776 6 chanx_left_in[8]
port 23 nsew default input
rlabel metal3 s 23520 10616 24000 10736 6 chanx_left_out[0]
port 24 nsew default tristate
rlabel metal2 s 10874 0 10930 480 6 chanx_left_out[1]
port 25 nsew default tristate
rlabel metal2 s 11978 23520 12034 24000 6 chanx_left_out[2]
port 26 nsew default tristate
rlabel metal2 s 12898 0 12954 480 6 chanx_left_out[3]
port 27 nsew default tristate
rlabel metal2 s 14922 0 14978 480 6 chanx_left_out[4]
port 28 nsew default tristate
rlabel metal2 s 16946 0 17002 480 6 chanx_left_out[5]
port 29 nsew default tristate
rlabel metal3 s 23520 11840 24000 11960 6 chanx_left_out[6]
port 30 nsew default tristate
rlabel metal3 s 0 14152 480 14272 6 chanx_left_out[7]
port 31 nsew default tristate
rlabel metal3 s 23520 13064 24000 13184 6 chanx_left_out[8]
port 32 nsew default tristate
rlabel metal3 s 0 15648 480 15768 6 chanx_right_in[0]
port 33 nsew default input
rlabel metal3 s 23520 14288 24000 14408 6 chanx_right_in[1]
port 34 nsew default input
rlabel metal3 s 0 17144 480 17264 6 chanx_right_in[2]
port 35 nsew default input
rlabel metal2 s 14646 23520 14702 24000 6 chanx_right_in[3]
port 36 nsew default input
rlabel metal2 s 18878 0 18934 480 6 chanx_right_in[4]
port 37 nsew default input
rlabel metal2 s 17314 23520 17370 24000 6 chanx_right_in[5]
port 38 nsew default input
rlabel metal3 s 23520 15648 24000 15768 6 chanx_right_in[6]
port 39 nsew default input
rlabel metal3 s 0 18640 480 18760 6 chanx_right_in[7]
port 40 nsew default input
rlabel metal3 s 23520 16872 24000 16992 6 chanx_right_in[8]
port 41 nsew default input
rlabel metal3 s 0 20136 480 20256 6 chanx_right_out[0]
port 42 nsew default tristate
rlabel metal2 s 20902 0 20958 480 6 chanx_right_out[1]
port 43 nsew default tristate
rlabel metal3 s 23520 18096 24000 18216 6 chanx_right_out[2]
port 44 nsew default tristate
rlabel metal2 s 19982 23520 20038 24000 6 chanx_right_out[3]
port 45 nsew default tristate
rlabel metal3 s 0 21632 480 21752 6 chanx_right_out[4]
port 46 nsew default tristate
rlabel metal3 s 23520 19320 24000 19440 6 chanx_right_out[5]
port 47 nsew default tristate
rlabel metal3 s 0 23128 480 23248 6 chanx_right_out[6]
port 48 nsew default tristate
rlabel metal2 s 22650 23520 22706 24000 6 chanx_right_out[7]
port 49 nsew default tristate
rlabel metal2 s 22926 0 22982 480 6 chanx_right_out[8]
port 50 nsew default tristate
rlabel metal2 s 2870 0 2926 480 6 data_in
port 51 nsew default input
rlabel metal2 s 938 0 994 480 6 enable
port 52 nsew default input
rlabel metal3 s 23520 23128 24000 23248 6 top_grid_pin_14_
port 53 nsew default tristate
rlabel metal3 s 23520 20680 24000 20800 6 top_grid_pin_2_
port 54 nsew default tristate
rlabel metal3 s 23520 21904 24000 22024 6 top_grid_pin_6_
port 55 nsew default tristate
rlabel metal4 s 4944 2128 5264 21808 6 vpwr
port 56 nsew default input
rlabel metal4 s 8944 2128 9264 21808 6 vgnd
port 57 nsew default input
<< end >>
