magic
tech sky130A
magscale 1 2
timestamp 1605199304
<< locali >>
rect 8401 11543 8435 11645
<< viali >>
rect 16773 20553 16807 20587
rect 18521 20553 18555 20587
rect 5273 20485 5307 20519
rect 15669 20485 15703 20519
rect 5917 20417 5951 20451
rect 10701 20417 10735 20451
rect 10885 20417 10919 20451
rect 2145 20349 2179 20383
rect 4077 20349 4111 20383
rect 6929 20349 6963 20383
rect 8401 20349 8435 20383
rect 12633 20349 12667 20383
rect 13737 20349 13771 20383
rect 15485 20349 15519 20383
rect 16589 20349 16623 20383
rect 18337 20349 18371 20383
rect 2421 20281 2455 20315
rect 8677 20281 8711 20315
rect 4261 20213 4295 20247
rect 5641 20213 5675 20247
rect 5733 20213 5767 20247
rect 7113 20213 7147 20247
rect 10241 20213 10275 20247
rect 10609 20213 10643 20247
rect 12817 20213 12851 20247
rect 13921 20213 13955 20247
rect 8125 20009 8159 20043
rect 17693 20009 17727 20043
rect 18797 20009 18831 20043
rect 2789 19941 2823 19975
rect 12142 19941 12176 19975
rect 1409 19873 1443 19907
rect 2513 19873 2547 19907
rect 4077 19873 4111 19907
rect 5540 19873 5574 19907
rect 8033 19873 8067 19907
rect 9945 19873 9979 19907
rect 14105 19873 14139 19907
rect 15301 19873 15335 19907
rect 16405 19873 16439 19907
rect 17509 19873 17543 19907
rect 18613 19873 18647 19907
rect 5273 19805 5307 19839
rect 8217 19805 8251 19839
rect 9689 19805 9723 19839
rect 11897 19805 11931 19839
rect 19717 19805 19751 19839
rect 14289 19737 14323 19771
rect 15485 19737 15519 19771
rect 1593 19669 1627 19703
rect 4261 19669 4295 19703
rect 6653 19669 6687 19703
rect 7665 19669 7699 19703
rect 11069 19669 11103 19703
rect 13277 19669 13311 19703
rect 16589 19669 16623 19703
rect 9137 19465 9171 19499
rect 10057 19465 10091 19499
rect 5825 19329 5859 19363
rect 10517 19329 10551 19363
rect 10701 19329 10735 19363
rect 19165 19329 19199 19363
rect 1777 19261 1811 19295
rect 2881 19261 2915 19295
rect 3148 19261 3182 19295
rect 5641 19261 5675 19295
rect 7757 19261 7791 19295
rect 13185 19261 13219 19295
rect 15393 19261 15427 19295
rect 18061 19261 18095 19295
rect 8024 19193 8058 19227
rect 10425 19193 10459 19227
rect 13452 19193 13486 19227
rect 15638 19193 15672 19227
rect 1961 19125 1995 19159
rect 4261 19125 4295 19159
rect 5181 19125 5215 19159
rect 5549 19125 5583 19159
rect 14565 19125 14599 19159
rect 16773 19125 16807 19159
rect 18245 19125 18279 19159
rect 2881 18921 2915 18955
rect 6837 18921 6871 18955
rect 8125 18921 8159 18955
rect 15485 18921 15519 18955
rect 16589 18921 16623 18955
rect 17693 18921 17727 18955
rect 4353 18853 4387 18887
rect 5724 18853 5758 18887
rect 9689 18853 9723 18887
rect 13277 18853 13311 18887
rect 2789 18785 2823 18819
rect 4077 18785 4111 18819
rect 8033 18785 8067 18819
rect 10957 18785 10991 18819
rect 15301 18785 15335 18819
rect 16405 18785 16439 18819
rect 17509 18785 17543 18819
rect 1409 18717 1443 18751
rect 3065 18717 3099 18751
rect 5457 18717 5491 18751
rect 8309 18717 8343 18751
rect 10701 18717 10735 18751
rect 13369 18717 13403 18751
rect 13553 18717 13587 18751
rect 7665 18649 7699 18683
rect 2421 18581 2455 18615
rect 12081 18581 12115 18615
rect 12909 18581 12943 18615
rect 2973 18377 3007 18411
rect 12541 18377 12575 18411
rect 15669 18377 15703 18411
rect 2881 18241 2915 18275
rect 3433 18241 3467 18275
rect 3617 18241 3651 18275
rect 5181 18241 5215 18275
rect 7481 18241 7515 18275
rect 9229 18241 9263 18275
rect 11253 18241 11287 18275
rect 11437 18241 11471 18275
rect 13185 18241 13219 18275
rect 1777 18173 1811 18207
rect 4997 18173 5031 18207
rect 7205 18173 7239 18207
rect 13001 18173 13035 18207
rect 14289 18173 14323 18207
rect 16497 18173 16531 18207
rect 3341 18105 3375 18139
rect 7297 18105 7331 18139
rect 11161 18105 11195 18139
rect 12909 18105 12943 18139
rect 14556 18105 14590 18139
rect 18061 18105 18095 18139
rect 18337 18105 18371 18139
rect 1961 18037 1995 18071
rect 4537 18037 4571 18071
rect 4905 18037 4939 18071
rect 6837 18037 6871 18071
rect 8585 18037 8619 18071
rect 8953 18037 8987 18071
rect 9045 18037 9079 18071
rect 10793 18037 10827 18071
rect 8217 17833 8251 17867
rect 9689 17833 9723 17867
rect 10149 17833 10183 17867
rect 11253 17833 11287 17867
rect 15577 17765 15611 17799
rect 2237 17697 2271 17731
rect 4333 17697 4367 17731
rect 7104 17697 7138 17731
rect 10057 17697 10091 17731
rect 11437 17697 11471 17731
rect 11529 17697 11563 17731
rect 11796 17697 11830 17731
rect 13737 17697 13771 17731
rect 15301 17697 15335 17731
rect 2421 17629 2455 17663
rect 4077 17629 4111 17663
rect 6837 17629 6871 17663
rect 10333 17629 10367 17663
rect 13921 17629 13955 17663
rect 16589 17629 16623 17663
rect 5457 17493 5491 17527
rect 12909 17493 12943 17527
rect 8217 17289 8251 17323
rect 11437 17289 11471 17323
rect 12449 17289 12483 17323
rect 15485 17289 15519 17323
rect 6193 17221 6227 17255
rect 2421 17153 2455 17187
rect 3985 17153 4019 17187
rect 9045 17153 9079 17187
rect 13001 17153 13035 17187
rect 14105 17153 14139 17187
rect 2145 17085 2179 17119
rect 4252 17085 4286 17119
rect 6377 17085 6411 17119
rect 6837 17085 6871 17119
rect 9312 17085 9346 17119
rect 11253 17085 11287 17119
rect 12817 17085 12851 17119
rect 7104 17017 7138 17051
rect 12909 17017 12943 17051
rect 14372 17017 14406 17051
rect 5365 16949 5399 16983
rect 10425 16949 10459 16983
rect 16313 16949 16347 16983
rect 4077 16745 4111 16779
rect 4537 16745 4571 16779
rect 6837 16745 6871 16779
rect 7297 16745 7331 16779
rect 8585 16745 8619 16779
rect 10977 16745 11011 16779
rect 12633 16745 12667 16779
rect 13645 16745 13679 16779
rect 15301 16745 15335 16779
rect 15669 16745 15703 16779
rect 4445 16677 4479 16711
rect 11520 16677 11554 16711
rect 15761 16677 15795 16711
rect 2145 16609 2179 16643
rect 2421 16609 2455 16643
rect 5641 16609 5675 16643
rect 7205 16609 7239 16643
rect 8401 16609 8435 16643
rect 9689 16609 9723 16643
rect 11161 16609 11195 16643
rect 11253 16609 11287 16643
rect 14013 16609 14047 16643
rect 14105 16609 14139 16643
rect 4721 16541 4755 16575
rect 7481 16541 7515 16575
rect 9873 16541 9907 16575
rect 14289 16541 14323 16575
rect 15853 16541 15887 16575
rect 5825 16405 5859 16439
rect 6837 16201 6871 16235
rect 15117 16201 15151 16235
rect 9873 16133 9907 16167
rect 3801 16065 3835 16099
rect 7481 16065 7515 16099
rect 8493 16065 8527 16099
rect 11437 16065 11471 16099
rect 12633 16065 12667 16099
rect 15945 16065 15979 16099
rect 2145 15997 2179 16031
rect 4068 15997 4102 16031
rect 8760 15997 8794 16031
rect 12449 15997 12483 16031
rect 13737 15997 13771 16031
rect 2421 15929 2455 15963
rect 14004 15929 14038 15963
rect 5181 15861 5215 15895
rect 7205 15861 7239 15895
rect 7297 15861 7331 15895
rect 10793 15861 10827 15895
rect 11161 15861 11195 15895
rect 11253 15861 11287 15895
rect 8493 15657 8527 15691
rect 9689 15657 9723 15691
rect 10149 15657 10183 15691
rect 11345 15657 11379 15691
rect 12081 15657 12115 15691
rect 13185 15657 13219 15691
rect 13553 15657 13587 15691
rect 15669 15657 15703 15691
rect 5172 15589 5206 15623
rect 2237 15521 2271 15555
rect 4905 15521 4939 15555
rect 7380 15521 7414 15555
rect 10057 15521 10091 15555
rect 11529 15521 11563 15555
rect 11989 15521 12023 15555
rect 15485 15521 15519 15555
rect 2513 15453 2547 15487
rect 7113 15453 7147 15487
rect 10241 15453 10275 15487
rect 12173 15453 12207 15487
rect 13645 15453 13679 15487
rect 13829 15453 13863 15487
rect 11621 15385 11655 15419
rect 6285 15317 6319 15351
rect 3065 15113 3099 15147
rect 9229 15113 9263 15147
rect 10793 15113 10827 15147
rect 13829 15113 13863 15147
rect 16037 15113 16071 15147
rect 3709 14977 3743 15011
rect 5181 14977 5215 15011
rect 7849 14977 7883 15011
rect 11253 14977 11287 15011
rect 11437 14977 11471 15011
rect 1777 14909 1811 14943
rect 5089 14909 5123 14943
rect 6377 14909 6411 14943
rect 8116 14909 8150 14943
rect 11161 14909 11195 14943
rect 12449 14909 12483 14943
rect 14657 14909 14691 14943
rect 16865 14909 16899 14943
rect 3433 14841 3467 14875
rect 12694 14841 12728 14875
rect 14902 14841 14936 14875
rect 1961 14773 1995 14807
rect 3525 14773 3559 14807
rect 4629 14773 4663 14807
rect 4997 14773 5031 14807
rect 6193 14773 6227 14807
rect 6837 14773 6871 14807
rect 4261 14569 4295 14603
rect 9689 14569 9723 14603
rect 12081 14569 12115 14603
rect 16773 14569 16807 14603
rect 8585 14501 8619 14535
rect 13737 14501 13771 14535
rect 15577 14501 15611 14535
rect 2789 14433 2823 14467
rect 4077 14433 4111 14467
rect 5181 14433 5215 14467
rect 6837 14433 6871 14467
rect 8309 14433 8343 14467
rect 10957 14433 10991 14467
rect 13461 14433 13495 14467
rect 15301 14433 15335 14467
rect 16589 14433 16623 14467
rect 1409 14365 1443 14399
rect 2881 14365 2915 14399
rect 3065 14365 3099 14399
rect 6929 14365 6963 14399
rect 7021 14365 7055 14399
rect 10701 14365 10735 14399
rect 5365 14297 5399 14331
rect 2421 14229 2455 14263
rect 6469 14229 6503 14263
rect 4077 14025 4111 14059
rect 6837 13957 6871 13991
rect 10609 13957 10643 13991
rect 12449 13957 12483 13991
rect 7389 13889 7423 13923
rect 9229 13889 9263 13923
rect 13001 13889 13035 13923
rect 15025 13889 15059 13923
rect 16313 13889 16347 13923
rect 1869 13821 1903 13855
rect 4261 13821 4295 13855
rect 4353 13821 4387 13855
rect 9496 13821 9530 13855
rect 12909 13821 12943 13855
rect 14749 13821 14783 13855
rect 16037 13821 16071 13855
rect 2136 13753 2170 13787
rect 4620 13753 4654 13787
rect 12817 13753 12851 13787
rect 3249 13685 3283 13719
rect 5733 13685 5767 13719
rect 7205 13685 7239 13719
rect 7297 13685 7331 13719
rect 2421 13481 2455 13515
rect 7021 13481 7055 13515
rect 7481 13481 7515 13515
rect 8585 13481 8619 13515
rect 5080 13413 5114 13447
rect 10149 13413 10183 13447
rect 15577 13413 15611 13447
rect 2789 13345 2823 13379
rect 4813 13345 4847 13379
rect 7389 13345 7423 13379
rect 10057 13345 10091 13379
rect 11437 13345 11471 13379
rect 11805 13345 11839 13379
rect 12072 13345 12106 13379
rect 15301 13345 15335 13379
rect 1409 13277 1443 13311
rect 2881 13277 2915 13311
rect 3065 13277 3099 13311
rect 7573 13277 7607 13311
rect 10333 13277 10367 13311
rect 14197 13277 14231 13311
rect 6193 13141 6227 13175
rect 9689 13141 9723 13175
rect 11253 13141 11287 13175
rect 13185 13141 13219 13175
rect 1593 12937 1627 12971
rect 4537 12937 4571 12971
rect 5549 12937 5583 12971
rect 6469 12937 6503 12971
rect 7021 12937 7055 12971
rect 15761 12937 15795 12971
rect 10609 12869 10643 12903
rect 14933 12869 14967 12903
rect 2237 12801 2271 12835
rect 7573 12801 7607 12835
rect 10333 12801 10367 12835
rect 11069 12801 11103 12835
rect 11253 12801 11287 12835
rect 16313 12801 16347 12835
rect 1961 12733 1995 12767
rect 3157 12733 3191 12767
rect 3413 12733 3447 12767
rect 5365 12733 5399 12767
rect 6653 12733 6687 12767
rect 7389 12733 7423 12767
rect 10977 12733 11011 12767
rect 13553 12733 13587 12767
rect 16129 12733 16163 12767
rect 8769 12665 8803 12699
rect 13820 12665 13854 12699
rect 2053 12597 2087 12631
rect 7481 12597 7515 12631
rect 12449 12597 12483 12631
rect 16221 12597 16255 12631
rect 3065 12393 3099 12427
rect 6653 12393 6687 12427
rect 8585 12393 8619 12427
rect 8953 12393 8987 12427
rect 11621 12393 11655 12427
rect 7021 12325 7055 12359
rect 11713 12325 11747 12359
rect 15568 12325 15602 12359
rect 17785 12325 17819 12359
rect 1685 12257 1719 12291
rect 1952 12257 1986 12291
rect 4445 12257 4479 12291
rect 5641 12257 5675 12291
rect 8309 12257 8343 12291
rect 9045 12257 9079 12291
rect 10057 12257 10091 12291
rect 13185 12257 13219 12291
rect 13277 12257 13311 12291
rect 14565 12257 14599 12291
rect 17509 12257 17543 12291
rect 4537 12189 4571 12223
rect 4721 12189 4755 12223
rect 7113 12189 7147 12223
rect 7297 12189 7331 12223
rect 9229 12189 9263 12223
rect 10149 12189 10183 12223
rect 10241 12189 10275 12223
rect 11805 12189 11839 12223
rect 13369 12189 13403 12223
rect 15301 12189 15335 12223
rect 4077 12121 4111 12155
rect 11253 12121 11287 12155
rect 14381 12121 14415 12155
rect 9689 12053 9723 12087
rect 12817 12053 12851 12087
rect 16681 12053 16715 12087
rect 1961 11849 1995 11883
rect 2973 11849 3007 11883
rect 6837 11849 6871 11883
rect 9873 11849 9907 11883
rect 14657 11849 14691 11883
rect 16221 11849 16255 11883
rect 10701 11781 10735 11815
rect 13829 11781 13863 11815
rect 3617 11713 3651 11747
rect 7297 11713 7331 11747
rect 7389 11713 7423 11747
rect 11161 11713 11195 11747
rect 11345 11713 11379 11747
rect 15209 11713 15243 11747
rect 16773 11713 16807 11747
rect 1777 11645 1811 11679
rect 4537 11645 4571 11679
rect 7205 11645 7239 11679
rect 8401 11645 8435 11679
rect 8493 11645 8527 11679
rect 12449 11645 12483 11679
rect 12716 11645 12750 11679
rect 15025 11645 15059 11679
rect 3341 11577 3375 11611
rect 4804 11577 4838 11611
rect 8760 11577 8794 11611
rect 11069 11577 11103 11611
rect 15117 11577 15151 11611
rect 16681 11577 16715 11611
rect 3433 11509 3467 11543
rect 5917 11509 5951 11543
rect 8401 11509 8435 11543
rect 16589 11509 16623 11543
rect 2881 11305 2915 11339
rect 4077 11305 4111 11339
rect 4537 11305 4571 11339
rect 8585 11305 8619 11339
rect 14197 11305 14231 11339
rect 16396 11237 16430 11271
rect 18613 11237 18647 11271
rect 2789 11169 2823 11203
rect 4445 11169 4479 11203
rect 6009 11169 6043 11203
rect 7205 11169 7239 11203
rect 7472 11169 7506 11203
rect 10692 11169 10726 11203
rect 13001 11169 13035 11203
rect 14381 11169 14415 11203
rect 18337 11169 18371 11203
rect 1409 11101 1443 11135
rect 2973 11101 3007 11135
rect 4721 11101 4755 11135
rect 6101 11101 6135 11135
rect 6285 11101 6319 11135
rect 10425 11101 10459 11135
rect 13093 11101 13127 11135
rect 13185 11101 13219 11135
rect 16129 11101 16163 11135
rect 2421 11033 2455 11067
rect 5641 10965 5675 10999
rect 11805 10965 11839 10999
rect 12633 10965 12667 10999
rect 17509 10965 17543 10999
rect 3341 10761 3375 10795
rect 8217 10761 8251 10795
rect 4905 10693 4939 10727
rect 2053 10625 2087 10659
rect 2145 10625 2179 10659
rect 3893 10625 3927 10659
rect 5365 10625 5399 10659
rect 5457 10625 5491 10659
rect 9045 10625 9079 10659
rect 14013 10625 14047 10659
rect 1961 10557 1995 10591
rect 3709 10557 3743 10591
rect 6653 10557 6687 10591
rect 6837 10557 6871 10591
rect 10057 10557 10091 10591
rect 10324 10557 10358 10591
rect 13829 10557 13863 10591
rect 14933 10557 14967 10591
rect 15200 10557 15234 10591
rect 5273 10489 5307 10523
rect 7082 10489 7116 10523
rect 13737 10489 13771 10523
rect 1593 10421 1627 10455
rect 3801 10421 3835 10455
rect 6469 10421 6503 10455
rect 11437 10421 11471 10455
rect 13369 10421 13403 10455
rect 16313 10421 16347 10455
rect 18061 10421 18095 10455
rect 3157 10217 3191 10251
rect 6377 10217 6411 10251
rect 7205 10217 7239 10251
rect 7573 10217 7607 10251
rect 10057 10217 10091 10251
rect 11621 10217 11655 10251
rect 13645 10217 13679 10251
rect 16221 10217 16255 10251
rect 2044 10149 2078 10183
rect 5264 10149 5298 10183
rect 11713 10149 11747 10183
rect 17693 10149 17727 10183
rect 1777 10081 1811 10115
rect 7665 10081 7699 10115
rect 14013 10081 14047 10115
rect 16313 10081 16347 10115
rect 17417 10081 17451 10115
rect 4997 10013 5031 10047
rect 7757 10013 7791 10047
rect 10149 10013 10183 10047
rect 10241 10013 10275 10047
rect 11897 10013 11931 10047
rect 14105 10013 14139 10047
rect 14289 10013 14323 10047
rect 16405 10013 16439 10047
rect 15853 9945 15887 9979
rect 9689 9877 9723 9911
rect 11253 9877 11287 9911
rect 4997 9673 5031 9707
rect 6469 9673 6503 9707
rect 6837 9605 6871 9639
rect 9965 9605 9999 9639
rect 10793 9605 10827 9639
rect 18429 9605 18463 9639
rect 1409 9537 1443 9571
rect 3617 9537 3651 9571
rect 7297 9537 7331 9571
rect 7481 9537 7515 9571
rect 11345 9537 11379 9571
rect 15761 9537 15795 9571
rect 1676 9469 1710 9503
rect 3884 9469 3918 9503
rect 6653 9469 6687 9503
rect 8585 9469 8619 9503
rect 8852 9469 8886 9503
rect 11161 9469 11195 9503
rect 13185 9469 13219 9503
rect 16028 9469 16062 9503
rect 18245 9469 18279 9503
rect 13452 9401 13486 9435
rect 2789 9333 2823 9367
rect 7205 9333 7239 9367
rect 11253 9333 11287 9367
rect 14565 9333 14599 9367
rect 17141 9333 17175 9367
rect 1961 9129 1995 9163
rect 6101 9129 6135 9163
rect 6929 9129 6963 9163
rect 8585 9129 8619 9163
rect 11069 9129 11103 9163
rect 11897 9129 11931 9163
rect 12633 9129 12667 9163
rect 18153 9061 18187 9095
rect 1777 8993 1811 9027
rect 4905 8993 4939 9027
rect 6285 8993 6319 9027
rect 7297 8993 7331 9027
rect 9689 8993 9723 9027
rect 9956 8993 9990 9027
rect 12081 8993 12115 9027
rect 13001 8993 13035 9027
rect 15301 8993 15335 9027
rect 16589 8993 16623 9027
rect 17877 8993 17911 9027
rect 2881 8925 2915 8959
rect 4997 8925 5031 8959
rect 5181 8925 5215 8959
rect 7389 8925 7423 8959
rect 7573 8925 7607 8959
rect 13093 8925 13127 8959
rect 13277 8925 13311 8959
rect 14197 8925 14231 8959
rect 15577 8925 15611 8959
rect 16865 8925 16899 8959
rect 4537 8857 4571 8891
rect 3709 8585 3743 8619
rect 7113 8585 7147 8619
rect 19533 8585 19567 8619
rect 8677 8517 8711 8551
rect 10793 8517 10827 8551
rect 2237 8449 2271 8483
rect 4169 8449 4203 8483
rect 4353 8449 4387 8483
rect 5273 8449 5307 8483
rect 7573 8449 7607 8483
rect 7757 8449 7791 8483
rect 9321 8449 9355 8483
rect 11437 8449 11471 8483
rect 12449 8449 12483 8483
rect 14657 8449 14691 8483
rect 18245 8449 18279 8483
rect 2053 8381 2087 8415
rect 18061 8381 18095 8415
rect 19349 8381 19383 8415
rect 7481 8313 7515 8347
rect 9137 8313 9171 8347
rect 11253 8313 11287 8347
rect 12716 8313 12750 8347
rect 14902 8313 14936 8347
rect 4077 8245 4111 8279
rect 9045 8245 9079 8279
rect 11161 8245 11195 8279
rect 13829 8245 13863 8279
rect 16037 8245 16071 8279
rect 2605 8041 2639 8075
rect 7205 8041 7239 8075
rect 9689 8041 9723 8075
rect 15301 8041 15335 8075
rect 5242 7973 5276 8007
rect 11529 7973 11563 8007
rect 18061 7973 18095 8007
rect 2697 7905 2731 7939
rect 7573 7905 7607 7939
rect 10057 7905 10091 7939
rect 11253 7905 11287 7939
rect 12808 7905 12842 7939
rect 17785 7905 17819 7939
rect 2789 7837 2823 7871
rect 4997 7837 5031 7871
rect 7665 7837 7699 7871
rect 7757 7837 7791 7871
rect 10149 7837 10183 7871
rect 10333 7837 10367 7871
rect 12541 7837 12575 7871
rect 6377 7769 6411 7803
rect 2237 7701 2271 7735
rect 13921 7701 13955 7735
rect 5273 7497 5307 7531
rect 8217 7497 8251 7531
rect 9873 7497 9907 7531
rect 12633 7497 12667 7531
rect 3893 7361 3927 7395
rect 6837 7361 6871 7395
rect 10425 7361 10459 7395
rect 13093 7361 13127 7395
rect 13277 7361 13311 7395
rect 1685 7293 1719 7327
rect 4160 7293 4194 7327
rect 10241 7293 10275 7327
rect 13001 7293 13035 7327
rect 1952 7225 1986 7259
rect 7104 7225 7138 7259
rect 3065 7157 3099 7191
rect 10333 7157 10367 7191
rect 1869 6953 1903 6987
rect 4905 6953 4939 6987
rect 11897 6953 11931 6987
rect 2237 6885 2271 6919
rect 7196 6885 7230 6919
rect 10762 6885 10796 6919
rect 2329 6817 2363 6851
rect 18981 6817 19015 6851
rect 2421 6749 2455 6783
rect 4997 6749 5031 6783
rect 5181 6749 5215 6783
rect 6929 6749 6963 6783
rect 10517 6749 10551 6783
rect 19165 6681 19199 6715
rect 4537 6613 4571 6647
rect 8309 6613 8343 6647
rect 10609 6409 10643 6443
rect 19717 6409 19751 6443
rect 5089 6273 5123 6307
rect 5273 6273 5307 6307
rect 9229 6273 9263 6307
rect 2421 6205 2455 6239
rect 2688 6205 2722 6239
rect 6837 6205 6871 6239
rect 7093 6205 7127 6239
rect 9496 6205 9530 6239
rect 19533 6205 19567 6239
rect 3801 6069 3835 6103
rect 4629 6069 4663 6103
rect 4997 6069 5031 6103
rect 8217 6069 8251 6103
rect 2421 5865 2455 5899
rect 6561 5865 6595 5899
rect 7389 5865 7423 5899
rect 10701 5865 10735 5899
rect 11161 5865 11195 5899
rect 19901 5865 19935 5899
rect 2329 5797 2363 5831
rect 2881 5797 2915 5831
rect 5426 5797 5460 5831
rect 10609 5797 10643 5831
rect 2789 5729 2823 5763
rect 11069 5729 11103 5763
rect 19717 5729 19751 5763
rect 3065 5661 3099 5695
rect 5181 5661 5215 5695
rect 9689 5661 9723 5695
rect 11253 5661 11287 5695
rect 5089 5321 5123 5355
rect 9413 5321 9447 5355
rect 10241 5321 10275 5355
rect 19625 5321 19659 5355
rect 20729 5321 20763 5355
rect 3709 5185 3743 5219
rect 8033 5185 8067 5219
rect 10793 5185 10827 5219
rect 2053 5117 2087 5151
rect 3965 5117 3999 5151
rect 8300 5117 8334 5151
rect 10609 5117 10643 5151
rect 19441 5117 19475 5151
rect 20545 5117 20579 5151
rect 2329 5049 2363 5083
rect 6837 4981 6871 5015
rect 10701 4981 10735 5015
rect 1961 4777 1995 4811
rect 4905 4777 4939 4811
rect 5273 4777 5307 4811
rect 1777 4641 1811 4675
rect 5365 4573 5399 4607
rect 5457 4573 5491 4607
rect 20545 4029 20579 4063
rect 20729 3893 20763 3927
<< metal1 >>
rect 3510 21088 3516 21140
rect 3568 21128 3574 21140
rect 6086 21128 6092 21140
rect 3568 21100 6092 21128
rect 3568 21088 3574 21100
rect 6086 21088 6092 21100
rect 6144 21088 6150 21140
rect 3786 20952 3792 21004
rect 3844 20992 3850 21004
rect 11238 20992 11244 21004
rect 3844 20964 11244 20992
rect 3844 20952 3850 20964
rect 11238 20952 11244 20964
rect 11296 20952 11302 21004
rect 4062 20748 4068 20800
rect 4120 20788 4126 20800
rect 15470 20788 15476 20800
rect 4120 20760 15476 20788
rect 4120 20748 4126 20760
rect 15470 20748 15476 20760
rect 15528 20748 15534 20800
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 3970 20544 3976 20596
rect 4028 20584 4034 20596
rect 8754 20584 8760 20596
rect 4028 20556 8760 20584
rect 4028 20544 4034 20556
rect 8754 20544 8760 20556
rect 8812 20544 8818 20596
rect 8938 20544 8944 20596
rect 8996 20584 9002 20596
rect 11790 20584 11796 20596
rect 8996 20556 11796 20584
rect 8996 20544 9002 20556
rect 11790 20544 11796 20556
rect 11848 20544 11854 20596
rect 13262 20544 13268 20596
rect 13320 20584 13326 20596
rect 13320 20556 14504 20584
rect 13320 20544 13326 20556
rect 4062 20476 4068 20528
rect 4120 20516 4126 20528
rect 5261 20519 5319 20525
rect 5261 20516 5273 20519
rect 4120 20488 5273 20516
rect 4120 20476 4126 20488
rect 5261 20485 5273 20488
rect 5307 20485 5319 20519
rect 5261 20479 5319 20485
rect 5442 20476 5448 20528
rect 5500 20516 5506 20528
rect 5500 20488 6040 20516
rect 5500 20476 5506 20488
rect 5902 20448 5908 20460
rect 5863 20420 5908 20448
rect 5902 20408 5908 20420
rect 5960 20408 5966 20460
rect 6012 20448 6040 20488
rect 6178 20476 6184 20528
rect 6236 20516 6242 20528
rect 8110 20516 8116 20528
rect 6236 20488 8116 20516
rect 6236 20476 6242 20488
rect 8110 20476 8116 20488
rect 8168 20476 8174 20528
rect 12710 20516 12716 20528
rect 8220 20488 12716 20516
rect 8220 20448 8248 20488
rect 12710 20476 12716 20488
rect 12768 20476 12774 20528
rect 14476 20516 14504 20556
rect 14734 20544 14740 20596
rect 14792 20584 14798 20596
rect 16761 20587 16819 20593
rect 16761 20584 16773 20587
rect 14792 20556 16773 20584
rect 14792 20544 14798 20556
rect 16761 20553 16773 20556
rect 16807 20553 16819 20587
rect 16761 20547 16819 20553
rect 18509 20587 18567 20593
rect 18509 20553 18521 20587
rect 18555 20584 18567 20587
rect 18598 20584 18604 20596
rect 18555 20556 18604 20584
rect 18555 20553 18567 20556
rect 18509 20547 18567 20553
rect 18598 20544 18604 20556
rect 18656 20544 18662 20596
rect 15657 20519 15715 20525
rect 15657 20516 15669 20519
rect 12820 20488 13860 20516
rect 14476 20488 15669 20516
rect 6012 20420 8248 20448
rect 8312 20420 10180 20448
rect 2130 20380 2136 20392
rect 2091 20352 2136 20380
rect 2130 20340 2136 20352
rect 2188 20340 2194 20392
rect 4065 20383 4123 20389
rect 4065 20349 4077 20383
rect 4111 20380 4123 20383
rect 6178 20380 6184 20392
rect 4111 20352 6184 20380
rect 4111 20349 4123 20352
rect 4065 20343 4123 20349
rect 6178 20340 6184 20352
rect 6236 20340 6242 20392
rect 6822 20340 6828 20392
rect 6880 20380 6886 20392
rect 6917 20383 6975 20389
rect 6917 20380 6929 20383
rect 6880 20352 6929 20380
rect 6880 20340 6886 20352
rect 6917 20349 6929 20352
rect 6963 20349 6975 20383
rect 6917 20343 6975 20349
rect 2409 20315 2467 20321
rect 2409 20281 2421 20315
rect 2455 20312 2467 20315
rect 8312 20312 8340 20420
rect 8389 20383 8447 20389
rect 8389 20349 8401 20383
rect 8435 20380 8447 20383
rect 10042 20380 10048 20392
rect 8435 20352 10048 20380
rect 8435 20349 8447 20352
rect 8389 20343 8447 20349
rect 10042 20340 10048 20352
rect 10100 20340 10106 20392
rect 10152 20380 10180 20420
rect 10502 20408 10508 20460
rect 10560 20448 10566 20460
rect 10689 20451 10747 20457
rect 10689 20448 10701 20451
rect 10560 20420 10701 20448
rect 10560 20408 10566 20420
rect 10689 20417 10701 20420
rect 10735 20417 10747 20451
rect 10689 20411 10747 20417
rect 10873 20451 10931 20457
rect 10873 20417 10885 20451
rect 10919 20448 10931 20451
rect 12066 20448 12072 20460
rect 10919 20420 12072 20448
rect 10919 20417 10931 20420
rect 10873 20411 10931 20417
rect 12066 20408 12072 20420
rect 12124 20408 12130 20460
rect 12158 20408 12164 20460
rect 12216 20448 12222 20460
rect 12820 20448 12848 20488
rect 12216 20420 12848 20448
rect 12216 20408 12222 20420
rect 12621 20383 12679 20389
rect 12621 20380 12633 20383
rect 10152 20352 12633 20380
rect 12621 20349 12633 20352
rect 12667 20349 12679 20383
rect 12621 20343 12679 20349
rect 12710 20340 12716 20392
rect 12768 20380 12774 20392
rect 13725 20383 13783 20389
rect 13725 20380 13737 20383
rect 12768 20352 13737 20380
rect 12768 20340 12774 20352
rect 13725 20349 13737 20352
rect 13771 20349 13783 20383
rect 13832 20380 13860 20488
rect 15657 20485 15669 20488
rect 15703 20485 15715 20519
rect 15657 20479 15715 20485
rect 15473 20383 15531 20389
rect 15473 20380 15485 20383
rect 13832 20352 15485 20380
rect 13725 20343 13783 20349
rect 15473 20349 15485 20352
rect 15519 20349 15531 20383
rect 15473 20343 15531 20349
rect 16577 20383 16635 20389
rect 16577 20349 16589 20383
rect 16623 20380 16635 20383
rect 16942 20380 16948 20392
rect 16623 20352 16948 20380
rect 16623 20349 16635 20352
rect 16577 20343 16635 20349
rect 16942 20340 16948 20352
rect 17000 20340 17006 20392
rect 18138 20340 18144 20392
rect 18196 20380 18202 20392
rect 18325 20383 18383 20389
rect 18325 20380 18337 20383
rect 18196 20352 18337 20380
rect 18196 20340 18202 20352
rect 18325 20349 18337 20352
rect 18371 20349 18383 20383
rect 18325 20343 18383 20349
rect 8662 20312 8668 20324
rect 2455 20284 8340 20312
rect 8623 20284 8668 20312
rect 2455 20281 2467 20284
rect 2409 20275 2467 20281
rect 8662 20272 8668 20284
rect 8720 20272 8726 20324
rect 8754 20272 8760 20324
rect 8812 20312 8818 20324
rect 8812 20284 13952 20312
rect 8812 20272 8818 20284
rect 3234 20204 3240 20256
rect 3292 20244 3298 20256
rect 4249 20247 4307 20253
rect 4249 20244 4261 20247
rect 3292 20216 4261 20244
rect 3292 20204 3298 20216
rect 4249 20213 4261 20216
rect 4295 20213 4307 20247
rect 5626 20244 5632 20256
rect 5587 20216 5632 20244
rect 4249 20207 4307 20213
rect 5626 20204 5632 20216
rect 5684 20204 5690 20256
rect 5718 20204 5724 20256
rect 5776 20244 5782 20256
rect 7098 20244 7104 20256
rect 5776 20216 5821 20244
rect 7059 20216 7104 20244
rect 5776 20204 5782 20216
rect 7098 20204 7104 20216
rect 7156 20204 7162 20256
rect 10229 20247 10287 20253
rect 10229 20213 10241 20247
rect 10275 20244 10287 20247
rect 10410 20244 10416 20256
rect 10275 20216 10416 20244
rect 10275 20213 10287 20216
rect 10229 20207 10287 20213
rect 10410 20204 10416 20216
rect 10468 20204 10474 20256
rect 10594 20244 10600 20256
rect 10555 20216 10600 20244
rect 10594 20204 10600 20216
rect 10652 20204 10658 20256
rect 12802 20244 12808 20256
rect 12763 20216 12808 20244
rect 12802 20204 12808 20216
rect 12860 20204 12866 20256
rect 13924 20253 13952 20284
rect 13909 20247 13967 20253
rect 13909 20213 13921 20247
rect 13955 20213 13967 20247
rect 13909 20207 13967 20213
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 4246 20000 4252 20052
rect 4304 20040 4310 20052
rect 7098 20040 7104 20052
rect 4304 20012 7104 20040
rect 4304 20000 4310 20012
rect 7098 20000 7104 20012
rect 7156 20000 7162 20052
rect 7190 20000 7196 20052
rect 7248 20040 7254 20052
rect 8113 20043 8171 20049
rect 8113 20040 8125 20043
rect 7248 20012 8125 20040
rect 7248 20000 7254 20012
rect 8113 20009 8125 20012
rect 8159 20009 8171 20043
rect 8113 20003 8171 20009
rect 9048 20012 15148 20040
rect 2777 19975 2835 19981
rect 2777 19941 2789 19975
rect 2823 19972 2835 19975
rect 5442 19972 5448 19984
rect 2823 19944 5448 19972
rect 2823 19941 2835 19944
rect 2777 19935 2835 19941
rect 5442 19932 5448 19944
rect 5500 19932 5506 19984
rect 5626 19932 5632 19984
rect 5684 19972 5690 19984
rect 9048 19972 9076 20012
rect 5684 19944 9076 19972
rect 5684 19932 5690 19944
rect 9490 19932 9496 19984
rect 9548 19972 9554 19984
rect 10594 19972 10600 19984
rect 9548 19944 10600 19972
rect 9548 19932 9554 19944
rect 10594 19932 10600 19944
rect 10652 19932 10658 19984
rect 12066 19932 12072 19984
rect 12124 19981 12130 19984
rect 12124 19975 12188 19981
rect 12124 19941 12142 19975
rect 12176 19941 12188 19975
rect 15120 19972 15148 20012
rect 15194 20000 15200 20052
rect 15252 20040 15258 20052
rect 17681 20043 17739 20049
rect 17681 20040 17693 20043
rect 15252 20012 17693 20040
rect 15252 20000 15258 20012
rect 17681 20009 17693 20012
rect 17727 20009 17739 20043
rect 17681 20003 17739 20009
rect 17954 20000 17960 20052
rect 18012 20040 18018 20052
rect 18785 20043 18843 20049
rect 18785 20040 18797 20043
rect 18012 20012 18797 20040
rect 18012 20000 18018 20012
rect 18785 20009 18797 20012
rect 18831 20009 18843 20043
rect 18785 20003 18843 20009
rect 19150 19972 19156 19984
rect 15120 19944 19156 19972
rect 12124 19935 12188 19941
rect 12124 19932 12130 19935
rect 19150 19932 19156 19944
rect 19208 19932 19214 19984
rect 1394 19904 1400 19916
rect 1355 19876 1400 19904
rect 1394 19864 1400 19876
rect 1452 19864 1458 19916
rect 2501 19907 2559 19913
rect 2501 19873 2513 19907
rect 2547 19904 2559 19907
rect 2958 19904 2964 19916
rect 2547 19876 2964 19904
rect 2547 19873 2559 19876
rect 2501 19867 2559 19873
rect 2958 19864 2964 19876
rect 3016 19864 3022 19916
rect 3602 19864 3608 19916
rect 3660 19904 3666 19916
rect 4065 19907 4123 19913
rect 4065 19904 4077 19907
rect 3660 19876 4077 19904
rect 3660 19864 3666 19876
rect 4065 19873 4077 19876
rect 4111 19873 4123 19907
rect 4065 19867 4123 19873
rect 5528 19907 5586 19913
rect 5528 19873 5540 19907
rect 5574 19904 5586 19907
rect 5902 19904 5908 19916
rect 5574 19876 5908 19904
rect 5574 19873 5586 19876
rect 5528 19867 5586 19873
rect 5902 19864 5908 19876
rect 5960 19904 5966 19916
rect 6822 19904 6828 19916
rect 5960 19876 6828 19904
rect 5960 19864 5966 19876
rect 6822 19864 6828 19876
rect 6880 19864 6886 19916
rect 8021 19907 8079 19913
rect 8021 19873 8033 19907
rect 8067 19904 8079 19907
rect 8938 19904 8944 19916
rect 8067 19876 8944 19904
rect 8067 19873 8079 19876
rect 8021 19867 8079 19873
rect 8938 19864 8944 19876
rect 8996 19864 9002 19916
rect 9122 19864 9128 19916
rect 9180 19904 9186 19916
rect 9933 19907 9991 19913
rect 9933 19904 9945 19907
rect 9180 19876 9945 19904
rect 9180 19864 9186 19876
rect 9933 19873 9945 19876
rect 9979 19873 9991 19907
rect 9933 19867 9991 19873
rect 12894 19864 12900 19916
rect 12952 19904 12958 19916
rect 14093 19907 14151 19913
rect 14093 19904 14105 19907
rect 12952 19876 14105 19904
rect 12952 19864 12958 19876
rect 14093 19873 14105 19876
rect 14139 19873 14151 19907
rect 15286 19904 15292 19916
rect 15247 19876 15292 19904
rect 14093 19867 14151 19873
rect 15286 19864 15292 19876
rect 15344 19864 15350 19916
rect 16390 19904 16396 19916
rect 16351 19876 16396 19904
rect 16390 19864 16396 19876
rect 16448 19864 16454 19916
rect 17402 19864 17408 19916
rect 17460 19904 17466 19916
rect 17497 19907 17555 19913
rect 17497 19904 17509 19907
rect 17460 19876 17509 19904
rect 17460 19864 17466 19876
rect 17497 19873 17509 19876
rect 17543 19873 17555 19907
rect 18598 19904 18604 19916
rect 18559 19876 18604 19904
rect 17497 19867 17555 19873
rect 18598 19864 18604 19876
rect 18656 19864 18662 19916
rect 4982 19796 4988 19848
rect 5040 19836 5046 19848
rect 5261 19839 5319 19845
rect 5261 19836 5273 19839
rect 5040 19808 5273 19836
rect 5040 19796 5046 19808
rect 5261 19805 5273 19808
rect 5307 19805 5319 19839
rect 8202 19836 8208 19848
rect 8163 19808 8208 19836
rect 5261 19799 5319 19805
rect 8202 19796 8208 19808
rect 8260 19796 8266 19848
rect 9674 19836 9680 19848
rect 9635 19808 9680 19836
rect 9674 19796 9680 19808
rect 9732 19796 9738 19848
rect 11882 19836 11888 19848
rect 11843 19808 11888 19836
rect 11882 19796 11888 19808
rect 11940 19796 11946 19848
rect 19702 19836 19708 19848
rect 19663 19808 19708 19836
rect 19702 19796 19708 19808
rect 19760 19796 19766 19848
rect 6362 19728 6368 19780
rect 6420 19768 6426 19780
rect 6420 19740 7788 19768
rect 6420 19728 6426 19740
rect 1578 19700 1584 19712
rect 1539 19672 1584 19700
rect 1578 19660 1584 19672
rect 1636 19660 1642 19712
rect 3510 19660 3516 19712
rect 3568 19700 3574 19712
rect 4249 19703 4307 19709
rect 4249 19700 4261 19703
rect 3568 19672 4261 19700
rect 3568 19660 3574 19672
rect 4249 19669 4261 19672
rect 4295 19669 4307 19703
rect 4249 19663 4307 19669
rect 4338 19660 4344 19712
rect 4396 19700 4402 19712
rect 6641 19703 6699 19709
rect 6641 19700 6653 19703
rect 4396 19672 6653 19700
rect 4396 19660 4402 19672
rect 6641 19669 6653 19672
rect 6687 19669 6699 19703
rect 7650 19700 7656 19712
rect 7611 19672 7656 19700
rect 6641 19663 6699 19669
rect 7650 19660 7656 19672
rect 7708 19660 7714 19712
rect 7760 19700 7788 19740
rect 7834 19728 7840 19780
rect 7892 19768 7898 19780
rect 9214 19768 9220 19780
rect 7892 19740 9220 19768
rect 7892 19728 7898 19740
rect 9214 19728 9220 19740
rect 9272 19768 9278 19780
rect 9490 19768 9496 19780
rect 9272 19740 9496 19768
rect 9272 19728 9278 19740
rect 9490 19728 9496 19740
rect 9548 19728 9554 19780
rect 10686 19728 10692 19780
rect 10744 19768 10750 19780
rect 10744 19740 11192 19768
rect 10744 19728 10750 19740
rect 11057 19703 11115 19709
rect 11057 19700 11069 19703
rect 7760 19672 11069 19700
rect 11057 19669 11069 19672
rect 11103 19669 11115 19703
rect 11164 19700 11192 19740
rect 12986 19728 12992 19780
rect 13044 19768 13050 19780
rect 14277 19771 14335 19777
rect 14277 19768 14289 19771
rect 13044 19740 14289 19768
rect 13044 19728 13050 19740
rect 14277 19737 14289 19740
rect 14323 19737 14335 19771
rect 15470 19768 15476 19780
rect 15431 19740 15476 19768
rect 14277 19731 14335 19737
rect 15470 19728 15476 19740
rect 15528 19728 15534 19780
rect 13265 19703 13323 19709
rect 13265 19700 13277 19703
rect 11164 19672 13277 19700
rect 11057 19663 11115 19669
rect 13265 19669 13277 19672
rect 13311 19669 13323 19703
rect 13265 19663 13323 19669
rect 16577 19703 16635 19709
rect 16577 19669 16589 19703
rect 16623 19700 16635 19703
rect 16666 19700 16672 19712
rect 16623 19672 16672 19700
rect 16623 19669 16635 19672
rect 16577 19663 16635 19669
rect 16666 19660 16672 19672
rect 16724 19660 16730 19712
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 3786 19456 3792 19508
rect 3844 19456 3850 19508
rect 3970 19456 3976 19508
rect 4028 19496 4034 19508
rect 9122 19496 9128 19508
rect 4028 19468 8708 19496
rect 9083 19468 9128 19496
rect 4028 19456 4034 19468
rect 3804 19428 3832 19456
rect 8680 19428 8708 19468
rect 9122 19456 9128 19468
rect 9180 19456 9186 19508
rect 10042 19496 10048 19508
rect 10003 19468 10048 19496
rect 10042 19456 10048 19468
rect 10100 19456 10106 19508
rect 9950 19428 9956 19440
rect 3804 19400 6500 19428
rect 8680 19400 9956 19428
rect 5813 19363 5871 19369
rect 5813 19329 5825 19363
rect 5859 19360 5871 19363
rect 5902 19360 5908 19372
rect 5859 19332 5908 19360
rect 5859 19329 5871 19332
rect 5813 19323 5871 19329
rect 5902 19320 5908 19332
rect 5960 19360 5966 19372
rect 6362 19360 6368 19372
rect 5960 19332 6368 19360
rect 5960 19320 5966 19332
rect 6362 19320 6368 19332
rect 6420 19320 6426 19372
rect 6472 19360 6500 19400
rect 9950 19388 9956 19400
rect 10008 19388 10014 19440
rect 12986 19428 12992 19440
rect 10336 19400 12992 19428
rect 10336 19360 10364 19400
rect 12986 19388 12992 19400
rect 13044 19388 13050 19440
rect 6472 19332 7880 19360
rect 1765 19295 1823 19301
rect 1765 19261 1777 19295
rect 1811 19292 1823 19295
rect 2866 19292 2872 19304
rect 1811 19264 2452 19292
rect 2827 19264 2872 19292
rect 1811 19261 1823 19264
rect 1765 19255 1823 19261
rect 1762 19116 1768 19168
rect 1820 19156 1826 19168
rect 1949 19159 2007 19165
rect 1949 19156 1961 19159
rect 1820 19128 1961 19156
rect 1820 19116 1826 19128
rect 1949 19125 1961 19128
rect 1995 19125 2007 19159
rect 2424 19156 2452 19264
rect 2866 19252 2872 19264
rect 2924 19252 2930 19304
rect 3136 19295 3194 19301
rect 3136 19261 3148 19295
rect 3182 19292 3194 19295
rect 4338 19292 4344 19304
rect 3182 19264 4344 19292
rect 3182 19261 3194 19264
rect 3136 19255 3194 19261
rect 4338 19252 4344 19264
rect 4396 19252 4402 19304
rect 5534 19292 5540 19304
rect 4448 19264 5540 19292
rect 2498 19184 2504 19236
rect 2556 19224 2562 19236
rect 3694 19224 3700 19236
rect 2556 19196 3700 19224
rect 2556 19184 2562 19196
rect 3694 19184 3700 19196
rect 3752 19184 3758 19236
rect 4448 19224 4476 19264
rect 5534 19252 5540 19264
rect 5592 19252 5598 19304
rect 5629 19295 5687 19301
rect 5629 19261 5641 19295
rect 5675 19292 5687 19295
rect 6730 19292 6736 19304
rect 5675 19264 6736 19292
rect 5675 19261 5687 19264
rect 5629 19255 5687 19261
rect 6730 19252 6736 19264
rect 6788 19252 6794 19304
rect 7742 19292 7748 19304
rect 7703 19264 7748 19292
rect 7742 19252 7748 19264
rect 7800 19252 7806 19304
rect 7852 19292 7880 19332
rect 8772 19332 10364 19360
rect 8772 19292 8800 19332
rect 10410 19320 10416 19372
rect 10468 19360 10474 19372
rect 10505 19363 10563 19369
rect 10505 19360 10517 19363
rect 10468 19332 10517 19360
rect 10468 19320 10474 19332
rect 10505 19329 10517 19332
rect 10551 19329 10563 19363
rect 10686 19360 10692 19372
rect 10647 19332 10692 19360
rect 10505 19323 10563 19329
rect 10686 19320 10692 19332
rect 10744 19320 10750 19372
rect 11882 19320 11888 19372
rect 11940 19360 11946 19372
rect 19150 19360 19156 19372
rect 11940 19332 13216 19360
rect 19111 19332 19156 19360
rect 11940 19320 11946 19332
rect 13188 19304 13216 19332
rect 19150 19320 19156 19332
rect 19208 19320 19214 19372
rect 7852 19264 8800 19292
rect 12342 19252 12348 19304
rect 12400 19292 12406 19304
rect 12710 19292 12716 19304
rect 12400 19264 12716 19292
rect 12400 19252 12406 19264
rect 12710 19252 12716 19264
rect 12768 19252 12774 19304
rect 13170 19292 13176 19304
rect 13131 19264 13176 19292
rect 13170 19252 13176 19264
rect 13228 19252 13234 19304
rect 15286 19292 15292 19304
rect 13280 19264 15292 19292
rect 5718 19224 5724 19236
rect 4080 19196 4476 19224
rect 5184 19196 5724 19224
rect 4080 19156 4108 19196
rect 2424 19128 4108 19156
rect 1949 19119 2007 19125
rect 4154 19116 4160 19168
rect 4212 19156 4218 19168
rect 5184 19165 5212 19196
rect 5718 19184 5724 19196
rect 5776 19184 5782 19236
rect 7834 19224 7840 19236
rect 5828 19196 7840 19224
rect 4249 19159 4307 19165
rect 4249 19156 4261 19159
rect 4212 19128 4261 19156
rect 4212 19116 4218 19128
rect 4249 19125 4261 19128
rect 4295 19125 4307 19159
rect 4249 19119 4307 19125
rect 5169 19159 5227 19165
rect 5169 19125 5181 19159
rect 5215 19125 5227 19159
rect 5169 19119 5227 19125
rect 5537 19159 5595 19165
rect 5537 19125 5549 19159
rect 5583 19156 5595 19159
rect 5828 19156 5856 19196
rect 7834 19184 7840 19196
rect 7892 19184 7898 19236
rect 8012 19227 8070 19233
rect 8012 19193 8024 19227
rect 8058 19224 8070 19227
rect 8202 19224 8208 19236
rect 8058 19196 8208 19224
rect 8058 19193 8070 19196
rect 8012 19187 8070 19193
rect 8202 19184 8208 19196
rect 8260 19184 8266 19236
rect 10413 19227 10471 19233
rect 10413 19193 10425 19227
rect 10459 19224 10471 19227
rect 10459 19196 12020 19224
rect 10459 19193 10471 19196
rect 10413 19187 10471 19193
rect 5583 19128 5856 19156
rect 5583 19125 5595 19128
rect 5537 19119 5595 19125
rect 5994 19116 6000 19168
rect 6052 19156 6058 19168
rect 8662 19156 8668 19168
rect 6052 19128 8668 19156
rect 6052 19116 6058 19128
rect 8662 19116 8668 19128
rect 8720 19116 8726 19168
rect 11992 19156 12020 19196
rect 12250 19184 12256 19236
rect 12308 19224 12314 19236
rect 13280 19224 13308 19264
rect 15286 19252 15292 19264
rect 15344 19252 15350 19304
rect 15378 19252 15384 19304
rect 15436 19292 15442 19304
rect 15436 19264 15481 19292
rect 15436 19252 15442 19264
rect 17862 19252 17868 19304
rect 17920 19292 17926 19304
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 17920 19264 18061 19292
rect 17920 19252 17926 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 13446 19233 13452 19236
rect 13440 19224 13452 19233
rect 12308 19196 13308 19224
rect 13407 19196 13452 19224
rect 12308 19184 12314 19196
rect 13440 19187 13452 19196
rect 13446 19184 13452 19187
rect 13504 19184 13510 19236
rect 15626 19227 15684 19233
rect 15626 19224 15638 19227
rect 14568 19196 15638 19224
rect 14568 19168 14596 19196
rect 15626 19193 15638 19196
rect 15672 19193 15684 19227
rect 15626 19187 15684 19193
rect 14182 19156 14188 19168
rect 11992 19128 14188 19156
rect 14182 19116 14188 19128
rect 14240 19116 14246 19168
rect 14550 19156 14556 19168
rect 14511 19128 14556 19156
rect 14550 19116 14556 19128
rect 14608 19116 14614 19168
rect 14642 19116 14648 19168
rect 14700 19156 14706 19168
rect 16761 19159 16819 19165
rect 16761 19156 16773 19159
rect 14700 19128 16773 19156
rect 14700 19116 14706 19128
rect 16761 19125 16773 19128
rect 16807 19125 16819 19159
rect 16761 19119 16819 19125
rect 17034 19116 17040 19168
rect 17092 19156 17098 19168
rect 18233 19159 18291 19165
rect 18233 19156 18245 19159
rect 17092 19128 18245 19156
rect 17092 19116 17098 19128
rect 18233 19125 18245 19128
rect 18279 19125 18291 19159
rect 18233 19119 18291 19125
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 2869 18955 2927 18961
rect 2869 18921 2881 18955
rect 2915 18952 2927 18955
rect 6270 18952 6276 18964
rect 2915 18924 6276 18952
rect 2915 18921 2927 18924
rect 2869 18915 2927 18921
rect 6270 18912 6276 18924
rect 6328 18912 6334 18964
rect 6822 18952 6828 18964
rect 6783 18924 6828 18952
rect 6822 18912 6828 18924
rect 6880 18912 6886 18964
rect 7650 18912 7656 18964
rect 7708 18952 7714 18964
rect 8113 18955 8171 18961
rect 8113 18952 8125 18955
rect 7708 18924 8125 18952
rect 7708 18912 7714 18924
rect 8113 18921 8125 18924
rect 8159 18921 8171 18955
rect 8113 18915 8171 18921
rect 8294 18912 8300 18964
rect 8352 18952 8358 18964
rect 12894 18952 12900 18964
rect 8352 18924 12900 18952
rect 8352 18912 8358 18924
rect 12894 18912 12900 18924
rect 12952 18912 12958 18964
rect 14366 18912 14372 18964
rect 14424 18952 14430 18964
rect 15473 18955 15531 18961
rect 15473 18952 15485 18955
rect 14424 18924 15485 18952
rect 14424 18912 14430 18924
rect 15473 18921 15485 18924
rect 15519 18921 15531 18955
rect 16574 18952 16580 18964
rect 16535 18924 16580 18952
rect 15473 18915 15531 18921
rect 16574 18912 16580 18924
rect 16632 18912 16638 18964
rect 17494 18912 17500 18964
rect 17552 18952 17558 18964
rect 17681 18955 17739 18961
rect 17681 18952 17693 18955
rect 17552 18924 17693 18952
rect 17552 18912 17558 18924
rect 17681 18921 17693 18924
rect 17727 18921 17739 18955
rect 17681 18915 17739 18921
rect 4341 18887 4399 18893
rect 4341 18853 4353 18887
rect 4387 18884 4399 18887
rect 4522 18884 4528 18896
rect 4387 18856 4528 18884
rect 4387 18853 4399 18856
rect 4341 18847 4399 18853
rect 4522 18844 4528 18856
rect 4580 18844 4586 18896
rect 5718 18893 5724 18896
rect 5712 18847 5724 18893
rect 5776 18884 5782 18896
rect 9677 18887 9735 18893
rect 5776 18856 5812 18884
rect 5718 18844 5724 18847
rect 5776 18844 5782 18856
rect 9677 18853 9689 18887
rect 9723 18884 9735 18887
rect 13265 18887 13323 18893
rect 13265 18884 13277 18887
rect 9723 18856 13277 18884
rect 9723 18853 9735 18856
rect 9677 18847 9735 18853
rect 13265 18853 13277 18856
rect 13311 18853 13323 18887
rect 13265 18847 13323 18853
rect 13722 18844 13728 18896
rect 13780 18884 13786 18896
rect 16666 18884 16672 18896
rect 13780 18856 16672 18884
rect 13780 18844 13786 18856
rect 16666 18844 16672 18856
rect 16724 18844 16730 18896
rect 2774 18776 2780 18828
rect 2832 18816 2838 18828
rect 4062 18816 4068 18828
rect 2832 18788 2877 18816
rect 4023 18788 4068 18816
rect 2832 18776 2838 18788
rect 4062 18776 4068 18788
rect 4120 18776 4126 18828
rect 6822 18776 6828 18828
rect 6880 18816 6886 18828
rect 7742 18816 7748 18828
rect 6880 18788 7748 18816
rect 6880 18776 6886 18788
rect 7742 18776 7748 18788
rect 7800 18776 7806 18828
rect 8021 18819 8079 18825
rect 8021 18785 8033 18819
rect 8067 18785 8079 18819
rect 8021 18779 8079 18785
rect 1397 18751 1455 18757
rect 1397 18717 1409 18751
rect 1443 18717 1455 18751
rect 1397 18711 1455 18717
rect 3053 18751 3111 18757
rect 3053 18717 3065 18751
rect 3099 18748 3111 18751
rect 4338 18748 4344 18760
rect 3099 18720 4344 18748
rect 3099 18717 3111 18720
rect 3053 18711 3111 18717
rect 1412 18680 1440 18711
rect 4338 18708 4344 18720
rect 4396 18708 4402 18760
rect 4982 18708 4988 18760
rect 5040 18748 5046 18760
rect 5445 18751 5503 18757
rect 5445 18748 5457 18751
rect 5040 18720 5457 18748
rect 5040 18708 5046 18720
rect 5445 18717 5457 18720
rect 5491 18717 5503 18751
rect 5445 18711 5503 18717
rect 1412 18652 5028 18680
rect 2409 18615 2467 18621
rect 2409 18581 2421 18615
rect 2455 18612 2467 18615
rect 3050 18612 3056 18624
rect 2455 18584 3056 18612
rect 2455 18581 2467 18584
rect 2409 18575 2467 18581
rect 3050 18572 3056 18584
rect 3108 18572 3114 18624
rect 5000 18612 5028 18652
rect 6914 18640 6920 18692
rect 6972 18680 6978 18692
rect 7653 18683 7711 18689
rect 7653 18680 7665 18683
rect 6972 18652 7665 18680
rect 6972 18640 6978 18652
rect 7653 18649 7665 18652
rect 7699 18649 7711 18683
rect 7653 18643 7711 18649
rect 7190 18612 7196 18624
rect 5000 18584 7196 18612
rect 7190 18572 7196 18584
rect 7248 18572 7254 18624
rect 8036 18612 8064 18779
rect 10778 18776 10784 18828
rect 10836 18816 10842 18828
rect 10945 18819 11003 18825
rect 10945 18816 10957 18819
rect 10836 18788 10957 18816
rect 10836 18776 10842 18788
rect 10945 18785 10957 18788
rect 10991 18785 11003 18819
rect 10945 18779 11003 18785
rect 12066 18776 12072 18828
rect 12124 18816 12130 18828
rect 14642 18816 14648 18828
rect 12124 18788 14648 18816
rect 12124 18776 12130 18788
rect 14642 18776 14648 18788
rect 14700 18776 14706 18828
rect 14734 18776 14740 18828
rect 14792 18816 14798 18828
rect 15289 18819 15347 18825
rect 15289 18816 15301 18819
rect 14792 18788 15301 18816
rect 14792 18776 14798 18788
rect 15289 18785 15301 18788
rect 15335 18785 15347 18819
rect 15289 18779 15347 18785
rect 15562 18776 15568 18828
rect 15620 18816 15626 18828
rect 16393 18819 16451 18825
rect 16393 18816 16405 18819
rect 15620 18788 16405 18816
rect 15620 18776 15626 18788
rect 16393 18785 16405 18788
rect 16439 18785 16451 18819
rect 17494 18816 17500 18828
rect 17455 18788 17500 18816
rect 16393 18779 16451 18785
rect 17494 18776 17500 18788
rect 17552 18776 17558 18828
rect 8297 18751 8355 18757
rect 8297 18717 8309 18751
rect 8343 18748 8355 18751
rect 9122 18748 9128 18760
rect 8343 18720 9128 18748
rect 8343 18717 8355 18720
rect 8297 18711 8355 18717
rect 9122 18708 9128 18720
rect 9180 18708 9186 18760
rect 9674 18708 9680 18760
rect 9732 18748 9738 18760
rect 9950 18748 9956 18760
rect 9732 18720 9956 18748
rect 9732 18708 9738 18720
rect 9950 18708 9956 18720
rect 10008 18748 10014 18760
rect 10689 18751 10747 18757
rect 10689 18748 10701 18751
rect 10008 18720 10701 18748
rect 10008 18708 10014 18720
rect 10689 18717 10701 18720
rect 10735 18717 10747 18751
rect 10689 18711 10747 18717
rect 12526 18708 12532 18760
rect 12584 18748 12590 18760
rect 13357 18751 13415 18757
rect 13357 18748 13369 18751
rect 12584 18720 13369 18748
rect 12584 18708 12590 18720
rect 13357 18717 13369 18720
rect 13403 18717 13415 18751
rect 13357 18711 13415 18717
rect 13541 18751 13599 18757
rect 13541 18717 13553 18751
rect 13587 18748 13599 18751
rect 14550 18748 14556 18760
rect 13587 18720 14556 18748
rect 13587 18717 13599 18720
rect 13541 18711 13599 18717
rect 14550 18708 14556 18720
rect 14608 18708 14614 18760
rect 19702 18680 19708 18692
rect 11624 18652 19708 18680
rect 11624 18612 11652 18652
rect 19702 18640 19708 18652
rect 19760 18640 19766 18692
rect 12066 18612 12072 18624
rect 8036 18584 11652 18612
rect 12027 18584 12072 18612
rect 12066 18572 12072 18584
rect 12124 18572 12130 18624
rect 12434 18572 12440 18624
rect 12492 18612 12498 18624
rect 12897 18615 12955 18621
rect 12897 18612 12909 18615
rect 12492 18584 12909 18612
rect 12492 18572 12498 18584
rect 12897 18581 12909 18584
rect 12943 18581 12955 18615
rect 12897 18575 12955 18581
rect 13078 18572 13084 18624
rect 13136 18612 13142 18624
rect 22646 18612 22652 18624
rect 13136 18584 22652 18612
rect 13136 18572 13142 18584
rect 22646 18572 22652 18584
rect 22704 18572 22710 18624
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 2958 18408 2964 18420
rect 2919 18380 2964 18408
rect 2958 18368 2964 18380
rect 3016 18368 3022 18420
rect 3142 18368 3148 18420
rect 3200 18408 3206 18420
rect 4062 18408 4068 18420
rect 3200 18380 4068 18408
rect 3200 18368 3206 18380
rect 4062 18368 4068 18380
rect 4120 18368 4126 18420
rect 4890 18368 4896 18420
rect 4948 18408 4954 18420
rect 12250 18408 12256 18420
rect 4948 18380 12256 18408
rect 4948 18368 4954 18380
rect 12250 18368 12256 18380
rect 12308 18368 12314 18420
rect 12526 18408 12532 18420
rect 12487 18380 12532 18408
rect 12526 18368 12532 18380
rect 12584 18368 12590 18420
rect 13446 18408 13452 18420
rect 13188 18380 13452 18408
rect 8570 18340 8576 18352
rect 1780 18312 8576 18340
rect 1780 18213 1808 18312
rect 8570 18300 8576 18312
rect 8628 18300 8634 18352
rect 13078 18340 13084 18352
rect 8680 18312 13084 18340
rect 1946 18232 1952 18284
rect 2004 18232 2010 18284
rect 2869 18275 2927 18281
rect 2869 18241 2881 18275
rect 2915 18272 2927 18275
rect 2958 18272 2964 18284
rect 2915 18244 2964 18272
rect 2915 18241 2927 18244
rect 2869 18235 2927 18241
rect 2958 18232 2964 18244
rect 3016 18232 3022 18284
rect 3050 18232 3056 18284
rect 3108 18272 3114 18284
rect 3421 18275 3479 18281
rect 3421 18272 3433 18275
rect 3108 18244 3433 18272
rect 3108 18232 3114 18244
rect 3421 18241 3433 18244
rect 3467 18241 3479 18275
rect 3421 18235 3479 18241
rect 3605 18275 3663 18281
rect 3605 18241 3617 18275
rect 3651 18272 3663 18275
rect 4154 18272 4160 18284
rect 3651 18244 4160 18272
rect 3651 18241 3663 18244
rect 3605 18235 3663 18241
rect 4154 18232 4160 18244
rect 4212 18232 4218 18284
rect 5169 18275 5227 18281
rect 5169 18241 5181 18275
rect 5215 18272 5227 18275
rect 5442 18272 5448 18284
rect 5215 18244 5448 18272
rect 5215 18241 5227 18244
rect 5169 18235 5227 18241
rect 5442 18232 5448 18244
rect 5500 18232 5506 18284
rect 7466 18272 7472 18284
rect 6840 18244 7328 18272
rect 7427 18244 7472 18272
rect 1765 18207 1823 18213
rect 1765 18173 1777 18207
rect 1811 18173 1823 18207
rect 1964 18204 1992 18232
rect 4890 18204 4896 18216
rect 1964 18176 4896 18204
rect 1765 18167 1823 18173
rect 4890 18164 4896 18176
rect 4948 18164 4954 18216
rect 4985 18207 5043 18213
rect 4985 18173 4997 18207
rect 5031 18204 5043 18207
rect 5626 18204 5632 18216
rect 5031 18176 5632 18204
rect 5031 18173 5043 18176
rect 4985 18167 5043 18173
rect 5626 18164 5632 18176
rect 5684 18164 5690 18216
rect 198 18096 204 18148
rect 256 18136 262 18148
rect 256 18108 2912 18136
rect 256 18096 262 18108
rect 1946 18068 1952 18080
rect 1907 18040 1952 18068
rect 1946 18028 1952 18040
rect 2004 18028 2010 18080
rect 2038 18028 2044 18080
rect 2096 18068 2102 18080
rect 2774 18068 2780 18080
rect 2096 18040 2780 18068
rect 2096 18028 2102 18040
rect 2774 18028 2780 18040
rect 2832 18028 2838 18080
rect 2884 18068 2912 18108
rect 2958 18096 2964 18148
rect 3016 18136 3022 18148
rect 3326 18136 3332 18148
rect 3016 18108 3332 18136
rect 3016 18096 3022 18108
rect 3326 18096 3332 18108
rect 3384 18096 3390 18148
rect 4706 18136 4712 18148
rect 4264 18108 4712 18136
rect 4264 18068 4292 18108
rect 4706 18096 4712 18108
rect 4764 18096 4770 18148
rect 4798 18096 4804 18148
rect 4856 18136 4862 18148
rect 6840 18136 6868 18244
rect 7190 18204 7196 18216
rect 7151 18176 7196 18204
rect 7190 18164 7196 18176
rect 7248 18164 7254 18216
rect 7300 18204 7328 18244
rect 7466 18232 7472 18244
rect 7524 18232 7530 18284
rect 8386 18232 8392 18284
rect 8444 18272 8450 18284
rect 8680 18272 8708 18312
rect 13078 18300 13084 18312
rect 13136 18300 13142 18352
rect 8444 18244 8708 18272
rect 9217 18275 9275 18281
rect 8444 18232 8450 18244
rect 9217 18241 9229 18275
rect 9263 18272 9275 18275
rect 9490 18272 9496 18284
rect 9263 18244 9496 18272
rect 9263 18241 9275 18244
rect 9217 18235 9275 18241
rect 9490 18232 9496 18244
rect 9548 18232 9554 18284
rect 10134 18232 10140 18284
rect 10192 18272 10198 18284
rect 11241 18275 11299 18281
rect 11241 18272 11253 18275
rect 10192 18244 11253 18272
rect 10192 18232 10198 18244
rect 11241 18241 11253 18244
rect 11287 18241 11299 18275
rect 11241 18235 11299 18241
rect 11425 18275 11483 18281
rect 11425 18241 11437 18275
rect 11471 18272 11483 18275
rect 12066 18272 12072 18284
rect 11471 18244 12072 18272
rect 11471 18241 11483 18244
rect 11425 18235 11483 18241
rect 12066 18232 12072 18244
rect 12124 18232 12130 18284
rect 13188 18281 13216 18380
rect 13446 18368 13452 18380
rect 13504 18408 13510 18420
rect 15657 18411 15715 18417
rect 15657 18408 15669 18411
rect 13504 18380 15669 18408
rect 13504 18368 13510 18380
rect 15657 18377 15669 18380
rect 15703 18377 15715 18411
rect 15657 18371 15715 18377
rect 13173 18275 13231 18281
rect 13173 18241 13185 18275
rect 13219 18241 13231 18275
rect 13173 18235 13231 18241
rect 14182 18232 14188 18284
rect 14240 18272 14246 18284
rect 14240 18244 14412 18272
rect 14240 18232 14246 18244
rect 7300 18176 8984 18204
rect 4856 18108 6868 18136
rect 4856 18096 4862 18108
rect 6914 18096 6920 18148
rect 6972 18136 6978 18148
rect 7285 18139 7343 18145
rect 7285 18136 7297 18139
rect 6972 18108 7297 18136
rect 6972 18096 6978 18108
rect 7285 18105 7297 18108
rect 7331 18105 7343 18139
rect 8956 18136 8984 18176
rect 9030 18164 9036 18216
rect 9088 18204 9094 18216
rect 10042 18204 10048 18216
rect 9088 18176 10048 18204
rect 9088 18164 9094 18176
rect 10042 18164 10048 18176
rect 10100 18164 10106 18216
rect 10962 18164 10968 18216
rect 11020 18204 11026 18216
rect 12989 18207 13047 18213
rect 12989 18204 13001 18207
rect 11020 18176 13001 18204
rect 11020 18164 11026 18176
rect 12989 18173 13001 18176
rect 13035 18173 13047 18207
rect 12989 18167 13047 18173
rect 13630 18164 13636 18216
rect 13688 18204 13694 18216
rect 14277 18207 14335 18213
rect 14277 18204 14289 18207
rect 13688 18176 14289 18204
rect 13688 18164 13694 18176
rect 14277 18173 14289 18176
rect 14323 18173 14335 18207
rect 14384 18204 14412 18244
rect 16485 18207 16543 18213
rect 16485 18204 16497 18207
rect 14384 18176 16497 18204
rect 14277 18167 14335 18173
rect 16485 18173 16497 18176
rect 16531 18173 16543 18207
rect 16485 18167 16543 18173
rect 10870 18136 10876 18148
rect 8956 18108 10876 18136
rect 7285 18099 7343 18105
rect 10870 18096 10876 18108
rect 10928 18096 10934 18148
rect 11146 18136 11152 18148
rect 11107 18108 11152 18136
rect 11146 18096 11152 18108
rect 11204 18096 11210 18148
rect 11882 18096 11888 18148
rect 11940 18136 11946 18148
rect 12897 18139 12955 18145
rect 12897 18136 12909 18139
rect 11940 18108 12909 18136
rect 11940 18096 11946 18108
rect 12897 18105 12909 18108
rect 12943 18105 12955 18139
rect 12897 18099 12955 18105
rect 2884 18040 4292 18068
rect 4338 18028 4344 18080
rect 4396 18068 4402 18080
rect 4525 18071 4583 18077
rect 4525 18068 4537 18071
rect 4396 18040 4537 18068
rect 4396 18028 4402 18040
rect 4525 18037 4537 18040
rect 4571 18037 4583 18071
rect 4525 18031 4583 18037
rect 4893 18071 4951 18077
rect 4893 18037 4905 18071
rect 4939 18068 4951 18071
rect 5258 18068 5264 18080
rect 4939 18040 5264 18068
rect 4939 18037 4951 18040
rect 4893 18031 4951 18037
rect 5258 18028 5264 18040
rect 5316 18028 5322 18080
rect 5534 18028 5540 18080
rect 5592 18068 5598 18080
rect 6825 18071 6883 18077
rect 6825 18068 6837 18071
rect 5592 18040 6837 18068
rect 5592 18028 5598 18040
rect 6825 18037 6837 18040
rect 6871 18037 6883 18071
rect 8570 18068 8576 18080
rect 8531 18040 8576 18068
rect 6825 18031 6883 18037
rect 8570 18028 8576 18040
rect 8628 18028 8634 18080
rect 8938 18068 8944 18080
rect 8899 18040 8944 18068
rect 8938 18028 8944 18040
rect 8996 18028 9002 18080
rect 9033 18071 9091 18077
rect 9033 18037 9045 18071
rect 9079 18068 9091 18071
rect 9674 18068 9680 18080
rect 9079 18040 9680 18068
rect 9079 18037 9091 18040
rect 9033 18031 9091 18037
rect 9674 18028 9680 18040
rect 9732 18028 9738 18080
rect 10781 18071 10839 18077
rect 10781 18037 10793 18071
rect 10827 18068 10839 18071
rect 11054 18068 11060 18080
rect 10827 18040 11060 18068
rect 10827 18037 10839 18040
rect 10781 18031 10839 18037
rect 11054 18028 11060 18040
rect 11112 18028 11118 18080
rect 11698 18028 11704 18080
rect 11756 18068 11762 18080
rect 13262 18068 13268 18080
rect 11756 18040 13268 18068
rect 11756 18028 11762 18040
rect 13262 18028 13268 18040
rect 13320 18028 13326 18080
rect 14292 18068 14320 18167
rect 19610 18164 19616 18216
rect 19668 18204 19674 18216
rect 21266 18204 21272 18216
rect 19668 18176 21272 18204
rect 19668 18164 19674 18176
rect 21266 18164 21272 18176
rect 21324 18164 21330 18216
rect 14544 18139 14602 18145
rect 14544 18105 14556 18139
rect 14590 18136 14602 18139
rect 15470 18136 15476 18148
rect 14590 18108 15476 18136
rect 14590 18105 14602 18108
rect 14544 18099 14602 18105
rect 15470 18096 15476 18108
rect 15528 18096 15534 18148
rect 15654 18096 15660 18148
rect 15712 18136 15718 18148
rect 16758 18136 16764 18148
rect 15712 18108 16764 18136
rect 15712 18096 15718 18108
rect 16758 18096 16764 18108
rect 16816 18096 16822 18148
rect 18046 18136 18052 18148
rect 18007 18108 18052 18136
rect 18046 18096 18052 18108
rect 18104 18136 18110 18148
rect 18325 18139 18383 18145
rect 18325 18136 18337 18139
rect 18104 18108 18337 18136
rect 18104 18096 18110 18108
rect 18325 18105 18337 18108
rect 18371 18105 18383 18139
rect 18325 18099 18383 18105
rect 21082 18096 21088 18148
rect 21140 18136 21146 18148
rect 22186 18136 22192 18148
rect 21140 18108 22192 18136
rect 21140 18096 21146 18108
rect 22186 18096 22192 18108
rect 22244 18096 22250 18148
rect 15378 18068 15384 18080
rect 14292 18040 15384 18068
rect 15378 18028 15384 18040
rect 15436 18028 15442 18080
rect 17954 18028 17960 18080
rect 18012 18068 18018 18080
rect 18966 18068 18972 18080
rect 18012 18040 18972 18068
rect 18012 18028 18018 18040
rect 18966 18028 18972 18040
rect 19024 18028 19030 18080
rect 19702 18028 19708 18080
rect 19760 18068 19766 18080
rect 20346 18068 20352 18080
rect 19760 18040 20352 18068
rect 19760 18028 19766 18040
rect 20346 18028 20352 18040
rect 20404 18028 20410 18080
rect 20714 18028 20720 18080
rect 20772 18068 20778 18080
rect 21726 18068 21732 18080
rect 20772 18040 21732 18068
rect 20772 18028 20778 18040
rect 21726 18028 21732 18040
rect 21784 18028 21790 18080
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 2498 17824 2504 17876
rect 2556 17864 2562 17876
rect 7006 17864 7012 17876
rect 2556 17836 7012 17864
rect 2556 17824 2562 17836
rect 7006 17824 7012 17836
rect 7064 17824 7070 17876
rect 8202 17864 8208 17876
rect 8163 17836 8208 17864
rect 8202 17824 8208 17836
rect 8260 17824 8266 17876
rect 9674 17864 9680 17876
rect 9635 17836 9680 17864
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 9766 17824 9772 17876
rect 9824 17864 9830 17876
rect 10137 17867 10195 17873
rect 10137 17864 10149 17867
rect 9824 17836 10149 17864
rect 9824 17824 9830 17836
rect 10137 17833 10149 17836
rect 10183 17833 10195 17867
rect 10137 17827 10195 17833
rect 11241 17867 11299 17873
rect 11241 17833 11253 17867
rect 11287 17864 11299 17867
rect 13170 17864 13176 17876
rect 11287 17836 13176 17864
rect 11287 17833 11299 17836
rect 11241 17827 11299 17833
rect 1394 17756 1400 17808
rect 1452 17796 1458 17808
rect 1452 17768 10732 17796
rect 1452 17756 1458 17768
rect 2222 17728 2228 17740
rect 2183 17700 2228 17728
rect 2222 17688 2228 17700
rect 2280 17688 2286 17740
rect 4154 17688 4160 17740
rect 4212 17728 4218 17740
rect 4321 17731 4379 17737
rect 4321 17728 4333 17731
rect 4212 17700 4333 17728
rect 4212 17688 4218 17700
rect 4321 17697 4333 17700
rect 4367 17697 4379 17731
rect 4321 17691 4379 17697
rect 7092 17731 7150 17737
rect 7092 17697 7104 17731
rect 7138 17728 7150 17731
rect 7466 17728 7472 17740
rect 7138 17700 7472 17728
rect 7138 17697 7150 17700
rect 7092 17691 7150 17697
rect 7466 17688 7472 17700
rect 7524 17728 7530 17740
rect 8202 17728 8208 17740
rect 7524 17700 8208 17728
rect 7524 17688 7530 17700
rect 8202 17688 8208 17700
rect 8260 17688 8266 17740
rect 10045 17731 10103 17737
rect 10045 17697 10057 17731
rect 10091 17728 10103 17731
rect 10134 17728 10140 17740
rect 10091 17700 10140 17728
rect 10091 17697 10103 17700
rect 10045 17691 10103 17697
rect 10134 17688 10140 17700
rect 10192 17688 10198 17740
rect 2406 17660 2412 17672
rect 2367 17632 2412 17660
rect 2406 17620 2412 17632
rect 2464 17620 2470 17672
rect 4065 17663 4123 17669
rect 4065 17629 4077 17663
rect 4111 17629 4123 17663
rect 6822 17660 6828 17672
rect 6783 17632 6828 17660
rect 4065 17623 4123 17629
rect 4080 17536 4108 17623
rect 6822 17620 6828 17632
rect 6880 17620 6886 17672
rect 10318 17660 10324 17672
rect 10231 17632 10324 17660
rect 10318 17620 10324 17632
rect 10376 17660 10382 17672
rect 10704 17660 10732 17768
rect 11146 17688 11152 17740
rect 11204 17728 11210 17740
rect 11532 17737 11560 17836
rect 13170 17824 13176 17836
rect 13228 17864 13234 17876
rect 13630 17864 13636 17876
rect 13228 17836 13636 17864
rect 13228 17824 13234 17836
rect 13630 17824 13636 17836
rect 13688 17824 13694 17876
rect 15565 17799 15623 17805
rect 15565 17796 15577 17799
rect 11624 17768 15577 17796
rect 11425 17731 11483 17737
rect 11425 17728 11437 17731
rect 11204 17700 11437 17728
rect 11204 17688 11210 17700
rect 11425 17697 11437 17700
rect 11471 17697 11483 17731
rect 11425 17691 11483 17697
rect 11517 17731 11575 17737
rect 11517 17697 11529 17731
rect 11563 17697 11575 17731
rect 11517 17691 11575 17697
rect 11624 17660 11652 17768
rect 15565 17765 15577 17768
rect 15611 17765 15623 17799
rect 15565 17759 15623 17765
rect 11784 17731 11842 17737
rect 11784 17697 11796 17731
rect 11830 17728 11842 17731
rect 12986 17728 12992 17740
rect 11830 17700 12992 17728
rect 11830 17697 11842 17700
rect 11784 17691 11842 17697
rect 12986 17688 12992 17700
rect 13044 17688 13050 17740
rect 13722 17728 13728 17740
rect 13683 17700 13728 17728
rect 13722 17688 13728 17700
rect 13780 17688 13786 17740
rect 15286 17728 15292 17740
rect 15247 17700 15292 17728
rect 15286 17688 15292 17700
rect 15344 17688 15350 17740
rect 13906 17660 13912 17672
rect 10376 17632 10640 17660
rect 10704 17632 11652 17660
rect 13867 17632 13912 17660
rect 10376 17620 10382 17632
rect 3142 17484 3148 17536
rect 3200 17524 3206 17536
rect 3878 17524 3884 17536
rect 3200 17496 3884 17524
rect 3200 17484 3206 17496
rect 3878 17484 3884 17496
rect 3936 17484 3942 17536
rect 4062 17524 4068 17536
rect 3975 17496 4068 17524
rect 4062 17484 4068 17496
rect 4120 17524 4126 17536
rect 4982 17524 4988 17536
rect 4120 17496 4988 17524
rect 4120 17484 4126 17496
rect 4982 17484 4988 17496
rect 5040 17484 5046 17536
rect 5442 17524 5448 17536
rect 5403 17496 5448 17524
rect 5442 17484 5448 17496
rect 5500 17484 5506 17536
rect 10612 17524 10640 17632
rect 13906 17620 13912 17632
rect 13964 17620 13970 17672
rect 13998 17620 14004 17672
rect 14056 17660 14062 17672
rect 16577 17663 16635 17669
rect 16577 17660 16589 17663
rect 14056 17632 16589 17660
rect 14056 17620 14062 17632
rect 16577 17629 16589 17632
rect 16623 17629 16635 17663
rect 16577 17623 16635 17629
rect 12897 17527 12955 17533
rect 12897 17524 12909 17527
rect 10612 17496 12909 17524
rect 12897 17493 12909 17496
rect 12943 17493 12955 17527
rect 12897 17487 12955 17493
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 3970 17280 3976 17332
rect 4028 17320 4034 17332
rect 7742 17320 7748 17332
rect 4028 17292 7748 17320
rect 4028 17280 4034 17292
rect 7742 17280 7748 17292
rect 7800 17280 7806 17332
rect 8202 17320 8208 17332
rect 8163 17292 8208 17320
rect 8202 17280 8208 17292
rect 8260 17280 8266 17332
rect 9950 17320 9956 17332
rect 9048 17292 9956 17320
rect 4982 17212 4988 17264
rect 5040 17252 5046 17264
rect 6181 17255 6239 17261
rect 6181 17252 6193 17255
rect 5040 17224 6193 17252
rect 5040 17212 5046 17224
rect 6181 17221 6193 17224
rect 6227 17252 6239 17255
rect 6822 17252 6828 17264
rect 6227 17224 6828 17252
rect 6227 17221 6239 17224
rect 6181 17215 6239 17221
rect 6822 17212 6828 17224
rect 6880 17212 6886 17264
rect 2409 17187 2467 17193
rect 2409 17153 2421 17187
rect 2455 17184 2467 17187
rect 2498 17184 2504 17196
rect 2455 17156 2504 17184
rect 2455 17153 2467 17156
rect 2409 17147 2467 17153
rect 2498 17144 2504 17156
rect 2556 17144 2562 17196
rect 3970 17184 3976 17196
rect 3931 17156 3976 17184
rect 3970 17144 3976 17156
rect 4028 17144 4034 17196
rect 8478 17144 8484 17196
rect 8536 17184 8542 17196
rect 9048 17193 9076 17292
rect 9950 17280 9956 17292
rect 10008 17280 10014 17332
rect 11238 17280 11244 17332
rect 11296 17320 11302 17332
rect 11425 17323 11483 17329
rect 11425 17320 11437 17323
rect 11296 17292 11437 17320
rect 11296 17280 11302 17292
rect 11425 17289 11437 17292
rect 11471 17289 11483 17323
rect 11425 17283 11483 17289
rect 12437 17323 12495 17329
rect 12437 17289 12449 17323
rect 12483 17320 12495 17323
rect 15286 17320 15292 17332
rect 12483 17292 15292 17320
rect 12483 17289 12495 17292
rect 12437 17283 12495 17289
rect 15286 17280 15292 17292
rect 15344 17280 15350 17332
rect 15470 17320 15476 17332
rect 15431 17292 15476 17320
rect 15470 17280 15476 17292
rect 15528 17280 15534 17332
rect 12618 17252 12624 17264
rect 10428 17224 12624 17252
rect 9033 17187 9091 17193
rect 9033 17184 9045 17187
rect 8536 17156 9045 17184
rect 8536 17144 8542 17156
rect 9033 17153 9045 17156
rect 9079 17153 9091 17187
rect 9033 17147 9091 17153
rect 2133 17119 2191 17125
rect 2133 17085 2145 17119
rect 2179 17085 2191 17119
rect 2133 17079 2191 17085
rect 4240 17119 4298 17125
rect 4240 17085 4252 17119
rect 4286 17116 4298 17119
rect 5442 17116 5448 17128
rect 4286 17088 5448 17116
rect 4286 17085 4298 17088
rect 4240 17079 4298 17085
rect 2148 17048 2176 17079
rect 5442 17076 5448 17088
rect 5500 17076 5506 17128
rect 6178 17076 6184 17128
rect 6236 17116 6242 17128
rect 6365 17119 6423 17125
rect 6365 17116 6377 17119
rect 6236 17088 6377 17116
rect 6236 17076 6242 17088
rect 6365 17085 6377 17088
rect 6411 17085 6423 17119
rect 6822 17116 6828 17128
rect 6783 17088 6828 17116
rect 6365 17079 6423 17085
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 8570 17116 8576 17128
rect 6932 17088 8576 17116
rect 5534 17048 5540 17060
rect 2148 17020 5540 17048
rect 5534 17008 5540 17020
rect 5592 17008 5598 17060
rect 6932 17048 6960 17088
rect 8570 17076 8576 17088
rect 8628 17076 8634 17128
rect 9300 17119 9358 17125
rect 9300 17085 9312 17119
rect 9346 17116 9358 17119
rect 10318 17116 10324 17128
rect 9346 17088 10324 17116
rect 9346 17085 9358 17088
rect 9300 17079 9358 17085
rect 10318 17076 10324 17088
rect 10376 17076 10382 17128
rect 5644 17020 6960 17048
rect 7092 17051 7150 17057
rect 4706 16940 4712 16992
rect 4764 16980 4770 16992
rect 5353 16983 5411 16989
rect 5353 16980 5365 16983
rect 4764 16952 5365 16980
rect 4764 16940 4770 16952
rect 5353 16949 5365 16952
rect 5399 16949 5411 16983
rect 5353 16943 5411 16949
rect 5442 16940 5448 16992
rect 5500 16980 5506 16992
rect 5644 16980 5672 17020
rect 7092 17017 7104 17051
rect 7138 17048 7150 17051
rect 7466 17048 7472 17060
rect 7138 17020 7472 17048
rect 7138 17017 7150 17020
rect 7092 17011 7150 17017
rect 7466 17008 7472 17020
rect 7524 17008 7530 17060
rect 10428 17048 10456 17224
rect 12618 17212 12624 17224
rect 12676 17212 12682 17264
rect 20806 17212 20812 17264
rect 20864 17252 20870 17264
rect 21082 17252 21088 17264
rect 20864 17224 21088 17252
rect 20864 17212 20870 17224
rect 21082 17212 21088 17224
rect 21140 17212 21146 17264
rect 12986 17184 12992 17196
rect 12947 17156 12992 17184
rect 12986 17144 12992 17156
rect 13044 17144 13050 17196
rect 13630 17144 13636 17196
rect 13688 17184 13694 17196
rect 14093 17187 14151 17193
rect 14093 17184 14105 17187
rect 13688 17156 14105 17184
rect 13688 17144 13694 17156
rect 14093 17153 14105 17156
rect 14139 17153 14151 17187
rect 14093 17147 14151 17153
rect 10870 17076 10876 17128
rect 10928 17116 10934 17128
rect 11241 17119 11299 17125
rect 11241 17116 11253 17119
rect 10928 17088 11253 17116
rect 10928 17076 10934 17088
rect 11241 17085 11253 17088
rect 11287 17085 11299 17119
rect 11241 17079 11299 17085
rect 12805 17119 12863 17125
rect 12805 17085 12817 17119
rect 12851 17116 12863 17119
rect 13998 17116 14004 17128
rect 12851 17088 14004 17116
rect 12851 17085 12863 17088
rect 12805 17079 12863 17085
rect 13998 17076 14004 17088
rect 14056 17076 14062 17128
rect 9416 17020 10456 17048
rect 5500 16952 5672 16980
rect 5500 16940 5506 16952
rect 7006 16940 7012 16992
rect 7064 16980 7070 16992
rect 9416 16980 9444 17020
rect 11054 17008 11060 17060
rect 11112 17048 11118 17060
rect 14366 17057 14372 17060
rect 12897 17051 12955 17057
rect 12897 17048 12909 17051
rect 11112 17020 12909 17048
rect 11112 17008 11118 17020
rect 12897 17017 12909 17020
rect 12943 17017 12955 17051
rect 14360 17048 14372 17057
rect 14327 17020 14372 17048
rect 12897 17011 12955 17017
rect 14360 17011 14372 17020
rect 14366 17008 14372 17011
rect 14424 17008 14430 17060
rect 7064 16952 9444 16980
rect 7064 16940 7070 16952
rect 9490 16940 9496 16992
rect 9548 16980 9554 16992
rect 10413 16983 10471 16989
rect 10413 16980 10425 16983
rect 9548 16952 10425 16980
rect 9548 16940 9554 16952
rect 10413 16949 10425 16952
rect 10459 16949 10471 16983
rect 10413 16943 10471 16949
rect 15654 16940 15660 16992
rect 15712 16980 15718 16992
rect 16301 16983 16359 16989
rect 16301 16980 16313 16983
rect 15712 16952 16313 16980
rect 15712 16940 15718 16952
rect 16301 16949 16313 16952
rect 16347 16949 16359 16983
rect 16301 16943 16359 16949
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 2222 16736 2228 16788
rect 2280 16776 2286 16788
rect 4065 16779 4123 16785
rect 4065 16776 4077 16779
rect 2280 16748 4077 16776
rect 2280 16736 2286 16748
rect 4065 16745 4077 16748
rect 4111 16745 4123 16779
rect 4065 16739 4123 16745
rect 4338 16736 4344 16788
rect 4396 16776 4402 16788
rect 4525 16779 4583 16785
rect 4525 16776 4537 16779
rect 4396 16748 4537 16776
rect 4396 16736 4402 16748
rect 4525 16745 4537 16748
rect 4571 16745 4583 16779
rect 4525 16739 4583 16745
rect 6825 16779 6883 16785
rect 6825 16745 6837 16779
rect 6871 16776 6883 16779
rect 6914 16776 6920 16788
rect 6871 16748 6920 16776
rect 6871 16745 6883 16748
rect 6825 16739 6883 16745
rect 6914 16736 6920 16748
rect 6972 16736 6978 16788
rect 7285 16779 7343 16785
rect 7285 16745 7297 16779
rect 7331 16776 7343 16779
rect 7558 16776 7564 16788
rect 7331 16748 7564 16776
rect 7331 16745 7343 16748
rect 7285 16739 7343 16745
rect 7558 16736 7564 16748
rect 7616 16736 7622 16788
rect 7742 16736 7748 16788
rect 7800 16776 7806 16788
rect 8573 16779 8631 16785
rect 8573 16776 8585 16779
rect 7800 16748 8585 16776
rect 7800 16736 7806 16748
rect 8573 16745 8585 16748
rect 8619 16745 8631 16779
rect 9674 16776 9680 16788
rect 8573 16739 8631 16745
rect 9508 16748 9680 16776
rect 4433 16711 4491 16717
rect 2148 16680 4384 16708
rect 2148 16649 2176 16680
rect 2133 16643 2191 16649
rect 2133 16609 2145 16643
rect 2179 16609 2191 16643
rect 2133 16603 2191 16609
rect 2409 16643 2467 16649
rect 2409 16609 2421 16643
rect 2455 16640 2467 16643
rect 3602 16640 3608 16652
rect 2455 16612 3608 16640
rect 2455 16609 2467 16612
rect 2409 16603 2467 16609
rect 3602 16600 3608 16612
rect 3660 16600 3666 16652
rect 4356 16640 4384 16680
rect 4433 16677 4445 16711
rect 4479 16708 4491 16711
rect 9508 16708 9536 16748
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 9950 16736 9956 16788
rect 10008 16776 10014 16788
rect 10965 16779 11023 16785
rect 10965 16776 10977 16779
rect 10008 16748 10977 16776
rect 10008 16736 10014 16748
rect 10965 16745 10977 16748
rect 11011 16776 11023 16779
rect 12621 16779 12679 16785
rect 11011 16748 11284 16776
rect 11011 16745 11023 16748
rect 10965 16739 11023 16745
rect 4479 16680 9536 16708
rect 4479 16677 4491 16680
rect 4433 16671 4491 16677
rect 5442 16640 5448 16652
rect 4356 16612 5448 16640
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 5629 16643 5687 16649
rect 5629 16609 5641 16643
rect 5675 16640 5687 16643
rect 7006 16640 7012 16652
rect 5675 16612 7012 16640
rect 5675 16609 5687 16612
rect 5629 16603 5687 16609
rect 7006 16600 7012 16612
rect 7064 16600 7070 16652
rect 7193 16643 7251 16649
rect 7193 16609 7205 16643
rect 7239 16609 7251 16643
rect 7193 16603 7251 16609
rect 4338 16532 4344 16584
rect 4396 16572 4402 16584
rect 4706 16572 4712 16584
rect 4396 16544 4712 16572
rect 4396 16532 4402 16544
rect 4706 16532 4712 16544
rect 4764 16532 4770 16584
rect 7208 16504 7236 16603
rect 7374 16600 7380 16652
rect 7432 16640 7438 16652
rect 8389 16643 8447 16649
rect 8389 16640 8401 16643
rect 7432 16612 8401 16640
rect 7432 16600 7438 16612
rect 8389 16609 8401 16612
rect 8435 16609 8447 16643
rect 9677 16643 9735 16649
rect 8389 16603 8447 16609
rect 8496 16612 9628 16640
rect 7466 16572 7472 16584
rect 7427 16544 7472 16572
rect 7466 16532 7472 16544
rect 7524 16532 7530 16584
rect 8202 16532 8208 16584
rect 8260 16572 8266 16584
rect 8496 16572 8524 16612
rect 8260 16544 8524 16572
rect 9600 16572 9628 16612
rect 9677 16609 9689 16643
rect 9723 16640 9735 16643
rect 11146 16640 11152 16652
rect 9723 16612 11008 16640
rect 11107 16612 11152 16640
rect 9723 16609 9735 16612
rect 9677 16603 9735 16609
rect 9861 16575 9919 16581
rect 9861 16572 9873 16575
rect 9600 16544 9873 16572
rect 8260 16532 8266 16544
rect 9861 16541 9873 16544
rect 9907 16541 9919 16575
rect 10980 16572 11008 16612
rect 11146 16600 11152 16612
rect 11204 16600 11210 16652
rect 11256 16649 11284 16748
rect 12621 16745 12633 16779
rect 12667 16776 12679 16779
rect 12986 16776 12992 16788
rect 12667 16748 12992 16776
rect 12667 16745 12679 16748
rect 12621 16739 12679 16745
rect 12986 16736 12992 16748
rect 13044 16736 13050 16788
rect 13633 16779 13691 16785
rect 13633 16745 13645 16779
rect 13679 16745 13691 16779
rect 13633 16739 13691 16745
rect 11508 16711 11566 16717
rect 11508 16677 11520 16711
rect 11554 16708 11566 16711
rect 12066 16708 12072 16720
rect 11554 16680 12072 16708
rect 11554 16677 11566 16680
rect 11508 16671 11566 16677
rect 12066 16668 12072 16680
rect 12124 16668 12130 16720
rect 13648 16708 13676 16739
rect 13722 16736 13728 16788
rect 13780 16776 13786 16788
rect 15289 16779 15347 16785
rect 15289 16776 15301 16779
rect 13780 16748 15301 16776
rect 13780 16736 13786 16748
rect 15289 16745 15301 16748
rect 15335 16745 15347 16779
rect 15654 16776 15660 16788
rect 15615 16748 15660 16776
rect 15289 16739 15347 16745
rect 15654 16736 15660 16748
rect 15712 16736 15718 16788
rect 15749 16711 15807 16717
rect 15749 16708 15761 16711
rect 13648 16680 15761 16708
rect 15749 16677 15761 16680
rect 15795 16677 15807 16711
rect 15749 16671 15807 16677
rect 11241 16643 11299 16649
rect 11241 16609 11253 16643
rect 11287 16609 11299 16643
rect 11241 16603 11299 16609
rect 13262 16600 13268 16652
rect 13320 16640 13326 16652
rect 13998 16640 14004 16652
rect 13320 16612 13860 16640
rect 13959 16612 14004 16640
rect 13320 16600 13326 16612
rect 13832 16572 13860 16612
rect 13998 16600 14004 16612
rect 14056 16600 14062 16652
rect 14093 16643 14151 16649
rect 14093 16609 14105 16643
rect 14139 16609 14151 16643
rect 14093 16603 14151 16609
rect 14108 16572 14136 16603
rect 10980 16544 11284 16572
rect 13832 16544 14136 16572
rect 14277 16575 14335 16581
rect 9861 16535 9919 16541
rect 7558 16504 7564 16516
rect 7208 16476 7564 16504
rect 7558 16464 7564 16476
rect 7616 16464 7622 16516
rect 4062 16396 4068 16448
rect 4120 16436 4126 16448
rect 5813 16439 5871 16445
rect 5813 16436 5825 16439
rect 4120 16408 5825 16436
rect 4120 16396 4126 16408
rect 5813 16405 5825 16408
rect 5859 16405 5871 16439
rect 11256 16436 11284 16544
rect 14277 16541 14289 16575
rect 14323 16572 14335 16575
rect 14366 16572 14372 16584
rect 14323 16544 14372 16572
rect 14323 16541 14335 16544
rect 14277 16535 14335 16541
rect 14366 16532 14372 16544
rect 14424 16572 14430 16584
rect 15102 16572 15108 16584
rect 14424 16544 15108 16572
rect 14424 16532 14430 16544
rect 15102 16532 15108 16544
rect 15160 16532 15166 16584
rect 15470 16532 15476 16584
rect 15528 16572 15534 16584
rect 15841 16575 15899 16581
rect 15841 16572 15853 16575
rect 15528 16544 15853 16572
rect 15528 16532 15534 16544
rect 15841 16541 15853 16544
rect 15887 16541 15899 16575
rect 15841 16535 15899 16541
rect 12158 16436 12164 16448
rect 11256 16408 12164 16436
rect 5813 16399 5871 16405
rect 12158 16396 12164 16408
rect 12216 16396 12222 16448
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 6825 16235 6883 16241
rect 6825 16232 6837 16235
rect 2148 16204 6837 16232
rect 2148 16037 2176 16204
rect 6825 16201 6837 16204
rect 6871 16201 6883 16235
rect 6825 16195 6883 16201
rect 9674 16192 9680 16244
rect 9732 16232 9738 16244
rect 15102 16232 15108 16244
rect 9732 16204 14688 16232
rect 15063 16204 15108 16232
rect 9732 16192 9738 16204
rect 9582 16124 9588 16176
rect 9640 16164 9646 16176
rect 9861 16167 9919 16173
rect 9861 16164 9873 16167
rect 9640 16136 9873 16164
rect 9640 16124 9646 16136
rect 9861 16133 9873 16136
rect 9907 16133 9919 16167
rect 14660 16164 14688 16204
rect 15102 16192 15108 16204
rect 15160 16192 15166 16244
rect 14660 16136 15976 16164
rect 9861 16127 9919 16133
rect 2866 16056 2872 16108
rect 2924 16096 2930 16108
rect 3786 16096 3792 16108
rect 2924 16068 3792 16096
rect 2924 16056 2930 16068
rect 3786 16056 3792 16068
rect 3844 16056 3850 16108
rect 7469 16099 7527 16105
rect 7469 16065 7481 16099
rect 7515 16096 7527 16099
rect 8294 16096 8300 16108
rect 7515 16068 8300 16096
rect 7515 16065 7527 16068
rect 7469 16059 7527 16065
rect 8294 16056 8300 16068
rect 8352 16056 8358 16108
rect 8478 16096 8484 16108
rect 8439 16068 8484 16096
rect 8478 16056 8484 16068
rect 8536 16056 8542 16108
rect 11425 16099 11483 16105
rect 11425 16065 11437 16099
rect 11471 16096 11483 16099
rect 11698 16096 11704 16108
rect 11471 16068 11704 16096
rect 11471 16065 11483 16068
rect 11425 16059 11483 16065
rect 11698 16056 11704 16068
rect 11756 16056 11762 16108
rect 12618 16096 12624 16108
rect 12579 16068 12624 16096
rect 12618 16056 12624 16068
rect 12676 16056 12682 16108
rect 15948 16105 15976 16136
rect 15933 16099 15991 16105
rect 15933 16065 15945 16099
rect 15979 16065 15991 16099
rect 15933 16059 15991 16065
rect 2133 16031 2191 16037
rect 2133 15997 2145 16031
rect 2179 15997 2191 16031
rect 2133 15991 2191 15997
rect 4056 16031 4114 16037
rect 4056 15997 4068 16031
rect 4102 16028 4114 16031
rect 4338 16028 4344 16040
rect 4102 16000 4344 16028
rect 4102 15997 4114 16000
rect 4056 15991 4114 15997
rect 4338 15988 4344 16000
rect 4396 15988 4402 16040
rect 8748 16031 8806 16037
rect 8748 15997 8760 16031
rect 8794 16028 8806 16031
rect 9490 16028 9496 16040
rect 8794 16000 9496 16028
rect 8794 15997 8806 16000
rect 8748 15991 8806 15997
rect 9490 15988 9496 16000
rect 9548 15988 9554 16040
rect 12434 15988 12440 16040
rect 12492 16028 12498 16040
rect 13722 16028 13728 16040
rect 12492 16000 12537 16028
rect 13683 16000 13728 16028
rect 12492 15988 12498 16000
rect 13722 15988 13728 16000
rect 13780 15988 13786 16040
rect 2409 15963 2467 15969
rect 2409 15929 2421 15963
rect 2455 15960 2467 15963
rect 7374 15960 7380 15972
rect 2455 15932 7380 15960
rect 2455 15929 2467 15932
rect 2409 15923 2467 15929
rect 7374 15920 7380 15932
rect 7432 15920 7438 15972
rect 13538 15960 13544 15972
rect 10796 15932 13544 15960
rect 5166 15892 5172 15904
rect 5127 15864 5172 15892
rect 5166 15852 5172 15864
rect 5224 15852 5230 15904
rect 6914 15852 6920 15904
rect 6972 15892 6978 15904
rect 7193 15895 7251 15901
rect 7193 15892 7205 15895
rect 6972 15864 7205 15892
rect 6972 15852 6978 15864
rect 7193 15861 7205 15864
rect 7239 15861 7251 15895
rect 7193 15855 7251 15861
rect 7285 15895 7343 15901
rect 7285 15861 7297 15895
rect 7331 15892 7343 15895
rect 9674 15892 9680 15904
rect 7331 15864 9680 15892
rect 7331 15861 7343 15864
rect 7285 15855 7343 15861
rect 9674 15852 9680 15864
rect 9732 15852 9738 15904
rect 10796 15901 10824 15932
rect 13538 15920 13544 15932
rect 13596 15920 13602 15972
rect 13998 15969 14004 15972
rect 13992 15960 14004 15969
rect 13959 15932 14004 15960
rect 13992 15923 14004 15932
rect 13998 15920 14004 15923
rect 14056 15920 14062 15972
rect 10781 15895 10839 15901
rect 10781 15861 10793 15895
rect 10827 15861 10839 15895
rect 10781 15855 10839 15861
rect 11054 15852 11060 15904
rect 11112 15892 11118 15904
rect 11149 15895 11207 15901
rect 11149 15892 11161 15895
rect 11112 15864 11161 15892
rect 11112 15852 11118 15864
rect 11149 15861 11161 15864
rect 11195 15861 11207 15895
rect 11149 15855 11207 15861
rect 11238 15852 11244 15904
rect 11296 15892 11302 15904
rect 11296 15864 11341 15892
rect 11296 15852 11302 15864
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 7466 15648 7472 15700
rect 7524 15688 7530 15700
rect 8481 15691 8539 15697
rect 8481 15688 8493 15691
rect 7524 15660 8493 15688
rect 7524 15648 7530 15660
rect 8481 15657 8493 15660
rect 8527 15657 8539 15691
rect 9674 15688 9680 15700
rect 9635 15660 9680 15688
rect 8481 15651 8539 15657
rect 9674 15648 9680 15660
rect 9732 15648 9738 15700
rect 10042 15648 10048 15700
rect 10100 15688 10106 15700
rect 10137 15691 10195 15697
rect 10137 15688 10149 15691
rect 10100 15660 10149 15688
rect 10100 15648 10106 15660
rect 10137 15657 10149 15660
rect 10183 15657 10195 15691
rect 10137 15651 10195 15657
rect 11146 15648 11152 15700
rect 11204 15688 11210 15700
rect 11333 15691 11391 15697
rect 11333 15688 11345 15691
rect 11204 15660 11345 15688
rect 11204 15648 11210 15660
rect 11333 15657 11345 15660
rect 11379 15657 11391 15691
rect 11333 15651 11391 15657
rect 11974 15648 11980 15700
rect 12032 15688 12038 15700
rect 12069 15691 12127 15697
rect 12069 15688 12081 15691
rect 12032 15660 12081 15688
rect 12032 15648 12038 15660
rect 12069 15657 12081 15660
rect 12115 15657 12127 15691
rect 12069 15651 12127 15657
rect 12158 15648 12164 15700
rect 12216 15688 12222 15700
rect 13173 15691 13231 15697
rect 13173 15688 13185 15691
rect 12216 15660 13185 15688
rect 12216 15648 12222 15660
rect 13173 15657 13185 15660
rect 13219 15657 13231 15691
rect 13538 15688 13544 15700
rect 13499 15660 13544 15688
rect 13173 15651 13231 15657
rect 13538 15648 13544 15660
rect 13596 15648 13602 15700
rect 15657 15691 15715 15697
rect 15657 15657 15669 15691
rect 15703 15688 15715 15691
rect 16114 15688 16120 15700
rect 15703 15660 16120 15688
rect 15703 15657 15715 15660
rect 15657 15651 15715 15657
rect 16114 15648 16120 15660
rect 16172 15648 16178 15700
rect 5166 15629 5172 15632
rect 5160 15620 5172 15629
rect 5127 15592 5172 15620
rect 5160 15583 5172 15592
rect 5166 15580 5172 15583
rect 5224 15580 5230 15632
rect 5534 15580 5540 15632
rect 5592 15620 5598 15632
rect 6546 15620 6552 15632
rect 5592 15592 6552 15620
rect 5592 15580 5598 15592
rect 6546 15580 6552 15592
rect 6604 15620 6610 15632
rect 6604 15592 10088 15620
rect 6604 15580 6610 15592
rect 2225 15555 2283 15561
rect 2225 15521 2237 15555
rect 2271 15552 2283 15555
rect 3050 15552 3056 15564
rect 2271 15524 3056 15552
rect 2271 15521 2283 15524
rect 2225 15515 2283 15521
rect 3050 15512 3056 15524
rect 3108 15512 3114 15564
rect 4893 15555 4951 15561
rect 4893 15521 4905 15555
rect 4939 15552 4951 15555
rect 7368 15555 7426 15561
rect 4939 15524 6868 15552
rect 4939 15521 4951 15524
rect 4893 15515 4951 15521
rect 6840 15496 6868 15524
rect 7368 15521 7380 15555
rect 7414 15552 7426 15555
rect 8294 15552 8300 15564
rect 7414 15524 8300 15552
rect 7414 15521 7426 15524
rect 7368 15515 7426 15521
rect 8294 15512 8300 15524
rect 8352 15552 8358 15564
rect 9214 15552 9220 15564
rect 8352 15524 9220 15552
rect 8352 15512 8358 15524
rect 9214 15512 9220 15524
rect 9272 15512 9278 15564
rect 10060 15561 10088 15592
rect 10045 15555 10103 15561
rect 10045 15521 10057 15555
rect 10091 15552 10103 15555
rect 11238 15552 11244 15564
rect 10091 15524 11244 15552
rect 10091 15521 10103 15524
rect 10045 15515 10103 15521
rect 11238 15512 11244 15524
rect 11296 15512 11302 15564
rect 11517 15555 11575 15561
rect 11517 15521 11529 15555
rect 11563 15552 11575 15555
rect 11790 15552 11796 15564
rect 11563 15524 11796 15552
rect 11563 15521 11575 15524
rect 11517 15515 11575 15521
rect 11790 15512 11796 15524
rect 11848 15512 11854 15564
rect 11882 15512 11888 15564
rect 11940 15552 11946 15564
rect 11977 15555 12035 15561
rect 11977 15552 11989 15555
rect 11940 15524 11989 15552
rect 11940 15512 11946 15524
rect 11977 15521 11989 15524
rect 12023 15521 12035 15555
rect 15470 15552 15476 15564
rect 15431 15524 15476 15552
rect 11977 15515 12035 15521
rect 15470 15512 15476 15524
rect 15528 15512 15534 15564
rect 2501 15487 2559 15493
rect 2501 15453 2513 15487
rect 2547 15484 2559 15487
rect 4246 15484 4252 15496
rect 2547 15456 4252 15484
rect 2547 15453 2559 15456
rect 2501 15447 2559 15453
rect 4246 15444 4252 15456
rect 4304 15444 4310 15496
rect 6822 15444 6828 15496
rect 6880 15484 6886 15496
rect 7098 15484 7104 15496
rect 6880 15456 7104 15484
rect 6880 15444 6886 15456
rect 7098 15444 7104 15456
rect 7156 15444 7162 15496
rect 10229 15487 10287 15493
rect 10229 15453 10241 15487
rect 10275 15453 10287 15487
rect 10229 15447 10287 15453
rect 9582 15376 9588 15428
rect 9640 15416 9646 15428
rect 10244 15416 10272 15447
rect 12066 15444 12072 15496
rect 12124 15484 12130 15496
rect 12161 15487 12219 15493
rect 12161 15484 12173 15487
rect 12124 15456 12173 15484
rect 12124 15444 12130 15456
rect 12161 15453 12173 15456
rect 12207 15453 12219 15487
rect 12161 15447 12219 15453
rect 12250 15444 12256 15496
rect 12308 15484 12314 15496
rect 13633 15487 13691 15493
rect 13633 15484 13645 15487
rect 12308 15456 13645 15484
rect 12308 15444 12314 15456
rect 13633 15453 13645 15456
rect 13679 15453 13691 15487
rect 13633 15447 13691 15453
rect 13817 15487 13875 15493
rect 13817 15453 13829 15487
rect 13863 15484 13875 15487
rect 13998 15484 14004 15496
rect 13863 15456 14004 15484
rect 13863 15453 13875 15456
rect 13817 15447 13875 15453
rect 13998 15444 14004 15456
rect 14056 15484 14062 15496
rect 14918 15484 14924 15496
rect 14056 15456 14924 15484
rect 14056 15444 14062 15456
rect 14918 15444 14924 15456
rect 14976 15444 14982 15496
rect 9640 15388 10272 15416
rect 9640 15376 9646 15388
rect 11238 15376 11244 15428
rect 11296 15416 11302 15428
rect 11609 15419 11667 15425
rect 11609 15416 11621 15419
rect 11296 15388 11621 15416
rect 11296 15376 11302 15388
rect 11609 15385 11621 15388
rect 11655 15385 11667 15419
rect 11609 15379 11667 15385
rect 6273 15351 6331 15357
rect 6273 15317 6285 15351
rect 6319 15348 6331 15351
rect 6454 15348 6460 15360
rect 6319 15320 6460 15348
rect 6319 15317 6331 15320
rect 6273 15311 6331 15317
rect 6454 15308 6460 15320
rect 6512 15308 6518 15360
rect 7742 15308 7748 15360
rect 7800 15348 7806 15360
rect 12802 15348 12808 15360
rect 7800 15320 12808 15348
rect 7800 15308 7806 15320
rect 12802 15308 12808 15320
rect 12860 15348 12866 15360
rect 14090 15348 14096 15360
rect 12860 15320 14096 15348
rect 12860 15308 12866 15320
rect 14090 15308 14096 15320
rect 14148 15308 14154 15360
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 3050 15144 3056 15156
rect 3011 15116 3056 15144
rect 3050 15104 3056 15116
rect 3108 15104 3114 15156
rect 4062 15104 4068 15156
rect 4120 15144 4126 15156
rect 8202 15144 8208 15156
rect 4120 15116 8208 15144
rect 4120 15104 4126 15116
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 9214 15144 9220 15156
rect 9175 15116 9220 15144
rect 9214 15104 9220 15116
rect 9272 15104 9278 15156
rect 10781 15147 10839 15153
rect 10781 15113 10793 15147
rect 10827 15144 10839 15147
rect 12250 15144 12256 15156
rect 10827 15116 12256 15144
rect 10827 15113 10839 15116
rect 10781 15107 10839 15113
rect 12250 15104 12256 15116
rect 12308 15104 12314 15156
rect 13817 15147 13875 15153
rect 13817 15144 13829 15147
rect 12452 15116 13829 15144
rect 6454 15076 6460 15088
rect 3712 15048 6460 15076
rect 3712 15017 3740 15048
rect 6454 15036 6460 15048
rect 6512 15036 6518 15088
rect 11698 15076 11704 15088
rect 11440 15048 11704 15076
rect 3697 15011 3755 15017
rect 3697 14977 3709 15011
rect 3743 14977 3755 15011
rect 5166 15008 5172 15020
rect 5127 14980 5172 15008
rect 3697 14971 3755 14977
rect 5166 14968 5172 14980
rect 5224 14968 5230 15020
rect 7098 14968 7104 15020
rect 7156 15008 7162 15020
rect 7837 15011 7895 15017
rect 7837 15008 7849 15011
rect 7156 14980 7849 15008
rect 7156 14968 7162 14980
rect 7837 14977 7849 14980
rect 7883 14977 7895 15011
rect 11238 15008 11244 15020
rect 11199 14980 11244 15008
rect 7837 14971 7895 14977
rect 11238 14968 11244 14980
rect 11296 14968 11302 15020
rect 11440 15017 11468 15048
rect 11698 15036 11704 15048
rect 11756 15076 11762 15088
rect 12452 15076 12480 15116
rect 13817 15113 13829 15116
rect 13863 15144 13875 15147
rect 14826 15144 14832 15156
rect 13863 15116 14832 15144
rect 13863 15113 13875 15116
rect 13817 15107 13875 15113
rect 14826 15104 14832 15116
rect 14884 15104 14890 15156
rect 14918 15104 14924 15156
rect 14976 15144 14982 15156
rect 16025 15147 16083 15153
rect 16025 15144 16037 15147
rect 14976 15116 16037 15144
rect 14976 15104 14982 15116
rect 16025 15113 16037 15116
rect 16071 15113 16083 15147
rect 16025 15107 16083 15113
rect 11756 15048 12480 15076
rect 11756 15036 11762 15048
rect 11425 15011 11483 15017
rect 11425 14977 11437 15011
rect 11471 14977 11483 15011
rect 11425 14971 11483 14977
rect 1765 14943 1823 14949
rect 1765 14909 1777 14943
rect 1811 14940 1823 14943
rect 4982 14940 4988 14952
rect 1811 14912 4988 14940
rect 1811 14909 1823 14912
rect 1765 14903 1823 14909
rect 4982 14900 4988 14912
rect 5040 14900 5046 14952
rect 5077 14943 5135 14949
rect 5077 14909 5089 14943
rect 5123 14940 5135 14943
rect 5350 14940 5356 14952
rect 5123 14912 5356 14940
rect 5123 14909 5135 14912
rect 5077 14903 5135 14909
rect 5350 14900 5356 14912
rect 5408 14900 5414 14952
rect 6362 14940 6368 14952
rect 6323 14912 6368 14940
rect 6362 14900 6368 14912
rect 6420 14900 6426 14952
rect 6454 14900 6460 14952
rect 6512 14940 6518 14952
rect 7282 14940 7288 14952
rect 6512 14912 7288 14940
rect 6512 14900 6518 14912
rect 7282 14900 7288 14912
rect 7340 14900 7346 14952
rect 8104 14943 8162 14949
rect 8104 14909 8116 14943
rect 8150 14940 8162 14943
rect 9582 14940 9588 14952
rect 8150 14912 9588 14940
rect 8150 14909 8162 14912
rect 8104 14903 8162 14909
rect 9582 14900 9588 14912
rect 9640 14900 9646 14952
rect 10778 14900 10784 14952
rect 10836 14940 10842 14952
rect 11149 14943 11207 14949
rect 11149 14940 11161 14943
rect 10836 14912 11161 14940
rect 10836 14900 10842 14912
rect 11149 14909 11161 14912
rect 11195 14909 11207 14943
rect 11149 14903 11207 14909
rect 12434 14900 12440 14952
rect 12492 14940 12498 14952
rect 13722 14940 13728 14952
rect 12492 14912 13728 14940
rect 12492 14900 12498 14912
rect 13722 14900 13728 14912
rect 13780 14940 13786 14952
rect 14645 14943 14703 14949
rect 14645 14940 14657 14943
rect 13780 14912 14657 14940
rect 13780 14900 13786 14912
rect 14645 14909 14657 14912
rect 14691 14909 14703 14943
rect 16853 14943 16911 14949
rect 16853 14940 16865 14943
rect 14645 14903 14703 14909
rect 14752 14912 16865 14940
rect 3421 14875 3479 14881
rect 3421 14841 3433 14875
rect 3467 14872 3479 14875
rect 3467 14844 11284 14872
rect 3467 14841 3479 14844
rect 3421 14835 3479 14841
rect 1946 14804 1952 14816
rect 1907 14776 1952 14804
rect 1946 14764 1952 14776
rect 2004 14764 2010 14816
rect 3513 14807 3571 14813
rect 3513 14773 3525 14807
rect 3559 14804 3571 14807
rect 4617 14807 4675 14813
rect 4617 14804 4629 14807
rect 3559 14776 4629 14804
rect 3559 14773 3571 14776
rect 3513 14767 3571 14773
rect 4617 14773 4629 14776
rect 4663 14773 4675 14807
rect 4617 14767 4675 14773
rect 4985 14807 5043 14813
rect 4985 14773 4997 14807
rect 5031 14804 5043 14807
rect 5534 14804 5540 14816
rect 5031 14776 5540 14804
rect 5031 14773 5043 14776
rect 4985 14767 5043 14773
rect 5534 14764 5540 14776
rect 5592 14764 5598 14816
rect 6178 14804 6184 14816
rect 6139 14776 6184 14804
rect 6178 14764 6184 14776
rect 6236 14764 6242 14816
rect 6825 14807 6883 14813
rect 6825 14773 6837 14807
rect 6871 14804 6883 14807
rect 8938 14804 8944 14816
rect 6871 14776 8944 14804
rect 6871 14773 6883 14776
rect 6825 14767 6883 14773
rect 8938 14764 8944 14776
rect 8996 14764 9002 14816
rect 11256 14804 11284 14844
rect 12066 14832 12072 14884
rect 12124 14872 12130 14884
rect 12682 14875 12740 14881
rect 12682 14872 12694 14875
rect 12124 14844 12694 14872
rect 12124 14832 12130 14844
rect 12682 14841 12694 14844
rect 12728 14841 12740 14875
rect 14752 14872 14780 14912
rect 16853 14909 16865 14912
rect 16899 14909 16911 14943
rect 16853 14903 16911 14909
rect 12682 14835 12740 14841
rect 13740 14844 14780 14872
rect 13740 14804 13768 14844
rect 14826 14832 14832 14884
rect 14884 14881 14890 14884
rect 14884 14875 14948 14881
rect 14884 14841 14902 14875
rect 14936 14841 14948 14875
rect 14884 14835 14948 14841
rect 14884 14832 14890 14835
rect 11256 14776 13768 14804
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 3510 14560 3516 14612
rect 3568 14600 3574 14612
rect 4249 14603 4307 14609
rect 4249 14600 4261 14603
rect 3568 14572 4261 14600
rect 3568 14560 3574 14572
rect 4249 14569 4261 14572
rect 4295 14569 4307 14603
rect 4249 14563 4307 14569
rect 4982 14560 4988 14612
rect 5040 14600 5046 14612
rect 9677 14603 9735 14609
rect 5040 14572 8616 14600
rect 5040 14560 5046 14572
rect 8588 14541 8616 14572
rect 9677 14569 9689 14603
rect 9723 14600 9735 14603
rect 11054 14600 11060 14612
rect 9723 14572 11060 14600
rect 9723 14569 9735 14572
rect 9677 14563 9735 14569
rect 11054 14560 11060 14572
rect 11112 14560 11118 14612
rect 12066 14600 12072 14612
rect 12027 14572 12072 14600
rect 12066 14560 12072 14572
rect 12124 14560 12130 14612
rect 16758 14600 16764 14612
rect 16719 14572 16764 14600
rect 16758 14560 16764 14572
rect 16816 14560 16822 14612
rect 8573 14535 8631 14541
rect 5184 14504 8524 14532
rect 2777 14467 2835 14473
rect 2777 14433 2789 14467
rect 2823 14464 2835 14467
rect 2958 14464 2964 14476
rect 2823 14436 2964 14464
rect 2823 14433 2835 14436
rect 2777 14427 2835 14433
rect 2958 14424 2964 14436
rect 3016 14424 3022 14476
rect 4062 14464 4068 14476
rect 4023 14436 4068 14464
rect 4062 14424 4068 14436
rect 4120 14424 4126 14476
rect 5184 14473 5212 14504
rect 5169 14467 5227 14473
rect 5169 14433 5181 14467
rect 5215 14433 5227 14467
rect 6730 14464 6736 14476
rect 5169 14427 5227 14433
rect 5276 14436 6736 14464
rect 1397 14399 1455 14405
rect 1397 14365 1409 14399
rect 1443 14365 1455 14399
rect 2866 14396 2872 14408
rect 2827 14368 2872 14396
rect 1397 14359 1455 14365
rect 1412 14328 1440 14359
rect 2866 14356 2872 14368
rect 2924 14356 2930 14408
rect 3053 14399 3111 14405
rect 3053 14365 3065 14399
rect 3099 14396 3111 14399
rect 3234 14396 3240 14408
rect 3099 14368 3240 14396
rect 3099 14365 3111 14368
rect 3053 14359 3111 14365
rect 3234 14356 3240 14368
rect 3292 14356 3298 14408
rect 5276 14396 5304 14436
rect 6730 14424 6736 14436
rect 6788 14424 6794 14476
rect 6825 14467 6883 14473
rect 6825 14433 6837 14467
rect 6871 14464 6883 14467
rect 7650 14464 7656 14476
rect 6871 14436 7656 14464
rect 6871 14433 6883 14436
rect 6825 14427 6883 14433
rect 7650 14424 7656 14436
rect 7708 14424 7714 14476
rect 8294 14464 8300 14476
rect 8255 14436 8300 14464
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 8496 14464 8524 14504
rect 8573 14501 8585 14535
rect 8619 14501 8631 14535
rect 13725 14535 13783 14541
rect 8573 14495 8631 14501
rect 10520 14504 11744 14532
rect 10520 14464 10548 14504
rect 8496 14436 10548 14464
rect 10594 14424 10600 14476
rect 10652 14464 10658 14476
rect 10945 14467 11003 14473
rect 10945 14464 10957 14467
rect 10652 14436 10957 14464
rect 10652 14424 10658 14436
rect 10945 14433 10957 14436
rect 10991 14433 11003 14467
rect 10945 14427 11003 14433
rect 3804 14368 5304 14396
rect 3804 14328 3832 14368
rect 6638 14356 6644 14408
rect 6696 14396 6702 14408
rect 6917 14399 6975 14405
rect 6917 14396 6929 14399
rect 6696 14368 6929 14396
rect 6696 14356 6702 14368
rect 6917 14365 6929 14368
rect 6963 14365 6975 14399
rect 6917 14359 6975 14365
rect 7009 14399 7067 14405
rect 7009 14365 7021 14399
rect 7055 14365 7067 14399
rect 7009 14359 7067 14365
rect 1412 14300 3832 14328
rect 3878 14288 3884 14340
rect 3936 14328 3942 14340
rect 5353 14331 5411 14337
rect 5353 14328 5365 14331
rect 3936 14300 5365 14328
rect 3936 14288 3942 14300
rect 5353 14297 5365 14300
rect 5399 14297 5411 14331
rect 5353 14291 5411 14297
rect 6730 14288 6736 14340
rect 6788 14328 6794 14340
rect 7024 14328 7052 14359
rect 8478 14356 8484 14408
rect 8536 14396 8542 14408
rect 9214 14396 9220 14408
rect 8536 14368 9220 14396
rect 8536 14356 8542 14368
rect 9214 14356 9220 14368
rect 9272 14396 9278 14408
rect 10689 14399 10747 14405
rect 10689 14396 10701 14399
rect 9272 14368 10701 14396
rect 9272 14356 9278 14368
rect 10689 14365 10701 14368
rect 10735 14365 10747 14399
rect 11716 14396 11744 14504
rect 13725 14501 13737 14535
rect 13771 14532 13783 14535
rect 14734 14532 14740 14544
rect 13771 14504 14740 14532
rect 13771 14501 13783 14504
rect 13725 14495 13783 14501
rect 14734 14492 14740 14504
rect 14792 14492 14798 14544
rect 15565 14535 15623 14541
rect 15565 14501 15577 14535
rect 15611 14532 15623 14535
rect 16390 14532 16396 14544
rect 15611 14504 16396 14532
rect 15611 14501 15623 14504
rect 15565 14495 15623 14501
rect 16390 14492 16396 14504
rect 16448 14492 16454 14544
rect 13446 14464 13452 14476
rect 13407 14436 13452 14464
rect 13446 14424 13452 14436
rect 13504 14424 13510 14476
rect 15286 14464 15292 14476
rect 15247 14436 15292 14464
rect 15286 14424 15292 14436
rect 15344 14424 15350 14476
rect 16298 14424 16304 14476
rect 16356 14464 16362 14476
rect 16577 14467 16635 14473
rect 16577 14464 16589 14467
rect 16356 14436 16589 14464
rect 16356 14424 16362 14436
rect 16577 14433 16589 14436
rect 16623 14433 16635 14467
rect 16577 14427 16635 14433
rect 13906 14396 13912 14408
rect 11716 14368 13912 14396
rect 10689 14359 10747 14365
rect 13906 14356 13912 14368
rect 13964 14356 13970 14408
rect 6788 14300 7052 14328
rect 6788 14288 6794 14300
rect 2409 14263 2467 14269
rect 2409 14229 2421 14263
rect 2455 14260 2467 14263
rect 4154 14260 4160 14272
rect 2455 14232 4160 14260
rect 2455 14229 2467 14232
rect 2409 14223 2467 14229
rect 4154 14220 4160 14232
rect 4212 14220 4218 14272
rect 6457 14263 6515 14269
rect 6457 14229 6469 14263
rect 6503 14260 6515 14263
rect 7190 14260 7196 14272
rect 6503 14232 7196 14260
rect 6503 14229 6515 14232
rect 6457 14223 6515 14229
rect 7190 14220 7196 14232
rect 7248 14220 7254 14272
rect 7282 14220 7288 14272
rect 7340 14260 7346 14272
rect 16758 14260 16764 14272
rect 7340 14232 16764 14260
rect 7340 14220 7346 14232
rect 16758 14220 16764 14232
rect 16816 14220 16822 14272
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 3786 14016 3792 14068
rect 3844 14056 3850 14068
rect 4065 14059 4123 14065
rect 4065 14056 4077 14059
rect 3844 14028 4077 14056
rect 3844 14016 3850 14028
rect 4065 14025 4077 14028
rect 4111 14025 4123 14059
rect 4065 14019 4123 14025
rect 4154 14016 4160 14068
rect 4212 14056 4218 14068
rect 15286 14056 15292 14068
rect 4212 14028 15292 14056
rect 4212 14016 4218 14028
rect 15286 14016 15292 14028
rect 15344 14016 15350 14068
rect 6825 13991 6883 13997
rect 6825 13957 6837 13991
rect 6871 13988 6883 13991
rect 7098 13988 7104 14000
rect 6871 13960 7104 13988
rect 6871 13957 6883 13960
rect 6825 13951 6883 13957
rect 7098 13948 7104 13960
rect 7156 13948 7162 14000
rect 10594 13988 10600 14000
rect 10555 13960 10600 13988
rect 10594 13948 10600 13960
rect 10652 13948 10658 14000
rect 11054 13948 11060 14000
rect 11112 13988 11118 14000
rect 12437 13991 12495 13997
rect 12437 13988 12449 13991
rect 11112 13960 12449 13988
rect 11112 13948 11118 13960
rect 12437 13957 12449 13960
rect 12483 13957 12495 13991
rect 12437 13951 12495 13957
rect 4264 13892 4476 13920
rect 1670 13812 1676 13864
rect 1728 13852 1734 13864
rect 1857 13855 1915 13861
rect 1857 13852 1869 13855
rect 1728 13824 1869 13852
rect 1728 13812 1734 13824
rect 1857 13821 1869 13824
rect 1903 13852 1915 13855
rect 3786 13852 3792 13864
rect 1903 13824 3792 13852
rect 1903 13821 1915 13824
rect 1857 13815 1915 13821
rect 3786 13812 3792 13824
rect 3844 13812 3850 13864
rect 4264 13861 4292 13892
rect 4249 13855 4307 13861
rect 4249 13821 4261 13855
rect 4295 13821 4307 13855
rect 4249 13815 4307 13821
rect 4341 13855 4399 13861
rect 4341 13821 4353 13855
rect 4387 13821 4399 13855
rect 4448 13852 4476 13892
rect 5718 13880 5724 13932
rect 5776 13920 5782 13932
rect 6730 13920 6736 13932
rect 5776 13892 6736 13920
rect 5776 13880 5782 13892
rect 6730 13880 6736 13892
rect 6788 13920 6794 13932
rect 7377 13923 7435 13929
rect 7377 13920 7389 13923
rect 6788 13892 7389 13920
rect 6788 13880 6794 13892
rect 7377 13889 7389 13892
rect 7423 13889 7435 13923
rect 9214 13920 9220 13932
rect 9175 13892 9220 13920
rect 7377 13883 7435 13889
rect 9214 13880 9220 13892
rect 9272 13880 9278 13932
rect 12066 13880 12072 13932
rect 12124 13920 12130 13932
rect 12989 13923 13047 13929
rect 12989 13920 13001 13923
rect 12124 13892 13001 13920
rect 12124 13880 12130 13892
rect 12989 13889 13001 13892
rect 13035 13889 13047 13923
rect 12989 13883 13047 13889
rect 15013 13923 15071 13929
rect 15013 13889 15025 13923
rect 15059 13920 15071 13923
rect 15470 13920 15476 13932
rect 15059 13892 15476 13920
rect 15059 13889 15071 13892
rect 15013 13883 15071 13889
rect 15470 13880 15476 13892
rect 15528 13880 15534 13932
rect 16298 13920 16304 13932
rect 16259 13892 16304 13920
rect 16298 13880 16304 13892
rect 16356 13880 16362 13932
rect 6178 13852 6184 13864
rect 4448 13824 6184 13852
rect 4341 13815 4399 13821
rect 2124 13787 2182 13793
rect 2124 13753 2136 13787
rect 2170 13784 2182 13787
rect 3050 13784 3056 13796
rect 2170 13756 3056 13784
rect 2170 13753 2182 13756
rect 2124 13747 2182 13753
rect 3050 13744 3056 13756
rect 3108 13744 3114 13796
rect 3804 13784 3832 13812
rect 4356 13784 4384 13815
rect 6178 13812 6184 13824
rect 6236 13812 6242 13864
rect 9484 13855 9542 13861
rect 9484 13821 9496 13855
rect 9530 13852 9542 13855
rect 10686 13852 10692 13864
rect 9530 13824 10692 13852
rect 9530 13821 9542 13824
rect 9484 13815 9542 13821
rect 10686 13812 10692 13824
rect 10744 13812 10750 13864
rect 12710 13812 12716 13864
rect 12768 13852 12774 13864
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 12768 13824 12909 13852
rect 12768 13812 12774 13824
rect 12897 13821 12909 13824
rect 12943 13821 12955 13855
rect 14734 13852 14740 13864
rect 14695 13824 14740 13852
rect 12897 13815 12955 13821
rect 14734 13812 14740 13824
rect 14792 13812 14798 13864
rect 16022 13852 16028 13864
rect 15983 13824 16028 13852
rect 16022 13812 16028 13824
rect 16080 13812 16086 13864
rect 3804 13756 4384 13784
rect 4608 13787 4666 13793
rect 4608 13753 4620 13787
rect 4654 13784 4666 13787
rect 4798 13784 4804 13796
rect 4654 13756 4804 13784
rect 4654 13753 4666 13756
rect 4608 13747 4666 13753
rect 4798 13744 4804 13756
rect 4856 13744 4862 13796
rect 12802 13784 12808 13796
rect 12763 13756 12808 13784
rect 12802 13744 12808 13756
rect 12860 13744 12866 13796
rect 3234 13716 3240 13728
rect 3195 13688 3240 13716
rect 3234 13676 3240 13688
rect 3292 13676 3298 13728
rect 5718 13716 5724 13728
rect 5679 13688 5724 13716
rect 5718 13676 5724 13688
rect 5776 13676 5782 13728
rect 7006 13676 7012 13728
rect 7064 13716 7070 13728
rect 7193 13719 7251 13725
rect 7193 13716 7205 13719
rect 7064 13688 7205 13716
rect 7064 13676 7070 13688
rect 7193 13685 7205 13688
rect 7239 13685 7251 13719
rect 7193 13679 7251 13685
rect 7282 13676 7288 13728
rect 7340 13716 7346 13728
rect 7340 13688 7385 13716
rect 7340 13676 7346 13688
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 2409 13515 2467 13521
rect 2409 13481 2421 13515
rect 2455 13512 2467 13515
rect 2866 13512 2872 13524
rect 2455 13484 2872 13512
rect 2455 13481 2467 13484
rect 2409 13475 2467 13481
rect 2866 13472 2872 13484
rect 2924 13472 2930 13524
rect 5258 13472 5264 13524
rect 5316 13512 5322 13524
rect 7009 13515 7067 13521
rect 5316 13484 6960 13512
rect 5316 13472 5322 13484
rect 1118 13404 1124 13456
rect 1176 13444 1182 13456
rect 5068 13447 5126 13453
rect 1176 13416 5028 13444
rect 1176 13404 1182 13416
rect 2774 13336 2780 13388
rect 2832 13376 2838 13388
rect 2832 13348 2877 13376
rect 2832 13336 2838 13348
rect 3786 13336 3792 13388
rect 3844 13376 3850 13388
rect 4801 13379 4859 13385
rect 4801 13376 4813 13379
rect 3844 13348 4813 13376
rect 3844 13336 3850 13348
rect 4801 13345 4813 13348
rect 4847 13345 4859 13379
rect 5000 13376 5028 13416
rect 5068 13413 5080 13447
rect 5114 13444 5126 13447
rect 5718 13444 5724 13456
rect 5114 13416 5724 13444
rect 5114 13413 5126 13416
rect 5068 13407 5126 13413
rect 5718 13404 5724 13416
rect 5776 13404 5782 13456
rect 6932 13444 6960 13484
rect 7009 13481 7021 13515
rect 7055 13512 7067 13515
rect 7282 13512 7288 13524
rect 7055 13484 7288 13512
rect 7055 13481 7067 13484
rect 7009 13475 7067 13481
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 7374 13472 7380 13524
rect 7432 13512 7438 13524
rect 7469 13515 7527 13521
rect 7469 13512 7481 13515
rect 7432 13484 7481 13512
rect 7432 13472 7438 13484
rect 7469 13481 7481 13484
rect 7515 13481 7527 13515
rect 7469 13475 7527 13481
rect 7650 13472 7656 13524
rect 7708 13512 7714 13524
rect 8573 13515 8631 13521
rect 8573 13512 8585 13515
rect 7708 13484 8585 13512
rect 7708 13472 7714 13484
rect 8573 13481 8585 13484
rect 8619 13481 8631 13515
rect 8573 13475 8631 13481
rect 10962 13472 10968 13524
rect 11020 13512 11026 13524
rect 13446 13512 13452 13524
rect 11020 13484 13452 13512
rect 11020 13472 11026 13484
rect 13446 13472 13452 13484
rect 13504 13472 13510 13524
rect 10134 13444 10140 13456
rect 6932 13416 10140 13444
rect 10134 13404 10140 13416
rect 10192 13404 10198 13456
rect 12434 13444 12440 13456
rect 11808 13416 12440 13444
rect 7377 13379 7435 13385
rect 7377 13376 7389 13379
rect 5000 13348 7389 13376
rect 4801 13339 4859 13345
rect 7377 13345 7389 13348
rect 7423 13376 7435 13379
rect 7742 13376 7748 13388
rect 7423 13348 7748 13376
rect 7423 13345 7435 13348
rect 7377 13339 7435 13345
rect 7742 13336 7748 13348
rect 7800 13336 7806 13388
rect 9122 13336 9128 13388
rect 9180 13376 9186 13388
rect 10045 13379 10103 13385
rect 10045 13376 10057 13379
rect 9180 13348 10057 13376
rect 9180 13336 9186 13348
rect 10045 13345 10057 13348
rect 10091 13345 10103 13379
rect 10045 13339 10103 13345
rect 10870 13336 10876 13388
rect 10928 13376 10934 13388
rect 11808 13385 11836 13416
rect 12434 13404 12440 13416
rect 12492 13404 12498 13456
rect 15562 13444 15568 13456
rect 15523 13416 15568 13444
rect 15562 13404 15568 13416
rect 15620 13404 15626 13456
rect 12066 13385 12072 13388
rect 11425 13379 11483 13385
rect 11425 13376 11437 13379
rect 10928 13348 11437 13376
rect 10928 13336 10934 13348
rect 11425 13345 11437 13348
rect 11471 13345 11483 13379
rect 11425 13339 11483 13345
rect 11793 13379 11851 13385
rect 11793 13345 11805 13379
rect 11839 13345 11851 13379
rect 12060 13376 12072 13385
rect 12027 13348 12072 13376
rect 11793 13339 11851 13345
rect 12060 13339 12072 13348
rect 12066 13336 12072 13339
rect 12124 13336 12130 13388
rect 15289 13379 15347 13385
rect 15289 13345 15301 13379
rect 15335 13376 15347 13379
rect 15746 13376 15752 13388
rect 15335 13348 15752 13376
rect 15335 13345 15347 13348
rect 15289 13339 15347 13345
rect 15746 13336 15752 13348
rect 15804 13336 15810 13388
rect 1397 13311 1455 13317
rect 1397 13277 1409 13311
rect 1443 13308 1455 13311
rect 1946 13308 1952 13320
rect 1443 13280 1952 13308
rect 1443 13277 1455 13280
rect 1397 13271 1455 13277
rect 1946 13268 1952 13280
rect 2004 13268 2010 13320
rect 2866 13308 2872 13320
rect 2827 13280 2872 13308
rect 2866 13268 2872 13280
rect 2924 13268 2930 13320
rect 3050 13308 3056 13320
rect 3011 13280 3056 13308
rect 3050 13268 3056 13280
rect 3108 13268 3114 13320
rect 7558 13308 7564 13320
rect 6012 13280 7564 13308
rect 4798 13132 4804 13184
rect 4856 13172 4862 13184
rect 6012 13172 6040 13280
rect 7558 13268 7564 13280
rect 7616 13268 7622 13320
rect 10321 13311 10379 13317
rect 10321 13277 10333 13311
rect 10367 13308 10379 13311
rect 10686 13308 10692 13320
rect 10367 13280 10692 13308
rect 10367 13277 10379 13280
rect 10321 13271 10379 13277
rect 10686 13268 10692 13280
rect 10744 13268 10750 13320
rect 14182 13308 14188 13320
rect 14143 13280 14188 13308
rect 14182 13268 14188 13280
rect 14240 13268 14246 13320
rect 13446 13240 13452 13252
rect 12719 13212 13452 13240
rect 6178 13172 6184 13184
rect 4856 13144 6040 13172
rect 6139 13144 6184 13172
rect 4856 13132 4862 13144
rect 6178 13132 6184 13144
rect 6236 13132 6242 13184
rect 8846 13132 8852 13184
rect 8904 13172 8910 13184
rect 9677 13175 9735 13181
rect 9677 13172 9689 13175
rect 8904 13144 9689 13172
rect 8904 13132 8910 13144
rect 9677 13141 9689 13144
rect 9723 13141 9735 13175
rect 9677 13135 9735 13141
rect 11241 13175 11299 13181
rect 11241 13141 11253 13175
rect 11287 13172 11299 13175
rect 11790 13172 11796 13184
rect 11287 13144 11796 13172
rect 11287 13141 11299 13144
rect 11241 13135 11299 13141
rect 11790 13132 11796 13144
rect 11848 13172 11854 13184
rect 12719 13172 12747 13212
rect 13446 13200 13452 13212
rect 13504 13200 13510 13252
rect 13170 13172 13176 13184
rect 11848 13144 12747 13172
rect 13131 13144 13176 13172
rect 11848 13132 11854 13144
rect 13170 13132 13176 13144
rect 13228 13132 13234 13184
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12968 1639 12971
rect 2958 12968 2964 12980
rect 1627 12940 2964 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 2958 12928 2964 12940
rect 3016 12928 3022 12980
rect 4525 12971 4583 12977
rect 4525 12937 4537 12971
rect 4571 12968 4583 12971
rect 4798 12968 4804 12980
rect 4571 12940 4804 12968
rect 4571 12937 4583 12940
rect 4525 12931 4583 12937
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 5537 12971 5595 12977
rect 5537 12937 5549 12971
rect 5583 12968 5595 12971
rect 6086 12968 6092 12980
rect 5583 12940 6092 12968
rect 5583 12937 5595 12940
rect 5537 12931 5595 12937
rect 6086 12928 6092 12940
rect 6144 12928 6150 12980
rect 6362 12928 6368 12980
rect 6420 12968 6426 12980
rect 6457 12971 6515 12977
rect 6457 12968 6469 12971
rect 6420 12940 6469 12968
rect 6420 12928 6426 12940
rect 6457 12937 6469 12940
rect 6503 12937 6515 12971
rect 7006 12968 7012 12980
rect 6967 12940 7012 12968
rect 6457 12931 6515 12937
rect 7006 12928 7012 12940
rect 7064 12928 7070 12980
rect 7282 12928 7288 12980
rect 7340 12968 7346 12980
rect 11238 12968 11244 12980
rect 7340 12940 11244 12968
rect 7340 12928 7346 12940
rect 11238 12928 11244 12940
rect 11296 12928 11302 12980
rect 15746 12968 15752 12980
rect 15707 12940 15752 12968
rect 15746 12928 15752 12940
rect 15804 12928 15810 12980
rect 6656 12872 8892 12900
rect 2225 12835 2283 12841
rect 2225 12801 2237 12835
rect 2271 12832 2283 12835
rect 3050 12832 3056 12844
rect 2271 12804 3056 12832
rect 2271 12801 2283 12804
rect 2225 12795 2283 12801
rect 3050 12792 3056 12804
rect 3108 12792 3114 12844
rect 1946 12764 1952 12776
rect 1907 12736 1952 12764
rect 1946 12724 1952 12736
rect 2004 12724 2010 12776
rect 2958 12724 2964 12776
rect 3016 12764 3022 12776
rect 3145 12767 3203 12773
rect 3145 12764 3157 12767
rect 3016 12736 3157 12764
rect 3016 12724 3022 12736
rect 3145 12733 3157 12736
rect 3191 12733 3203 12767
rect 3145 12727 3203 12733
rect 3234 12724 3240 12776
rect 3292 12764 3298 12776
rect 3401 12767 3459 12773
rect 3401 12764 3413 12767
rect 3292 12736 3413 12764
rect 3292 12724 3298 12736
rect 3401 12733 3413 12736
rect 3447 12733 3459 12767
rect 3401 12727 3459 12733
rect 4246 12724 4252 12776
rect 4304 12764 4310 12776
rect 6656 12773 6684 12872
rect 7558 12832 7564 12844
rect 7519 12804 7564 12832
rect 7558 12792 7564 12804
rect 7616 12792 7622 12844
rect 8864 12832 8892 12872
rect 8938 12860 8944 12912
rect 8996 12900 9002 12912
rect 10597 12903 10655 12909
rect 10597 12900 10609 12903
rect 8996 12872 10609 12900
rect 8996 12860 9002 12872
rect 10597 12869 10609 12872
rect 10643 12869 10655 12903
rect 10597 12863 10655 12869
rect 10686 12860 10692 12912
rect 10744 12900 10750 12912
rect 14921 12903 14979 12909
rect 10744 12872 11284 12900
rect 10744 12860 10750 12872
rect 10321 12835 10379 12841
rect 10321 12832 10333 12835
rect 8864 12804 10333 12832
rect 10321 12801 10333 12804
rect 10367 12832 10379 12835
rect 10870 12832 10876 12844
rect 10367 12804 10876 12832
rect 10367 12801 10379 12804
rect 10321 12795 10379 12801
rect 10870 12792 10876 12804
rect 10928 12792 10934 12844
rect 11054 12832 11060 12844
rect 11015 12804 11060 12832
rect 11054 12792 11060 12804
rect 11112 12792 11118 12844
rect 11256 12841 11284 12872
rect 14921 12869 14933 12903
rect 14967 12900 14979 12903
rect 14967 12872 16344 12900
rect 14967 12869 14979 12872
rect 14921 12863 14979 12869
rect 16316 12844 16344 12872
rect 11241 12835 11299 12841
rect 11241 12801 11253 12835
rect 11287 12832 11299 12835
rect 13170 12832 13176 12844
rect 11287 12804 13176 12832
rect 11287 12801 11299 12804
rect 11241 12795 11299 12801
rect 13170 12792 13176 12804
rect 13228 12792 13234 12844
rect 16298 12832 16304 12844
rect 16211 12804 16304 12832
rect 16298 12792 16304 12804
rect 16356 12792 16362 12844
rect 5353 12767 5411 12773
rect 5353 12764 5365 12767
rect 4304 12736 5365 12764
rect 4304 12724 4310 12736
rect 5353 12733 5365 12736
rect 5399 12733 5411 12767
rect 5353 12727 5411 12733
rect 6641 12767 6699 12773
rect 6641 12733 6653 12767
rect 6687 12733 6699 12767
rect 6641 12727 6699 12733
rect 6914 12724 6920 12776
rect 6972 12764 6978 12776
rect 7282 12764 7288 12776
rect 6972 12736 7288 12764
rect 6972 12724 6978 12736
rect 7282 12724 7288 12736
rect 7340 12764 7346 12776
rect 7377 12767 7435 12773
rect 7377 12764 7389 12767
rect 7340 12736 7389 12764
rect 7340 12724 7346 12736
rect 7377 12733 7389 12736
rect 7423 12733 7435 12767
rect 7377 12727 7435 12733
rect 9030 12724 9036 12776
rect 9088 12764 9094 12776
rect 10965 12767 11023 12773
rect 10965 12764 10977 12767
rect 9088 12736 10977 12764
rect 9088 12724 9094 12736
rect 10965 12733 10977 12736
rect 11011 12733 11023 12767
rect 10965 12727 11023 12733
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 13538 12764 13544 12776
rect 12492 12736 13544 12764
rect 12492 12724 12498 12736
rect 13538 12724 13544 12736
rect 13596 12724 13602 12776
rect 14182 12724 14188 12776
rect 14240 12764 14246 12776
rect 16117 12767 16175 12773
rect 16117 12764 16129 12767
rect 14240 12736 16129 12764
rect 14240 12724 14246 12736
rect 16117 12733 16129 12736
rect 16163 12733 16175 12767
rect 16117 12727 16175 12733
rect 658 12656 664 12708
rect 716 12696 722 12708
rect 2314 12696 2320 12708
rect 716 12668 2320 12696
rect 716 12656 722 12668
rect 2314 12656 2320 12668
rect 2372 12656 2378 12708
rect 6730 12656 6736 12708
rect 6788 12696 6794 12708
rect 8757 12699 8815 12705
rect 8757 12696 8769 12699
rect 6788 12668 8769 12696
rect 6788 12656 6794 12668
rect 8757 12665 8769 12668
rect 8803 12665 8815 12699
rect 12250 12696 12256 12708
rect 8757 12659 8815 12665
rect 8956 12668 12256 12696
rect 2038 12628 2044 12640
rect 1999 12600 2044 12628
rect 2038 12588 2044 12600
rect 2096 12588 2102 12640
rect 5626 12588 5632 12640
rect 5684 12628 5690 12640
rect 7469 12631 7527 12637
rect 7469 12628 7481 12631
rect 5684 12600 7481 12628
rect 5684 12588 5690 12600
rect 7469 12597 7481 12600
rect 7515 12628 7527 12631
rect 8956 12628 8984 12668
rect 12250 12656 12256 12668
rect 12308 12656 12314 12708
rect 13814 12705 13820 12708
rect 13808 12659 13820 12705
rect 13872 12696 13878 12708
rect 13872 12668 13908 12696
rect 13814 12656 13820 12659
rect 13872 12656 13878 12668
rect 7515 12600 8984 12628
rect 12437 12631 12495 12637
rect 7515 12597 7527 12600
rect 7469 12591 7527 12597
rect 12437 12597 12449 12631
rect 12483 12628 12495 12631
rect 14642 12628 14648 12640
rect 12483 12600 14648 12628
rect 12483 12597 12495 12600
rect 12437 12591 12495 12597
rect 14642 12588 14648 12600
rect 14700 12588 14706 12640
rect 16206 12628 16212 12640
rect 16167 12600 16212 12628
rect 16206 12588 16212 12600
rect 16264 12588 16270 12640
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 3050 12424 3056 12436
rect 3011 12396 3056 12424
rect 3050 12384 3056 12396
rect 3108 12384 3114 12436
rect 6638 12424 6644 12436
rect 6599 12396 6644 12424
rect 6638 12384 6644 12396
rect 6696 12384 6702 12436
rect 8294 12384 8300 12436
rect 8352 12424 8358 12436
rect 8573 12427 8631 12433
rect 8573 12424 8585 12427
rect 8352 12396 8585 12424
rect 8352 12384 8358 12396
rect 8573 12393 8585 12396
rect 8619 12393 8631 12427
rect 8573 12387 8631 12393
rect 8846 12384 8852 12436
rect 8904 12424 8910 12436
rect 8941 12427 8999 12433
rect 8941 12424 8953 12427
rect 8904 12396 8953 12424
rect 8904 12384 8910 12396
rect 8941 12393 8953 12396
rect 8987 12393 8999 12427
rect 11609 12427 11667 12433
rect 11609 12424 11621 12427
rect 8941 12387 8999 12393
rect 9140 12396 11621 12424
rect 2958 12356 2964 12368
rect 1688 12328 2964 12356
rect 1688 12300 1716 12328
rect 2958 12316 2964 12328
rect 3016 12316 3022 12368
rect 4062 12316 4068 12368
rect 4120 12356 4126 12368
rect 7009 12359 7067 12365
rect 7009 12356 7021 12359
rect 4120 12328 7021 12356
rect 4120 12316 4126 12328
rect 7009 12325 7021 12328
rect 7055 12325 7067 12359
rect 9140 12356 9168 12396
rect 11609 12393 11621 12396
rect 11655 12393 11667 12427
rect 16022 12424 16028 12436
rect 11609 12387 11667 12393
rect 11900 12396 16028 12424
rect 11900 12368 11928 12396
rect 16022 12384 16028 12396
rect 16080 12384 16086 12436
rect 10594 12356 10600 12368
rect 7009 12319 7067 12325
rect 8312 12328 9168 12356
rect 9232 12328 10600 12356
rect 1670 12288 1676 12300
rect 1631 12260 1676 12288
rect 1670 12248 1676 12260
rect 1728 12248 1734 12300
rect 1940 12291 1998 12297
rect 1940 12257 1952 12291
rect 1986 12288 1998 12291
rect 3602 12288 3608 12300
rect 1986 12260 3608 12288
rect 1986 12257 1998 12260
rect 1940 12251 1998 12257
rect 3602 12248 3608 12260
rect 3660 12248 3666 12300
rect 4338 12248 4344 12300
rect 4396 12288 4402 12300
rect 4433 12291 4491 12297
rect 4433 12288 4445 12291
rect 4396 12260 4445 12288
rect 4396 12248 4402 12260
rect 4433 12257 4445 12260
rect 4479 12288 4491 12291
rect 4890 12288 4896 12300
rect 4479 12260 4896 12288
rect 4479 12257 4491 12260
rect 4433 12251 4491 12257
rect 4890 12248 4896 12260
rect 4948 12248 4954 12300
rect 5629 12291 5687 12297
rect 5629 12257 5641 12291
rect 5675 12288 5687 12291
rect 7466 12288 7472 12300
rect 5675 12260 7472 12288
rect 5675 12257 5687 12260
rect 5629 12251 5687 12257
rect 7466 12248 7472 12260
rect 7524 12248 7530 12300
rect 8312 12297 8340 12328
rect 8297 12291 8355 12297
rect 8297 12257 8309 12291
rect 8343 12257 8355 12291
rect 8297 12251 8355 12257
rect 8938 12248 8944 12300
rect 8996 12288 9002 12300
rect 9033 12291 9091 12297
rect 9033 12288 9045 12291
rect 8996 12260 9045 12288
rect 8996 12248 9002 12260
rect 9033 12257 9045 12260
rect 9079 12257 9091 12291
rect 9033 12251 9091 12257
rect 4525 12223 4583 12229
rect 4525 12189 4537 12223
rect 4571 12189 4583 12223
rect 4525 12183 4583 12189
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12220 4767 12223
rect 5534 12220 5540 12232
rect 4755 12192 5540 12220
rect 4755 12189 4767 12192
rect 4709 12183 4767 12189
rect 2866 12112 2872 12164
rect 2924 12152 2930 12164
rect 4065 12155 4123 12161
rect 4065 12152 4077 12155
rect 2924 12124 4077 12152
rect 2924 12112 2930 12124
rect 4065 12121 4077 12124
rect 4111 12121 4123 12155
rect 4540 12152 4568 12183
rect 5534 12180 5540 12192
rect 5592 12220 5598 12232
rect 6546 12220 6552 12232
rect 5592 12192 6552 12220
rect 5592 12180 5598 12192
rect 6546 12180 6552 12192
rect 6604 12180 6610 12232
rect 7101 12223 7159 12229
rect 7101 12189 7113 12223
rect 7147 12189 7159 12223
rect 7101 12183 7159 12189
rect 7285 12223 7343 12229
rect 7285 12189 7297 12223
rect 7331 12220 7343 12223
rect 7558 12220 7564 12232
rect 7331 12192 7564 12220
rect 7331 12189 7343 12192
rect 7285 12183 7343 12189
rect 4798 12152 4804 12164
rect 4540 12124 4804 12152
rect 4065 12115 4123 12121
rect 4798 12112 4804 12124
rect 4856 12112 4862 12164
rect 7116 12152 7144 12183
rect 7558 12180 7564 12192
rect 7616 12180 7622 12232
rect 9232 12229 9260 12328
rect 10594 12316 10600 12328
rect 10652 12316 10658 12368
rect 11698 12356 11704 12368
rect 11659 12328 11704 12356
rect 11698 12316 11704 12328
rect 11756 12316 11762 12368
rect 11882 12316 11888 12368
rect 11940 12316 11946 12368
rect 15556 12359 15614 12365
rect 15556 12325 15568 12359
rect 15602 12356 15614 12359
rect 16298 12356 16304 12368
rect 15602 12328 16304 12356
rect 15602 12325 15614 12328
rect 15556 12319 15614 12325
rect 16298 12316 16304 12328
rect 16356 12316 16362 12368
rect 17773 12359 17831 12365
rect 17773 12325 17785 12359
rect 17819 12356 17831 12359
rect 17862 12356 17868 12368
rect 17819 12328 17868 12356
rect 17819 12325 17831 12328
rect 17773 12319 17831 12325
rect 17862 12316 17868 12328
rect 17920 12316 17926 12368
rect 9306 12248 9312 12300
rect 9364 12288 9370 12300
rect 10045 12291 10103 12297
rect 10045 12288 10057 12291
rect 9364 12260 10057 12288
rect 9364 12248 9370 12260
rect 10045 12257 10057 12260
rect 10091 12257 10103 12291
rect 10045 12251 10103 12257
rect 12618 12248 12624 12300
rect 12676 12288 12682 12300
rect 13173 12291 13231 12297
rect 13173 12288 13185 12291
rect 12676 12260 13185 12288
rect 12676 12248 12682 12260
rect 13173 12257 13185 12260
rect 13219 12257 13231 12291
rect 13173 12251 13231 12257
rect 13262 12248 13268 12300
rect 13320 12288 13326 12300
rect 13320 12260 13365 12288
rect 13320 12248 13326 12260
rect 14182 12248 14188 12300
rect 14240 12288 14246 12300
rect 14553 12291 14611 12297
rect 14553 12288 14565 12291
rect 14240 12260 14565 12288
rect 14240 12248 14246 12260
rect 14553 12257 14565 12260
rect 14599 12257 14611 12291
rect 14553 12251 14611 12257
rect 16574 12248 16580 12300
rect 16632 12288 16638 12300
rect 17497 12291 17555 12297
rect 17497 12288 17509 12291
rect 16632 12260 17509 12288
rect 16632 12248 16638 12260
rect 17497 12257 17509 12260
rect 17543 12257 17555 12291
rect 17497 12251 17555 12257
rect 9217 12223 9275 12229
rect 9217 12189 9229 12223
rect 9263 12189 9275 12223
rect 9217 12183 9275 12189
rect 9398 12180 9404 12232
rect 9456 12220 9462 12232
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 9456 12192 10149 12220
rect 9456 12180 9462 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 10226 12180 10232 12232
rect 10284 12220 10290 12232
rect 10284 12192 10329 12220
rect 10284 12180 10290 12192
rect 10410 12180 10416 12232
rect 10468 12220 10474 12232
rect 11793 12223 11851 12229
rect 11793 12220 11805 12223
rect 10468 12192 11805 12220
rect 10468 12180 10474 12192
rect 11793 12189 11805 12192
rect 11839 12189 11851 12223
rect 11793 12183 11851 12189
rect 12710 12180 12716 12232
rect 12768 12220 12774 12232
rect 13357 12223 13415 12229
rect 13357 12220 13369 12223
rect 12768 12192 13369 12220
rect 12768 12180 12774 12192
rect 13357 12189 13369 12192
rect 13403 12189 13415 12223
rect 13357 12183 13415 12189
rect 15289 12223 15347 12229
rect 15289 12189 15301 12223
rect 15335 12189 15347 12223
rect 15289 12183 15347 12189
rect 8386 12152 8392 12164
rect 7116 12124 8392 12152
rect 8386 12112 8392 12124
rect 8444 12112 8450 12164
rect 10594 12152 10600 12164
rect 8496 12124 10600 12152
rect 5626 12044 5632 12096
rect 5684 12084 5690 12096
rect 8496 12084 8524 12124
rect 10594 12112 10600 12124
rect 10652 12112 10658 12164
rect 11241 12155 11299 12161
rect 11241 12121 11253 12155
rect 11287 12152 11299 12155
rect 11882 12152 11888 12164
rect 11287 12124 11888 12152
rect 11287 12121 11299 12124
rect 11241 12115 11299 12121
rect 11882 12112 11888 12124
rect 11940 12112 11946 12164
rect 13538 12112 13544 12164
rect 13596 12152 13602 12164
rect 14369 12155 14427 12161
rect 14369 12152 14381 12155
rect 13596 12124 14381 12152
rect 13596 12112 13602 12124
rect 14369 12121 14381 12124
rect 14415 12152 14427 12155
rect 14550 12152 14556 12164
rect 14415 12124 14556 12152
rect 14415 12121 14427 12124
rect 14369 12115 14427 12121
rect 14550 12112 14556 12124
rect 14608 12152 14614 12164
rect 15304 12152 15332 12183
rect 14608 12124 15332 12152
rect 14608 12112 14614 12124
rect 5684 12056 8524 12084
rect 9677 12087 9735 12093
rect 5684 12044 5690 12056
rect 9677 12053 9689 12087
rect 9723 12084 9735 12087
rect 10686 12084 10692 12096
rect 9723 12056 10692 12084
rect 9723 12053 9735 12056
rect 9677 12047 9735 12053
rect 10686 12044 10692 12056
rect 10744 12044 10750 12096
rect 12802 12044 12808 12096
rect 12860 12084 12866 12096
rect 12860 12056 12905 12084
rect 12860 12044 12866 12056
rect 14458 12044 14464 12096
rect 14516 12084 14522 12096
rect 16298 12084 16304 12096
rect 14516 12056 16304 12084
rect 14516 12044 14522 12056
rect 16298 12044 16304 12056
rect 16356 12044 16362 12096
rect 16666 12084 16672 12096
rect 16627 12056 16672 12084
rect 16666 12044 16672 12056
rect 16724 12044 16730 12096
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 1854 11840 1860 11892
rect 1912 11880 1918 11892
rect 1949 11883 2007 11889
rect 1949 11880 1961 11883
rect 1912 11852 1961 11880
rect 1912 11840 1918 11852
rect 1949 11849 1961 11852
rect 1995 11849 2007 11883
rect 1949 11843 2007 11849
rect 2774 11840 2780 11892
rect 2832 11880 2838 11892
rect 2961 11883 3019 11889
rect 2961 11880 2973 11883
rect 2832 11852 2973 11880
rect 2832 11840 2838 11852
rect 2961 11849 2973 11852
rect 3007 11849 3019 11883
rect 5534 11880 5540 11892
rect 2961 11843 3019 11849
rect 4264 11852 5540 11880
rect 3602 11744 3608 11756
rect 3515 11716 3608 11744
rect 3602 11704 3608 11716
rect 3660 11744 3666 11756
rect 4264 11744 4292 11852
rect 5534 11840 5540 11852
rect 5592 11840 5598 11892
rect 6825 11883 6883 11889
rect 6825 11849 6837 11883
rect 6871 11880 6883 11883
rect 9861 11883 9919 11889
rect 6871 11852 9536 11880
rect 6871 11849 6883 11852
rect 6825 11843 6883 11849
rect 3660 11716 4292 11744
rect 5552 11784 7512 11812
rect 3660 11704 3666 11716
rect 1765 11679 1823 11685
rect 1765 11645 1777 11679
rect 1811 11676 1823 11679
rect 2406 11676 2412 11688
rect 1811 11648 2412 11676
rect 1811 11645 1823 11648
rect 1765 11639 1823 11645
rect 2406 11636 2412 11648
rect 2464 11636 2470 11688
rect 3418 11636 3424 11688
rect 3476 11636 3482 11688
rect 4525 11679 4583 11685
rect 4525 11645 4537 11679
rect 4571 11645 4583 11679
rect 4525 11639 4583 11645
rect 3329 11611 3387 11617
rect 3329 11577 3341 11611
rect 3375 11608 3387 11611
rect 3436 11608 3464 11636
rect 3786 11608 3792 11620
rect 3375 11580 3792 11608
rect 3375 11577 3387 11580
rect 3329 11571 3387 11577
rect 3786 11568 3792 11580
rect 3844 11568 3850 11620
rect 4338 11568 4344 11620
rect 4396 11608 4402 11620
rect 4540 11608 4568 11639
rect 4614 11636 4620 11688
rect 4672 11676 4678 11688
rect 5552 11676 5580 11784
rect 7098 11704 7104 11756
rect 7156 11744 7162 11756
rect 7285 11747 7343 11753
rect 7285 11744 7297 11747
rect 7156 11716 7297 11744
rect 7156 11704 7162 11716
rect 7285 11713 7297 11716
rect 7331 11713 7343 11747
rect 7285 11707 7343 11713
rect 7377 11747 7435 11753
rect 7377 11713 7389 11747
rect 7423 11713 7435 11747
rect 7377 11707 7435 11713
rect 7190 11676 7196 11688
rect 4672 11648 5580 11676
rect 7151 11648 7196 11676
rect 4672 11636 4678 11648
rect 7190 11636 7196 11648
rect 7248 11636 7254 11688
rect 7392 11676 7420 11707
rect 7300 11648 7420 11676
rect 4396 11580 4568 11608
rect 4792 11611 4850 11617
rect 4396 11568 4402 11580
rect 4792 11577 4804 11611
rect 4838 11608 4850 11611
rect 6178 11608 6184 11620
rect 4838 11580 6184 11608
rect 4838 11577 4850 11580
rect 4792 11571 4850 11577
rect 6178 11568 6184 11580
rect 6236 11608 6242 11620
rect 7300 11608 7328 11648
rect 6236 11580 7328 11608
rect 7484 11608 7512 11784
rect 7742 11704 7748 11756
rect 7800 11744 7806 11756
rect 9508 11744 9536 11852
rect 9861 11849 9873 11883
rect 9907 11880 9919 11883
rect 12710 11880 12716 11892
rect 9907 11852 12716 11880
rect 9907 11849 9919 11852
rect 9861 11843 9919 11849
rect 12710 11840 12716 11852
rect 12768 11840 12774 11892
rect 14645 11883 14703 11889
rect 14645 11849 14657 11883
rect 14691 11880 14703 11883
rect 14734 11880 14740 11892
rect 14691 11852 14740 11880
rect 14691 11849 14703 11852
rect 14645 11843 14703 11849
rect 14734 11840 14740 11852
rect 14792 11840 14798 11892
rect 16206 11880 16212 11892
rect 16167 11852 16212 11880
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 16298 11840 16304 11892
rect 16356 11880 16362 11892
rect 16356 11852 16804 11880
rect 16356 11840 16362 11852
rect 10689 11815 10747 11821
rect 10689 11781 10701 11815
rect 10735 11812 10747 11815
rect 11882 11812 11888 11824
rect 10735 11784 11888 11812
rect 10735 11781 10747 11784
rect 10689 11775 10747 11781
rect 11882 11772 11888 11784
rect 11940 11772 11946 11824
rect 13814 11812 13820 11824
rect 13727 11784 13820 11812
rect 13814 11772 13820 11784
rect 13872 11812 13878 11824
rect 14366 11812 14372 11824
rect 13872 11784 14372 11812
rect 13872 11772 13878 11784
rect 14366 11772 14372 11784
rect 14424 11772 14430 11824
rect 10962 11744 10968 11756
rect 7800 11716 8616 11744
rect 9508 11716 10968 11744
rect 7800 11704 7806 11716
rect 8389 11679 8447 11685
rect 8389 11645 8401 11679
rect 8435 11676 8447 11679
rect 8481 11679 8539 11685
rect 8481 11676 8493 11679
rect 8435 11648 8493 11676
rect 8435 11645 8447 11648
rect 8389 11639 8447 11645
rect 8481 11645 8493 11648
rect 8527 11645 8539 11679
rect 8588 11676 8616 11716
rect 10962 11704 10968 11716
rect 11020 11704 11026 11756
rect 11146 11744 11152 11756
rect 11107 11716 11152 11744
rect 11146 11704 11152 11716
rect 11204 11704 11210 11756
rect 11330 11744 11336 11756
rect 11291 11716 11336 11744
rect 11330 11704 11336 11716
rect 11388 11704 11394 11756
rect 16776 11753 16804 11852
rect 15197 11747 15255 11753
rect 15197 11744 15209 11747
rect 13455 11716 15209 11744
rect 10318 11676 10324 11688
rect 8588 11648 10324 11676
rect 8481 11639 8539 11645
rect 10318 11636 10324 11648
rect 10376 11636 10382 11688
rect 12434 11636 12440 11688
rect 12492 11676 12498 11688
rect 12704 11679 12762 11685
rect 12492 11648 12537 11676
rect 12492 11636 12498 11648
rect 12704 11645 12716 11679
rect 12750 11676 12762 11679
rect 13455 11676 13483 11716
rect 15197 11713 15209 11716
rect 15243 11713 15255 11747
rect 15197 11707 15255 11713
rect 16761 11747 16819 11753
rect 16761 11713 16773 11747
rect 16807 11713 16819 11747
rect 16761 11707 16819 11713
rect 12750 11648 13483 11676
rect 12750 11645 12762 11648
rect 12704 11639 12762 11645
rect 7484 11580 8524 11608
rect 6236 11568 6242 11580
rect 3418 11540 3424 11552
rect 3379 11512 3424 11540
rect 3418 11500 3424 11512
rect 3476 11540 3482 11552
rect 3694 11540 3700 11552
rect 3476 11512 3700 11540
rect 3476 11500 3482 11512
rect 3694 11500 3700 11512
rect 3752 11500 3758 11552
rect 5902 11540 5908 11552
rect 5863 11512 5908 11540
rect 5902 11500 5908 11512
rect 5960 11500 5966 11552
rect 7190 11500 7196 11552
rect 7248 11540 7254 11552
rect 8389 11543 8447 11549
rect 8389 11540 8401 11543
rect 7248 11512 8401 11540
rect 7248 11500 7254 11512
rect 8389 11509 8401 11512
rect 8435 11509 8447 11543
rect 8496 11540 8524 11580
rect 8570 11568 8576 11620
rect 8628 11608 8634 11620
rect 8748 11611 8806 11617
rect 8748 11608 8760 11611
rect 8628 11580 8760 11608
rect 8628 11568 8634 11580
rect 8748 11577 8760 11580
rect 8794 11608 8806 11611
rect 10410 11608 10416 11620
rect 8794 11580 10416 11608
rect 8794 11577 8806 11580
rect 8748 11571 8806 11577
rect 10410 11568 10416 11580
rect 10468 11568 10474 11620
rect 10686 11568 10692 11620
rect 10744 11608 10750 11620
rect 11057 11611 11115 11617
rect 11057 11608 11069 11611
rect 10744 11580 11069 11608
rect 10744 11568 10750 11580
rect 11057 11577 11069 11580
rect 11103 11577 11115 11611
rect 11057 11571 11115 11577
rect 12158 11568 12164 11620
rect 12216 11608 12222 11620
rect 12719 11608 12747 11639
rect 14642 11636 14648 11688
rect 14700 11676 14706 11688
rect 15013 11679 15071 11685
rect 15013 11676 15025 11679
rect 14700 11648 15025 11676
rect 14700 11636 14706 11648
rect 15013 11645 15025 11648
rect 15059 11645 15071 11679
rect 15013 11639 15071 11645
rect 12216 11580 12747 11608
rect 12216 11568 12222 11580
rect 12802 11568 12808 11620
rect 12860 11608 12866 11620
rect 15105 11611 15163 11617
rect 15105 11608 15117 11611
rect 12860 11580 15117 11608
rect 12860 11568 12866 11580
rect 15105 11577 15117 11580
rect 15151 11577 15163 11611
rect 16669 11611 16727 11617
rect 16669 11608 16681 11611
rect 15105 11571 15163 11577
rect 15212 11580 16681 11608
rect 15212 11540 15240 11580
rect 16669 11577 16681 11580
rect 16715 11577 16727 11611
rect 16669 11571 16727 11577
rect 8496 11512 15240 11540
rect 8389 11503 8447 11509
rect 15286 11500 15292 11552
rect 15344 11540 15350 11552
rect 16577 11543 16635 11549
rect 16577 11540 16589 11543
rect 15344 11512 16589 11540
rect 15344 11500 15350 11512
rect 16577 11509 16589 11512
rect 16623 11509 16635 11543
rect 16577 11503 16635 11509
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 2869 11339 2927 11345
rect 2869 11305 2881 11339
rect 2915 11336 2927 11339
rect 4065 11339 4123 11345
rect 4065 11336 4077 11339
rect 2915 11308 4077 11336
rect 2915 11305 2927 11308
rect 2869 11299 2927 11305
rect 4065 11305 4077 11308
rect 4111 11305 4123 11339
rect 4525 11339 4583 11345
rect 4525 11336 4537 11339
rect 4065 11299 4123 11305
rect 4172 11308 4537 11336
rect 2314 11228 2320 11280
rect 2372 11268 2378 11280
rect 4172 11268 4200 11308
rect 4525 11305 4537 11308
rect 4571 11336 4583 11339
rect 4798 11336 4804 11348
rect 4571 11308 4804 11336
rect 4571 11305 4583 11308
rect 4525 11299 4583 11305
rect 4798 11296 4804 11308
rect 4856 11336 4862 11348
rect 8294 11336 8300 11348
rect 4856 11308 8300 11336
rect 4856 11296 4862 11308
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 8570 11336 8576 11348
rect 8531 11308 8576 11336
rect 8570 11296 8576 11308
rect 8628 11296 8634 11348
rect 8662 11296 8668 11348
rect 8720 11336 8726 11348
rect 11514 11336 11520 11348
rect 8720 11308 11520 11336
rect 8720 11296 8726 11308
rect 11514 11296 11520 11308
rect 11572 11296 11578 11348
rect 12526 11336 12532 11348
rect 12084 11308 12532 11336
rect 2372 11240 4200 11268
rect 2372 11228 2378 11240
rect 4246 11228 4252 11280
rect 4304 11268 4310 11280
rect 5534 11268 5540 11280
rect 4304 11240 5540 11268
rect 4304 11228 4310 11240
rect 5534 11228 5540 11240
rect 5592 11228 5598 11280
rect 10962 11268 10968 11280
rect 8763 11240 10968 11268
rect 2774 11160 2780 11212
rect 2832 11200 2838 11212
rect 4433 11203 4491 11209
rect 2832 11172 2877 11200
rect 2832 11160 2838 11172
rect 4433 11169 4445 11203
rect 4479 11200 4491 11203
rect 4522 11200 4528 11212
rect 4479 11172 4528 11200
rect 4479 11169 4491 11172
rect 4433 11163 4491 11169
rect 4522 11160 4528 11172
rect 4580 11160 4586 11212
rect 5997 11203 6055 11209
rect 5997 11169 6009 11203
rect 6043 11200 6055 11203
rect 7098 11200 7104 11212
rect 6043 11172 7104 11200
rect 6043 11169 6055 11172
rect 5997 11163 6055 11169
rect 7098 11160 7104 11172
rect 7156 11160 7162 11212
rect 7190 11160 7196 11212
rect 7248 11200 7254 11212
rect 7460 11203 7518 11209
rect 7248 11172 7293 11200
rect 7248 11160 7254 11172
rect 7460 11169 7472 11203
rect 7506 11200 7518 11203
rect 7506 11172 8248 11200
rect 7506 11169 7518 11172
rect 7460 11163 7518 11169
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11092 1458 11144
rect 2130 11092 2136 11144
rect 2188 11132 2194 11144
rect 2961 11135 3019 11141
rect 2961 11132 2973 11135
rect 2188 11104 2973 11132
rect 2188 11092 2194 11104
rect 2961 11101 2973 11104
rect 3007 11101 3019 11135
rect 2961 11095 3019 11101
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11132 4767 11135
rect 5902 11132 5908 11144
rect 4755 11104 5908 11132
rect 4755 11101 4767 11104
rect 4709 11095 4767 11101
rect 2409 11067 2467 11073
rect 2409 11033 2421 11067
rect 2455 11064 2467 11067
rect 4154 11064 4160 11076
rect 2455 11036 4160 11064
rect 2455 11033 2467 11036
rect 2409 11027 2467 11033
rect 4154 11024 4160 11036
rect 4212 11024 4218 11076
rect 3878 10956 3884 11008
rect 3936 10996 3942 11008
rect 4724 10996 4752 11095
rect 5902 11092 5908 11104
rect 5960 11092 5966 11144
rect 6086 11132 6092 11144
rect 6047 11104 6092 11132
rect 6086 11092 6092 11104
rect 6144 11092 6150 11144
rect 6270 11132 6276 11144
rect 6231 11104 6276 11132
rect 6270 11092 6276 11104
rect 6328 11092 6334 11144
rect 6914 11092 6920 11144
rect 6972 11132 6978 11144
rect 7208 11132 7236 11160
rect 6972 11104 7236 11132
rect 6972 11092 6978 11104
rect 8220 11076 8248 11172
rect 8294 11160 8300 11212
rect 8352 11200 8358 11212
rect 8763 11200 8791 11240
rect 10962 11228 10968 11240
rect 11020 11228 11026 11280
rect 11054 11228 11060 11280
rect 11112 11268 11118 11280
rect 11330 11268 11336 11280
rect 11112 11240 11336 11268
rect 11112 11228 11118 11240
rect 11330 11228 11336 11240
rect 11388 11228 11394 11280
rect 11698 11228 11704 11280
rect 11756 11268 11762 11280
rect 12084 11268 12112 11308
rect 12526 11296 12532 11308
rect 12584 11296 12590 11348
rect 14182 11336 14188 11348
rect 14143 11308 14188 11336
rect 14182 11296 14188 11308
rect 14240 11296 14246 11348
rect 17034 11296 17040 11348
rect 17092 11336 17098 11348
rect 17092 11308 18644 11336
rect 17092 11296 17098 11308
rect 11756 11240 12112 11268
rect 16384 11271 16442 11277
rect 11756 11228 11762 11240
rect 16384 11237 16396 11271
rect 16430 11268 16442 11271
rect 17954 11268 17960 11280
rect 16430 11240 17960 11268
rect 16430 11237 16442 11240
rect 16384 11231 16442 11237
rect 17954 11228 17960 11240
rect 18012 11228 18018 11280
rect 18616 11277 18644 11308
rect 18601 11271 18659 11277
rect 18601 11237 18613 11271
rect 18647 11237 18659 11271
rect 18601 11231 18659 11237
rect 8352 11172 8791 11200
rect 8352 11160 8358 11172
rect 8846 11160 8852 11212
rect 8904 11200 8910 11212
rect 10502 11200 10508 11212
rect 8904 11172 10508 11200
rect 8904 11160 8910 11172
rect 10502 11160 10508 11172
rect 10560 11160 10566 11212
rect 10680 11203 10738 11209
rect 10680 11169 10692 11203
rect 10726 11200 10738 11203
rect 12710 11200 12716 11212
rect 10726 11172 12716 11200
rect 10726 11169 10738 11172
rect 10680 11163 10738 11169
rect 12710 11160 12716 11172
rect 12768 11160 12774 11212
rect 12989 11203 13047 11209
rect 12989 11200 13001 11203
rect 12820 11172 13001 11200
rect 9674 11092 9680 11144
rect 9732 11132 9738 11144
rect 10413 11135 10471 11141
rect 10413 11132 10425 11135
rect 9732 11104 10425 11132
rect 9732 11092 9738 11104
rect 10413 11101 10425 11104
rect 10459 11101 10471 11135
rect 10413 11095 10471 11101
rect 8202 11024 8208 11076
rect 8260 11064 8266 11076
rect 10042 11064 10048 11076
rect 8260 11036 10048 11064
rect 8260 11024 8266 11036
rect 10042 11024 10048 11036
rect 10100 11024 10106 11076
rect 12820 11064 12848 11172
rect 12989 11169 13001 11172
rect 13035 11169 13047 11203
rect 12989 11163 13047 11169
rect 13446 11160 13452 11212
rect 13504 11200 13510 11212
rect 14369 11203 14427 11209
rect 14369 11200 14381 11203
rect 13504 11172 14381 11200
rect 13504 11160 13510 11172
rect 14369 11169 14381 11172
rect 14415 11169 14427 11203
rect 14369 11163 14427 11169
rect 14458 11160 14464 11212
rect 14516 11200 14522 11212
rect 18325 11203 18383 11209
rect 18325 11200 18337 11203
rect 14516 11172 18337 11200
rect 14516 11160 14522 11172
rect 18325 11169 18337 11172
rect 18371 11169 18383 11203
rect 18325 11163 18383 11169
rect 13078 11132 13084 11144
rect 13039 11104 13084 11132
rect 13078 11092 13084 11104
rect 13136 11092 13142 11144
rect 13170 11092 13176 11144
rect 13228 11132 13234 11144
rect 13228 11104 13273 11132
rect 13228 11092 13234 11104
rect 14550 11092 14556 11144
rect 14608 11132 14614 11144
rect 16117 11135 16175 11141
rect 16117 11132 16129 11135
rect 14608 11104 16129 11132
rect 14608 11092 14614 11104
rect 16117 11101 16129 11104
rect 16163 11101 16175 11135
rect 16117 11095 16175 11101
rect 11348 11036 12848 11064
rect 5626 10996 5632 11008
rect 3936 10968 4752 10996
rect 5587 10968 5632 10996
rect 3936 10956 3942 10968
rect 5626 10956 5632 10968
rect 5684 10956 5690 11008
rect 9950 10956 9956 11008
rect 10008 10996 10014 11008
rect 11348 10996 11376 11036
rect 10008 10968 11376 10996
rect 11793 10999 11851 11005
rect 10008 10956 10014 10968
rect 11793 10965 11805 10999
rect 11839 10996 11851 10999
rect 12158 10996 12164 11008
rect 11839 10968 12164 10996
rect 11839 10965 11851 10968
rect 11793 10959 11851 10965
rect 12158 10956 12164 10968
rect 12216 10956 12222 11008
rect 12526 10956 12532 11008
rect 12584 10996 12590 11008
rect 12621 10999 12679 11005
rect 12621 10996 12633 10999
rect 12584 10968 12633 10996
rect 12584 10956 12590 10968
rect 12621 10965 12633 10968
rect 12667 10965 12679 10999
rect 12621 10959 12679 10965
rect 12710 10956 12716 11008
rect 12768 10996 12774 11008
rect 17497 10999 17555 11005
rect 17497 10996 17509 10999
rect 12768 10968 17509 10996
rect 12768 10956 12774 10968
rect 17497 10965 17509 10968
rect 17543 10965 17555 10999
rect 17497 10959 17555 10965
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 2774 10752 2780 10804
rect 2832 10792 2838 10804
rect 3329 10795 3387 10801
rect 3329 10792 3341 10795
rect 2832 10764 3341 10792
rect 2832 10752 2838 10764
rect 3329 10761 3341 10764
rect 3375 10761 3387 10795
rect 8202 10792 8208 10804
rect 8163 10764 8208 10792
rect 3329 10755 3387 10761
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 9950 10792 9956 10804
rect 9600 10764 9956 10792
rect 9600 10736 9628 10764
rect 9950 10752 9956 10764
rect 10008 10752 10014 10804
rect 10042 10752 10048 10804
rect 10100 10792 10106 10804
rect 13170 10792 13176 10804
rect 10100 10764 13176 10792
rect 10100 10752 10106 10764
rect 13170 10752 13176 10764
rect 13228 10752 13234 10804
rect 4890 10724 4896 10736
rect 4851 10696 4896 10724
rect 4890 10684 4896 10696
rect 4948 10684 4954 10736
rect 9582 10684 9588 10736
rect 9640 10684 9646 10736
rect 2038 10656 2044 10668
rect 1999 10628 2044 10656
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 2130 10616 2136 10668
rect 2188 10656 2194 10668
rect 3878 10656 3884 10668
rect 2188 10628 2233 10656
rect 3839 10628 3884 10656
rect 2188 10616 2194 10628
rect 3878 10616 3884 10628
rect 3936 10616 3942 10668
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 5353 10659 5411 10665
rect 5353 10656 5365 10659
rect 4212 10628 5365 10656
rect 4212 10616 4218 10628
rect 5353 10625 5365 10628
rect 5399 10625 5411 10659
rect 5353 10619 5411 10625
rect 5442 10616 5448 10668
rect 5500 10656 5506 10668
rect 9033 10659 9091 10665
rect 5500 10628 5545 10656
rect 5644 10628 6960 10656
rect 5500 10616 5506 10628
rect 1394 10548 1400 10600
rect 1452 10588 1458 10600
rect 1949 10591 2007 10597
rect 1949 10588 1961 10591
rect 1452 10560 1961 10588
rect 1452 10548 1458 10560
rect 1949 10557 1961 10560
rect 1995 10557 2007 10591
rect 1949 10551 2007 10557
rect 3697 10591 3755 10597
rect 3697 10557 3709 10591
rect 3743 10588 3755 10591
rect 3786 10588 3792 10600
rect 3743 10560 3792 10588
rect 3743 10557 3755 10560
rect 3697 10551 3755 10557
rect 3786 10548 3792 10560
rect 3844 10548 3850 10600
rect 4062 10548 4068 10600
rect 4120 10588 4126 10600
rect 5644 10588 5672 10628
rect 4120 10560 5672 10588
rect 4120 10548 4126 10560
rect 6362 10548 6368 10600
rect 6420 10588 6426 10600
rect 6641 10591 6699 10597
rect 6641 10588 6653 10591
rect 6420 10560 6653 10588
rect 6420 10548 6426 10560
rect 6641 10557 6653 10560
rect 6687 10557 6699 10591
rect 6822 10588 6828 10600
rect 6783 10560 6828 10588
rect 6641 10551 6699 10557
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 6932 10588 6960 10628
rect 9033 10625 9045 10659
rect 9079 10656 9091 10659
rect 9122 10656 9128 10668
rect 9079 10628 9128 10656
rect 9079 10625 9091 10628
rect 9033 10619 9091 10625
rect 9122 10616 9128 10628
rect 9180 10616 9186 10668
rect 14001 10659 14059 10665
rect 14001 10625 14013 10659
rect 14047 10656 14059 10659
rect 14047 10628 15056 10656
rect 14047 10625 14059 10628
rect 14001 10619 14059 10625
rect 6932 10560 7236 10588
rect 5261 10523 5319 10529
rect 5261 10520 5273 10523
rect 1596 10492 5273 10520
rect 1596 10461 1624 10492
rect 5261 10489 5273 10492
rect 5307 10489 5319 10523
rect 5261 10483 5319 10489
rect 6270 10480 6276 10532
rect 6328 10520 6334 10532
rect 7070 10523 7128 10529
rect 7070 10520 7082 10523
rect 6328 10492 7082 10520
rect 6328 10480 6334 10492
rect 7070 10489 7082 10492
rect 7116 10489 7128 10523
rect 7208 10520 7236 10560
rect 9674 10548 9680 10600
rect 9732 10588 9738 10600
rect 10045 10591 10103 10597
rect 10045 10588 10057 10591
rect 9732 10560 10057 10588
rect 9732 10548 9738 10560
rect 10045 10557 10057 10560
rect 10091 10557 10103 10591
rect 10045 10551 10103 10557
rect 10312 10591 10370 10597
rect 10312 10557 10324 10591
rect 10358 10588 10370 10591
rect 11054 10588 11060 10600
rect 10358 10560 11060 10588
rect 10358 10557 10370 10560
rect 10312 10551 10370 10557
rect 11054 10548 11060 10560
rect 11112 10548 11118 10600
rect 12250 10548 12256 10600
rect 12308 10588 12314 10600
rect 13817 10591 13875 10597
rect 13817 10588 13829 10591
rect 12308 10560 13829 10588
rect 12308 10548 12314 10560
rect 13817 10557 13829 10560
rect 13863 10557 13875 10591
rect 13817 10551 13875 10557
rect 14550 10548 14556 10600
rect 14608 10588 14614 10600
rect 14921 10591 14979 10597
rect 14921 10588 14933 10591
rect 14608 10560 14933 10588
rect 14608 10548 14614 10560
rect 14921 10557 14933 10560
rect 14967 10557 14979 10591
rect 15028 10588 15056 10628
rect 15188 10591 15246 10597
rect 15188 10588 15200 10591
rect 15028 10560 15200 10588
rect 14921 10551 14979 10557
rect 15188 10557 15200 10560
rect 15234 10588 15246 10591
rect 16666 10588 16672 10600
rect 15234 10560 16672 10588
rect 15234 10557 15246 10560
rect 15188 10551 15246 10557
rect 16666 10548 16672 10560
rect 16724 10548 16730 10600
rect 12618 10520 12624 10532
rect 7208 10492 12624 10520
rect 7070 10483 7128 10489
rect 12618 10480 12624 10492
rect 12676 10480 12682 10532
rect 12894 10480 12900 10532
rect 12952 10520 12958 10532
rect 13725 10523 13783 10529
rect 13725 10520 13737 10523
rect 12952 10492 13737 10520
rect 12952 10480 12958 10492
rect 13725 10489 13737 10492
rect 13771 10489 13783 10523
rect 13725 10483 13783 10489
rect 1581 10455 1639 10461
rect 1581 10421 1593 10455
rect 1627 10421 1639 10455
rect 1581 10415 1639 10421
rect 3418 10412 3424 10464
rect 3476 10452 3482 10464
rect 3789 10455 3847 10461
rect 3789 10452 3801 10455
rect 3476 10424 3801 10452
rect 3476 10412 3482 10424
rect 3789 10421 3801 10424
rect 3835 10452 3847 10455
rect 3970 10452 3976 10464
rect 3835 10424 3976 10452
rect 3835 10421 3847 10424
rect 3789 10415 3847 10421
rect 3970 10412 3976 10424
rect 4028 10412 4034 10464
rect 6454 10452 6460 10464
rect 6415 10424 6460 10452
rect 6454 10412 6460 10424
rect 6512 10412 6518 10464
rect 6546 10412 6552 10464
rect 6604 10452 6610 10464
rect 11425 10455 11483 10461
rect 11425 10452 11437 10455
rect 6604 10424 11437 10452
rect 6604 10412 6610 10424
rect 11425 10421 11437 10424
rect 11471 10421 11483 10455
rect 11425 10415 11483 10421
rect 13357 10455 13415 10461
rect 13357 10421 13369 10455
rect 13403 10452 13415 10455
rect 16206 10452 16212 10464
rect 13403 10424 16212 10452
rect 13403 10421 13415 10424
rect 13357 10415 13415 10421
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 16301 10455 16359 10461
rect 16301 10421 16313 10455
rect 16347 10452 16359 10455
rect 16390 10452 16396 10464
rect 16347 10424 16396 10452
rect 16347 10421 16359 10424
rect 16301 10415 16359 10421
rect 16390 10412 16396 10424
rect 16448 10412 16454 10464
rect 18046 10452 18052 10464
rect 18007 10424 18052 10452
rect 18046 10412 18052 10424
rect 18104 10412 18110 10464
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 2130 10208 2136 10260
rect 2188 10248 2194 10260
rect 3145 10251 3203 10257
rect 3145 10248 3157 10251
rect 2188 10220 3157 10248
rect 2188 10208 2194 10220
rect 3145 10217 3157 10220
rect 3191 10217 3203 10251
rect 3145 10211 3203 10217
rect 6270 10208 6276 10260
rect 6328 10248 6334 10260
rect 6365 10251 6423 10257
rect 6365 10248 6377 10251
rect 6328 10220 6377 10248
rect 6328 10208 6334 10220
rect 6365 10217 6377 10220
rect 6411 10217 6423 10251
rect 6365 10211 6423 10217
rect 7098 10208 7104 10260
rect 7156 10248 7162 10260
rect 7193 10251 7251 10257
rect 7193 10248 7205 10251
rect 7156 10220 7205 10248
rect 7156 10208 7162 10220
rect 7193 10217 7205 10220
rect 7239 10217 7251 10251
rect 7193 10211 7251 10217
rect 7466 10208 7472 10260
rect 7524 10248 7530 10260
rect 7561 10251 7619 10257
rect 7561 10248 7573 10251
rect 7524 10220 7573 10248
rect 7524 10208 7530 10220
rect 7561 10217 7573 10220
rect 7607 10217 7619 10251
rect 7561 10211 7619 10217
rect 10045 10251 10103 10257
rect 10045 10217 10057 10251
rect 10091 10248 10103 10251
rect 10318 10248 10324 10260
rect 10091 10220 10324 10248
rect 10091 10217 10103 10220
rect 10045 10211 10103 10217
rect 10318 10208 10324 10220
rect 10376 10208 10382 10260
rect 11238 10208 11244 10260
rect 11296 10248 11302 10260
rect 11609 10251 11667 10257
rect 11609 10248 11621 10251
rect 11296 10220 11621 10248
rect 11296 10208 11302 10220
rect 11609 10217 11621 10220
rect 11655 10248 11667 10251
rect 11790 10248 11796 10260
rect 11655 10220 11796 10248
rect 11655 10217 11667 10220
rect 11609 10211 11667 10217
rect 11790 10208 11796 10220
rect 11848 10208 11854 10260
rect 13633 10251 13691 10257
rect 13633 10217 13645 10251
rect 13679 10217 13691 10251
rect 13633 10211 13691 10217
rect 16209 10251 16267 10257
rect 16209 10217 16221 10251
rect 16255 10248 16267 10251
rect 18046 10248 18052 10260
rect 16255 10220 18052 10248
rect 16255 10217 16267 10220
rect 16209 10211 16267 10217
rect 2032 10183 2090 10189
rect 2032 10149 2044 10183
rect 2078 10180 2090 10183
rect 3878 10180 3884 10192
rect 2078 10152 3884 10180
rect 2078 10149 2090 10152
rect 2032 10143 2090 10149
rect 3878 10140 3884 10152
rect 3936 10140 3942 10192
rect 4982 10140 4988 10192
rect 5040 10180 5046 10192
rect 5252 10183 5310 10189
rect 5252 10180 5264 10183
rect 5040 10152 5264 10180
rect 5040 10140 5046 10152
rect 5252 10149 5264 10152
rect 5298 10180 5310 10183
rect 11701 10183 11759 10189
rect 5298 10152 7788 10180
rect 5298 10149 5310 10152
rect 5252 10143 5310 10149
rect 1765 10115 1823 10121
rect 1765 10081 1777 10115
rect 1811 10112 1823 10115
rect 2406 10112 2412 10124
rect 1811 10084 2412 10112
rect 1811 10081 1823 10084
rect 1765 10075 1823 10081
rect 2406 10072 2412 10084
rect 2464 10072 2470 10124
rect 5534 10072 5540 10124
rect 5592 10112 5598 10124
rect 7653 10115 7711 10121
rect 7653 10112 7665 10115
rect 5592 10084 7665 10112
rect 5592 10072 5598 10084
rect 7653 10081 7665 10084
rect 7699 10081 7711 10115
rect 7653 10075 7711 10081
rect 7760 10056 7788 10152
rect 11701 10149 11713 10183
rect 11747 10180 11759 10183
rect 12250 10180 12256 10192
rect 11747 10152 12256 10180
rect 11747 10149 11759 10152
rect 11701 10143 11759 10149
rect 12250 10140 12256 10152
rect 12308 10140 12314 10192
rect 13648 10180 13676 10211
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 13648 10152 17448 10180
rect 10318 10112 10324 10124
rect 10231 10084 10324 10112
rect 4338 10004 4344 10056
rect 4396 10044 4402 10056
rect 4985 10047 5043 10053
rect 4985 10044 4997 10047
rect 4396 10016 4997 10044
rect 4396 10004 4402 10016
rect 4985 10013 4997 10016
rect 5031 10013 5043 10047
rect 4985 10007 5043 10013
rect 7742 10004 7748 10056
rect 7800 10044 7806 10056
rect 10244 10053 10272 10084
rect 10318 10072 10324 10084
rect 10376 10112 10382 10124
rect 14001 10115 14059 10121
rect 10376 10084 11928 10112
rect 10376 10072 10382 10084
rect 11900 10053 11928 10084
rect 14001 10081 14013 10115
rect 14047 10112 14059 10115
rect 15286 10112 15292 10124
rect 14047 10084 15292 10112
rect 14047 10081 14059 10084
rect 14001 10075 14059 10081
rect 15286 10072 15292 10084
rect 15344 10072 15350 10124
rect 16206 10072 16212 10124
rect 16264 10112 16270 10124
rect 17420 10121 17448 10152
rect 17494 10140 17500 10192
rect 17552 10180 17558 10192
rect 17681 10183 17739 10189
rect 17681 10180 17693 10183
rect 17552 10152 17693 10180
rect 17552 10140 17558 10152
rect 17681 10149 17693 10152
rect 17727 10149 17739 10183
rect 17681 10143 17739 10149
rect 16301 10115 16359 10121
rect 16301 10112 16313 10115
rect 16264 10084 16313 10112
rect 16264 10072 16270 10084
rect 16301 10081 16313 10084
rect 16347 10081 16359 10115
rect 16301 10075 16359 10081
rect 17405 10115 17463 10121
rect 17405 10081 17417 10115
rect 17451 10081 17463 10115
rect 17405 10075 17463 10081
rect 10137 10047 10195 10053
rect 7800 10016 7845 10044
rect 7800 10004 7806 10016
rect 10137 10013 10149 10047
rect 10183 10013 10195 10047
rect 10137 10007 10195 10013
rect 10229 10047 10287 10053
rect 10229 10013 10241 10047
rect 10275 10013 10287 10047
rect 10229 10007 10287 10013
rect 11885 10047 11943 10053
rect 11885 10013 11897 10047
rect 11931 10013 11943 10047
rect 14090 10044 14096 10056
rect 14051 10016 14096 10044
rect 11885 10007 11943 10013
rect 7374 9936 7380 9988
rect 7432 9976 7438 9988
rect 10152 9976 10180 10007
rect 7432 9948 10180 9976
rect 11900 9976 11928 10007
rect 14090 10004 14096 10016
rect 14148 10004 14154 10056
rect 14277 10047 14335 10053
rect 14277 10013 14289 10047
rect 14323 10044 14335 10047
rect 14734 10044 14740 10056
rect 14323 10016 14740 10044
rect 14323 10013 14335 10016
rect 14277 10007 14335 10013
rect 14734 10004 14740 10016
rect 14792 10004 14798 10056
rect 16390 10004 16396 10056
rect 16448 10044 16454 10056
rect 16448 10016 16493 10044
rect 16448 10004 16454 10016
rect 12710 9976 12716 9988
rect 11900 9948 12716 9976
rect 7432 9936 7438 9948
rect 12710 9936 12716 9948
rect 12768 9936 12774 9988
rect 15841 9979 15899 9985
rect 15841 9945 15853 9979
rect 15887 9976 15899 9979
rect 16574 9976 16580 9988
rect 15887 9948 16580 9976
rect 15887 9945 15899 9948
rect 15841 9939 15899 9945
rect 16574 9936 16580 9948
rect 16632 9936 16638 9988
rect 3694 9868 3700 9920
rect 3752 9908 3758 9920
rect 8846 9908 8852 9920
rect 3752 9880 8852 9908
rect 3752 9868 3758 9880
rect 8846 9868 8852 9880
rect 8904 9868 8910 9920
rect 9677 9911 9735 9917
rect 9677 9877 9689 9911
rect 9723 9908 9735 9911
rect 11054 9908 11060 9920
rect 9723 9880 11060 9908
rect 9723 9877 9735 9880
rect 9677 9871 9735 9877
rect 11054 9868 11060 9880
rect 11112 9868 11118 9920
rect 11238 9908 11244 9920
rect 11199 9880 11244 9908
rect 11238 9868 11244 9880
rect 11296 9868 11302 9920
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 4338 9704 4344 9716
rect 1412 9676 2452 9704
rect 1412 9577 1440 9676
rect 2424 9648 2452 9676
rect 3620 9676 4344 9704
rect 2406 9596 2412 9648
rect 2464 9636 2470 9648
rect 3620 9636 3648 9676
rect 4338 9664 4344 9676
rect 4396 9664 4402 9716
rect 4982 9704 4988 9716
rect 4943 9676 4988 9704
rect 4982 9664 4988 9676
rect 5040 9664 5046 9716
rect 6457 9707 6515 9713
rect 6457 9673 6469 9707
rect 6503 9704 6515 9707
rect 6914 9704 6920 9716
rect 6503 9676 6920 9704
rect 6503 9673 6515 9676
rect 6457 9667 6515 9673
rect 6914 9664 6920 9676
rect 6972 9664 6978 9716
rect 10594 9664 10600 9716
rect 10652 9704 10658 9716
rect 15194 9704 15200 9716
rect 10652 9676 15200 9704
rect 10652 9664 10658 9676
rect 15194 9664 15200 9676
rect 15252 9664 15258 9716
rect 2464 9608 3648 9636
rect 2464 9596 2470 9608
rect 3620 9577 3648 9608
rect 6086 9596 6092 9648
rect 6144 9636 6150 9648
rect 6825 9639 6883 9645
rect 6825 9636 6837 9639
rect 6144 9608 6837 9636
rect 6144 9596 6150 9608
rect 6825 9605 6837 9608
rect 6871 9605 6883 9639
rect 6825 9599 6883 9605
rect 7190 9596 7196 9648
rect 7248 9636 7254 9648
rect 8386 9636 8392 9648
rect 7248 9608 8392 9636
rect 7248 9596 7254 9608
rect 8386 9596 8392 9608
rect 8444 9596 8450 9648
rect 9953 9639 10011 9645
rect 9953 9605 9965 9639
rect 9999 9636 10011 9639
rect 10226 9636 10232 9648
rect 9999 9608 10232 9636
rect 9999 9605 10011 9608
rect 9953 9599 10011 9605
rect 10226 9596 10232 9608
rect 10284 9596 10290 9648
rect 10781 9639 10839 9645
rect 10781 9605 10793 9639
rect 10827 9636 10839 9639
rect 11146 9636 11152 9648
rect 10827 9608 11152 9636
rect 10827 9605 10839 9608
rect 10781 9599 10839 9605
rect 11146 9596 11152 9608
rect 11204 9596 11210 9648
rect 17954 9596 17960 9648
rect 18012 9636 18018 9648
rect 18417 9639 18475 9645
rect 18417 9636 18429 9639
rect 18012 9608 18429 9636
rect 18012 9596 18018 9608
rect 18417 9605 18429 9608
rect 18463 9605 18475 9639
rect 18417 9599 18475 9605
rect 1397 9571 1455 9577
rect 1397 9537 1409 9571
rect 1443 9537 1455 9571
rect 1397 9531 1455 9537
rect 3605 9571 3663 9577
rect 3605 9537 3617 9571
rect 3651 9537 3663 9571
rect 3605 9531 3663 9537
rect 7285 9571 7343 9577
rect 7285 9537 7297 9571
rect 7331 9568 7343 9571
rect 7374 9568 7380 9580
rect 7331 9540 7380 9568
rect 7331 9537 7343 9540
rect 7285 9531 7343 9537
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9568 7527 9571
rect 7742 9568 7748 9580
rect 7515 9540 7748 9568
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 7742 9528 7748 9540
rect 7800 9528 7806 9580
rect 10244 9568 10272 9596
rect 11333 9571 11391 9577
rect 11333 9568 11345 9571
rect 10244 9540 11345 9568
rect 11333 9537 11345 9540
rect 11379 9537 11391 9571
rect 11333 9531 11391 9537
rect 14550 9528 14556 9580
rect 14608 9568 14614 9580
rect 15749 9571 15807 9577
rect 15749 9568 15761 9571
rect 14608 9540 15761 9568
rect 14608 9528 14614 9540
rect 15749 9537 15761 9540
rect 15795 9537 15807 9571
rect 15749 9531 15807 9537
rect 1664 9503 1722 9509
rect 1664 9469 1676 9503
rect 1710 9500 1722 9503
rect 2130 9500 2136 9512
rect 1710 9472 2136 9500
rect 1710 9469 1722 9472
rect 1664 9463 1722 9469
rect 2130 9460 2136 9472
rect 2188 9460 2194 9512
rect 3872 9503 3930 9509
rect 3872 9500 3884 9503
rect 3804 9472 3884 9500
rect 2777 9367 2835 9373
rect 2777 9333 2789 9367
rect 2823 9364 2835 9367
rect 3804 9364 3832 9472
rect 3872 9469 3884 9472
rect 3918 9500 3930 9503
rect 5442 9500 5448 9512
rect 3918 9472 5448 9500
rect 3918 9469 3930 9472
rect 3872 9463 3930 9469
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 6454 9460 6460 9512
rect 6512 9500 6518 9512
rect 6641 9503 6699 9509
rect 6641 9500 6653 9503
rect 6512 9472 6653 9500
rect 6512 9460 6518 9472
rect 6641 9469 6653 9472
rect 6687 9469 6699 9503
rect 6641 9463 6699 9469
rect 6914 9460 6920 9512
rect 6972 9500 6978 9512
rect 8573 9503 8631 9509
rect 8573 9500 8585 9503
rect 6972 9472 8585 9500
rect 6972 9460 6978 9472
rect 8573 9469 8585 9472
rect 8619 9469 8631 9503
rect 8573 9463 8631 9469
rect 8840 9503 8898 9509
rect 8840 9469 8852 9503
rect 8886 9500 8898 9503
rect 9766 9500 9772 9512
rect 8886 9472 9772 9500
rect 8886 9469 8898 9472
rect 8840 9463 8898 9469
rect 9766 9460 9772 9472
rect 9824 9500 9830 9512
rect 10318 9500 10324 9512
rect 9824 9472 10324 9500
rect 9824 9460 9830 9472
rect 10318 9460 10324 9472
rect 10376 9460 10382 9512
rect 11149 9503 11207 9509
rect 11149 9469 11161 9503
rect 11195 9500 11207 9503
rect 11238 9500 11244 9512
rect 11195 9472 11244 9500
rect 11195 9469 11207 9472
rect 11149 9463 11207 9469
rect 11238 9460 11244 9472
rect 11296 9460 11302 9512
rect 12066 9460 12072 9512
rect 12124 9500 12130 9512
rect 12250 9500 12256 9512
rect 12124 9472 12256 9500
rect 12124 9460 12130 9472
rect 12250 9460 12256 9472
rect 12308 9460 12314 9512
rect 13173 9503 13231 9509
rect 13173 9469 13185 9503
rect 13219 9500 13231 9503
rect 14568 9500 14596 9528
rect 13219 9472 14596 9500
rect 16016 9503 16074 9509
rect 13219 9469 13231 9472
rect 13173 9463 13231 9469
rect 16016 9469 16028 9503
rect 16062 9500 16074 9503
rect 16390 9500 16396 9512
rect 16062 9472 16396 9500
rect 16062 9469 16074 9472
rect 16016 9463 16074 9469
rect 16390 9460 16396 9472
rect 16448 9460 16454 9512
rect 18138 9460 18144 9512
rect 18196 9500 18202 9512
rect 18233 9503 18291 9509
rect 18233 9500 18245 9503
rect 18196 9472 18245 9500
rect 18196 9460 18202 9472
rect 18233 9469 18245 9472
rect 18279 9469 18291 9503
rect 18233 9463 18291 9469
rect 4062 9392 4068 9444
rect 4120 9432 4126 9444
rect 12894 9432 12900 9444
rect 4120 9404 7420 9432
rect 4120 9392 4126 9404
rect 7190 9364 7196 9376
rect 2823 9336 3832 9364
rect 7151 9336 7196 9364
rect 2823 9333 2835 9336
rect 2777 9327 2835 9333
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 7392 9364 7420 9404
rect 8956 9404 12900 9432
rect 8956 9364 8984 9404
rect 12894 9392 12900 9404
rect 12952 9392 12958 9444
rect 13262 9392 13268 9444
rect 13320 9432 13326 9444
rect 13440 9435 13498 9441
rect 13440 9432 13452 9435
rect 13320 9404 13452 9432
rect 13320 9392 13326 9404
rect 13440 9401 13452 9404
rect 13486 9432 13498 9435
rect 13486 9404 17172 9432
rect 13486 9401 13498 9404
rect 13440 9395 13498 9401
rect 7392 9336 8984 9364
rect 11054 9324 11060 9376
rect 11112 9364 11118 9376
rect 11241 9367 11299 9373
rect 11241 9364 11253 9367
rect 11112 9336 11253 9364
rect 11112 9324 11118 9336
rect 11241 9333 11253 9336
rect 11287 9333 11299 9367
rect 11241 9327 11299 9333
rect 12066 9324 12072 9376
rect 12124 9364 12130 9376
rect 14182 9364 14188 9376
rect 12124 9336 14188 9364
rect 12124 9324 12130 9336
rect 14182 9324 14188 9336
rect 14240 9324 14246 9376
rect 14553 9367 14611 9373
rect 14553 9333 14565 9367
rect 14599 9364 14611 9367
rect 14734 9364 14740 9376
rect 14599 9336 14740 9364
rect 14599 9333 14611 9336
rect 14553 9327 14611 9333
rect 14734 9324 14740 9336
rect 14792 9324 14798 9376
rect 17144 9373 17172 9404
rect 17129 9367 17187 9373
rect 17129 9333 17141 9367
rect 17175 9333 17187 9367
rect 17129 9327 17187 9333
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 1949 9163 2007 9169
rect 1949 9129 1961 9163
rect 1995 9160 2007 9163
rect 3326 9160 3332 9172
rect 1995 9132 3332 9160
rect 1995 9129 2007 9132
rect 1949 9123 2007 9129
rect 3326 9120 3332 9132
rect 3384 9120 3390 9172
rect 4338 9120 4344 9172
rect 4396 9160 4402 9172
rect 4982 9160 4988 9172
rect 4396 9132 4988 9160
rect 4396 9120 4402 9132
rect 4982 9120 4988 9132
rect 5040 9160 5046 9172
rect 6089 9163 6147 9169
rect 6089 9160 6101 9163
rect 5040 9132 6101 9160
rect 5040 9120 5046 9132
rect 6089 9129 6101 9132
rect 6135 9129 6147 9163
rect 6089 9123 6147 9129
rect 6917 9163 6975 9169
rect 6917 9129 6929 9163
rect 6963 9129 6975 9163
rect 6917 9123 6975 9129
rect 8573 9163 8631 9169
rect 8573 9129 8585 9163
rect 8619 9160 8631 9163
rect 9306 9160 9312 9172
rect 8619 9132 9312 9160
rect 8619 9129 8631 9132
rect 8573 9123 8631 9129
rect 6932 9092 6960 9123
rect 9306 9120 9312 9132
rect 9364 9120 9370 9172
rect 11054 9160 11060 9172
rect 11015 9132 11060 9160
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 11606 9120 11612 9172
rect 11664 9160 11670 9172
rect 11885 9163 11943 9169
rect 11885 9160 11897 9163
rect 11664 9132 11897 9160
rect 11664 9120 11670 9132
rect 11885 9129 11897 9132
rect 11931 9160 11943 9163
rect 11974 9160 11980 9172
rect 11931 9132 11980 9160
rect 11931 9129 11943 9132
rect 11885 9123 11943 9129
rect 11974 9120 11980 9132
rect 12032 9120 12038 9172
rect 12621 9163 12679 9169
rect 12621 9129 12633 9163
rect 12667 9160 12679 9163
rect 14090 9160 14096 9172
rect 12667 9132 14096 9160
rect 12667 9129 12679 9132
rect 12621 9123 12679 9129
rect 14090 9120 14096 9132
rect 14148 9120 14154 9172
rect 12158 9092 12164 9104
rect 6932 9064 12164 9092
rect 12158 9052 12164 9064
rect 12216 9052 12222 9104
rect 18138 9092 18144 9104
rect 18099 9064 18144 9092
rect 18138 9052 18144 9064
rect 18196 9052 18202 9104
rect 1765 9027 1823 9033
rect 1765 8993 1777 9027
rect 1811 9024 1823 9027
rect 2222 9024 2228 9036
rect 1811 8996 2228 9024
rect 1811 8993 1823 8996
rect 1765 8987 1823 8993
rect 2222 8984 2228 8996
rect 2280 8984 2286 9036
rect 4893 9027 4951 9033
rect 4893 8993 4905 9027
rect 4939 9024 4951 9027
rect 5258 9024 5264 9036
rect 4939 8996 5264 9024
rect 4939 8993 4951 8996
rect 4893 8987 4951 8993
rect 5258 8984 5264 8996
rect 5316 8984 5322 9036
rect 6273 9027 6331 9033
rect 6273 8993 6285 9027
rect 6319 9024 6331 9027
rect 6454 9024 6460 9036
rect 6319 8996 6460 9024
rect 6319 8993 6331 8996
rect 6273 8987 6331 8993
rect 6454 8984 6460 8996
rect 6512 8984 6518 9036
rect 7282 9024 7288 9036
rect 7243 8996 7288 9024
rect 7282 8984 7288 8996
rect 7340 8984 7346 9036
rect 9674 8984 9680 9036
rect 9732 9024 9738 9036
rect 9944 9027 10002 9033
rect 9732 8996 9777 9024
rect 9732 8984 9738 8996
rect 9944 8993 9956 9027
rect 9990 9024 10002 9027
rect 10226 9024 10232 9036
rect 9990 8996 10232 9024
rect 9990 8993 10002 8996
rect 9944 8987 10002 8993
rect 10226 8984 10232 8996
rect 10284 8984 10290 9036
rect 12066 9024 12072 9036
rect 12027 8996 12072 9024
rect 12066 8984 12072 8996
rect 12124 8984 12130 9036
rect 12989 9027 13047 9033
rect 12989 8993 13001 9027
rect 13035 8993 13047 9027
rect 12989 8987 13047 8993
rect 2866 8956 2872 8968
rect 2827 8928 2872 8956
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 3694 8916 3700 8968
rect 3752 8956 3758 8968
rect 4985 8959 5043 8965
rect 4985 8956 4997 8959
rect 3752 8928 4997 8956
rect 3752 8916 3758 8928
rect 4985 8925 4997 8928
rect 5031 8925 5043 8959
rect 5166 8956 5172 8968
rect 5127 8928 5172 8956
rect 4985 8919 5043 8925
rect 5166 8916 5172 8928
rect 5224 8916 5230 8968
rect 7098 8916 7104 8968
rect 7156 8956 7162 8968
rect 7377 8959 7435 8965
rect 7377 8956 7389 8959
rect 7156 8928 7389 8956
rect 7156 8916 7162 8928
rect 7377 8925 7389 8928
rect 7423 8925 7435 8959
rect 7377 8919 7435 8925
rect 7561 8959 7619 8965
rect 7561 8925 7573 8959
rect 7607 8956 7619 8959
rect 8202 8956 8208 8968
rect 7607 8928 8208 8956
rect 7607 8925 7619 8928
rect 7561 8919 7619 8925
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 13004 8956 13032 8987
rect 15194 8984 15200 9036
rect 15252 9024 15258 9036
rect 15289 9027 15347 9033
rect 15289 9024 15301 9027
rect 15252 8996 15301 9024
rect 15252 8984 15258 8996
rect 15289 8993 15301 8996
rect 15335 8993 15347 9027
rect 16574 9024 16580 9036
rect 16535 8996 16580 9024
rect 15289 8987 15347 8993
rect 16574 8984 16580 8996
rect 16632 8984 16638 9036
rect 17402 9024 17408 9036
rect 16684 8996 17408 9024
rect 10796 8928 13032 8956
rect 13081 8959 13139 8965
rect 4525 8891 4583 8897
rect 4525 8857 4537 8891
rect 4571 8888 4583 8891
rect 8478 8888 8484 8900
rect 4571 8860 8484 8888
rect 4571 8857 4583 8860
rect 4525 8851 4583 8857
rect 8478 8848 8484 8860
rect 8536 8848 8542 8900
rect 3510 8780 3516 8832
rect 3568 8820 3574 8832
rect 10796 8820 10824 8928
rect 13081 8925 13093 8959
rect 13127 8925 13139 8959
rect 13262 8956 13268 8968
rect 13223 8928 13268 8956
rect 13081 8919 13139 8925
rect 10870 8848 10876 8900
rect 10928 8888 10934 8900
rect 13096 8888 13124 8919
rect 13262 8916 13268 8928
rect 13320 8916 13326 8968
rect 14182 8956 14188 8968
rect 14143 8928 14188 8956
rect 14182 8916 14188 8928
rect 14240 8916 14246 8968
rect 15565 8959 15623 8965
rect 15565 8925 15577 8959
rect 15611 8956 15623 8959
rect 16684 8956 16712 8996
rect 17402 8984 17408 8996
rect 17460 8984 17466 9036
rect 17862 9024 17868 9036
rect 17823 8996 17868 9024
rect 17862 8984 17868 8996
rect 17920 8984 17926 9036
rect 15611 8928 16712 8956
rect 16853 8959 16911 8965
rect 15611 8925 15623 8928
rect 15565 8919 15623 8925
rect 16853 8925 16865 8959
rect 16899 8956 16911 8959
rect 18598 8956 18604 8968
rect 16899 8928 18604 8956
rect 16899 8925 16911 8928
rect 16853 8919 16911 8925
rect 18598 8916 18604 8928
rect 18656 8916 18662 8968
rect 10928 8860 13124 8888
rect 10928 8848 10934 8860
rect 3568 8792 10824 8820
rect 3568 8780 3574 8792
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 3694 8616 3700 8628
rect 3655 8588 3700 8616
rect 3694 8576 3700 8588
rect 3752 8576 3758 8628
rect 7098 8616 7104 8628
rect 7059 8588 7104 8616
rect 7098 8576 7104 8588
rect 7156 8576 7162 8628
rect 8478 8576 8484 8628
rect 8536 8616 8542 8628
rect 8536 8588 15700 8616
rect 8536 8576 8542 8588
rect 3970 8508 3976 8560
rect 4028 8548 4034 8560
rect 8665 8551 8723 8557
rect 4028 8520 7880 8548
rect 4028 8508 4034 8520
rect 2222 8480 2228 8492
rect 2183 8452 2228 8480
rect 2222 8440 2228 8452
rect 2280 8440 2286 8492
rect 3786 8440 3792 8492
rect 3844 8480 3850 8492
rect 4157 8483 4215 8489
rect 4157 8480 4169 8483
rect 3844 8452 4169 8480
rect 3844 8440 3850 8452
rect 4157 8449 4169 8452
rect 4203 8449 4215 8483
rect 4338 8480 4344 8492
rect 4299 8452 4344 8480
rect 4157 8443 4215 8449
rect 4338 8440 4344 8452
rect 4396 8440 4402 8492
rect 5258 8480 5264 8492
rect 5219 8452 5264 8480
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 7374 8440 7380 8492
rect 7432 8480 7438 8492
rect 7561 8483 7619 8489
rect 7561 8480 7573 8483
rect 7432 8452 7573 8480
rect 7432 8440 7438 8452
rect 7561 8449 7573 8452
rect 7607 8449 7619 8483
rect 7742 8480 7748 8492
rect 7703 8452 7748 8480
rect 7561 8443 7619 8449
rect 7742 8440 7748 8452
rect 7800 8440 7806 8492
rect 7852 8480 7880 8520
rect 8665 8517 8677 8551
rect 8711 8548 8723 8551
rect 9398 8548 9404 8560
rect 8711 8520 9404 8548
rect 8711 8517 8723 8520
rect 8665 8511 8723 8517
rect 9398 8508 9404 8520
rect 9456 8508 9462 8560
rect 10781 8551 10839 8557
rect 10781 8517 10793 8551
rect 10827 8548 10839 8551
rect 11698 8548 11704 8560
rect 10827 8520 11704 8548
rect 10827 8517 10839 8520
rect 10781 8511 10839 8517
rect 11698 8508 11704 8520
rect 11756 8508 11762 8560
rect 11974 8508 11980 8560
rect 12032 8548 12038 8560
rect 12032 8520 12480 8548
rect 12032 8508 12038 8520
rect 9309 8483 9367 8489
rect 7852 8452 9076 8480
rect 2041 8415 2099 8421
rect 2041 8381 2053 8415
rect 2087 8412 2099 8415
rect 8938 8412 8944 8424
rect 2087 8384 8944 8412
rect 2087 8381 2099 8384
rect 2041 8375 2099 8381
rect 8938 8372 8944 8384
rect 8996 8372 9002 8424
rect 9048 8412 9076 8452
rect 9309 8449 9321 8483
rect 9355 8480 9367 8483
rect 9766 8480 9772 8492
rect 9355 8452 9772 8480
rect 9355 8449 9367 8452
rect 9309 8443 9367 8449
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 12452 8489 12480 8520
rect 11425 8483 11483 8489
rect 11425 8449 11437 8483
rect 11471 8480 11483 8483
rect 12437 8483 12495 8489
rect 11471 8452 12296 8480
rect 11471 8449 11483 8452
rect 11425 8443 11483 8449
rect 10870 8412 10876 8424
rect 9048 8384 10876 8412
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 7469 8347 7527 8353
rect 7469 8313 7481 8347
rect 7515 8344 7527 8347
rect 8386 8344 8392 8356
rect 7515 8316 8392 8344
rect 7515 8313 7527 8316
rect 7469 8307 7527 8313
rect 8386 8304 8392 8316
rect 8444 8344 8450 8356
rect 9125 8347 9183 8353
rect 9125 8344 9137 8347
rect 8444 8316 9137 8344
rect 8444 8304 8450 8316
rect 9125 8313 9137 8316
rect 9171 8313 9183 8347
rect 9125 8307 9183 8313
rect 11241 8347 11299 8353
rect 11241 8313 11253 8347
rect 11287 8344 11299 8347
rect 11790 8344 11796 8356
rect 11287 8316 11796 8344
rect 11287 8313 11299 8316
rect 11241 8307 11299 8313
rect 11790 8304 11796 8316
rect 11848 8304 11854 8356
rect 12268 8344 12296 8452
rect 12437 8449 12449 8483
rect 12483 8449 12495 8483
rect 12437 8443 12495 8449
rect 14550 8440 14556 8492
rect 14608 8480 14614 8492
rect 14645 8483 14703 8489
rect 14645 8480 14657 8483
rect 14608 8452 14657 8480
rect 14608 8440 14614 8452
rect 14645 8449 14657 8452
rect 14691 8449 14703 8483
rect 14645 8443 14703 8449
rect 15672 8412 15700 8588
rect 19426 8576 19432 8628
rect 19484 8616 19490 8628
rect 19521 8619 19579 8625
rect 19521 8616 19533 8619
rect 19484 8588 19533 8616
rect 19484 8576 19490 8588
rect 19521 8585 19533 8588
rect 19567 8585 19579 8619
rect 19521 8579 19579 8585
rect 18046 8508 18052 8560
rect 18104 8548 18110 8560
rect 18104 8520 18276 8548
rect 18104 8508 18110 8520
rect 18248 8489 18276 8520
rect 18233 8483 18291 8489
rect 18233 8449 18245 8483
rect 18279 8449 18291 8483
rect 18233 8443 18291 8449
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 15672 8384 18061 8412
rect 18049 8381 18061 8384
rect 18095 8381 18107 8415
rect 19334 8412 19340 8424
rect 19295 8384 19340 8412
rect 18049 8375 18107 8381
rect 19334 8372 19340 8384
rect 19392 8372 19398 8424
rect 12704 8347 12762 8353
rect 12704 8344 12716 8347
rect 12268 8316 12716 8344
rect 12704 8313 12716 8316
rect 12750 8344 12762 8347
rect 12750 8316 13952 8344
rect 12750 8313 12762 8316
rect 12704 8307 12762 8313
rect 4062 8276 4068 8288
rect 4023 8248 4068 8276
rect 4062 8236 4068 8248
rect 4120 8236 4126 8288
rect 7650 8236 7656 8288
rect 7708 8276 7714 8288
rect 9033 8279 9091 8285
rect 9033 8276 9045 8279
rect 7708 8248 9045 8276
rect 7708 8236 7714 8248
rect 9033 8245 9045 8248
rect 9079 8245 9091 8279
rect 11146 8276 11152 8288
rect 11107 8248 11152 8276
rect 9033 8239 9091 8245
rect 11146 8236 11152 8248
rect 11204 8236 11210 8288
rect 13814 8276 13820 8288
rect 13775 8248 13820 8276
rect 13814 8236 13820 8248
rect 13872 8236 13878 8288
rect 13924 8276 13952 8316
rect 14826 8304 14832 8356
rect 14884 8353 14890 8356
rect 14884 8347 14948 8353
rect 14884 8313 14902 8347
rect 14936 8313 14948 8347
rect 14884 8307 14948 8313
rect 14884 8304 14890 8307
rect 16025 8279 16083 8285
rect 16025 8276 16037 8279
rect 13924 8248 16037 8276
rect 16025 8245 16037 8248
rect 16071 8245 16083 8279
rect 16025 8239 16083 8245
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 2593 8075 2651 8081
rect 2593 8041 2605 8075
rect 2639 8072 2651 8075
rect 2866 8072 2872 8084
rect 2639 8044 2872 8072
rect 2639 8041 2651 8044
rect 2593 8035 2651 8041
rect 2866 8032 2872 8044
rect 2924 8032 2930 8084
rect 3970 8032 3976 8084
rect 4028 8072 4034 8084
rect 7193 8075 7251 8081
rect 4028 8044 5396 8072
rect 4028 8032 4034 8044
rect 5166 7964 5172 8016
rect 5224 8013 5230 8016
rect 5224 8007 5288 8013
rect 5224 7973 5242 8007
rect 5276 7973 5288 8007
rect 5368 8004 5396 8044
rect 7193 8041 7205 8075
rect 7239 8072 7251 8075
rect 7282 8072 7288 8084
rect 7239 8044 7288 8072
rect 7239 8041 7251 8044
rect 7193 8035 7251 8041
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 8938 8032 8944 8084
rect 8996 8072 9002 8084
rect 9677 8075 9735 8081
rect 9677 8072 9689 8075
rect 8996 8044 9689 8072
rect 8996 8032 9002 8044
rect 9677 8041 9689 8044
rect 9723 8041 9735 8075
rect 15286 8072 15292 8084
rect 15247 8044 15292 8072
rect 9677 8035 9735 8041
rect 15286 8032 15292 8044
rect 15344 8032 15350 8084
rect 11146 8004 11152 8016
rect 5368 7976 11152 8004
rect 5224 7967 5288 7973
rect 5224 7964 5230 7967
rect 11146 7964 11152 7976
rect 11204 7964 11210 8016
rect 11517 8007 11575 8013
rect 11517 7973 11529 8007
rect 11563 8004 11575 8007
rect 12342 8004 12348 8016
rect 11563 7976 12348 8004
rect 11563 7973 11575 7976
rect 11517 7967 11575 7973
rect 12342 7964 12348 7976
rect 12400 7964 12406 8016
rect 18049 8007 18107 8013
rect 12728 7976 17816 8004
rect 1854 7896 1860 7948
rect 1912 7936 1918 7948
rect 2685 7939 2743 7945
rect 2685 7936 2697 7939
rect 1912 7908 2697 7936
rect 1912 7896 1918 7908
rect 2685 7905 2697 7908
rect 2731 7905 2743 7939
rect 7558 7936 7564 7948
rect 7519 7908 7564 7936
rect 2685 7899 2743 7905
rect 7558 7896 7564 7908
rect 7616 7896 7622 7948
rect 10042 7936 10048 7948
rect 10003 7908 10048 7936
rect 10042 7896 10048 7908
rect 10100 7896 10106 7948
rect 11241 7939 11299 7945
rect 11241 7905 11253 7939
rect 11287 7936 11299 7939
rect 11882 7936 11888 7948
rect 11287 7908 11888 7936
rect 11287 7905 11299 7908
rect 11241 7899 11299 7905
rect 11882 7896 11888 7908
rect 11940 7896 11946 7948
rect 12728 7936 12756 7976
rect 11992 7908 12756 7936
rect 12796 7939 12854 7945
rect 2774 7828 2780 7880
rect 2832 7868 2838 7880
rect 4982 7868 4988 7880
rect 2832 7840 2877 7868
rect 4943 7840 4988 7868
rect 2832 7828 2838 7840
rect 4982 7828 4988 7840
rect 5040 7828 5046 7880
rect 6086 7828 6092 7880
rect 6144 7868 6150 7880
rect 7653 7871 7711 7877
rect 7653 7868 7665 7871
rect 6144 7840 7665 7868
rect 6144 7828 6150 7840
rect 7653 7837 7665 7840
rect 7699 7837 7711 7871
rect 7653 7831 7711 7837
rect 7742 7828 7748 7880
rect 7800 7868 7806 7880
rect 7800 7840 7845 7868
rect 7800 7828 7806 7840
rect 9858 7828 9864 7880
rect 9916 7868 9922 7880
rect 10137 7871 10195 7877
rect 10137 7868 10149 7871
rect 9916 7840 10149 7868
rect 9916 7828 9922 7840
rect 10137 7837 10149 7840
rect 10183 7837 10195 7871
rect 10137 7831 10195 7837
rect 10321 7871 10379 7877
rect 10321 7837 10333 7871
rect 10367 7868 10379 7871
rect 10686 7868 10692 7880
rect 10367 7840 10692 7868
rect 10367 7837 10379 7840
rect 10321 7831 10379 7837
rect 10686 7828 10692 7840
rect 10744 7828 10750 7880
rect 6365 7803 6423 7809
rect 6365 7769 6377 7803
rect 6411 7800 6423 7803
rect 7760 7800 7788 7828
rect 11992 7800 12020 7908
rect 12796 7905 12808 7939
rect 12842 7936 12854 7939
rect 13814 7936 13820 7948
rect 12842 7908 13820 7936
rect 12842 7905 12854 7908
rect 12796 7899 12854 7905
rect 13814 7896 13820 7908
rect 13872 7896 13878 7948
rect 17788 7945 17816 7976
rect 18049 7973 18061 8007
rect 18095 8004 18107 8007
rect 19334 8004 19340 8016
rect 18095 7976 19340 8004
rect 18095 7973 18107 7976
rect 18049 7967 18107 7973
rect 19334 7964 19340 7976
rect 19392 7964 19398 8016
rect 17773 7939 17831 7945
rect 17773 7905 17785 7939
rect 17819 7905 17831 7939
rect 17773 7899 17831 7905
rect 12066 7828 12072 7880
rect 12124 7868 12130 7880
rect 12529 7871 12587 7877
rect 12529 7868 12541 7871
rect 12124 7840 12541 7868
rect 12124 7828 12130 7840
rect 12529 7837 12541 7840
rect 12575 7837 12587 7871
rect 12529 7831 12587 7837
rect 6411 7772 7788 7800
rect 7852 7772 12020 7800
rect 6411 7769 6423 7772
rect 6365 7763 6423 7769
rect 2225 7735 2283 7741
rect 2225 7701 2237 7735
rect 2271 7732 2283 7735
rect 7852 7732 7880 7772
rect 2271 7704 7880 7732
rect 2271 7701 2283 7704
rect 2225 7695 2283 7701
rect 7926 7692 7932 7744
rect 7984 7732 7990 7744
rect 13909 7735 13967 7741
rect 13909 7732 13921 7735
rect 7984 7704 13921 7732
rect 7984 7692 7990 7704
rect 13909 7701 13921 7704
rect 13955 7701 13967 7735
rect 13909 7695 13967 7701
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 4982 7528 4988 7540
rect 3896 7500 4988 7528
rect 3896 7401 3924 7500
rect 4982 7488 4988 7500
rect 5040 7488 5046 7540
rect 5166 7488 5172 7540
rect 5224 7528 5230 7540
rect 5261 7531 5319 7537
rect 5261 7528 5273 7531
rect 5224 7500 5273 7528
rect 5224 7488 5230 7500
rect 5261 7497 5273 7500
rect 5307 7497 5319 7531
rect 8202 7528 8208 7540
rect 8163 7500 8208 7528
rect 5261 7491 5319 7497
rect 8202 7488 8208 7500
rect 8260 7488 8266 7540
rect 9858 7528 9864 7540
rect 9819 7500 9864 7528
rect 9858 7488 9864 7500
rect 9916 7488 9922 7540
rect 12621 7531 12679 7537
rect 12621 7497 12633 7531
rect 12667 7528 12679 7531
rect 16574 7528 16580 7540
rect 12667 7500 16580 7528
rect 12667 7497 12679 7500
rect 12621 7491 12679 7497
rect 16574 7488 16580 7500
rect 16632 7488 16638 7540
rect 3881 7395 3939 7401
rect 3881 7361 3893 7395
rect 3927 7361 3939 7395
rect 6822 7392 6828 7404
rect 6783 7364 6828 7392
rect 3881 7355 3939 7361
rect 1673 7327 1731 7333
rect 1673 7293 1685 7327
rect 1719 7324 1731 7327
rect 2774 7324 2780 7336
rect 1719 7296 2780 7324
rect 1719 7293 1731 7296
rect 1673 7287 1731 7293
rect 2774 7284 2780 7296
rect 2832 7324 2838 7336
rect 3896 7324 3924 7355
rect 6822 7352 6828 7364
rect 6880 7352 6886 7404
rect 9490 7352 9496 7404
rect 9548 7392 9554 7404
rect 10413 7395 10471 7401
rect 10413 7392 10425 7395
rect 9548 7364 10425 7392
rect 9548 7352 9554 7364
rect 10413 7361 10425 7364
rect 10459 7361 10471 7395
rect 10413 7355 10471 7361
rect 11698 7352 11704 7404
rect 11756 7392 11762 7404
rect 13081 7395 13139 7401
rect 13081 7392 13093 7395
rect 11756 7364 13093 7392
rect 11756 7352 11762 7364
rect 13081 7361 13093 7364
rect 13127 7361 13139 7395
rect 13081 7355 13139 7361
rect 13265 7395 13323 7401
rect 13265 7361 13277 7395
rect 13311 7392 13323 7395
rect 13814 7392 13820 7404
rect 13311 7364 13820 7392
rect 13311 7361 13323 7364
rect 13265 7355 13323 7361
rect 13814 7352 13820 7364
rect 13872 7352 13878 7404
rect 2832 7296 3924 7324
rect 4148 7327 4206 7333
rect 2832 7284 2838 7296
rect 4148 7293 4160 7327
rect 4194 7324 4206 7327
rect 7926 7324 7932 7336
rect 4194 7296 7932 7324
rect 4194 7293 4206 7296
rect 4148 7287 4206 7293
rect 4356 7268 4384 7296
rect 7926 7284 7932 7296
rect 7984 7284 7990 7336
rect 10226 7324 10232 7336
rect 10139 7296 10232 7324
rect 10226 7284 10232 7296
rect 10284 7324 10290 7336
rect 10778 7324 10784 7336
rect 10284 7296 10784 7324
rect 10284 7284 10290 7296
rect 10778 7284 10784 7296
rect 10836 7284 10842 7336
rect 12989 7327 13047 7333
rect 12989 7293 13001 7327
rect 13035 7324 13047 7327
rect 14182 7324 14188 7336
rect 13035 7296 14188 7324
rect 13035 7293 13047 7296
rect 12989 7287 13047 7293
rect 14182 7284 14188 7296
rect 14240 7284 14246 7336
rect 1940 7259 1998 7265
rect 1940 7225 1952 7259
rect 1986 7256 1998 7259
rect 2406 7256 2412 7268
rect 1986 7228 2412 7256
rect 1986 7225 1998 7228
rect 1940 7219 1998 7225
rect 2406 7216 2412 7228
rect 2464 7216 2470 7268
rect 4338 7216 4344 7268
rect 4396 7216 4402 7268
rect 7092 7259 7150 7265
rect 7092 7225 7104 7259
rect 7138 7256 7150 7259
rect 7742 7256 7748 7268
rect 7138 7228 7748 7256
rect 7138 7225 7150 7228
rect 7092 7219 7150 7225
rect 7742 7216 7748 7228
rect 7800 7216 7806 7268
rect 2682 7148 2688 7200
rect 2740 7188 2746 7200
rect 3053 7191 3111 7197
rect 3053 7188 3065 7191
rect 2740 7160 3065 7188
rect 2740 7148 2746 7160
rect 3053 7157 3065 7160
rect 3099 7157 3111 7191
rect 3053 7151 3111 7157
rect 10318 7148 10324 7200
rect 10376 7188 10382 7200
rect 10376 7160 10421 7188
rect 10376 7148 10382 7160
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 1854 6984 1860 6996
rect 1815 6956 1860 6984
rect 1854 6944 1860 6956
rect 1912 6944 1918 6996
rect 3878 6944 3884 6996
rect 3936 6984 3942 6996
rect 4893 6987 4951 6993
rect 4893 6984 4905 6987
rect 3936 6956 4905 6984
rect 3936 6944 3942 6956
rect 4893 6953 4905 6956
rect 4939 6984 4951 6987
rect 9030 6984 9036 6996
rect 4939 6956 9036 6984
rect 4939 6953 4951 6956
rect 4893 6947 4951 6953
rect 9030 6944 9036 6956
rect 9088 6944 9094 6996
rect 11885 6987 11943 6993
rect 11885 6953 11897 6987
rect 11931 6984 11943 6987
rect 12250 6984 12256 6996
rect 11931 6956 12256 6984
rect 11931 6953 11943 6956
rect 11885 6947 11943 6953
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 2222 6916 2228 6928
rect 2183 6888 2228 6916
rect 2222 6876 2228 6888
rect 2280 6876 2286 6928
rect 7184 6919 7242 6925
rect 7184 6885 7196 6919
rect 7230 6916 7242 6919
rect 8202 6916 8208 6928
rect 7230 6888 8208 6916
rect 7230 6885 7242 6888
rect 7184 6879 7242 6885
rect 8202 6876 8208 6888
rect 8260 6876 8266 6928
rect 10686 6876 10692 6928
rect 10744 6925 10750 6928
rect 10744 6919 10808 6925
rect 10744 6885 10762 6919
rect 10796 6885 10808 6919
rect 10744 6879 10808 6885
rect 10744 6876 10750 6879
rect 2314 6848 2320 6860
rect 2275 6820 2320 6848
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 18969 6851 19027 6857
rect 18969 6848 18981 6851
rect 5276 6820 18981 6848
rect 2406 6780 2412 6792
rect 2367 6752 2412 6780
rect 2406 6740 2412 6752
rect 2464 6740 2470 6792
rect 2498 6740 2504 6792
rect 2556 6780 2562 6792
rect 4985 6783 5043 6789
rect 4985 6780 4997 6783
rect 2556 6752 4997 6780
rect 2556 6740 2562 6752
rect 4985 6749 4997 6752
rect 5031 6749 5043 6783
rect 5166 6780 5172 6792
rect 5127 6752 5172 6780
rect 4985 6743 5043 6749
rect 5166 6740 5172 6752
rect 5224 6740 5230 6792
rect 4062 6672 4068 6724
rect 4120 6712 4126 6724
rect 5276 6712 5304 6820
rect 18969 6817 18981 6820
rect 19015 6817 19027 6851
rect 18969 6811 19027 6817
rect 6822 6740 6828 6792
rect 6880 6780 6886 6792
rect 6917 6783 6975 6789
rect 6917 6780 6929 6783
rect 6880 6752 6929 6780
rect 6880 6740 6886 6752
rect 6917 6749 6929 6752
rect 6963 6749 6975 6783
rect 10502 6780 10508 6792
rect 10463 6752 10508 6780
rect 6917 6743 6975 6749
rect 10502 6740 10508 6752
rect 10560 6740 10566 6792
rect 4120 6684 5304 6712
rect 19153 6715 19211 6721
rect 4120 6672 4126 6684
rect 19153 6681 19165 6715
rect 19199 6712 19211 6715
rect 19886 6712 19892 6724
rect 19199 6684 19892 6712
rect 19199 6681 19211 6684
rect 19153 6675 19211 6681
rect 19886 6672 19892 6684
rect 19944 6672 19950 6724
rect 4525 6647 4583 6653
rect 4525 6613 4537 6647
rect 4571 6644 4583 6647
rect 5074 6644 5080 6656
rect 4571 6616 5080 6644
rect 4571 6613 4583 6616
rect 4525 6607 4583 6613
rect 5074 6604 5080 6616
rect 5132 6604 5138 6656
rect 8294 6644 8300 6656
rect 8255 6616 8300 6644
rect 8294 6604 8300 6616
rect 8352 6604 8358 6656
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 2406 6400 2412 6452
rect 2464 6440 2470 6452
rect 8294 6440 8300 6452
rect 2464 6412 8300 6440
rect 2464 6400 2470 6412
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 10502 6440 10508 6452
rect 9232 6412 10508 6440
rect 5074 6304 5080 6316
rect 5035 6276 5080 6304
rect 5074 6264 5080 6276
rect 5132 6264 5138 6316
rect 5261 6307 5319 6313
rect 5261 6273 5273 6307
rect 5307 6304 5319 6307
rect 6546 6304 6552 6316
rect 5307 6276 6552 6304
rect 5307 6273 5319 6276
rect 5261 6267 5319 6273
rect 6546 6264 6552 6276
rect 6604 6304 6610 6316
rect 9232 6313 9260 6412
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 10597 6443 10655 6449
rect 10597 6409 10609 6443
rect 10643 6440 10655 6443
rect 10686 6440 10692 6452
rect 10643 6412 10692 6440
rect 10643 6409 10655 6412
rect 10597 6403 10655 6409
rect 10686 6400 10692 6412
rect 10744 6400 10750 6452
rect 19702 6440 19708 6452
rect 12452 6412 19564 6440
rect 19663 6412 19708 6440
rect 12342 6332 12348 6384
rect 12400 6372 12406 6384
rect 12452 6372 12480 6412
rect 12400 6344 12480 6372
rect 12400 6332 12406 6344
rect 9217 6307 9275 6313
rect 6604 6276 6960 6304
rect 6604 6264 6610 6276
rect 2682 6245 2688 6248
rect 2409 6239 2467 6245
rect 2409 6205 2421 6239
rect 2455 6205 2467 6239
rect 2409 6199 2467 6205
rect 2676 6199 2688 6245
rect 2740 6236 2746 6248
rect 6822 6236 6828 6248
rect 2740 6208 2776 6236
rect 6783 6208 6828 6236
rect 2424 6168 2452 6199
rect 2682 6196 2688 6199
rect 2740 6196 2746 6208
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 6932 6236 6960 6276
rect 9217 6273 9229 6307
rect 9263 6273 9275 6307
rect 9217 6267 9275 6273
rect 9490 6245 9496 6248
rect 7081 6239 7139 6245
rect 7081 6236 7093 6239
rect 6932 6208 7093 6236
rect 7081 6205 7093 6208
rect 7127 6205 7139 6239
rect 9484 6236 9496 6245
rect 9451 6208 9496 6236
rect 7081 6199 7139 6205
rect 9484 6199 9496 6208
rect 9490 6196 9496 6199
rect 9548 6196 9554 6248
rect 19536 6245 19564 6412
rect 19702 6400 19708 6412
rect 19760 6400 19766 6452
rect 19521 6239 19579 6245
rect 19521 6205 19533 6239
rect 19567 6205 19579 6239
rect 19521 6199 19579 6205
rect 2774 6168 2780 6180
rect 2424 6140 2780 6168
rect 2774 6128 2780 6140
rect 2832 6128 2838 6180
rect 3970 6128 3976 6180
rect 4028 6168 4034 6180
rect 12342 6168 12348 6180
rect 4028 6140 12348 6168
rect 4028 6128 4034 6140
rect 12342 6128 12348 6140
rect 12400 6128 12406 6180
rect 3786 6100 3792 6112
rect 3747 6072 3792 6100
rect 3786 6060 3792 6072
rect 3844 6060 3850 6112
rect 4338 6060 4344 6112
rect 4396 6100 4402 6112
rect 4617 6103 4675 6109
rect 4617 6100 4629 6103
rect 4396 6072 4629 6100
rect 4396 6060 4402 6072
rect 4617 6069 4629 6072
rect 4663 6069 4675 6103
rect 4982 6100 4988 6112
rect 4943 6072 4988 6100
rect 4617 6063 4675 6069
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 8205 6103 8263 6109
rect 8205 6069 8217 6103
rect 8251 6100 8263 6103
rect 8294 6100 8300 6112
rect 8251 6072 8300 6100
rect 8251 6069 8263 6072
rect 8205 6063 8263 6069
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 2409 5899 2467 5905
rect 2409 5865 2421 5899
rect 2455 5896 2467 5899
rect 2498 5896 2504 5908
rect 2455 5868 2504 5896
rect 2455 5865 2467 5868
rect 2409 5859 2467 5865
rect 2498 5856 2504 5868
rect 2556 5856 2562 5908
rect 6546 5896 6552 5908
rect 6507 5868 6552 5896
rect 6546 5856 6552 5868
rect 6604 5856 6610 5908
rect 7377 5899 7435 5905
rect 7377 5865 7389 5899
rect 7423 5896 7435 5899
rect 7558 5896 7564 5908
rect 7423 5868 7564 5896
rect 7423 5865 7435 5868
rect 7377 5859 7435 5865
rect 7558 5856 7564 5868
rect 7616 5856 7622 5908
rect 10318 5856 10324 5908
rect 10376 5896 10382 5908
rect 10689 5899 10747 5905
rect 10689 5896 10701 5899
rect 10376 5868 10701 5896
rect 10376 5856 10382 5868
rect 10689 5865 10701 5868
rect 10735 5865 10747 5899
rect 10689 5859 10747 5865
rect 11149 5899 11207 5905
rect 11149 5865 11161 5899
rect 11195 5896 11207 5899
rect 13354 5896 13360 5908
rect 11195 5868 13360 5896
rect 11195 5865 11207 5868
rect 11149 5859 11207 5865
rect 2317 5831 2375 5837
rect 2317 5797 2329 5831
rect 2363 5828 2375 5831
rect 2869 5831 2927 5837
rect 2869 5828 2881 5831
rect 2363 5800 2881 5828
rect 2363 5797 2375 5800
rect 2317 5791 2375 5797
rect 2869 5797 2881 5800
rect 2915 5828 2927 5831
rect 3142 5828 3148 5840
rect 2915 5800 3148 5828
rect 2915 5797 2927 5800
rect 2869 5791 2927 5797
rect 3142 5788 3148 5800
rect 3200 5788 3206 5840
rect 5166 5788 5172 5840
rect 5224 5828 5230 5840
rect 5414 5831 5472 5837
rect 5414 5828 5426 5831
rect 5224 5800 5426 5828
rect 5224 5788 5230 5800
rect 5414 5797 5426 5800
rect 5460 5797 5472 5831
rect 5414 5791 5472 5797
rect 10597 5831 10655 5837
rect 10597 5797 10609 5831
rect 10643 5828 10655 5831
rect 11164 5828 11192 5859
rect 13354 5856 13360 5868
rect 13412 5856 13418 5908
rect 19889 5899 19947 5905
rect 19889 5865 19901 5899
rect 19935 5896 19947 5899
rect 20990 5896 20996 5908
rect 19935 5868 20996 5896
rect 19935 5865 19947 5868
rect 19889 5859 19947 5865
rect 20990 5856 20996 5868
rect 21048 5856 21054 5908
rect 10643 5800 11192 5828
rect 10643 5797 10655 5800
rect 10597 5791 10655 5797
rect 11238 5788 11244 5840
rect 11296 5788 11302 5840
rect 12452 5800 19748 5828
rect 2682 5720 2688 5772
rect 2740 5760 2746 5772
rect 2777 5763 2835 5769
rect 2777 5760 2789 5763
rect 2740 5732 2789 5760
rect 2740 5720 2746 5732
rect 2777 5729 2789 5732
rect 2823 5760 2835 5763
rect 7466 5760 7472 5772
rect 2823 5732 7472 5760
rect 2823 5729 2835 5732
rect 2777 5723 2835 5729
rect 7466 5720 7472 5732
rect 7524 5720 7530 5772
rect 8294 5720 8300 5772
rect 8352 5760 8358 5772
rect 11054 5760 11060 5772
rect 8352 5732 9812 5760
rect 10967 5732 11060 5760
rect 8352 5720 8358 5732
rect 3053 5695 3111 5701
rect 3053 5661 3065 5695
rect 3099 5692 3111 5695
rect 3786 5692 3792 5704
rect 3099 5664 3792 5692
rect 3099 5661 3111 5664
rect 3053 5655 3111 5661
rect 3786 5652 3792 5664
rect 3844 5652 3850 5704
rect 5169 5695 5227 5701
rect 5169 5661 5181 5695
rect 5215 5661 5227 5695
rect 9674 5692 9680 5704
rect 9635 5664 9680 5692
rect 5169 5655 5227 5661
rect 2774 5584 2780 5636
rect 2832 5624 2838 5636
rect 3694 5624 3700 5636
rect 2832 5596 3700 5624
rect 2832 5584 2838 5596
rect 3694 5584 3700 5596
rect 3752 5624 3758 5636
rect 5184 5624 5212 5655
rect 9674 5652 9680 5664
rect 9732 5652 9738 5704
rect 9784 5692 9812 5732
rect 11054 5720 11060 5732
rect 11112 5760 11118 5772
rect 11256 5760 11284 5788
rect 11112 5732 11284 5760
rect 11112 5720 11118 5732
rect 12342 5720 12348 5772
rect 12400 5760 12406 5772
rect 12452 5760 12480 5800
rect 19720 5769 19748 5800
rect 12400 5732 12480 5760
rect 19705 5763 19763 5769
rect 12400 5720 12406 5732
rect 19705 5729 19717 5763
rect 19751 5729 19763 5763
rect 19705 5723 19763 5729
rect 11241 5695 11299 5701
rect 11241 5692 11253 5695
rect 9784 5664 11253 5692
rect 11241 5661 11253 5664
rect 11287 5661 11299 5695
rect 11241 5655 11299 5661
rect 3752 5596 5212 5624
rect 3752 5584 3758 5596
rect 4062 5516 4068 5568
rect 4120 5556 4126 5568
rect 12342 5556 12348 5568
rect 4120 5528 12348 5556
rect 4120 5516 4126 5528
rect 12342 5516 12348 5528
rect 12400 5516 12406 5568
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 4338 5352 4344 5364
rect 2516 5324 4344 5352
rect 2041 5151 2099 5157
rect 2041 5117 2053 5151
rect 2087 5148 2099 5151
rect 2516 5148 2544 5324
rect 4338 5312 4344 5324
rect 4396 5312 4402 5364
rect 5077 5355 5135 5361
rect 5077 5321 5089 5355
rect 5123 5352 5135 5355
rect 5166 5352 5172 5364
rect 5123 5324 5172 5352
rect 5123 5321 5135 5324
rect 5077 5315 5135 5321
rect 5166 5312 5172 5324
rect 5224 5312 5230 5364
rect 9401 5355 9459 5361
rect 5276 5324 9076 5352
rect 3694 5216 3700 5228
rect 3655 5188 3700 5216
rect 3694 5176 3700 5188
rect 3752 5176 3758 5228
rect 2087 5120 2544 5148
rect 2087 5117 2099 5120
rect 2041 5111 2099 5117
rect 3786 5108 3792 5160
rect 3844 5148 3850 5160
rect 3953 5151 4011 5157
rect 3953 5148 3965 5151
rect 3844 5120 3965 5148
rect 3844 5108 3850 5120
rect 3953 5117 3965 5120
rect 3999 5117 4011 5151
rect 3953 5111 4011 5117
rect 1762 5040 1768 5092
rect 1820 5080 1826 5092
rect 2317 5083 2375 5089
rect 2317 5080 2329 5083
rect 1820 5052 2329 5080
rect 1820 5040 1826 5052
rect 2317 5049 2329 5052
rect 2363 5049 2375 5083
rect 2317 5043 2375 5049
rect 3234 5040 3240 5092
rect 3292 5080 3298 5092
rect 5276 5080 5304 5324
rect 5534 5176 5540 5228
rect 5592 5216 5598 5228
rect 6638 5216 6644 5228
rect 5592 5188 6644 5216
rect 5592 5176 5598 5188
rect 6638 5176 6644 5188
rect 6696 5176 6702 5228
rect 6822 5176 6828 5228
rect 6880 5216 6886 5228
rect 8021 5219 8079 5225
rect 8021 5216 8033 5219
rect 6880 5188 8033 5216
rect 6880 5176 6886 5188
rect 8021 5185 8033 5188
rect 8067 5185 8079 5219
rect 8021 5179 8079 5185
rect 6656 5148 6684 5176
rect 8294 5157 8300 5160
rect 8288 5148 8300 5157
rect 6656 5120 7696 5148
rect 8255 5120 8300 5148
rect 3292 5052 5304 5080
rect 3292 5040 3298 5052
rect 5258 4972 5264 5024
rect 5316 5012 5322 5024
rect 6825 5015 6883 5021
rect 6825 5012 6837 5015
rect 5316 4984 6837 5012
rect 5316 4972 5322 4984
rect 6825 4981 6837 4984
rect 6871 4981 6883 5015
rect 7668 5012 7696 5120
rect 8288 5111 8300 5120
rect 8294 5108 8300 5111
rect 8352 5108 8358 5160
rect 9048 5080 9076 5324
rect 9401 5321 9413 5355
rect 9447 5352 9459 5355
rect 9490 5352 9496 5364
rect 9447 5324 9496 5352
rect 9447 5321 9459 5324
rect 9401 5315 9459 5321
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 10042 5312 10048 5364
rect 10100 5352 10106 5364
rect 10229 5355 10287 5361
rect 10229 5352 10241 5355
rect 10100 5324 10241 5352
rect 10100 5312 10106 5324
rect 10229 5321 10241 5324
rect 10275 5321 10287 5355
rect 19610 5352 19616 5364
rect 19571 5324 19616 5352
rect 10229 5315 10287 5321
rect 19610 5312 19616 5324
rect 19668 5312 19674 5364
rect 20717 5355 20775 5361
rect 20717 5321 20729 5355
rect 20763 5352 20775 5355
rect 20898 5352 20904 5364
rect 20763 5324 20904 5352
rect 20763 5321 20775 5324
rect 20717 5315 20775 5321
rect 20898 5312 20904 5324
rect 20956 5312 20962 5364
rect 9508 5216 9536 5312
rect 10781 5219 10839 5225
rect 10781 5216 10793 5219
rect 9508 5188 10793 5216
rect 10781 5185 10793 5188
rect 10827 5185 10839 5219
rect 10781 5179 10839 5185
rect 9674 5108 9680 5160
rect 9732 5148 9738 5160
rect 10597 5151 10655 5157
rect 10597 5148 10609 5151
rect 9732 5120 10609 5148
rect 9732 5108 9738 5120
rect 10597 5117 10609 5120
rect 10643 5117 10655 5151
rect 10597 5111 10655 5117
rect 19429 5151 19487 5157
rect 19429 5117 19441 5151
rect 19475 5117 19487 5151
rect 20530 5148 20536 5160
rect 20491 5120 20536 5148
rect 19429 5111 19487 5117
rect 19444 5080 19472 5111
rect 20530 5108 20536 5120
rect 20588 5108 20594 5160
rect 9048 5052 19472 5080
rect 10689 5015 10747 5021
rect 10689 5012 10701 5015
rect 7668 4984 10701 5012
rect 6825 4975 6883 4981
rect 10689 4981 10701 4984
rect 10735 4981 10747 5015
rect 10689 4975 10747 4981
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 1578 4768 1584 4820
rect 1636 4808 1642 4820
rect 1949 4811 2007 4817
rect 1949 4808 1961 4811
rect 1636 4780 1961 4808
rect 1636 4768 1642 4780
rect 1949 4777 1961 4780
rect 1995 4777 2007 4811
rect 1949 4771 2007 4777
rect 4893 4811 4951 4817
rect 4893 4777 4905 4811
rect 4939 4808 4951 4811
rect 4982 4808 4988 4820
rect 4939 4780 4988 4808
rect 4939 4777 4951 4780
rect 4893 4771 4951 4777
rect 4982 4768 4988 4780
rect 5040 4768 5046 4820
rect 5258 4808 5264 4820
rect 5219 4780 5264 4808
rect 5258 4768 5264 4780
rect 5316 4768 5322 4820
rect 12434 4768 12440 4820
rect 12492 4808 12498 4820
rect 20530 4808 20536 4820
rect 12492 4780 20536 4808
rect 12492 4768 12498 4780
rect 20530 4768 20536 4780
rect 20588 4768 20594 4820
rect 4062 4700 4068 4752
rect 4120 4740 4126 4752
rect 12342 4740 12348 4752
rect 4120 4712 12348 4740
rect 4120 4700 4126 4712
rect 12342 4700 12348 4712
rect 12400 4700 12406 4752
rect 1762 4672 1768 4684
rect 1723 4644 1768 4672
rect 1762 4632 1768 4644
rect 1820 4632 1826 4684
rect 5166 4632 5172 4684
rect 5224 4672 5230 4684
rect 5224 4644 5488 4672
rect 5224 4632 5230 4644
rect 4154 4564 4160 4616
rect 4212 4604 4218 4616
rect 5350 4604 5356 4616
rect 4212 4576 5356 4604
rect 4212 4564 4218 4576
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 5460 4613 5488 4644
rect 5445 4607 5503 4613
rect 5445 4573 5457 4607
rect 5491 4573 5503 4607
rect 5445 4567 5503 4573
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 3510 4088 3516 4140
rect 3568 4128 3574 4140
rect 7650 4128 7656 4140
rect 3568 4100 7656 4128
rect 3568 4088 3574 4100
rect 7650 4088 7656 4100
rect 7708 4088 7714 4140
rect 4062 4020 4068 4072
rect 4120 4060 4126 4072
rect 20533 4063 20591 4069
rect 20533 4060 20545 4063
rect 4120 4032 20545 4060
rect 4120 4020 4126 4032
rect 20533 4029 20545 4032
rect 20579 4029 20591 4063
rect 20533 4023 20591 4029
rect 5718 3952 5724 4004
rect 5776 3992 5782 4004
rect 6730 3992 6736 4004
rect 5776 3964 6736 3992
rect 5776 3952 5782 3964
rect 6730 3952 6736 3964
rect 6788 3952 6794 4004
rect 20717 3927 20775 3933
rect 20717 3893 20729 3927
rect 20763 3924 20775 3927
rect 20806 3924 20812 3936
rect 20763 3896 20812 3924
rect 20763 3893 20775 3896
rect 20717 3887 20775 3893
rect 20806 3884 20812 3896
rect 20864 3884 20870 3936
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 4062 2592 4068 2644
rect 4120 2632 4126 2644
rect 5534 2632 5540 2644
rect 4120 2604 5540 2632
rect 4120 2592 4126 2604
rect 5534 2592 5540 2604
rect 5592 2592 5598 2644
rect 3050 2456 3056 2508
rect 3108 2496 3114 2508
rect 10226 2496 10232 2508
rect 3108 2468 10232 2496
rect 3108 2456 3114 2468
rect 10226 2456 10232 2468
rect 10284 2456 10290 2508
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 3418 1300 3424 1352
rect 3476 1340 3482 1352
rect 11054 1340 11060 1352
rect 3476 1312 11060 1340
rect 3476 1300 3482 1312
rect 11054 1300 11060 1312
rect 11112 1300 11118 1352
<< via1 >>
rect 3516 21088 3568 21140
rect 6092 21088 6144 21140
rect 3792 20952 3844 21004
rect 11244 20952 11296 21004
rect 4068 20748 4120 20800
rect 15476 20748 15528 20800
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 3976 20544 4028 20596
rect 8760 20544 8812 20596
rect 8944 20544 8996 20596
rect 11796 20544 11848 20596
rect 13268 20544 13320 20596
rect 4068 20476 4120 20528
rect 5448 20476 5500 20528
rect 5908 20451 5960 20460
rect 5908 20417 5917 20451
rect 5917 20417 5951 20451
rect 5951 20417 5960 20451
rect 5908 20408 5960 20417
rect 6184 20476 6236 20528
rect 8116 20476 8168 20528
rect 12716 20476 12768 20528
rect 14740 20544 14792 20596
rect 18604 20544 18656 20596
rect 2136 20383 2188 20392
rect 2136 20349 2145 20383
rect 2145 20349 2179 20383
rect 2179 20349 2188 20383
rect 2136 20340 2188 20349
rect 6184 20340 6236 20392
rect 6828 20340 6880 20392
rect 10048 20340 10100 20392
rect 10508 20408 10560 20460
rect 12072 20408 12124 20460
rect 12164 20408 12216 20460
rect 12716 20340 12768 20392
rect 16948 20340 17000 20392
rect 18144 20340 18196 20392
rect 8668 20315 8720 20324
rect 8668 20281 8677 20315
rect 8677 20281 8711 20315
rect 8711 20281 8720 20315
rect 8668 20272 8720 20281
rect 8760 20272 8812 20324
rect 3240 20204 3292 20256
rect 5632 20247 5684 20256
rect 5632 20213 5641 20247
rect 5641 20213 5675 20247
rect 5675 20213 5684 20247
rect 5632 20204 5684 20213
rect 5724 20247 5776 20256
rect 5724 20213 5733 20247
rect 5733 20213 5767 20247
rect 5767 20213 5776 20247
rect 7104 20247 7156 20256
rect 5724 20204 5776 20213
rect 7104 20213 7113 20247
rect 7113 20213 7147 20247
rect 7147 20213 7156 20247
rect 7104 20204 7156 20213
rect 10416 20204 10468 20256
rect 10600 20247 10652 20256
rect 10600 20213 10609 20247
rect 10609 20213 10643 20247
rect 10643 20213 10652 20247
rect 10600 20204 10652 20213
rect 12808 20247 12860 20256
rect 12808 20213 12817 20247
rect 12817 20213 12851 20247
rect 12851 20213 12860 20247
rect 12808 20204 12860 20213
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 4252 20000 4304 20052
rect 7104 20000 7156 20052
rect 7196 20000 7248 20052
rect 5448 19932 5500 19984
rect 5632 19932 5684 19984
rect 9496 19932 9548 19984
rect 10600 19932 10652 19984
rect 12072 19932 12124 19984
rect 15200 20000 15252 20052
rect 17960 20000 18012 20052
rect 19156 19932 19208 19984
rect 1400 19907 1452 19916
rect 1400 19873 1409 19907
rect 1409 19873 1443 19907
rect 1443 19873 1452 19907
rect 1400 19864 1452 19873
rect 2964 19864 3016 19916
rect 3608 19864 3660 19916
rect 5908 19864 5960 19916
rect 6828 19864 6880 19916
rect 8944 19864 8996 19916
rect 9128 19864 9180 19916
rect 12900 19864 12952 19916
rect 15292 19907 15344 19916
rect 15292 19873 15301 19907
rect 15301 19873 15335 19907
rect 15335 19873 15344 19907
rect 15292 19864 15344 19873
rect 16396 19907 16448 19916
rect 16396 19873 16405 19907
rect 16405 19873 16439 19907
rect 16439 19873 16448 19907
rect 16396 19864 16448 19873
rect 17408 19864 17460 19916
rect 18604 19907 18656 19916
rect 18604 19873 18613 19907
rect 18613 19873 18647 19907
rect 18647 19873 18656 19907
rect 18604 19864 18656 19873
rect 4988 19796 5040 19848
rect 8208 19839 8260 19848
rect 8208 19805 8217 19839
rect 8217 19805 8251 19839
rect 8251 19805 8260 19839
rect 8208 19796 8260 19805
rect 9680 19839 9732 19848
rect 9680 19805 9689 19839
rect 9689 19805 9723 19839
rect 9723 19805 9732 19839
rect 9680 19796 9732 19805
rect 11888 19839 11940 19848
rect 11888 19805 11897 19839
rect 11897 19805 11931 19839
rect 11931 19805 11940 19839
rect 11888 19796 11940 19805
rect 19708 19839 19760 19848
rect 19708 19805 19717 19839
rect 19717 19805 19751 19839
rect 19751 19805 19760 19839
rect 19708 19796 19760 19805
rect 6368 19728 6420 19780
rect 1584 19703 1636 19712
rect 1584 19669 1593 19703
rect 1593 19669 1627 19703
rect 1627 19669 1636 19703
rect 1584 19660 1636 19669
rect 3516 19660 3568 19712
rect 4344 19660 4396 19712
rect 7656 19703 7708 19712
rect 7656 19669 7665 19703
rect 7665 19669 7699 19703
rect 7699 19669 7708 19703
rect 7656 19660 7708 19669
rect 7840 19728 7892 19780
rect 9220 19728 9272 19780
rect 9496 19728 9548 19780
rect 10692 19728 10744 19780
rect 12992 19728 13044 19780
rect 15476 19771 15528 19780
rect 15476 19737 15485 19771
rect 15485 19737 15519 19771
rect 15519 19737 15528 19771
rect 15476 19728 15528 19737
rect 16672 19660 16724 19712
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 3792 19456 3844 19508
rect 3976 19456 4028 19508
rect 9128 19499 9180 19508
rect 9128 19465 9137 19499
rect 9137 19465 9171 19499
rect 9171 19465 9180 19499
rect 9128 19456 9180 19465
rect 10048 19499 10100 19508
rect 10048 19465 10057 19499
rect 10057 19465 10091 19499
rect 10091 19465 10100 19499
rect 10048 19456 10100 19465
rect 5908 19320 5960 19372
rect 6368 19320 6420 19372
rect 9956 19388 10008 19440
rect 12992 19388 13044 19440
rect 2872 19295 2924 19304
rect 1768 19116 1820 19168
rect 2872 19261 2881 19295
rect 2881 19261 2915 19295
rect 2915 19261 2924 19295
rect 2872 19252 2924 19261
rect 4344 19252 4396 19304
rect 2504 19184 2556 19236
rect 3700 19184 3752 19236
rect 5540 19252 5592 19304
rect 6736 19252 6788 19304
rect 7748 19295 7800 19304
rect 7748 19261 7757 19295
rect 7757 19261 7791 19295
rect 7791 19261 7800 19295
rect 7748 19252 7800 19261
rect 10416 19320 10468 19372
rect 10692 19363 10744 19372
rect 10692 19329 10701 19363
rect 10701 19329 10735 19363
rect 10735 19329 10744 19363
rect 10692 19320 10744 19329
rect 11888 19320 11940 19372
rect 19156 19363 19208 19372
rect 19156 19329 19165 19363
rect 19165 19329 19199 19363
rect 19199 19329 19208 19363
rect 19156 19320 19208 19329
rect 12348 19252 12400 19304
rect 12716 19252 12768 19304
rect 13176 19295 13228 19304
rect 13176 19261 13185 19295
rect 13185 19261 13219 19295
rect 13219 19261 13228 19295
rect 13176 19252 13228 19261
rect 4160 19116 4212 19168
rect 5724 19184 5776 19236
rect 7840 19184 7892 19236
rect 8208 19184 8260 19236
rect 6000 19116 6052 19168
rect 8668 19116 8720 19168
rect 12256 19184 12308 19236
rect 15292 19252 15344 19304
rect 15384 19295 15436 19304
rect 15384 19261 15393 19295
rect 15393 19261 15427 19295
rect 15427 19261 15436 19295
rect 15384 19252 15436 19261
rect 17868 19252 17920 19304
rect 13452 19227 13504 19236
rect 13452 19193 13486 19227
rect 13486 19193 13504 19227
rect 13452 19184 13504 19193
rect 14188 19116 14240 19168
rect 14556 19159 14608 19168
rect 14556 19125 14565 19159
rect 14565 19125 14599 19159
rect 14599 19125 14608 19159
rect 14556 19116 14608 19125
rect 14648 19116 14700 19168
rect 17040 19116 17092 19168
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 6276 18912 6328 18964
rect 6828 18955 6880 18964
rect 6828 18921 6837 18955
rect 6837 18921 6871 18955
rect 6871 18921 6880 18955
rect 6828 18912 6880 18921
rect 7656 18912 7708 18964
rect 8300 18912 8352 18964
rect 12900 18912 12952 18964
rect 14372 18912 14424 18964
rect 16580 18955 16632 18964
rect 16580 18921 16589 18955
rect 16589 18921 16623 18955
rect 16623 18921 16632 18955
rect 16580 18912 16632 18921
rect 17500 18912 17552 18964
rect 4528 18844 4580 18896
rect 5724 18887 5776 18896
rect 5724 18853 5758 18887
rect 5758 18853 5776 18887
rect 5724 18844 5776 18853
rect 13728 18844 13780 18896
rect 16672 18844 16724 18896
rect 2780 18819 2832 18828
rect 2780 18785 2789 18819
rect 2789 18785 2823 18819
rect 2823 18785 2832 18819
rect 4068 18819 4120 18828
rect 2780 18776 2832 18785
rect 4068 18785 4077 18819
rect 4077 18785 4111 18819
rect 4111 18785 4120 18819
rect 4068 18776 4120 18785
rect 6828 18776 6880 18828
rect 7748 18776 7800 18828
rect 4344 18708 4396 18760
rect 4988 18708 5040 18760
rect 3056 18572 3108 18624
rect 6920 18640 6972 18692
rect 7196 18572 7248 18624
rect 10784 18776 10836 18828
rect 12072 18776 12124 18828
rect 14648 18776 14700 18828
rect 14740 18776 14792 18828
rect 15568 18776 15620 18828
rect 17500 18819 17552 18828
rect 17500 18785 17509 18819
rect 17509 18785 17543 18819
rect 17543 18785 17552 18819
rect 17500 18776 17552 18785
rect 9128 18708 9180 18760
rect 9680 18708 9732 18760
rect 9956 18708 10008 18760
rect 12532 18708 12584 18760
rect 14556 18708 14608 18760
rect 19708 18640 19760 18692
rect 12072 18615 12124 18624
rect 12072 18581 12081 18615
rect 12081 18581 12115 18615
rect 12115 18581 12124 18615
rect 12072 18572 12124 18581
rect 12440 18572 12492 18624
rect 13084 18572 13136 18624
rect 22652 18572 22704 18624
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 2964 18411 3016 18420
rect 2964 18377 2973 18411
rect 2973 18377 3007 18411
rect 3007 18377 3016 18411
rect 2964 18368 3016 18377
rect 3148 18368 3200 18420
rect 4068 18368 4120 18420
rect 4896 18368 4948 18420
rect 12256 18368 12308 18420
rect 12532 18411 12584 18420
rect 12532 18377 12541 18411
rect 12541 18377 12575 18411
rect 12575 18377 12584 18411
rect 12532 18368 12584 18377
rect 8576 18300 8628 18352
rect 1952 18232 2004 18284
rect 2964 18232 3016 18284
rect 3056 18232 3108 18284
rect 4160 18232 4212 18284
rect 5448 18232 5500 18284
rect 7472 18275 7524 18284
rect 4896 18164 4948 18216
rect 5632 18164 5684 18216
rect 204 18096 256 18148
rect 1952 18071 2004 18080
rect 1952 18037 1961 18071
rect 1961 18037 1995 18071
rect 1995 18037 2004 18071
rect 1952 18028 2004 18037
rect 2044 18028 2096 18080
rect 2780 18028 2832 18080
rect 2964 18096 3016 18148
rect 3332 18139 3384 18148
rect 3332 18105 3341 18139
rect 3341 18105 3375 18139
rect 3375 18105 3384 18139
rect 3332 18096 3384 18105
rect 4712 18096 4764 18148
rect 4804 18096 4856 18148
rect 7196 18207 7248 18216
rect 7196 18173 7205 18207
rect 7205 18173 7239 18207
rect 7239 18173 7248 18207
rect 7196 18164 7248 18173
rect 7472 18241 7481 18275
rect 7481 18241 7515 18275
rect 7515 18241 7524 18275
rect 7472 18232 7524 18241
rect 8392 18232 8444 18284
rect 13084 18300 13136 18352
rect 9496 18232 9548 18284
rect 10140 18232 10192 18284
rect 12072 18232 12124 18284
rect 13452 18368 13504 18420
rect 14188 18232 14240 18284
rect 6920 18096 6972 18148
rect 9036 18164 9088 18216
rect 10048 18164 10100 18216
rect 10968 18164 11020 18216
rect 13636 18164 13688 18216
rect 10876 18096 10928 18148
rect 11152 18139 11204 18148
rect 11152 18105 11161 18139
rect 11161 18105 11195 18139
rect 11195 18105 11204 18139
rect 11152 18096 11204 18105
rect 11888 18096 11940 18148
rect 4344 18028 4396 18080
rect 5264 18028 5316 18080
rect 5540 18028 5592 18080
rect 8576 18071 8628 18080
rect 8576 18037 8585 18071
rect 8585 18037 8619 18071
rect 8619 18037 8628 18071
rect 8576 18028 8628 18037
rect 8944 18071 8996 18080
rect 8944 18037 8953 18071
rect 8953 18037 8987 18071
rect 8987 18037 8996 18071
rect 8944 18028 8996 18037
rect 9680 18028 9732 18080
rect 11060 18028 11112 18080
rect 11704 18028 11756 18080
rect 13268 18028 13320 18080
rect 19616 18164 19668 18216
rect 21272 18164 21324 18216
rect 15476 18096 15528 18148
rect 15660 18096 15712 18148
rect 16764 18096 16816 18148
rect 18052 18139 18104 18148
rect 18052 18105 18061 18139
rect 18061 18105 18095 18139
rect 18095 18105 18104 18139
rect 18052 18096 18104 18105
rect 21088 18096 21140 18148
rect 22192 18096 22244 18148
rect 15384 18028 15436 18080
rect 17960 18028 18012 18080
rect 18972 18028 19024 18080
rect 19708 18028 19760 18080
rect 20352 18028 20404 18080
rect 20720 18028 20772 18080
rect 21732 18028 21784 18080
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 2504 17824 2556 17876
rect 7012 17824 7064 17876
rect 8208 17867 8260 17876
rect 8208 17833 8217 17867
rect 8217 17833 8251 17867
rect 8251 17833 8260 17867
rect 8208 17824 8260 17833
rect 9680 17867 9732 17876
rect 9680 17833 9689 17867
rect 9689 17833 9723 17867
rect 9723 17833 9732 17867
rect 9680 17824 9732 17833
rect 9772 17824 9824 17876
rect 1400 17756 1452 17808
rect 2228 17731 2280 17740
rect 2228 17697 2237 17731
rect 2237 17697 2271 17731
rect 2271 17697 2280 17731
rect 2228 17688 2280 17697
rect 4160 17688 4212 17740
rect 7472 17688 7524 17740
rect 8208 17688 8260 17740
rect 10140 17688 10192 17740
rect 2412 17663 2464 17672
rect 2412 17629 2421 17663
rect 2421 17629 2455 17663
rect 2455 17629 2464 17663
rect 2412 17620 2464 17629
rect 6828 17663 6880 17672
rect 6828 17629 6837 17663
rect 6837 17629 6871 17663
rect 6871 17629 6880 17663
rect 6828 17620 6880 17629
rect 10324 17663 10376 17672
rect 10324 17629 10333 17663
rect 10333 17629 10367 17663
rect 10367 17629 10376 17663
rect 11152 17688 11204 17740
rect 13176 17824 13228 17876
rect 13636 17824 13688 17876
rect 12992 17688 13044 17740
rect 13728 17731 13780 17740
rect 13728 17697 13737 17731
rect 13737 17697 13771 17731
rect 13771 17697 13780 17731
rect 13728 17688 13780 17697
rect 15292 17731 15344 17740
rect 15292 17697 15301 17731
rect 15301 17697 15335 17731
rect 15335 17697 15344 17731
rect 15292 17688 15344 17697
rect 13912 17663 13964 17672
rect 10324 17620 10376 17629
rect 3148 17484 3200 17536
rect 3884 17484 3936 17536
rect 4068 17484 4120 17536
rect 4988 17484 5040 17536
rect 5448 17527 5500 17536
rect 5448 17493 5457 17527
rect 5457 17493 5491 17527
rect 5491 17493 5500 17527
rect 5448 17484 5500 17493
rect 13912 17629 13921 17663
rect 13921 17629 13955 17663
rect 13955 17629 13964 17663
rect 13912 17620 13964 17629
rect 14004 17620 14056 17672
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 3976 17280 4028 17332
rect 7748 17280 7800 17332
rect 8208 17323 8260 17332
rect 8208 17289 8217 17323
rect 8217 17289 8251 17323
rect 8251 17289 8260 17323
rect 8208 17280 8260 17289
rect 4988 17212 5040 17264
rect 6828 17212 6880 17264
rect 2504 17144 2556 17196
rect 3976 17187 4028 17196
rect 3976 17153 3985 17187
rect 3985 17153 4019 17187
rect 4019 17153 4028 17187
rect 3976 17144 4028 17153
rect 8484 17144 8536 17196
rect 9956 17280 10008 17332
rect 11244 17280 11296 17332
rect 15292 17280 15344 17332
rect 15476 17323 15528 17332
rect 15476 17289 15485 17323
rect 15485 17289 15519 17323
rect 15519 17289 15528 17323
rect 15476 17280 15528 17289
rect 5448 17076 5500 17128
rect 6184 17076 6236 17128
rect 6828 17119 6880 17128
rect 6828 17085 6837 17119
rect 6837 17085 6871 17119
rect 6871 17085 6880 17119
rect 6828 17076 6880 17085
rect 5540 17008 5592 17060
rect 8576 17076 8628 17128
rect 10324 17076 10376 17128
rect 4712 16940 4764 16992
rect 5448 16940 5500 16992
rect 7472 17008 7524 17060
rect 12624 17212 12676 17264
rect 20812 17212 20864 17264
rect 21088 17212 21140 17264
rect 12992 17187 13044 17196
rect 12992 17153 13001 17187
rect 13001 17153 13035 17187
rect 13035 17153 13044 17187
rect 12992 17144 13044 17153
rect 13636 17144 13688 17196
rect 10876 17076 10928 17128
rect 14004 17076 14056 17128
rect 7012 16940 7064 16992
rect 11060 17008 11112 17060
rect 14372 17051 14424 17060
rect 14372 17017 14406 17051
rect 14406 17017 14424 17051
rect 14372 17008 14424 17017
rect 9496 16940 9548 16992
rect 15660 16940 15712 16992
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 2228 16736 2280 16788
rect 4344 16736 4396 16788
rect 6920 16736 6972 16788
rect 7564 16736 7616 16788
rect 7748 16736 7800 16788
rect 3608 16600 3660 16652
rect 9680 16736 9732 16788
rect 9956 16736 10008 16788
rect 5448 16600 5500 16652
rect 7012 16600 7064 16652
rect 4344 16532 4396 16584
rect 4712 16575 4764 16584
rect 4712 16541 4721 16575
rect 4721 16541 4755 16575
rect 4755 16541 4764 16575
rect 4712 16532 4764 16541
rect 7380 16600 7432 16652
rect 7472 16575 7524 16584
rect 7472 16541 7481 16575
rect 7481 16541 7515 16575
rect 7515 16541 7524 16575
rect 7472 16532 7524 16541
rect 8208 16532 8260 16584
rect 11152 16643 11204 16652
rect 11152 16609 11161 16643
rect 11161 16609 11195 16643
rect 11195 16609 11204 16643
rect 11152 16600 11204 16609
rect 12992 16736 13044 16788
rect 12072 16668 12124 16720
rect 13728 16736 13780 16788
rect 15660 16779 15712 16788
rect 15660 16745 15669 16779
rect 15669 16745 15703 16779
rect 15703 16745 15712 16779
rect 15660 16736 15712 16745
rect 13268 16600 13320 16652
rect 14004 16643 14056 16652
rect 14004 16609 14013 16643
rect 14013 16609 14047 16643
rect 14047 16609 14056 16643
rect 14004 16600 14056 16609
rect 7564 16464 7616 16516
rect 4068 16396 4120 16448
rect 14372 16532 14424 16584
rect 15108 16532 15160 16584
rect 15476 16532 15528 16584
rect 12164 16396 12216 16448
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 9680 16192 9732 16244
rect 15108 16235 15160 16244
rect 9588 16124 9640 16176
rect 15108 16201 15117 16235
rect 15117 16201 15151 16235
rect 15151 16201 15160 16235
rect 15108 16192 15160 16201
rect 2872 16056 2924 16108
rect 3792 16099 3844 16108
rect 3792 16065 3801 16099
rect 3801 16065 3835 16099
rect 3835 16065 3844 16099
rect 3792 16056 3844 16065
rect 8300 16056 8352 16108
rect 8484 16099 8536 16108
rect 8484 16065 8493 16099
rect 8493 16065 8527 16099
rect 8527 16065 8536 16099
rect 8484 16056 8536 16065
rect 11704 16056 11756 16108
rect 12624 16099 12676 16108
rect 12624 16065 12633 16099
rect 12633 16065 12667 16099
rect 12667 16065 12676 16099
rect 12624 16056 12676 16065
rect 4344 15988 4396 16040
rect 9496 15988 9548 16040
rect 12440 16031 12492 16040
rect 12440 15997 12449 16031
rect 12449 15997 12483 16031
rect 12483 15997 12492 16031
rect 13728 16031 13780 16040
rect 12440 15988 12492 15997
rect 13728 15997 13737 16031
rect 13737 15997 13771 16031
rect 13771 15997 13780 16031
rect 13728 15988 13780 15997
rect 7380 15920 7432 15972
rect 5172 15895 5224 15904
rect 5172 15861 5181 15895
rect 5181 15861 5215 15895
rect 5215 15861 5224 15895
rect 5172 15852 5224 15861
rect 6920 15852 6972 15904
rect 9680 15852 9732 15904
rect 13544 15920 13596 15972
rect 14004 15963 14056 15972
rect 14004 15929 14038 15963
rect 14038 15929 14056 15963
rect 14004 15920 14056 15929
rect 11060 15852 11112 15904
rect 11244 15895 11296 15904
rect 11244 15861 11253 15895
rect 11253 15861 11287 15895
rect 11287 15861 11296 15895
rect 11244 15852 11296 15861
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 7472 15648 7524 15700
rect 9680 15691 9732 15700
rect 9680 15657 9689 15691
rect 9689 15657 9723 15691
rect 9723 15657 9732 15691
rect 9680 15648 9732 15657
rect 10048 15648 10100 15700
rect 11152 15648 11204 15700
rect 11980 15648 12032 15700
rect 12164 15648 12216 15700
rect 13544 15691 13596 15700
rect 13544 15657 13553 15691
rect 13553 15657 13587 15691
rect 13587 15657 13596 15691
rect 13544 15648 13596 15657
rect 16120 15648 16172 15700
rect 5172 15623 5224 15632
rect 5172 15589 5206 15623
rect 5206 15589 5224 15623
rect 5172 15580 5224 15589
rect 5540 15580 5592 15632
rect 6552 15580 6604 15632
rect 3056 15512 3108 15564
rect 8300 15512 8352 15564
rect 9220 15512 9272 15564
rect 11244 15512 11296 15564
rect 11796 15512 11848 15564
rect 11888 15512 11940 15564
rect 15476 15555 15528 15564
rect 15476 15521 15485 15555
rect 15485 15521 15519 15555
rect 15519 15521 15528 15555
rect 15476 15512 15528 15521
rect 4252 15444 4304 15496
rect 6828 15444 6880 15496
rect 7104 15487 7156 15496
rect 7104 15453 7113 15487
rect 7113 15453 7147 15487
rect 7147 15453 7156 15487
rect 7104 15444 7156 15453
rect 9588 15376 9640 15428
rect 12072 15444 12124 15496
rect 12256 15444 12308 15496
rect 14004 15444 14056 15496
rect 14924 15444 14976 15496
rect 11244 15376 11296 15428
rect 6460 15308 6512 15360
rect 7748 15308 7800 15360
rect 12808 15308 12860 15360
rect 14096 15308 14148 15360
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 3056 15147 3108 15156
rect 3056 15113 3065 15147
rect 3065 15113 3099 15147
rect 3099 15113 3108 15147
rect 3056 15104 3108 15113
rect 4068 15104 4120 15156
rect 8208 15104 8260 15156
rect 9220 15147 9272 15156
rect 9220 15113 9229 15147
rect 9229 15113 9263 15147
rect 9263 15113 9272 15147
rect 9220 15104 9272 15113
rect 12256 15104 12308 15156
rect 6460 15036 6512 15088
rect 5172 15011 5224 15020
rect 5172 14977 5181 15011
rect 5181 14977 5215 15011
rect 5215 14977 5224 15011
rect 5172 14968 5224 14977
rect 7104 14968 7156 15020
rect 11244 15011 11296 15020
rect 11244 14977 11253 15011
rect 11253 14977 11287 15011
rect 11287 14977 11296 15011
rect 11244 14968 11296 14977
rect 11704 15036 11756 15088
rect 14832 15104 14884 15156
rect 14924 15104 14976 15156
rect 4988 14900 5040 14952
rect 5356 14900 5408 14952
rect 6368 14943 6420 14952
rect 6368 14909 6377 14943
rect 6377 14909 6411 14943
rect 6411 14909 6420 14943
rect 6368 14900 6420 14909
rect 6460 14900 6512 14952
rect 7288 14900 7340 14952
rect 9588 14900 9640 14952
rect 10784 14900 10836 14952
rect 12440 14943 12492 14952
rect 12440 14909 12449 14943
rect 12449 14909 12483 14943
rect 12483 14909 12492 14943
rect 12440 14900 12492 14909
rect 13728 14900 13780 14952
rect 1952 14807 2004 14816
rect 1952 14773 1961 14807
rect 1961 14773 1995 14807
rect 1995 14773 2004 14807
rect 1952 14764 2004 14773
rect 5540 14764 5592 14816
rect 6184 14807 6236 14816
rect 6184 14773 6193 14807
rect 6193 14773 6227 14807
rect 6227 14773 6236 14807
rect 6184 14764 6236 14773
rect 8944 14764 8996 14816
rect 12072 14832 12124 14884
rect 14832 14832 14884 14884
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 3516 14560 3568 14612
rect 4988 14560 5040 14612
rect 11060 14560 11112 14612
rect 12072 14603 12124 14612
rect 12072 14569 12081 14603
rect 12081 14569 12115 14603
rect 12115 14569 12124 14603
rect 12072 14560 12124 14569
rect 16764 14603 16816 14612
rect 16764 14569 16773 14603
rect 16773 14569 16807 14603
rect 16807 14569 16816 14603
rect 16764 14560 16816 14569
rect 2964 14424 3016 14476
rect 4068 14467 4120 14476
rect 4068 14433 4077 14467
rect 4077 14433 4111 14467
rect 4111 14433 4120 14467
rect 4068 14424 4120 14433
rect 2872 14399 2924 14408
rect 2872 14365 2881 14399
rect 2881 14365 2915 14399
rect 2915 14365 2924 14399
rect 2872 14356 2924 14365
rect 3240 14356 3292 14408
rect 6736 14424 6788 14476
rect 7656 14424 7708 14476
rect 8300 14467 8352 14476
rect 8300 14433 8309 14467
rect 8309 14433 8343 14467
rect 8343 14433 8352 14467
rect 8300 14424 8352 14433
rect 10600 14424 10652 14476
rect 6644 14356 6696 14408
rect 3884 14288 3936 14340
rect 6736 14288 6788 14340
rect 8484 14356 8536 14408
rect 9220 14356 9272 14408
rect 14740 14492 14792 14544
rect 16396 14492 16448 14544
rect 13452 14467 13504 14476
rect 13452 14433 13461 14467
rect 13461 14433 13495 14467
rect 13495 14433 13504 14467
rect 13452 14424 13504 14433
rect 15292 14467 15344 14476
rect 15292 14433 15301 14467
rect 15301 14433 15335 14467
rect 15335 14433 15344 14467
rect 15292 14424 15344 14433
rect 16304 14424 16356 14476
rect 13912 14356 13964 14408
rect 4160 14220 4212 14272
rect 7196 14220 7248 14272
rect 7288 14220 7340 14272
rect 16764 14220 16816 14272
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 3792 14016 3844 14068
rect 4160 14016 4212 14068
rect 15292 14016 15344 14068
rect 7104 13948 7156 14000
rect 10600 13991 10652 14000
rect 10600 13957 10609 13991
rect 10609 13957 10643 13991
rect 10643 13957 10652 13991
rect 10600 13948 10652 13957
rect 11060 13948 11112 14000
rect 1676 13812 1728 13864
rect 3792 13812 3844 13864
rect 5724 13880 5776 13932
rect 6736 13880 6788 13932
rect 9220 13923 9272 13932
rect 9220 13889 9229 13923
rect 9229 13889 9263 13923
rect 9263 13889 9272 13923
rect 9220 13880 9272 13889
rect 12072 13880 12124 13932
rect 15476 13880 15528 13932
rect 16304 13923 16356 13932
rect 16304 13889 16313 13923
rect 16313 13889 16347 13923
rect 16347 13889 16356 13923
rect 16304 13880 16356 13889
rect 3056 13744 3108 13796
rect 6184 13812 6236 13864
rect 10692 13812 10744 13864
rect 12716 13812 12768 13864
rect 14740 13855 14792 13864
rect 14740 13821 14749 13855
rect 14749 13821 14783 13855
rect 14783 13821 14792 13855
rect 14740 13812 14792 13821
rect 16028 13855 16080 13864
rect 16028 13821 16037 13855
rect 16037 13821 16071 13855
rect 16071 13821 16080 13855
rect 16028 13812 16080 13821
rect 4804 13744 4856 13796
rect 12808 13787 12860 13796
rect 12808 13753 12817 13787
rect 12817 13753 12851 13787
rect 12851 13753 12860 13787
rect 12808 13744 12860 13753
rect 3240 13719 3292 13728
rect 3240 13685 3249 13719
rect 3249 13685 3283 13719
rect 3283 13685 3292 13719
rect 3240 13676 3292 13685
rect 5724 13719 5776 13728
rect 5724 13685 5733 13719
rect 5733 13685 5767 13719
rect 5767 13685 5776 13719
rect 5724 13676 5776 13685
rect 7012 13676 7064 13728
rect 7288 13719 7340 13728
rect 7288 13685 7297 13719
rect 7297 13685 7331 13719
rect 7331 13685 7340 13719
rect 7288 13676 7340 13685
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 2872 13472 2924 13524
rect 5264 13472 5316 13524
rect 1124 13404 1176 13456
rect 2780 13379 2832 13388
rect 2780 13345 2789 13379
rect 2789 13345 2823 13379
rect 2823 13345 2832 13379
rect 2780 13336 2832 13345
rect 3792 13336 3844 13388
rect 5724 13404 5776 13456
rect 7288 13472 7340 13524
rect 7380 13472 7432 13524
rect 7656 13472 7708 13524
rect 10968 13472 11020 13524
rect 13452 13472 13504 13524
rect 10140 13447 10192 13456
rect 10140 13413 10149 13447
rect 10149 13413 10183 13447
rect 10183 13413 10192 13447
rect 10140 13404 10192 13413
rect 7748 13336 7800 13388
rect 9128 13336 9180 13388
rect 10876 13336 10928 13388
rect 12440 13404 12492 13456
rect 15568 13447 15620 13456
rect 15568 13413 15577 13447
rect 15577 13413 15611 13447
rect 15611 13413 15620 13447
rect 15568 13404 15620 13413
rect 12072 13379 12124 13388
rect 12072 13345 12106 13379
rect 12106 13345 12124 13379
rect 12072 13336 12124 13345
rect 15752 13336 15804 13388
rect 1952 13268 2004 13320
rect 2872 13311 2924 13320
rect 2872 13277 2881 13311
rect 2881 13277 2915 13311
rect 2915 13277 2924 13311
rect 2872 13268 2924 13277
rect 3056 13311 3108 13320
rect 3056 13277 3065 13311
rect 3065 13277 3099 13311
rect 3099 13277 3108 13311
rect 3056 13268 3108 13277
rect 7564 13311 7616 13320
rect 4804 13132 4856 13184
rect 7564 13277 7573 13311
rect 7573 13277 7607 13311
rect 7607 13277 7616 13311
rect 7564 13268 7616 13277
rect 10692 13268 10744 13320
rect 14188 13311 14240 13320
rect 14188 13277 14197 13311
rect 14197 13277 14231 13311
rect 14231 13277 14240 13311
rect 14188 13268 14240 13277
rect 6184 13175 6236 13184
rect 6184 13141 6193 13175
rect 6193 13141 6227 13175
rect 6227 13141 6236 13175
rect 6184 13132 6236 13141
rect 8852 13132 8904 13184
rect 11796 13132 11848 13184
rect 13452 13200 13504 13252
rect 13176 13175 13228 13184
rect 13176 13141 13185 13175
rect 13185 13141 13219 13175
rect 13219 13141 13228 13175
rect 13176 13132 13228 13141
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 2964 12928 3016 12980
rect 4804 12928 4856 12980
rect 6092 12928 6144 12980
rect 6368 12928 6420 12980
rect 7012 12971 7064 12980
rect 7012 12937 7021 12971
rect 7021 12937 7055 12971
rect 7055 12937 7064 12971
rect 7012 12928 7064 12937
rect 7288 12928 7340 12980
rect 11244 12928 11296 12980
rect 15752 12971 15804 12980
rect 15752 12937 15761 12971
rect 15761 12937 15795 12971
rect 15795 12937 15804 12971
rect 15752 12928 15804 12937
rect 3056 12792 3108 12844
rect 1952 12767 2004 12776
rect 1952 12733 1961 12767
rect 1961 12733 1995 12767
rect 1995 12733 2004 12767
rect 1952 12724 2004 12733
rect 2964 12724 3016 12776
rect 3240 12724 3292 12776
rect 4252 12724 4304 12776
rect 7564 12835 7616 12844
rect 7564 12801 7573 12835
rect 7573 12801 7607 12835
rect 7607 12801 7616 12835
rect 7564 12792 7616 12801
rect 8944 12860 8996 12912
rect 10692 12860 10744 12912
rect 10876 12792 10928 12844
rect 11060 12835 11112 12844
rect 11060 12801 11069 12835
rect 11069 12801 11103 12835
rect 11103 12801 11112 12835
rect 11060 12792 11112 12801
rect 13176 12792 13228 12844
rect 16304 12835 16356 12844
rect 16304 12801 16313 12835
rect 16313 12801 16347 12835
rect 16347 12801 16356 12835
rect 16304 12792 16356 12801
rect 6920 12724 6972 12776
rect 7288 12724 7340 12776
rect 9036 12724 9088 12776
rect 12440 12724 12492 12776
rect 13544 12767 13596 12776
rect 13544 12733 13553 12767
rect 13553 12733 13587 12767
rect 13587 12733 13596 12767
rect 13544 12724 13596 12733
rect 14188 12724 14240 12776
rect 664 12656 716 12708
rect 2320 12656 2372 12708
rect 6736 12656 6788 12708
rect 2044 12631 2096 12640
rect 2044 12597 2053 12631
rect 2053 12597 2087 12631
rect 2087 12597 2096 12631
rect 2044 12588 2096 12597
rect 5632 12588 5684 12640
rect 12256 12656 12308 12708
rect 13820 12699 13872 12708
rect 13820 12665 13854 12699
rect 13854 12665 13872 12699
rect 13820 12656 13872 12665
rect 14648 12588 14700 12640
rect 16212 12631 16264 12640
rect 16212 12597 16221 12631
rect 16221 12597 16255 12631
rect 16255 12597 16264 12631
rect 16212 12588 16264 12597
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 3056 12427 3108 12436
rect 3056 12393 3065 12427
rect 3065 12393 3099 12427
rect 3099 12393 3108 12427
rect 3056 12384 3108 12393
rect 6644 12427 6696 12436
rect 6644 12393 6653 12427
rect 6653 12393 6687 12427
rect 6687 12393 6696 12427
rect 6644 12384 6696 12393
rect 8300 12384 8352 12436
rect 8852 12384 8904 12436
rect 2964 12316 3016 12368
rect 4068 12316 4120 12368
rect 16028 12384 16080 12436
rect 1676 12291 1728 12300
rect 1676 12257 1685 12291
rect 1685 12257 1719 12291
rect 1719 12257 1728 12291
rect 1676 12248 1728 12257
rect 3608 12248 3660 12300
rect 4344 12248 4396 12300
rect 4896 12248 4948 12300
rect 7472 12248 7524 12300
rect 8944 12248 8996 12300
rect 2872 12112 2924 12164
rect 5540 12180 5592 12232
rect 6552 12180 6604 12232
rect 4804 12112 4856 12164
rect 7564 12180 7616 12232
rect 10600 12316 10652 12368
rect 11704 12359 11756 12368
rect 11704 12325 11713 12359
rect 11713 12325 11747 12359
rect 11747 12325 11756 12359
rect 11704 12316 11756 12325
rect 11888 12316 11940 12368
rect 16304 12316 16356 12368
rect 17868 12316 17920 12368
rect 9312 12248 9364 12300
rect 12624 12248 12676 12300
rect 13268 12291 13320 12300
rect 13268 12257 13277 12291
rect 13277 12257 13311 12291
rect 13311 12257 13320 12291
rect 13268 12248 13320 12257
rect 14188 12248 14240 12300
rect 16580 12248 16632 12300
rect 9404 12180 9456 12232
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 10416 12180 10468 12232
rect 12716 12180 12768 12232
rect 8392 12112 8444 12164
rect 5632 12044 5684 12096
rect 10600 12112 10652 12164
rect 11888 12112 11940 12164
rect 13544 12112 13596 12164
rect 14556 12112 14608 12164
rect 10692 12044 10744 12096
rect 12808 12087 12860 12096
rect 12808 12053 12817 12087
rect 12817 12053 12851 12087
rect 12851 12053 12860 12087
rect 12808 12044 12860 12053
rect 14464 12044 14516 12096
rect 16304 12044 16356 12096
rect 16672 12087 16724 12096
rect 16672 12053 16681 12087
rect 16681 12053 16715 12087
rect 16715 12053 16724 12087
rect 16672 12044 16724 12053
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 1860 11840 1912 11892
rect 2780 11840 2832 11892
rect 3608 11747 3660 11756
rect 3608 11713 3617 11747
rect 3617 11713 3651 11747
rect 3651 11713 3660 11747
rect 5540 11840 5592 11892
rect 3608 11704 3660 11713
rect 2412 11636 2464 11688
rect 3424 11636 3476 11688
rect 3792 11568 3844 11620
rect 4344 11568 4396 11620
rect 4620 11636 4672 11688
rect 7104 11704 7156 11756
rect 7196 11679 7248 11688
rect 7196 11645 7205 11679
rect 7205 11645 7239 11679
rect 7239 11645 7248 11679
rect 7196 11636 7248 11645
rect 6184 11568 6236 11620
rect 7748 11704 7800 11756
rect 12716 11840 12768 11892
rect 14740 11840 14792 11892
rect 16212 11883 16264 11892
rect 16212 11849 16221 11883
rect 16221 11849 16255 11883
rect 16255 11849 16264 11883
rect 16212 11840 16264 11849
rect 16304 11840 16356 11892
rect 11888 11772 11940 11824
rect 13820 11815 13872 11824
rect 13820 11781 13829 11815
rect 13829 11781 13863 11815
rect 13863 11781 13872 11815
rect 13820 11772 13872 11781
rect 14372 11772 14424 11824
rect 10968 11704 11020 11756
rect 11152 11747 11204 11756
rect 11152 11713 11161 11747
rect 11161 11713 11195 11747
rect 11195 11713 11204 11747
rect 11152 11704 11204 11713
rect 11336 11747 11388 11756
rect 11336 11713 11345 11747
rect 11345 11713 11379 11747
rect 11379 11713 11388 11747
rect 11336 11704 11388 11713
rect 10324 11636 10376 11688
rect 12440 11679 12492 11688
rect 12440 11645 12449 11679
rect 12449 11645 12483 11679
rect 12483 11645 12492 11679
rect 12440 11636 12492 11645
rect 3424 11543 3476 11552
rect 3424 11509 3433 11543
rect 3433 11509 3467 11543
rect 3467 11509 3476 11543
rect 3424 11500 3476 11509
rect 3700 11500 3752 11552
rect 5908 11543 5960 11552
rect 5908 11509 5917 11543
rect 5917 11509 5951 11543
rect 5951 11509 5960 11543
rect 5908 11500 5960 11509
rect 7196 11500 7248 11552
rect 8576 11568 8628 11620
rect 10416 11568 10468 11620
rect 10692 11568 10744 11620
rect 12164 11568 12216 11620
rect 14648 11636 14700 11688
rect 12808 11568 12860 11620
rect 15292 11500 15344 11552
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 2320 11228 2372 11280
rect 4804 11296 4856 11348
rect 8300 11296 8352 11348
rect 8576 11339 8628 11348
rect 8576 11305 8585 11339
rect 8585 11305 8619 11339
rect 8619 11305 8628 11339
rect 8576 11296 8628 11305
rect 8668 11296 8720 11348
rect 11520 11296 11572 11348
rect 4252 11228 4304 11280
rect 5540 11228 5592 11280
rect 2780 11203 2832 11212
rect 2780 11169 2789 11203
rect 2789 11169 2823 11203
rect 2823 11169 2832 11203
rect 2780 11160 2832 11169
rect 4528 11160 4580 11212
rect 7104 11160 7156 11212
rect 7196 11203 7248 11212
rect 7196 11169 7205 11203
rect 7205 11169 7239 11203
rect 7239 11169 7248 11203
rect 7196 11160 7248 11169
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 2136 11092 2188 11144
rect 4160 11024 4212 11076
rect 3884 10956 3936 11008
rect 5908 11092 5960 11144
rect 6092 11135 6144 11144
rect 6092 11101 6101 11135
rect 6101 11101 6135 11135
rect 6135 11101 6144 11135
rect 6092 11092 6144 11101
rect 6276 11135 6328 11144
rect 6276 11101 6285 11135
rect 6285 11101 6319 11135
rect 6319 11101 6328 11135
rect 6276 11092 6328 11101
rect 6920 11092 6972 11144
rect 8300 11160 8352 11212
rect 10968 11228 11020 11280
rect 11060 11228 11112 11280
rect 11336 11228 11388 11280
rect 11704 11228 11756 11280
rect 12532 11296 12584 11348
rect 14188 11339 14240 11348
rect 14188 11305 14197 11339
rect 14197 11305 14231 11339
rect 14231 11305 14240 11339
rect 14188 11296 14240 11305
rect 17040 11296 17092 11348
rect 17960 11228 18012 11280
rect 8852 11160 8904 11212
rect 10508 11160 10560 11212
rect 12716 11160 12768 11212
rect 9680 11092 9732 11144
rect 8208 11024 8260 11076
rect 10048 11024 10100 11076
rect 13452 11160 13504 11212
rect 14464 11160 14516 11212
rect 13084 11135 13136 11144
rect 13084 11101 13093 11135
rect 13093 11101 13127 11135
rect 13127 11101 13136 11135
rect 13084 11092 13136 11101
rect 13176 11135 13228 11144
rect 13176 11101 13185 11135
rect 13185 11101 13219 11135
rect 13219 11101 13228 11135
rect 13176 11092 13228 11101
rect 14556 11092 14608 11144
rect 5632 10999 5684 11008
rect 5632 10965 5641 10999
rect 5641 10965 5675 10999
rect 5675 10965 5684 10999
rect 5632 10956 5684 10965
rect 9956 10956 10008 11008
rect 12164 10956 12216 11008
rect 12532 10956 12584 11008
rect 12716 10956 12768 11008
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 2780 10752 2832 10804
rect 8208 10795 8260 10804
rect 8208 10761 8217 10795
rect 8217 10761 8251 10795
rect 8251 10761 8260 10795
rect 8208 10752 8260 10761
rect 9956 10752 10008 10804
rect 10048 10752 10100 10804
rect 13176 10752 13228 10804
rect 4896 10727 4948 10736
rect 4896 10693 4905 10727
rect 4905 10693 4939 10727
rect 4939 10693 4948 10727
rect 4896 10684 4948 10693
rect 9588 10684 9640 10736
rect 2044 10659 2096 10668
rect 2044 10625 2053 10659
rect 2053 10625 2087 10659
rect 2087 10625 2096 10659
rect 2044 10616 2096 10625
rect 2136 10659 2188 10668
rect 2136 10625 2145 10659
rect 2145 10625 2179 10659
rect 2179 10625 2188 10659
rect 3884 10659 3936 10668
rect 2136 10616 2188 10625
rect 3884 10625 3893 10659
rect 3893 10625 3927 10659
rect 3927 10625 3936 10659
rect 3884 10616 3936 10625
rect 4160 10616 4212 10668
rect 5448 10659 5500 10668
rect 5448 10625 5457 10659
rect 5457 10625 5491 10659
rect 5491 10625 5500 10659
rect 5448 10616 5500 10625
rect 1400 10548 1452 10600
rect 3792 10548 3844 10600
rect 4068 10548 4120 10600
rect 6368 10548 6420 10600
rect 6828 10591 6880 10600
rect 6828 10557 6837 10591
rect 6837 10557 6871 10591
rect 6871 10557 6880 10591
rect 6828 10548 6880 10557
rect 9128 10616 9180 10668
rect 6276 10480 6328 10532
rect 9680 10548 9732 10600
rect 11060 10548 11112 10600
rect 12256 10548 12308 10600
rect 14556 10548 14608 10600
rect 16672 10548 16724 10600
rect 12624 10480 12676 10532
rect 12900 10480 12952 10532
rect 3424 10412 3476 10464
rect 3976 10412 4028 10464
rect 6460 10455 6512 10464
rect 6460 10421 6469 10455
rect 6469 10421 6503 10455
rect 6503 10421 6512 10455
rect 6460 10412 6512 10421
rect 6552 10412 6604 10464
rect 16212 10412 16264 10464
rect 16396 10412 16448 10464
rect 18052 10455 18104 10464
rect 18052 10421 18061 10455
rect 18061 10421 18095 10455
rect 18095 10421 18104 10455
rect 18052 10412 18104 10421
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 2136 10208 2188 10260
rect 6276 10208 6328 10260
rect 7104 10208 7156 10260
rect 7472 10208 7524 10260
rect 10324 10208 10376 10260
rect 11244 10208 11296 10260
rect 11796 10208 11848 10260
rect 3884 10140 3936 10192
rect 4988 10140 5040 10192
rect 2412 10072 2464 10124
rect 5540 10072 5592 10124
rect 12256 10140 12308 10192
rect 18052 10208 18104 10260
rect 4344 10004 4396 10056
rect 7748 10047 7800 10056
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 10324 10072 10376 10124
rect 15292 10072 15344 10124
rect 16212 10072 16264 10124
rect 17500 10140 17552 10192
rect 7748 10004 7800 10013
rect 14096 10047 14148 10056
rect 7380 9936 7432 9988
rect 14096 10013 14105 10047
rect 14105 10013 14139 10047
rect 14139 10013 14148 10047
rect 14096 10004 14148 10013
rect 14740 10004 14792 10056
rect 16396 10047 16448 10056
rect 16396 10013 16405 10047
rect 16405 10013 16439 10047
rect 16439 10013 16448 10047
rect 16396 10004 16448 10013
rect 12716 9936 12768 9988
rect 16580 9936 16632 9988
rect 3700 9868 3752 9920
rect 8852 9868 8904 9920
rect 11060 9868 11112 9920
rect 11244 9911 11296 9920
rect 11244 9877 11253 9911
rect 11253 9877 11287 9911
rect 11287 9877 11296 9911
rect 11244 9868 11296 9877
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 2412 9596 2464 9648
rect 4344 9664 4396 9716
rect 4988 9707 5040 9716
rect 4988 9673 4997 9707
rect 4997 9673 5031 9707
rect 5031 9673 5040 9707
rect 4988 9664 5040 9673
rect 6920 9664 6972 9716
rect 10600 9664 10652 9716
rect 15200 9664 15252 9716
rect 6092 9596 6144 9648
rect 7196 9596 7248 9648
rect 8392 9596 8444 9648
rect 10232 9596 10284 9648
rect 11152 9596 11204 9648
rect 17960 9596 18012 9648
rect 7380 9528 7432 9580
rect 7748 9528 7800 9580
rect 14556 9528 14608 9580
rect 2136 9460 2188 9512
rect 5448 9460 5500 9512
rect 6460 9460 6512 9512
rect 6920 9460 6972 9512
rect 9772 9460 9824 9512
rect 10324 9460 10376 9512
rect 11244 9460 11296 9512
rect 12072 9460 12124 9512
rect 12256 9460 12308 9512
rect 16396 9460 16448 9512
rect 18144 9460 18196 9512
rect 4068 9392 4120 9444
rect 7196 9367 7248 9376
rect 7196 9333 7205 9367
rect 7205 9333 7239 9367
rect 7239 9333 7248 9367
rect 7196 9324 7248 9333
rect 12900 9392 12952 9444
rect 13268 9392 13320 9444
rect 11060 9324 11112 9376
rect 12072 9324 12124 9376
rect 14188 9324 14240 9376
rect 14740 9324 14792 9376
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 3332 9120 3384 9172
rect 4344 9120 4396 9172
rect 4988 9120 5040 9172
rect 9312 9120 9364 9172
rect 11060 9163 11112 9172
rect 11060 9129 11069 9163
rect 11069 9129 11103 9163
rect 11103 9129 11112 9163
rect 11060 9120 11112 9129
rect 11612 9120 11664 9172
rect 11980 9120 12032 9172
rect 14096 9120 14148 9172
rect 12164 9052 12216 9104
rect 18144 9095 18196 9104
rect 18144 9061 18153 9095
rect 18153 9061 18187 9095
rect 18187 9061 18196 9095
rect 18144 9052 18196 9061
rect 2228 8984 2280 9036
rect 5264 8984 5316 9036
rect 6460 8984 6512 9036
rect 7288 9027 7340 9036
rect 7288 8993 7297 9027
rect 7297 8993 7331 9027
rect 7331 8993 7340 9027
rect 7288 8984 7340 8993
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 10232 8984 10284 9036
rect 12072 9027 12124 9036
rect 12072 8993 12081 9027
rect 12081 8993 12115 9027
rect 12115 8993 12124 9027
rect 12072 8984 12124 8993
rect 2872 8959 2924 8968
rect 2872 8925 2881 8959
rect 2881 8925 2915 8959
rect 2915 8925 2924 8959
rect 2872 8916 2924 8925
rect 3700 8916 3752 8968
rect 5172 8959 5224 8968
rect 5172 8925 5181 8959
rect 5181 8925 5215 8959
rect 5215 8925 5224 8959
rect 5172 8916 5224 8925
rect 7104 8916 7156 8968
rect 8208 8916 8260 8968
rect 15200 8984 15252 9036
rect 16580 9027 16632 9036
rect 16580 8993 16589 9027
rect 16589 8993 16623 9027
rect 16623 8993 16632 9027
rect 16580 8984 16632 8993
rect 8484 8848 8536 8900
rect 3516 8780 3568 8832
rect 13268 8959 13320 8968
rect 10876 8848 10928 8900
rect 13268 8925 13277 8959
rect 13277 8925 13311 8959
rect 13311 8925 13320 8959
rect 13268 8916 13320 8925
rect 14188 8959 14240 8968
rect 14188 8925 14197 8959
rect 14197 8925 14231 8959
rect 14231 8925 14240 8959
rect 14188 8916 14240 8925
rect 17408 8984 17460 9036
rect 17868 9027 17920 9036
rect 17868 8993 17877 9027
rect 17877 8993 17911 9027
rect 17911 8993 17920 9027
rect 17868 8984 17920 8993
rect 18604 8916 18656 8968
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 3700 8619 3752 8628
rect 3700 8585 3709 8619
rect 3709 8585 3743 8619
rect 3743 8585 3752 8619
rect 3700 8576 3752 8585
rect 7104 8619 7156 8628
rect 7104 8585 7113 8619
rect 7113 8585 7147 8619
rect 7147 8585 7156 8619
rect 7104 8576 7156 8585
rect 8484 8576 8536 8628
rect 3976 8508 4028 8560
rect 2228 8483 2280 8492
rect 2228 8449 2237 8483
rect 2237 8449 2271 8483
rect 2271 8449 2280 8483
rect 2228 8440 2280 8449
rect 3792 8440 3844 8492
rect 4344 8483 4396 8492
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 5264 8483 5316 8492
rect 5264 8449 5273 8483
rect 5273 8449 5307 8483
rect 5307 8449 5316 8483
rect 5264 8440 5316 8449
rect 7380 8440 7432 8492
rect 7748 8483 7800 8492
rect 7748 8449 7757 8483
rect 7757 8449 7791 8483
rect 7791 8449 7800 8483
rect 7748 8440 7800 8449
rect 9404 8508 9456 8560
rect 11704 8508 11756 8560
rect 11980 8508 12032 8560
rect 8944 8372 8996 8424
rect 9772 8440 9824 8492
rect 10876 8372 10928 8424
rect 8392 8304 8444 8356
rect 11796 8304 11848 8356
rect 14556 8440 14608 8492
rect 19432 8576 19484 8628
rect 18052 8508 18104 8560
rect 19340 8415 19392 8424
rect 19340 8381 19349 8415
rect 19349 8381 19383 8415
rect 19383 8381 19392 8415
rect 19340 8372 19392 8381
rect 4068 8279 4120 8288
rect 4068 8245 4077 8279
rect 4077 8245 4111 8279
rect 4111 8245 4120 8279
rect 4068 8236 4120 8245
rect 7656 8236 7708 8288
rect 11152 8279 11204 8288
rect 11152 8245 11161 8279
rect 11161 8245 11195 8279
rect 11195 8245 11204 8279
rect 11152 8236 11204 8245
rect 13820 8279 13872 8288
rect 13820 8245 13829 8279
rect 13829 8245 13863 8279
rect 13863 8245 13872 8279
rect 13820 8236 13872 8245
rect 14832 8304 14884 8356
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 2872 8032 2924 8084
rect 3976 8032 4028 8084
rect 5172 7964 5224 8016
rect 7288 8032 7340 8084
rect 8944 8032 8996 8084
rect 15292 8075 15344 8084
rect 15292 8041 15301 8075
rect 15301 8041 15335 8075
rect 15335 8041 15344 8075
rect 15292 8032 15344 8041
rect 11152 7964 11204 8016
rect 12348 7964 12400 8016
rect 1860 7896 1912 7948
rect 7564 7939 7616 7948
rect 7564 7905 7573 7939
rect 7573 7905 7607 7939
rect 7607 7905 7616 7939
rect 7564 7896 7616 7905
rect 10048 7939 10100 7948
rect 10048 7905 10057 7939
rect 10057 7905 10091 7939
rect 10091 7905 10100 7939
rect 10048 7896 10100 7905
rect 11888 7896 11940 7948
rect 2780 7871 2832 7880
rect 2780 7837 2789 7871
rect 2789 7837 2823 7871
rect 2823 7837 2832 7871
rect 4988 7871 5040 7880
rect 2780 7828 2832 7837
rect 4988 7837 4997 7871
rect 4997 7837 5031 7871
rect 5031 7837 5040 7871
rect 4988 7828 5040 7837
rect 6092 7828 6144 7880
rect 7748 7871 7800 7880
rect 7748 7837 7757 7871
rect 7757 7837 7791 7871
rect 7791 7837 7800 7871
rect 7748 7828 7800 7837
rect 9864 7828 9916 7880
rect 10692 7828 10744 7880
rect 13820 7896 13872 7948
rect 19340 7964 19392 8016
rect 12072 7828 12124 7880
rect 7932 7692 7984 7744
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 4988 7488 5040 7540
rect 5172 7488 5224 7540
rect 8208 7531 8260 7540
rect 8208 7497 8217 7531
rect 8217 7497 8251 7531
rect 8251 7497 8260 7531
rect 8208 7488 8260 7497
rect 9864 7531 9916 7540
rect 9864 7497 9873 7531
rect 9873 7497 9907 7531
rect 9907 7497 9916 7531
rect 9864 7488 9916 7497
rect 16580 7488 16632 7540
rect 6828 7395 6880 7404
rect 2780 7284 2832 7336
rect 6828 7361 6837 7395
rect 6837 7361 6871 7395
rect 6871 7361 6880 7395
rect 6828 7352 6880 7361
rect 9496 7352 9548 7404
rect 11704 7352 11756 7404
rect 13820 7352 13872 7404
rect 7932 7284 7984 7336
rect 10232 7327 10284 7336
rect 10232 7293 10241 7327
rect 10241 7293 10275 7327
rect 10275 7293 10284 7327
rect 10232 7284 10284 7293
rect 10784 7284 10836 7336
rect 14188 7284 14240 7336
rect 2412 7216 2464 7268
rect 4344 7216 4396 7268
rect 7748 7216 7800 7268
rect 2688 7148 2740 7200
rect 10324 7191 10376 7200
rect 10324 7157 10333 7191
rect 10333 7157 10367 7191
rect 10367 7157 10376 7191
rect 10324 7148 10376 7157
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 1860 6987 1912 6996
rect 1860 6953 1869 6987
rect 1869 6953 1903 6987
rect 1903 6953 1912 6987
rect 1860 6944 1912 6953
rect 3884 6944 3936 6996
rect 9036 6944 9088 6996
rect 12256 6944 12308 6996
rect 2228 6919 2280 6928
rect 2228 6885 2237 6919
rect 2237 6885 2271 6919
rect 2271 6885 2280 6919
rect 2228 6876 2280 6885
rect 8208 6876 8260 6928
rect 10692 6876 10744 6928
rect 2320 6851 2372 6860
rect 2320 6817 2329 6851
rect 2329 6817 2363 6851
rect 2363 6817 2372 6851
rect 2320 6808 2372 6817
rect 2412 6783 2464 6792
rect 2412 6749 2421 6783
rect 2421 6749 2455 6783
rect 2455 6749 2464 6783
rect 2412 6740 2464 6749
rect 2504 6740 2556 6792
rect 5172 6783 5224 6792
rect 5172 6749 5181 6783
rect 5181 6749 5215 6783
rect 5215 6749 5224 6783
rect 5172 6740 5224 6749
rect 4068 6672 4120 6724
rect 6828 6740 6880 6792
rect 10508 6783 10560 6792
rect 10508 6749 10517 6783
rect 10517 6749 10551 6783
rect 10551 6749 10560 6783
rect 10508 6740 10560 6749
rect 19892 6672 19944 6724
rect 5080 6604 5132 6656
rect 8300 6647 8352 6656
rect 8300 6613 8309 6647
rect 8309 6613 8343 6647
rect 8343 6613 8352 6647
rect 8300 6604 8352 6613
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 2412 6400 2464 6452
rect 8300 6400 8352 6452
rect 5080 6307 5132 6316
rect 5080 6273 5089 6307
rect 5089 6273 5123 6307
rect 5123 6273 5132 6307
rect 5080 6264 5132 6273
rect 6552 6264 6604 6316
rect 10508 6400 10560 6452
rect 10692 6400 10744 6452
rect 19708 6443 19760 6452
rect 12348 6332 12400 6384
rect 2688 6239 2740 6248
rect 2688 6205 2722 6239
rect 2722 6205 2740 6239
rect 6828 6239 6880 6248
rect 2688 6196 2740 6205
rect 6828 6205 6837 6239
rect 6837 6205 6871 6239
rect 6871 6205 6880 6239
rect 6828 6196 6880 6205
rect 9496 6239 9548 6248
rect 9496 6205 9530 6239
rect 9530 6205 9548 6239
rect 9496 6196 9548 6205
rect 19708 6409 19717 6443
rect 19717 6409 19751 6443
rect 19751 6409 19760 6443
rect 19708 6400 19760 6409
rect 2780 6128 2832 6180
rect 3976 6128 4028 6180
rect 12348 6128 12400 6180
rect 3792 6103 3844 6112
rect 3792 6069 3801 6103
rect 3801 6069 3835 6103
rect 3835 6069 3844 6103
rect 3792 6060 3844 6069
rect 4344 6060 4396 6112
rect 4988 6103 5040 6112
rect 4988 6069 4997 6103
rect 4997 6069 5031 6103
rect 5031 6069 5040 6103
rect 4988 6060 5040 6069
rect 8300 6060 8352 6112
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 2504 5856 2556 5908
rect 6552 5899 6604 5908
rect 6552 5865 6561 5899
rect 6561 5865 6595 5899
rect 6595 5865 6604 5899
rect 6552 5856 6604 5865
rect 7564 5856 7616 5908
rect 10324 5856 10376 5908
rect 3148 5788 3200 5840
rect 5172 5788 5224 5840
rect 13360 5856 13412 5908
rect 20996 5856 21048 5908
rect 11244 5788 11296 5840
rect 2688 5720 2740 5772
rect 7472 5720 7524 5772
rect 8300 5720 8352 5772
rect 11060 5763 11112 5772
rect 3792 5652 3844 5704
rect 9680 5695 9732 5704
rect 2780 5584 2832 5636
rect 3700 5584 3752 5636
rect 9680 5661 9689 5695
rect 9689 5661 9723 5695
rect 9723 5661 9732 5695
rect 9680 5652 9732 5661
rect 11060 5729 11069 5763
rect 11069 5729 11103 5763
rect 11103 5729 11112 5763
rect 11060 5720 11112 5729
rect 12348 5720 12400 5772
rect 4068 5516 4120 5568
rect 12348 5516 12400 5568
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 4344 5312 4396 5364
rect 5172 5312 5224 5364
rect 3700 5219 3752 5228
rect 3700 5185 3709 5219
rect 3709 5185 3743 5219
rect 3743 5185 3752 5219
rect 3700 5176 3752 5185
rect 3792 5108 3844 5160
rect 1768 5040 1820 5092
rect 3240 5040 3292 5092
rect 5540 5176 5592 5228
rect 6644 5176 6696 5228
rect 6828 5176 6880 5228
rect 8300 5151 8352 5160
rect 5264 4972 5316 5024
rect 8300 5117 8334 5151
rect 8334 5117 8352 5151
rect 8300 5108 8352 5117
rect 9496 5312 9548 5364
rect 10048 5312 10100 5364
rect 19616 5355 19668 5364
rect 19616 5321 19625 5355
rect 19625 5321 19659 5355
rect 19659 5321 19668 5355
rect 19616 5312 19668 5321
rect 20904 5312 20956 5364
rect 9680 5108 9732 5160
rect 20536 5151 20588 5160
rect 20536 5117 20545 5151
rect 20545 5117 20579 5151
rect 20579 5117 20588 5151
rect 20536 5108 20588 5117
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 1584 4768 1636 4820
rect 4988 4768 5040 4820
rect 5264 4811 5316 4820
rect 5264 4777 5273 4811
rect 5273 4777 5307 4811
rect 5307 4777 5316 4811
rect 5264 4768 5316 4777
rect 12440 4768 12492 4820
rect 20536 4768 20588 4820
rect 4068 4700 4120 4752
rect 12348 4700 12400 4752
rect 1768 4675 1820 4684
rect 1768 4641 1777 4675
rect 1777 4641 1811 4675
rect 1811 4641 1820 4675
rect 1768 4632 1820 4641
rect 5172 4632 5224 4684
rect 4160 4564 4212 4616
rect 5356 4607 5408 4616
rect 5356 4573 5365 4607
rect 5365 4573 5399 4607
rect 5399 4573 5408 4607
rect 5356 4564 5408 4573
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 3516 4088 3568 4140
rect 7656 4088 7708 4140
rect 4068 4020 4120 4072
rect 5724 3952 5776 4004
rect 6736 3952 6788 4004
rect 20812 3884 20864 3936
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 4068 2592 4120 2644
rect 5540 2592 5592 2644
rect 3056 2456 3108 2508
rect 10232 2456 10284 2508
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 3424 1300 3476 1352
rect 11060 1300 11112 1352
<< metal2 >>
rect 202 22520 258 23000
rect 662 22520 718 23000
rect 1122 22520 1178 23000
rect 1582 22520 1638 23000
rect 2042 22520 2098 23000
rect 2502 22520 2558 23000
rect 2962 22520 3018 23000
rect 3422 22520 3478 23000
rect 3790 22672 3846 22681
rect 3790 22607 3846 22616
rect 216 18154 244 22520
rect 204 18148 256 18154
rect 204 18090 256 18096
rect 676 12714 704 22520
rect 1136 13462 1164 22520
rect 1596 21298 1624 22520
rect 1596 21270 1992 21298
rect 1858 21176 1914 21185
rect 1858 21111 1914 21120
rect 1400 19916 1452 19922
rect 1400 19858 1452 19864
rect 1412 17814 1440 19858
rect 1584 19712 1636 19718
rect 1584 19654 1636 19660
rect 1400 17808 1452 17814
rect 1400 17750 1452 17756
rect 1596 16697 1624 19654
rect 1768 19168 1820 19174
rect 1768 19110 1820 19116
rect 1582 16688 1638 16697
rect 1582 16623 1638 16632
rect 1780 16153 1808 19110
rect 1766 16144 1822 16153
rect 1766 16079 1822 16088
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 1124 13456 1176 13462
rect 1124 13398 1176 13404
rect 1582 13152 1638 13161
rect 1582 13087 1638 13096
rect 664 12708 716 12714
rect 664 12650 716 12656
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10606 1440 11086
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1596 4826 1624 13087
rect 1688 12306 1716 13806
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 1872 11898 1900 21111
rect 1964 18290 1992 21270
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 1950 18184 2006 18193
rect 1950 18119 2006 18128
rect 1964 18086 1992 18119
rect 2056 18086 2084 22520
rect 2136 20392 2188 20398
rect 2136 20334 2188 20340
rect 2148 19825 2176 20334
rect 2134 19816 2190 19825
rect 2134 19751 2190 19760
rect 2516 19242 2544 22520
rect 2976 20074 3004 22520
rect 3240 20256 3292 20262
rect 3240 20198 3292 20204
rect 2976 20046 3188 20074
rect 2964 19916 3016 19922
rect 2964 19858 3016 19864
rect 2872 19304 2924 19310
rect 2872 19246 2924 19252
rect 2504 19236 2556 19242
rect 2504 19178 2556 19184
rect 2780 18828 2832 18834
rect 2780 18770 2832 18776
rect 2792 18329 2820 18770
rect 2778 18320 2834 18329
rect 2778 18255 2834 18264
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 2044 18080 2096 18086
rect 2044 18022 2096 18028
rect 2780 18080 2832 18086
rect 2780 18022 2832 18028
rect 2792 17921 2820 18022
rect 2778 17912 2834 17921
rect 2504 17876 2556 17882
rect 2778 17847 2834 17856
rect 2504 17818 2556 17824
rect 2228 17740 2280 17746
rect 2228 17682 2280 17688
rect 2240 16794 2268 17682
rect 2412 17672 2464 17678
rect 2412 17614 2464 17620
rect 2228 16788 2280 16794
rect 2228 16730 2280 16736
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1964 14113 1992 14758
rect 1950 14104 2006 14113
rect 1950 14039 2006 14048
rect 1952 13320 2004 13326
rect 1952 13262 2004 13268
rect 1964 12782 1992 13262
rect 1952 12776 2004 12782
rect 1952 12718 2004 12724
rect 2320 12708 2372 12714
rect 2320 12650 2372 12656
rect 2044 12640 2096 12646
rect 2042 12608 2044 12617
rect 2096 12608 2098 12617
rect 2042 12543 2098 12552
rect 1860 11892 1912 11898
rect 1860 11834 1912 11840
rect 2042 11656 2098 11665
rect 2042 11591 2098 11600
rect 2056 10674 2084 11591
rect 2332 11286 2360 12650
rect 2424 11694 2452 17614
rect 2516 17202 2544 17818
rect 2504 17196 2556 17202
rect 2504 17138 2556 17144
rect 2884 16114 2912 19246
rect 2976 18426 3004 19858
rect 3056 18624 3108 18630
rect 3056 18566 3108 18572
rect 2964 18420 3016 18426
rect 2964 18362 3016 18368
rect 3068 18290 3096 18566
rect 3160 18426 3188 20046
rect 3252 18601 3280 20198
rect 3238 18592 3294 18601
rect 3238 18527 3294 18536
rect 3148 18420 3200 18426
rect 3148 18362 3200 18368
rect 2964 18284 3016 18290
rect 2964 18226 3016 18232
rect 3056 18284 3108 18290
rect 3056 18226 3108 18232
rect 2976 18154 3004 18226
rect 3330 18184 3386 18193
rect 2964 18148 3016 18154
rect 3330 18119 3332 18128
rect 2964 18090 3016 18096
rect 3384 18119 3386 18128
rect 3332 18090 3384 18096
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 2872 16108 2924 16114
rect 2872 16050 2924 16056
rect 3056 15564 3108 15570
rect 3056 15506 3108 15512
rect 3068 15162 3096 15506
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 2964 14476 3016 14482
rect 2964 14418 3016 14424
rect 2872 14408 2924 14414
rect 2872 14350 2924 14356
rect 2884 13530 2912 14350
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2792 11898 2820 13330
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 2884 12170 2912 13262
rect 2976 12986 3004 14418
rect 3056 13796 3108 13802
rect 3056 13738 3108 13744
rect 3068 13326 3096 13738
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 3068 12850 3096 13262
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 2964 12776 3016 12782
rect 2964 12718 3016 12724
rect 2976 12374 3004 12718
rect 3068 12442 3096 12786
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 2964 12368 3016 12374
rect 2964 12310 3016 12316
rect 2872 12164 2924 12170
rect 2872 12106 2924 12112
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2320 11280 2372 11286
rect 2320 11222 2372 11228
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 2148 10674 2176 11086
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2148 10266 2176 10610
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 2148 9518 2176 10202
rect 2136 9512 2188 9518
rect 2136 9454 2188 9460
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 2240 8498 2268 8978
rect 2228 8492 2280 8498
rect 2228 8434 2280 8440
rect 1860 7948 1912 7954
rect 1860 7890 1912 7896
rect 1872 7002 1900 7890
rect 1860 6996 1912 7002
rect 1860 6938 1912 6944
rect 2228 6928 2280 6934
rect 2228 6870 2280 6876
rect 2240 6633 2268 6870
rect 2332 6866 2360 11222
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2792 10810 2820 11154
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2412 10124 2464 10130
rect 2412 10066 2464 10072
rect 2424 9654 2452 10066
rect 2412 9648 2464 9654
rect 2412 9590 2464 9596
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2884 8090 2912 8910
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 2780 7880 2832 7886
rect 2700 7828 2780 7834
rect 2700 7822 2832 7828
rect 2700 7806 2820 7822
rect 2412 7268 2464 7274
rect 2412 7210 2464 7216
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2424 6798 2452 7210
rect 2700 7206 2728 7806
rect 2780 7336 2832 7342
rect 2780 7278 2832 7284
rect 2688 7200 2740 7206
rect 2688 7142 2740 7148
rect 2412 6792 2464 6798
rect 2412 6734 2464 6740
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2226 6624 2282 6633
rect 2226 6559 2282 6568
rect 2424 6458 2452 6734
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2516 5914 2544 6734
rect 2700 6254 2728 7142
rect 2688 6248 2740 6254
rect 2688 6190 2740 6196
rect 2792 6186 2820 7278
rect 2780 6180 2832 6186
rect 2780 6122 2832 6128
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 1768 5092 1820 5098
rect 1768 5034 1820 5040
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 1780 4690 1808 5034
rect 1768 4684 1820 4690
rect 1768 4626 1820 4632
rect 2700 241 2728 5714
rect 2792 5642 2820 6122
rect 3160 5846 3188 17478
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3252 13734 3280 14350
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3330 13696 3386 13705
rect 3252 12782 3280 13670
rect 3330 13631 3386 13640
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 3344 9178 3372 13631
rect 3436 11694 3464 22520
rect 3514 21584 3570 21593
rect 3514 21519 3570 21528
rect 3528 21146 3556 21519
rect 3516 21140 3568 21146
rect 3516 21082 3568 21088
rect 3804 21010 3832 22607
rect 3882 22520 3938 23000
rect 4342 22520 4398 23000
rect 4894 22520 4950 23000
rect 5354 22520 5410 23000
rect 5814 22520 5870 23000
rect 6274 22520 6330 23000
rect 6734 22520 6790 23000
rect 7194 22520 7250 23000
rect 7654 22520 7710 23000
rect 8114 22520 8170 23000
rect 8574 22520 8630 23000
rect 9034 22520 9090 23000
rect 9586 22520 9642 23000
rect 10046 22520 10102 23000
rect 10506 22520 10562 23000
rect 10966 22520 11022 23000
rect 11426 22520 11482 23000
rect 11886 22520 11942 23000
rect 12346 22520 12402 23000
rect 12806 22520 12862 23000
rect 13266 22520 13322 23000
rect 13726 22520 13782 23000
rect 14278 22520 14334 23000
rect 14738 22520 14794 23000
rect 15198 22520 15254 23000
rect 15658 22520 15714 23000
rect 16118 22520 16174 23000
rect 16578 22520 16634 23000
rect 17038 22520 17094 23000
rect 17498 22520 17554 23000
rect 17958 22520 18014 23000
rect 18418 22520 18474 23000
rect 18970 22520 19026 23000
rect 19430 22520 19486 23000
rect 19890 22520 19946 23000
rect 20350 22520 20406 23000
rect 20810 22520 20866 23000
rect 21270 22520 21326 23000
rect 21730 22520 21786 23000
rect 22190 22520 22246 23000
rect 22650 22520 22706 23000
rect 3792 21004 3844 21010
rect 3792 20946 3844 20952
rect 3790 20088 3846 20097
rect 3790 20023 3846 20032
rect 3608 19916 3660 19922
rect 3608 19858 3660 19864
rect 3516 19712 3568 19718
rect 3516 19654 3568 19660
rect 3528 17105 3556 19654
rect 3514 17096 3570 17105
rect 3514 17031 3570 17040
rect 3620 16658 3648 19858
rect 3804 19514 3832 20023
rect 3792 19508 3844 19514
rect 3792 19450 3844 19456
rect 3700 19236 3752 19242
rect 3700 19178 3752 19184
rect 3608 16652 3660 16658
rect 3608 16594 3660 16600
rect 3514 14648 3570 14657
rect 3514 14583 3516 14592
rect 3568 14583 3570 14592
rect 3516 14554 3568 14560
rect 3608 12300 3660 12306
rect 3608 12242 3660 12248
rect 3620 11762 3648 12242
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3712 11558 3740 19178
rect 3896 17542 3924 22520
rect 4066 22128 4122 22137
rect 4066 22063 4122 22072
rect 4080 20806 4108 22063
rect 4068 20800 4120 20806
rect 4068 20742 4120 20748
rect 3974 20632 4030 20641
rect 3974 20567 3976 20576
rect 4028 20567 4030 20576
rect 3976 20538 4028 20544
rect 4068 20528 4120 20534
rect 4068 20470 4120 20476
rect 3974 19680 4030 19689
rect 3974 19615 4030 19624
rect 3988 19514 4016 19615
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 4080 18834 4108 20470
rect 4252 20052 4304 20058
rect 4252 19994 4304 20000
rect 4160 19168 4212 19174
rect 4264 19145 4292 19994
rect 4356 19938 4384 22520
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 4356 19910 4844 19938
rect 4344 19712 4396 19718
rect 4344 19654 4396 19660
rect 4356 19310 4384 19654
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 4344 19304 4396 19310
rect 4344 19246 4396 19252
rect 4160 19110 4212 19116
rect 4250 19136 4306 19145
rect 4068 18828 4120 18834
rect 4068 18770 4120 18776
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 4080 17785 4108 18362
rect 4172 18290 4200 19110
rect 4250 19071 4306 19080
rect 4356 18766 4384 19246
rect 4528 18896 4580 18902
rect 4526 18864 4528 18873
rect 4580 18864 4582 18873
rect 4526 18799 4582 18808
rect 4344 18760 4396 18766
rect 4344 18702 4396 18708
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 4160 18284 4212 18290
rect 4160 18226 4212 18232
rect 4066 17776 4122 17785
rect 4172 17746 4200 18226
rect 4816 18154 4844 19910
rect 4908 18426 4936 22520
rect 4988 19848 5040 19854
rect 4988 19790 5040 19796
rect 5000 18766 5028 19790
rect 4988 18760 5040 18766
rect 4988 18702 5040 18708
rect 4896 18420 4948 18426
rect 4896 18362 4948 18368
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 4712 18148 4764 18154
rect 4712 18090 4764 18096
rect 4804 18148 4856 18154
rect 4804 18090 4856 18096
rect 4344 18080 4396 18086
rect 4724 18057 4752 18090
rect 4344 18022 4396 18028
rect 4710 18048 4766 18057
rect 4066 17711 4122 17720
rect 4160 17740 4212 17746
rect 4160 17682 4212 17688
rect 3974 17640 4030 17649
rect 3974 17575 4030 17584
rect 3884 17536 3936 17542
rect 3884 17478 3936 17484
rect 3988 17338 4016 17575
rect 4068 17536 4120 17542
rect 4068 17478 4120 17484
rect 3976 17332 4028 17338
rect 3976 17274 4028 17280
rect 4080 17218 4108 17478
rect 3988 17202 4108 17218
rect 3976 17196 4108 17202
rect 4028 17190 4108 17196
rect 3976 17138 4028 17144
rect 4356 16794 4384 18022
rect 4710 17983 4766 17992
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4344 16788 4396 16794
rect 4344 16730 4396 16736
rect 4724 16590 4752 16934
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 4712 16584 4764 16590
rect 4712 16526 4764 16532
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 3792 16108 3844 16114
rect 3792 16050 3844 16056
rect 3804 14074 3832 16050
rect 4080 15609 4108 16390
rect 4356 16046 4384 16526
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 4344 16040 4396 16046
rect 4344 15982 4396 15988
rect 4066 15600 4122 15609
rect 4066 15535 4122 15544
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 3882 15192 3938 15201
rect 3882 15127 3938 15136
rect 4068 15156 4120 15162
rect 3896 14346 3924 15127
rect 4068 15098 4120 15104
rect 4080 14482 4108 15098
rect 4068 14476 4120 14482
rect 4068 14418 4120 14424
rect 3884 14340 3936 14346
rect 3884 14282 3936 14288
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4172 14074 4200 14214
rect 3792 14068 3844 14074
rect 3792 14010 3844 14016
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 3804 13870 3832 14010
rect 3792 13864 3844 13870
rect 3792 13806 3844 13812
rect 3804 13394 3832 13806
rect 3792 13388 3844 13394
rect 3792 13330 3844 13336
rect 4264 12782 4292 15438
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 4804 13796 4856 13802
rect 4804 13738 4856 13744
rect 4816 13190 4844 13738
rect 4804 13184 4856 13190
rect 4804 13126 4856 13132
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 4816 12986 4844 13126
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4252 12776 4304 12782
rect 4252 12718 4304 12724
rect 4068 12368 4120 12374
rect 4068 12310 4120 12316
rect 4080 12209 4108 12310
rect 4908 12306 4936 18158
rect 5000 17542 5028 18702
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 4988 17536 5040 17542
rect 4988 17478 5040 17484
rect 5000 17270 5028 17478
rect 4988 17264 5040 17270
rect 4988 17206 5040 17212
rect 5172 15904 5224 15910
rect 5172 15846 5224 15852
rect 5184 15638 5212 15846
rect 5172 15632 5224 15638
rect 5172 15574 5224 15580
rect 5184 15026 5212 15574
rect 5172 15020 5224 15026
rect 5172 14962 5224 14968
rect 4988 14952 5040 14958
rect 4988 14894 5040 14900
rect 5000 14618 5028 14894
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 5276 13530 5304 18022
rect 5368 14958 5396 22520
rect 5448 20528 5500 20534
rect 5448 20470 5500 20476
rect 5460 19990 5488 20470
rect 5632 20256 5684 20262
rect 5632 20198 5684 20204
rect 5724 20256 5776 20262
rect 5724 20198 5776 20204
rect 5644 19990 5672 20198
rect 5448 19984 5500 19990
rect 5448 19926 5500 19932
rect 5632 19984 5684 19990
rect 5632 19926 5684 19932
rect 5540 19304 5592 19310
rect 5538 19272 5540 19281
rect 5592 19272 5594 19281
rect 5736 19242 5764 20198
rect 5538 19207 5594 19216
rect 5724 19236 5776 19242
rect 5724 19178 5776 19184
rect 5828 18986 5856 22520
rect 6092 21140 6144 21146
rect 6092 21082 6144 21088
rect 5908 20460 5960 20466
rect 5908 20402 5960 20408
rect 5920 19922 5948 20402
rect 5908 19916 5960 19922
rect 5908 19858 5960 19864
rect 5908 19372 5960 19378
rect 5908 19314 5960 19320
rect 5644 18958 5856 18986
rect 5448 18284 5500 18290
rect 5448 18226 5500 18232
rect 5460 17542 5488 18226
rect 5644 18222 5672 18958
rect 5724 18896 5776 18902
rect 5920 18850 5948 19314
rect 5998 19272 6054 19281
rect 5998 19207 6054 19216
rect 6012 19174 6040 19207
rect 6000 19168 6052 19174
rect 6000 19110 6052 19116
rect 5776 18844 5948 18850
rect 5724 18838 5948 18844
rect 5736 18822 5948 18838
rect 5632 18216 5684 18222
rect 5632 18158 5684 18164
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 5460 17134 5488 17478
rect 5448 17128 5500 17134
rect 5448 17070 5500 17076
rect 5552 17066 5580 18022
rect 5630 17912 5686 17921
rect 5630 17847 5686 17856
rect 5540 17060 5592 17066
rect 5540 17002 5592 17008
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5460 16658 5488 16934
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5540 15632 5592 15638
rect 5540 15574 5592 15580
rect 5356 14952 5408 14958
rect 5356 14894 5408 14900
rect 5552 14822 5580 15574
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 4344 12300 4396 12306
rect 4344 12242 4396 12248
rect 4896 12300 4948 12306
rect 4896 12242 4948 12248
rect 4066 12200 4122 12209
rect 4066 12135 4122 12144
rect 4356 11778 4384 12242
rect 4804 12164 4856 12170
rect 4804 12106 4856 12112
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 4356 11750 4476 11778
rect 4448 11676 4476 11750
rect 4620 11688 4672 11694
rect 4448 11648 4620 11676
rect 3792 11620 3844 11626
rect 3792 11562 3844 11568
rect 4344 11620 4396 11626
rect 4344 11562 4396 11568
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3436 10470 3464 11494
rect 3804 10606 3832 11562
rect 4252 11280 4304 11286
rect 4080 11240 4252 11268
rect 4080 11121 4108 11240
rect 4252 11222 4304 11228
rect 4066 11112 4122 11121
rect 4066 11047 4122 11056
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 3884 11008 3936 11014
rect 3884 10950 3936 10956
rect 3896 10674 3924 10950
rect 4172 10674 4200 11018
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 3792 10600 3844 10606
rect 3792 10542 3844 10548
rect 3424 10464 3476 10470
rect 3424 10406 3476 10412
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3712 9625 3740 9862
rect 3698 9616 3754 9625
rect 3698 9551 3754 9560
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3700 8968 3752 8974
rect 3700 8910 3752 8916
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3528 8673 3556 8774
rect 3514 8664 3570 8673
rect 3712 8634 3740 8910
rect 3514 8599 3570 8608
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 3804 8498 3832 10542
rect 3896 10198 3924 10610
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3884 10192 3936 10198
rect 3884 10134 3936 10140
rect 3988 8566 4016 10406
rect 4080 10169 4108 10542
rect 4066 10160 4122 10169
rect 4066 10095 4122 10104
rect 4356 10062 4384 11562
rect 4540 11218 4568 11648
rect 4620 11630 4672 11636
rect 4816 11354 4844 12106
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 4894 10840 4950 10849
rect 4894 10775 4950 10784
rect 4908 10742 4936 10775
rect 4896 10736 4948 10742
rect 4896 10678 4948 10684
rect 4988 10192 5040 10198
rect 4988 10134 5040 10140
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4356 9722 4384 9998
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 5000 9722 5028 10134
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4988 9716 5040 9722
rect 4988 9658 5040 9664
rect 4068 9444 4120 9450
rect 4068 9386 4120 9392
rect 4080 9217 4108 9386
rect 4066 9208 4122 9217
rect 4356 9178 4384 9658
rect 5276 9194 5304 13466
rect 5644 12646 5672 17847
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5736 13734 5764 13874
rect 5724 13728 5776 13734
rect 5724 13670 5776 13676
rect 5736 13462 5764 13670
rect 5724 13456 5776 13462
rect 5724 13398 5776 13404
rect 6104 12986 6132 21082
rect 6184 20528 6236 20534
rect 6184 20470 6236 20476
rect 6196 20398 6224 20470
rect 6184 20392 6236 20398
rect 6184 20334 6236 20340
rect 6288 18970 6316 22520
rect 6368 19780 6420 19786
rect 6368 19722 6420 19728
rect 6380 19378 6408 19722
rect 6368 19372 6420 19378
rect 6368 19314 6420 19320
rect 6748 19310 6776 22520
rect 6840 20454 7052 20482
rect 6840 20398 6868 20454
rect 6828 20392 6880 20398
rect 6828 20334 6880 20340
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 6736 19304 6788 19310
rect 6736 19246 6788 19252
rect 6840 18970 6868 19858
rect 6918 19816 6974 19825
rect 6918 19751 6974 19760
rect 6276 18964 6328 18970
rect 6276 18906 6328 18912
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 6828 18828 6880 18834
rect 6828 18770 6880 18776
rect 6840 17678 6868 18770
rect 6932 18698 6960 19751
rect 6920 18692 6972 18698
rect 6920 18634 6972 18640
rect 6920 18148 6972 18154
rect 6920 18090 6972 18096
rect 6828 17672 6880 17678
rect 6828 17614 6880 17620
rect 6840 17270 6868 17614
rect 6828 17264 6880 17270
rect 6828 17206 6880 17212
rect 6840 17134 6868 17206
rect 6184 17128 6236 17134
rect 6184 17070 6236 17076
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6196 14822 6224 17070
rect 6552 15632 6604 15638
rect 6552 15574 6604 15580
rect 6460 15360 6512 15366
rect 6460 15302 6512 15308
rect 6472 15094 6500 15302
rect 6460 15088 6512 15094
rect 6460 15030 6512 15036
rect 6472 14958 6500 15030
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 6460 14952 6512 14958
rect 6460 14894 6512 14900
rect 6184 14816 6236 14822
rect 6184 14758 6236 14764
rect 6196 13870 6224 14758
rect 6184 13864 6236 13870
rect 6184 13806 6236 13812
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5552 11898 5580 12174
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5540 11280 5592 11286
rect 5540 11222 5592 11228
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5460 9518 5488 10610
rect 5552 10130 5580 11222
rect 5644 11014 5672 12038
rect 6196 11626 6224 13126
rect 6380 12986 6408 14894
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 6184 11620 6236 11626
rect 6184 11562 6236 11568
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5920 11150 5948 11494
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 6104 9654 6132 11086
rect 6288 10538 6316 11086
rect 6380 10606 6408 12922
rect 6564 12322 6592 15574
rect 6840 15502 6868 17070
rect 6932 16794 6960 18090
rect 7024 17882 7052 20454
rect 7104 20256 7156 20262
rect 7104 20198 7156 20204
rect 7116 20058 7144 20198
rect 7208 20058 7236 22520
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 7196 20052 7248 20058
rect 7196 19994 7248 20000
rect 7668 19802 7696 22520
rect 8128 20534 8156 22520
rect 8116 20528 8168 20534
rect 8116 20470 8168 20476
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 7576 19774 7696 19802
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 7840 19780 7892 19786
rect 7196 18624 7248 18630
rect 7196 18566 7248 18572
rect 7208 18222 7236 18566
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 7196 18216 7248 18222
rect 7196 18158 7248 18164
rect 7286 18048 7342 18057
rect 7286 17983 7342 17992
rect 7012 17876 7064 17882
rect 7012 17818 7064 17824
rect 7194 17776 7250 17785
rect 7194 17711 7250 17720
rect 7012 16992 7064 16998
rect 7012 16934 7064 16940
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 7024 16658 7052 16934
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6828 15496 6880 15502
rect 6828 15438 6880 15444
rect 6932 14498 6960 15846
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 7116 15026 7144 15438
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 6748 14482 6960 14498
rect 6736 14476 6960 14482
rect 6788 14470 6960 14476
rect 6736 14418 6788 14424
rect 6644 14408 6696 14414
rect 7208 14362 7236 17711
rect 7300 15042 7328 17983
rect 7484 17746 7512 18226
rect 7472 17740 7524 17746
rect 7472 17682 7524 17688
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 7380 16652 7432 16658
rect 7380 16594 7432 16600
rect 7392 15978 7420 16594
rect 7484 16590 7512 17002
rect 7576 16794 7604 19774
rect 7840 19722 7892 19728
rect 7656 19712 7708 19718
rect 7656 19654 7708 19660
rect 7668 18970 7696 19654
rect 7748 19304 7800 19310
rect 7748 19246 7800 19252
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 7760 18834 7788 19246
rect 7852 19242 7880 19722
rect 8220 19242 8248 19790
rect 7840 19236 7892 19242
rect 7840 19178 7892 19184
rect 8208 19236 8260 19242
rect 8208 19178 8260 19184
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 8220 17882 8248 19178
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 8312 18873 8340 18906
rect 8298 18864 8354 18873
rect 8298 18799 8354 18808
rect 8588 18358 8616 22520
rect 8760 20596 8812 20602
rect 8760 20538 8812 20544
rect 8944 20596 8996 20602
rect 8944 20538 8996 20544
rect 8772 20330 8800 20538
rect 8668 20324 8720 20330
rect 8668 20266 8720 20272
rect 8760 20324 8812 20330
rect 8760 20266 8812 20272
rect 8680 19174 8708 20266
rect 8956 19922 8984 20538
rect 8944 19916 8996 19922
rect 8944 19858 8996 19864
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 8576 18352 8628 18358
rect 8576 18294 8628 18300
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 8208 17876 8260 17882
rect 8208 17818 8260 17824
rect 8208 17740 8260 17746
rect 8208 17682 8260 17688
rect 8220 17338 8248 17682
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 7760 16794 7788 17274
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 7380 15972 7432 15978
rect 7380 15914 7432 15920
rect 7484 15706 7512 16526
rect 7564 16516 7616 16522
rect 7564 16458 7616 16464
rect 7472 15700 7524 15706
rect 7472 15642 7524 15648
rect 7576 15314 7604 16458
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 7748 15360 7800 15366
rect 7576 15308 7748 15314
rect 7576 15302 7800 15308
rect 7576 15286 7788 15302
rect 7300 15014 7420 15042
rect 7288 14952 7340 14958
rect 7288 14894 7340 14900
rect 6644 14350 6696 14356
rect 6656 12442 6684 14350
rect 6736 14340 6788 14346
rect 6736 14282 6788 14288
rect 6932 14334 7236 14362
rect 6748 13938 6776 14282
rect 6736 13932 6788 13938
rect 6736 13874 6788 13880
rect 6932 12782 6960 14334
rect 7300 14278 7328 14894
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7104 14000 7156 14006
rect 7104 13942 7156 13948
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 7024 12986 7052 13670
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 6736 12708 6788 12714
rect 6736 12650 6788 12656
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6564 12294 6684 12322
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6276 10532 6328 10538
rect 6276 10474 6328 10480
rect 6288 10266 6316 10474
rect 6564 10470 6592 12174
rect 6460 10464 6512 10470
rect 6460 10406 6512 10412
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 6092 9648 6144 9654
rect 6092 9590 6144 9596
rect 6472 9518 6500 10406
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 4066 9143 4122 9152
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4988 9172 5040 9178
rect 5276 9166 5396 9194
rect 4988 9114 5040 9120
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 3976 8560 4028 8566
rect 3976 8502 4028 8508
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 3974 8120 4030 8129
rect 3974 8055 3976 8064
rect 4028 8055 4030 8064
rect 3976 8026 4028 8032
rect 4080 7721 4108 8230
rect 4066 7712 4122 7721
rect 4066 7647 4122 7656
rect 4356 7274 4384 8434
rect 5000 7886 5028 9114
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 5184 8022 5212 8910
rect 5276 8498 5304 8978
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5172 8016 5224 8022
rect 5172 7958 5224 7964
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 5000 7546 5028 7822
rect 5184 7546 5212 7958
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 4344 7268 4396 7274
rect 4344 7210 4396 7216
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3148 5840 3200 5846
rect 3148 5782 3200 5788
rect 3804 5710 3832 6054
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 2780 5636 2832 5642
rect 2780 5578 2832 5584
rect 3700 5636 3752 5642
rect 3700 5578 3752 5584
rect 3712 5234 3740 5578
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 3804 5166 3832 5646
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3240 5092 3292 5098
rect 3240 5034 3292 5040
rect 3252 4729 3280 5034
rect 3238 4720 3294 4729
rect 3238 4655 3294 4664
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3528 3233 3556 4082
rect 3514 3224 3570 3233
rect 3514 3159 3570 3168
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 3068 1737 3096 2450
rect 3054 1728 3110 1737
rect 3054 1663 3110 1672
rect 3424 1352 3476 1358
rect 3424 1294 3476 1300
rect 3436 649 3464 1294
rect 3896 1193 3924 6938
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 4068 6724 4120 6730
rect 4068 6666 4120 6672
rect 4080 6225 4108 6666
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 5092 6322 5120 6598
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 4066 6216 4122 6225
rect 3976 6180 4028 6186
rect 4066 6151 4122 6160
rect 3976 6122 4028 6128
rect 3988 5681 4016 6122
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 3974 5672 4030 5681
rect 3974 5607 4030 5616
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4080 5137 4108 5510
rect 4356 5370 4384 6054
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4066 5128 4122 5137
rect 4066 5063 4122 5072
rect 5000 4826 5028 6054
rect 5184 5846 5212 6734
rect 5172 5840 5224 5846
rect 5172 5782 5224 5788
rect 5184 5370 5212 5782
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4068 4752 4120 4758
rect 4068 4694 4120 4700
rect 4080 4185 4108 4694
rect 5184 4690 5212 5306
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5276 4826 5304 4966
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5368 4622 5396 9166
rect 6472 9042 6500 9454
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 6104 7177 6132 7822
rect 6090 7168 6146 7177
rect 6090 7103 6146 7112
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6564 5914 6592 6258
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6656 5234 6684 12294
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 4066 4176 4122 4185
rect 4066 4111 4122 4120
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 4080 3641 4108 4014
rect 4066 3632 4122 3641
rect 4066 3567 4122 3576
rect 4066 2680 4122 2689
rect 4066 2615 4068 2624
rect 4120 2615 4122 2624
rect 4068 2586 4120 2592
rect 4172 2145 4200 4558
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 5552 2650 5580 5170
rect 6748 4010 6776 12650
rect 7116 11762 7144 13942
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7208 11694 7236 14214
rect 7288 13728 7340 13734
rect 7288 13670 7340 13676
rect 7300 13530 7328 13670
rect 7392 13530 7420 15014
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7300 12782 7328 12922
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 7208 11218 7236 11494
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6932 10690 6960 11086
rect 6840 10662 6960 10690
rect 6840 10606 6868 10662
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6932 9722 6960 10662
rect 7116 10266 7144 11154
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 7392 9994 7420 13466
rect 7576 13410 7604 15286
rect 8220 15162 8248 16526
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 8312 15570 8340 16050
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 7668 13530 7696 14418
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 7576 13382 7696 13410
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7576 12850 7604 13262
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7484 10266 7512 12242
rect 7576 12238 7604 12786
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7472 10260 7524 10266
rect 7472 10202 7524 10208
rect 7380 9988 7432 9994
rect 7380 9930 7432 9936
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 6932 9518 6960 9658
rect 7196 9648 7248 9654
rect 7196 9590 7248 9596
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6932 8480 6960 9454
rect 7208 9382 7236 9590
rect 7392 9586 7420 9930
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7288 9036 7340 9042
rect 7288 8978 7340 8984
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7116 8634 7144 8910
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 6840 8452 6960 8480
rect 6840 7410 6868 8452
rect 7300 8090 7328 8978
rect 7392 8498 7420 9522
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7668 8378 7696 13382
rect 7748 13388 7800 13394
rect 7748 13330 7800 13336
rect 7760 11762 7788 13330
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 8312 12442 8340 14418
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 8404 12170 8432 18226
rect 9048 18222 9076 22520
rect 9496 19984 9548 19990
rect 9496 19926 9548 19932
rect 9128 19916 9180 19922
rect 9128 19858 9180 19864
rect 9140 19514 9168 19858
rect 9508 19786 9536 19926
rect 9220 19780 9272 19786
rect 9220 19722 9272 19728
rect 9496 19780 9548 19786
rect 9496 19722 9548 19728
rect 9128 19508 9180 19514
rect 9128 19450 9180 19456
rect 9140 18766 9168 19450
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 9036 18216 9088 18222
rect 9036 18158 9088 18164
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8944 18080 8996 18086
rect 8944 18022 8996 18028
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8496 16114 8524 17138
rect 8588 17134 8616 18022
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8484 16108 8536 16114
rect 8484 16050 8536 16056
rect 8496 14414 8524 16050
rect 8956 14822 8984 18022
rect 9232 16130 9260 19722
rect 9496 18284 9548 18290
rect 9496 18226 9548 18232
rect 9508 16998 9536 18226
rect 9600 18170 9628 22520
rect 10060 20482 10088 22520
rect 10060 20454 10180 20482
rect 10520 20466 10548 22520
rect 10048 20392 10100 20398
rect 10048 20334 10100 20340
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9954 19816 10010 19825
rect 9692 18766 9720 19790
rect 9954 19751 10010 19760
rect 9968 19446 9996 19751
rect 10060 19514 10088 20334
rect 10048 19508 10100 19514
rect 10048 19450 10100 19456
rect 9956 19440 10008 19446
rect 9956 19382 10008 19388
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 9600 18142 9812 18170
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9692 17882 9720 18022
rect 9784 17882 9812 18142
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9968 17338 9996 18702
rect 10152 18290 10180 20454
rect 10508 20460 10560 20466
rect 10508 20402 10560 20408
rect 10416 20256 10468 20262
rect 10416 20198 10468 20204
rect 10600 20256 10652 20262
rect 10600 20198 10652 20204
rect 10428 19378 10456 20198
rect 10612 19990 10640 20198
rect 10600 19984 10652 19990
rect 10600 19926 10652 19932
rect 10692 19780 10744 19786
rect 10692 19722 10744 19728
rect 10704 19378 10732 19722
rect 10416 19372 10468 19378
rect 10416 19314 10468 19320
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10704 18850 10732 19314
rect 10704 18834 10824 18850
rect 10704 18828 10836 18834
rect 10704 18822 10784 18828
rect 10784 18770 10836 18776
rect 10782 18320 10838 18329
rect 10140 18284 10192 18290
rect 10782 18255 10838 18264
rect 10140 18226 10192 18232
rect 10048 18216 10100 18222
rect 10048 18158 10100 18164
rect 9956 17332 10008 17338
rect 9956 17274 10008 17280
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9048 16102 9260 16130
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8852 13184 8904 13190
rect 8852 13126 8904 13132
rect 8864 12442 8892 13126
rect 8944 12912 8996 12918
rect 8944 12854 8996 12860
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8956 12306 8984 12854
rect 9048 12782 9076 16102
rect 9508 16046 9536 16934
rect 9968 16794 9996 17274
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9692 16250 9720 16730
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9588 16176 9640 16182
rect 9588 16118 9640 16124
rect 9496 16040 9548 16046
rect 9496 15982 9548 15988
rect 9220 15564 9272 15570
rect 9220 15506 9272 15512
rect 9232 15162 9260 15506
rect 9600 15434 9628 16118
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 9692 15706 9720 15846
rect 10060 15706 10088 18158
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 9588 15428 9640 15434
rect 9588 15370 9640 15376
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9600 14958 9628 15370
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 9232 13938 9260 14350
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 10152 13462 10180 17682
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 10336 17134 10364 17614
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10796 14958 10824 18255
rect 10980 18222 11008 22520
rect 11244 21004 11296 21010
rect 11244 20946 11296 20952
rect 11150 18320 11206 18329
rect 11150 18255 11206 18264
rect 10968 18216 11020 18222
rect 10968 18158 11020 18164
rect 11164 18154 11192 18255
rect 10876 18148 10928 18154
rect 10876 18090 10928 18096
rect 11152 18148 11204 18154
rect 11152 18090 11204 18096
rect 10888 17134 10916 18090
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 11072 17066 11100 18022
rect 11152 17740 11204 17746
rect 11152 17682 11204 17688
rect 11060 17060 11112 17066
rect 11060 17002 11112 17008
rect 11164 16658 11192 17682
rect 11256 17338 11284 20946
rect 11440 20890 11468 22520
rect 11440 20862 11744 20890
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 11716 18086 11744 20862
rect 11796 20596 11848 20602
rect 11796 20538 11848 20544
rect 11808 18136 11836 20538
rect 11900 19938 11928 22520
rect 12072 20460 12124 20466
rect 12072 20402 12124 20408
rect 12164 20460 12216 20466
rect 12164 20402 12216 20408
rect 12084 19990 12112 20402
rect 12072 19984 12124 19990
rect 11900 19910 12020 19938
rect 12072 19926 12124 19932
rect 11888 19848 11940 19854
rect 11888 19790 11940 19796
rect 11900 19378 11928 19790
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 11888 18148 11940 18154
rect 11808 18108 11888 18136
rect 11888 18090 11940 18096
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11244 17332 11296 17338
rect 11244 17274 11296 17280
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10612 14006 10640 14418
rect 10600 14000 10652 14006
rect 10600 13942 10652 13948
rect 10140 13456 10192 13462
rect 10140 13398 10192 13404
rect 9128 13388 9180 13394
rect 9128 13330 9180 13336
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 8392 12164 8444 12170
rect 8392 12106 8444 12112
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8312 11218 8340 11290
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 8208 11076 8260 11082
rect 8208 11018 8260 11024
rect 8220 10810 8248 11018
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7886 10288 8182 10308
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 7760 9586 7788 9998
rect 8404 9654 8432 12106
rect 8576 11620 8628 11626
rect 8576 11562 8628 11568
rect 8588 11354 8616 11562
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8680 10849 8708 11290
rect 8852 11212 8904 11218
rect 8852 11154 8904 11160
rect 8666 10840 8722 10849
rect 8666 10775 8722 10784
rect 8864 9926 8892 11154
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 7484 8350 7696 8378
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6840 6798 6868 7346
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6840 6254 6868 6734
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6840 5234 6868 6190
rect 7484 5778 7512 8350
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7576 5914 7604 7890
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 7668 4146 7696 8230
rect 7760 7886 7788 8434
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 7760 7274 7788 7822
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7944 7342 7972 7686
rect 8220 7546 8248 8910
rect 8404 8362 8432 9590
rect 8484 8900 8536 8906
rect 8484 8842 8536 8848
rect 8496 8634 8524 8842
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8944 8424 8996 8430
rect 8944 8366 8996 8372
rect 8392 8356 8444 8362
rect 8392 8298 8444 8304
rect 8956 8090 8984 8366
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 7748 7268 7800 7274
rect 7748 7210 7800 7216
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 8220 6934 8248 7482
rect 9048 7002 9076 12718
rect 9140 10674 9168 13330
rect 10612 12374 10640 13942
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10704 13326 10732 13806
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10704 12918 10732 13262
rect 10692 12912 10744 12918
rect 10692 12854 10744 12860
rect 10600 12368 10652 12374
rect 10600 12310 10652 12316
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9324 9178 9352 12242
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9416 8566 9444 12174
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9588 10736 9640 10742
rect 9586 10704 9588 10713
rect 9640 10704 9642 10713
rect 9586 10639 9642 10648
rect 9692 10606 9720 11086
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 9968 10810 9996 10950
rect 10060 10810 10088 11018
rect 9956 10804 10008 10810
rect 9956 10746 10008 10752
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9692 9217 9720 10542
rect 10244 9654 10272 12174
rect 10322 11792 10378 11801
rect 10322 11727 10378 11736
rect 10336 11694 10364 11727
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10336 10266 10364 11630
rect 10428 11626 10456 12174
rect 10600 12164 10652 12170
rect 10600 12106 10652 12112
rect 10416 11620 10468 11626
rect 10416 11562 10468 11568
rect 10506 11248 10562 11257
rect 10506 11183 10508 11192
rect 10560 11183 10562 11192
rect 10508 11154 10560 11160
rect 10324 10260 10376 10266
rect 10324 10202 10376 10208
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9678 9208 9734 9217
rect 9678 9143 9734 9152
rect 9692 9042 9720 9143
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9404 8560 9456 8566
rect 9404 8502 9456 8508
rect 9784 8498 9812 9454
rect 10244 9042 10272 9590
rect 10336 9518 10364 10066
rect 10612 9722 10640 12106
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10704 11626 10732 12038
rect 10692 11620 10744 11626
rect 10692 11562 10744 11568
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 10506 9208 10562 9217
rect 10506 9143 10562 9152
rect 10232 9036 10284 9042
rect 10232 8978 10284 8984
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 10048 7948 10100 7954
rect 10048 7890 10100 7896
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 9876 7546 9904 7822
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8312 6458 8340 6598
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 9508 6254 9536 7346
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 8312 5778 8340 6054
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8312 5166 8340 5714
rect 9508 5370 9536 6190
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9692 5166 9720 5646
rect 10060 5370 10088 7890
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 7656 4140 7708 4146
rect 7656 4082 7708 4088
rect 5724 4004 5776 4010
rect 5724 3946 5776 3952
rect 6736 4004 6788 4010
rect 6736 3946 6788 3952
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4158 2136 4214 2145
rect 4421 2128 4717 2148
rect 4158 2071 4214 2080
rect 3882 1184 3938 1193
rect 3882 1119 3938 1128
rect 3422 640 3478 649
rect 3422 575 3478 584
rect 5736 480 5764 3946
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 10244 2514 10272 7278
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 10336 5914 10364 7142
rect 10520 6798 10548 9143
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10704 6934 10732 7822
rect 10796 7342 10824 14894
rect 11072 14618 11100 15846
rect 11164 15706 11192 16594
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11244 15904 11296 15910
rect 11244 15846 11296 15852
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11256 15570 11284 15846
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11244 15428 11296 15434
rect 11244 15370 11296 15376
rect 11256 15026 11284 15370
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11716 15094 11744 16050
rect 11900 15570 11928 18090
rect 11992 15706 12020 19910
rect 12084 18834 12112 19926
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 12084 18290 12112 18566
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 12084 16726 12112 18226
rect 12176 16810 12204 20402
rect 12360 19310 12388 22520
rect 12716 20528 12768 20534
rect 12716 20470 12768 20476
rect 12728 20398 12756 20470
rect 12716 20392 12768 20398
rect 12716 20334 12768 20340
rect 12820 20346 12848 22520
rect 13280 20602 13308 22520
rect 13268 20596 13320 20602
rect 13268 20538 13320 20544
rect 12820 20318 13400 20346
rect 12808 20256 12860 20262
rect 12808 20198 12860 20204
rect 12820 19825 12848 20198
rect 12900 19916 12952 19922
rect 12900 19858 12952 19864
rect 12806 19816 12862 19825
rect 12806 19751 12862 19760
rect 12348 19304 12400 19310
rect 12348 19246 12400 19252
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 12256 19236 12308 19242
rect 12256 19178 12308 19184
rect 12268 18426 12296 19178
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12440 18624 12492 18630
rect 12440 18566 12492 18572
rect 12256 18420 12308 18426
rect 12256 18362 12308 18368
rect 12176 16782 12388 16810
rect 12072 16720 12124 16726
rect 12072 16662 12124 16668
rect 12164 16448 12216 16454
rect 12164 16390 12216 16396
rect 12176 15706 12204 16390
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 12164 15700 12216 15706
rect 12164 15642 12216 15648
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 11704 15088 11756 15094
rect 11704 15030 11756 15036
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11060 14000 11112 14006
rect 11060 13942 11112 13948
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10888 12850 10916 13330
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10980 11762 11008 13466
rect 11072 12850 11100 13942
rect 11808 13190 11836 15506
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11900 13002 11928 15506
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 12256 15496 12308 15502
rect 12256 15438 12308 15444
rect 12084 14890 12112 15438
rect 12268 15162 12296 15438
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12072 14884 12124 14890
rect 12072 14826 12124 14832
rect 12084 14618 12112 14826
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 12072 13932 12124 13938
rect 12072 13874 12124 13880
rect 12084 13394 12112 13874
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 11808 12974 11928 13002
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 10968 11756 11020 11762
rect 10968 11698 11020 11704
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 10968 11280 11020 11286
rect 10968 11222 11020 11228
rect 11060 11280 11112 11286
rect 11060 11222 11112 11228
rect 10980 11121 11008 11222
rect 10966 11112 11022 11121
rect 10966 11047 11022 11056
rect 11072 10606 11100 11222
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 11072 10010 11100 10542
rect 10980 9982 11100 10010
rect 10980 9194 11008 9982
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11072 9382 11100 9862
rect 11164 9654 11192 11698
rect 11256 10266 11284 12922
rect 11704 12368 11756 12374
rect 11704 12310 11756 12316
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 11348 11286 11376 11698
rect 11518 11384 11574 11393
rect 11518 11319 11520 11328
rect 11572 11319 11574 11328
rect 11520 11290 11572 11296
rect 11716 11286 11744 12310
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 11704 11280 11756 11286
rect 11704 11222 11756 11228
rect 11808 11132 11836 12974
rect 11888 12368 11940 12374
rect 11888 12310 11940 12316
rect 11900 12170 11928 12310
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 11888 11824 11940 11830
rect 11888 11766 11940 11772
rect 11716 11104 11836 11132
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11152 9648 11204 9654
rect 11152 9590 11204 9596
rect 11256 9518 11284 9862
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 11610 9208 11666 9217
rect 10980 9178 11100 9194
rect 10980 9172 11112 9178
rect 10980 9166 11060 9172
rect 11610 9143 11612 9152
rect 11060 9114 11112 9120
rect 11664 9143 11666 9152
rect 11612 9114 11664 9120
rect 10876 8900 10928 8906
rect 10876 8842 10928 8848
rect 10888 8430 10916 8842
rect 11716 8820 11744 11104
rect 11796 10260 11848 10266
rect 11796 10202 11848 10208
rect 11256 8792 11744 8820
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11164 8022 11192 8230
rect 11152 8016 11204 8022
rect 11152 7958 11204 7964
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10520 6458 10548 6734
rect 10704 6458 10732 6870
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 11256 5846 11284 8792
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11704 8560 11756 8566
rect 11704 8502 11756 8508
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11716 7410 11744 8502
rect 11808 8362 11836 10202
rect 11796 8356 11848 8362
rect 11796 8298 11848 8304
rect 11900 7954 11928 11766
rect 12084 9518 12112 13330
rect 12256 12708 12308 12714
rect 12256 12650 12308 12656
rect 12164 11620 12216 11626
rect 12164 11562 12216 11568
rect 12176 11014 12204 11562
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 12268 10606 12296 12650
rect 12256 10600 12308 10606
rect 12256 10542 12308 10548
rect 12268 10198 12296 10542
rect 12256 10192 12308 10198
rect 12256 10134 12308 10140
rect 12072 9512 12124 9518
rect 12072 9454 12124 9460
rect 12256 9512 12308 9518
rect 12256 9454 12308 9460
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11992 8566 12020 9114
rect 12084 9042 12112 9318
rect 12164 9104 12216 9110
rect 12162 9072 12164 9081
rect 12216 9072 12218 9081
rect 12072 9036 12124 9042
rect 12162 9007 12218 9016
rect 12072 8978 12124 8984
rect 11980 8560 12032 8566
rect 11980 8502 12032 8508
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11992 7868 12020 8502
rect 12072 7880 12124 7886
rect 11992 7840 12072 7868
rect 12072 7822 12124 7828
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 12268 7002 12296 9454
rect 12360 8022 12388 16782
rect 12452 16046 12480 18566
rect 12544 18426 12572 18702
rect 12532 18420 12584 18426
rect 12532 18362 12584 18368
rect 12624 17264 12676 17270
rect 12624 17206 12676 17212
rect 12636 16114 12664 17206
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12452 13462 12480 14894
rect 12728 13870 12756 19246
rect 12912 18970 12940 19858
rect 12992 19780 13044 19786
rect 12992 19722 13044 19728
rect 13004 19446 13032 19722
rect 12992 19440 13044 19446
rect 12992 19382 13044 19388
rect 13176 19304 13228 19310
rect 13176 19246 13228 19252
rect 12900 18964 12952 18970
rect 12900 18906 12952 18912
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 13096 18358 13124 18566
rect 13084 18352 13136 18358
rect 13084 18294 13136 18300
rect 13188 17882 13216 19246
rect 13268 18080 13320 18086
rect 13268 18022 13320 18028
rect 13176 17876 13228 17882
rect 13176 17818 13228 17824
rect 12992 17740 13044 17746
rect 12992 17682 13044 17688
rect 13004 17202 13032 17682
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 13004 16794 13032 17138
rect 12992 16788 13044 16794
rect 12992 16730 13044 16736
rect 13280 16658 13308 18022
rect 13268 16652 13320 16658
rect 13268 16594 13320 16600
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12716 13864 12768 13870
rect 12716 13806 12768 13812
rect 12820 13802 12848 15302
rect 12808 13796 12860 13802
rect 12808 13738 12860 13744
rect 12440 13456 12492 13462
rect 12440 13398 12492 13404
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 13188 12850 13216 13126
rect 13176 12844 13228 12850
rect 13176 12786 13228 12792
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12452 11694 12480 12718
rect 12624 12300 12676 12306
rect 12624 12242 12676 12248
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12544 11014 12572 11290
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12636 10538 12664 12242
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12728 11898 12756 12174
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12728 11218 12756 11834
rect 12820 11626 12848 12038
rect 13280 11801 13308 12242
rect 13266 11792 13322 11801
rect 13266 11727 13322 11736
rect 12808 11620 12860 11626
rect 12808 11562 12860 11568
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 13084 11144 13136 11150
rect 13082 11112 13084 11121
rect 13176 11144 13228 11150
rect 13136 11112 13138 11121
rect 13176 11086 13228 11092
rect 13082 11047 13138 11056
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12624 10532 12676 10538
rect 12624 10474 12676 10480
rect 12728 9994 12756 10950
rect 13188 10810 13216 11086
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 12900 10532 12952 10538
rect 12900 10474 12952 10480
rect 12716 9988 12768 9994
rect 12716 9930 12768 9936
rect 12912 9450 12940 10474
rect 12900 9444 12952 9450
rect 12900 9386 12952 9392
rect 13268 9444 13320 9450
rect 13268 9386 13320 9392
rect 13280 8974 13308 9386
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 12348 8016 12400 8022
rect 12348 7958 12400 7964
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 12348 6384 12400 6390
rect 12348 6326 12400 6332
rect 12360 6186 12388 6326
rect 12348 6180 12400 6186
rect 12348 6122 12400 6128
rect 13372 5914 13400 20318
rect 13452 19236 13504 19242
rect 13452 19178 13504 19184
rect 13464 18426 13492 19178
rect 13740 18902 13768 22520
rect 14292 19802 14320 22520
rect 14752 20602 14780 22520
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 15212 20058 15240 22520
rect 15476 20800 15528 20806
rect 15476 20742 15528 20748
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 14292 19774 14412 19802
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 13728 18896 13780 18902
rect 13728 18838 13780 18844
rect 13452 18420 13504 18426
rect 13452 18362 13504 18368
rect 14200 18290 14228 19110
rect 14384 18970 14412 19774
rect 15304 19310 15332 19858
rect 15488 19786 15516 20742
rect 15476 19780 15528 19786
rect 15476 19722 15528 19728
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15384 19304 15436 19310
rect 15384 19246 15436 19252
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 14648 19168 14700 19174
rect 14648 19110 14700 19116
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14568 18766 14596 19110
rect 14660 18834 14688 19110
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 14648 18828 14700 18834
rect 14648 18770 14700 18776
rect 14740 18828 14792 18834
rect 14740 18770 14792 18776
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 13636 18216 13688 18222
rect 13636 18158 13688 18164
rect 13648 17882 13676 18158
rect 13636 17876 13688 17882
rect 13636 17818 13688 17824
rect 13648 17202 13676 17818
rect 13728 17740 13780 17746
rect 13728 17682 13780 17688
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13648 16674 13676 17138
rect 13740 16794 13768 17682
rect 13912 17672 13964 17678
rect 13912 17614 13964 17620
rect 14004 17672 14056 17678
rect 14004 17614 14056 17620
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13648 16646 13768 16674
rect 13740 16046 13768 16646
rect 13728 16040 13780 16046
rect 13728 15982 13780 15988
rect 13544 15972 13596 15978
rect 13544 15914 13596 15920
rect 13556 15706 13584 15914
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13740 14958 13768 15982
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13464 13530 13492 14418
rect 13924 14414 13952 17614
rect 14016 17134 14044 17614
rect 14004 17128 14056 17134
rect 14004 17070 14056 17076
rect 14372 17060 14424 17066
rect 14372 17002 14424 17008
rect 14004 16652 14056 16658
rect 14004 16594 14056 16600
rect 14016 16130 14044 16594
rect 14384 16590 14412 17002
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14016 16102 14136 16130
rect 14004 15972 14056 15978
rect 14004 15914 14056 15920
rect 14016 15502 14044 15914
rect 14004 15496 14056 15502
rect 14004 15438 14056 15444
rect 14108 15366 14136 16102
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 14752 14550 14780 18770
rect 15396 18086 15424 19246
rect 15568 18828 15620 18834
rect 15568 18770 15620 18776
rect 15476 18148 15528 18154
rect 15476 18090 15528 18096
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 15292 17740 15344 17746
rect 15292 17682 15344 17688
rect 15304 17338 15332 17682
rect 15488 17338 15516 18090
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15476 17332 15528 17338
rect 15476 17274 15528 17280
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 15488 16590 15516 17274
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 15476 16584 15528 16590
rect 15476 16526 15528 16532
rect 15120 16250 15148 16526
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 14924 15496 14976 15502
rect 14924 15438 14976 15444
rect 14936 15162 14964 15438
rect 14832 15156 14884 15162
rect 14832 15098 14884 15104
rect 14924 15156 14976 15162
rect 14924 15098 14976 15104
rect 14844 14890 14872 15098
rect 14832 14884 14884 14890
rect 14832 14826 14884 14832
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 14740 14544 14792 14550
rect 14740 14486 14792 14492
rect 15292 14476 15344 14482
rect 15292 14418 15344 14424
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 15304 14074 15332 14418
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15488 13938 15516 15506
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 13452 13252 13504 13258
rect 13452 13194 13504 13200
rect 13464 11218 13492 13194
rect 14200 12782 14228 13262
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 13556 12170 13584 12718
rect 13820 12708 13872 12714
rect 13820 12650 13872 12656
rect 13544 12164 13596 12170
rect 13544 12106 13596 12112
rect 13832 11830 13860 12650
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14188 12300 14240 12306
rect 14188 12242 14240 12248
rect 13820 11824 13872 11830
rect 13820 11766 13872 11772
rect 14200 11354 14228 12242
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14476 11914 14504 12038
rect 14384 11886 14504 11914
rect 14384 11830 14412 11886
rect 14372 11824 14424 11830
rect 14372 11766 14424 11772
rect 14462 11384 14518 11393
rect 14188 11348 14240 11354
rect 14462 11319 14518 11328
rect 14188 11290 14240 11296
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 14108 9178 14136 9998
rect 14200 9382 14228 11290
rect 14476 11218 14504 11319
rect 14464 11212 14516 11218
rect 14464 11154 14516 11160
rect 14568 11150 14596 12106
rect 14660 11694 14688 12582
rect 14752 11898 14780 13806
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 15580 13462 15608 18770
rect 15672 18154 15700 22520
rect 15660 18148 15712 18154
rect 15660 18090 15712 18096
rect 15660 16992 15712 16998
rect 15660 16934 15712 16940
rect 15672 16794 15700 16934
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 16132 15706 16160 22520
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 16408 14550 16436 19858
rect 16592 18970 16620 22520
rect 16948 20392 17000 20398
rect 16948 20334 17000 20340
rect 16672 19712 16724 19718
rect 16672 19654 16724 19660
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 16684 18902 16712 19654
rect 16672 18896 16724 18902
rect 16672 18838 16724 18844
rect 16764 18148 16816 18154
rect 16764 18090 16816 18096
rect 16776 14618 16804 18090
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16396 14544 16448 14550
rect 16396 14486 16448 14492
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 16316 13938 16344 14418
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 16028 13864 16080 13870
rect 16028 13806 16080 13812
rect 15568 13456 15620 13462
rect 15568 13398 15620 13404
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15764 12986 15792 13330
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 16040 12442 16068 13806
rect 16304 12844 16356 12850
rect 16304 12786 16356 12792
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16028 12436 16080 12442
rect 16028 12378 16080 12384
rect 16224 11898 16252 12582
rect 16316 12374 16344 12786
rect 16304 12368 16356 12374
rect 16304 12310 16356 12316
rect 16580 12300 16632 12306
rect 16580 12242 16632 12248
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 16316 11898 16344 12038
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16304 11892 16356 11898
rect 16304 11834 16356 11840
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 15304 11257 15332 11494
rect 15290 11248 15346 11257
rect 15290 11183 15346 11192
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14568 10606 14596 11086
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14568 9586 14596 10542
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 16224 10130 16252 10406
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13832 7954 13860 8230
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 13832 7410 13860 7890
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 14200 7342 14228 8910
rect 14568 8498 14596 9522
rect 14752 9382 14780 9998
rect 15200 9716 15252 9722
rect 15200 9658 15252 9664
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14752 9058 14780 9318
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 14752 9030 14872 9058
rect 15212 9042 15240 9658
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14844 8362 14872 9030
rect 15200 9036 15252 9042
rect 15200 8978 15252 8984
rect 14832 8356 14884 8362
rect 14832 8298 14884 8304
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 15304 8090 15332 10066
rect 16408 10062 16436 10406
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 16408 9518 16436 9998
rect 16592 9994 16620 12242
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16684 10606 16712 12038
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16580 9988 16632 9994
rect 16580 9930 16632 9936
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 16592 7546 16620 8978
rect 16776 7562 16804 14214
rect 16960 13376 16988 20334
rect 17052 19174 17080 22520
rect 17408 19916 17460 19922
rect 17408 19858 17460 19864
rect 17040 19168 17092 19174
rect 17040 19110 17092 19116
rect 16960 13348 17080 13376
rect 17052 11354 17080 13348
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 17420 9042 17448 19858
rect 17512 18970 17540 22520
rect 17972 20058 18000 22520
rect 18432 21434 18460 22520
rect 18432 21406 18644 21434
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 18616 20602 18644 21406
rect 18604 20596 18656 20602
rect 18604 20538 18656 20544
rect 18144 20392 18196 20398
rect 18144 20334 18196 20340
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17500 18964 17552 18970
rect 17500 18906 17552 18912
rect 17500 18828 17552 18834
rect 17500 18770 17552 18776
rect 17512 10198 17540 18770
rect 17880 12374 17908 19246
rect 18050 18184 18106 18193
rect 18050 18119 18052 18128
rect 18104 18119 18106 18128
rect 18052 18090 18104 18096
rect 17960 18080 18012 18086
rect 17960 18022 18012 18028
rect 17868 12368 17920 12374
rect 17868 12310 17920 12316
rect 17972 11642 18000 18022
rect 17972 11614 18092 11642
rect 17958 11520 18014 11529
rect 17958 11455 18014 11464
rect 17972 11286 18000 11455
rect 17960 11280 18012 11286
rect 17960 11222 18012 11228
rect 18064 10588 18092 11614
rect 17972 10560 18092 10588
rect 17500 10192 17552 10198
rect 17500 10134 17552 10140
rect 17972 9654 18000 10560
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 18064 10266 18092 10406
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 18156 9738 18184 20334
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18282 14096 18578 14116
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 18064 9710 18184 9738
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 17866 9072 17922 9081
rect 17408 9036 17460 9042
rect 17866 9007 17868 9016
rect 17408 8978 17460 8984
rect 17920 9007 17922 9016
rect 17868 8978 17920 8984
rect 18064 8566 18092 9710
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 18156 9110 18184 9454
rect 18144 9104 18196 9110
rect 18144 9046 18196 9052
rect 18616 8974 18644 19858
rect 18984 18086 19012 22520
rect 19156 19984 19208 19990
rect 19156 19926 19208 19932
rect 19168 19378 19196 19926
rect 19156 19372 19208 19378
rect 19156 19314 19208 19320
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 18604 8968 18656 8974
rect 18604 8910 18656 8916
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 19444 8634 19472 22520
rect 19708 19848 19760 19854
rect 19708 19790 19760 19796
rect 19720 18698 19748 19790
rect 19708 18692 19760 18698
rect 19708 18634 19760 18640
rect 19616 18216 19668 18222
rect 19616 18158 19668 18164
rect 19432 8628 19484 8634
rect 19432 8570 19484 8576
rect 18052 8560 18104 8566
rect 18052 8502 18104 8508
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19352 8022 19380 8366
rect 19340 8016 19392 8022
rect 19340 7958 19392 7964
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 16580 7540 16632 7546
rect 16776 7534 17264 7562
rect 16580 7482 16632 7488
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 14817 7100 15113 7120
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 13360 5908 13412 5914
rect 13360 5850 13412 5856
rect 11244 5840 11296 5846
rect 11244 5782 11296 5788
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 10232 2508 10284 2514
rect 10232 2450 10284 2456
rect 11072 1358 11100 5714
rect 12360 5574 12388 5714
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12348 4752 12400 4758
rect 12452 4706 12480 4762
rect 12400 4700 12480 4706
rect 12348 4694 12480 4700
rect 12360 4678 12480 4694
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 11060 1352 11112 1358
rect 11060 1294 11112 1300
rect 17236 480 17264 7534
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 19628 5370 19656 18158
rect 19708 18080 19760 18086
rect 19708 18022 19760 18028
rect 19720 6458 19748 18022
rect 19904 6730 19932 22520
rect 20364 18086 20392 22520
rect 20352 18080 20404 18086
rect 20352 18022 20404 18028
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20732 17354 20760 18022
rect 20824 17490 20852 22520
rect 21284 18222 21312 22520
rect 21272 18216 21324 18222
rect 21272 18158 21324 18164
rect 21088 18148 21140 18154
rect 21088 18090 21140 18096
rect 20824 17462 21036 17490
rect 20732 17326 20944 17354
rect 20812 17264 20864 17270
rect 20812 17206 20864 17212
rect 19892 6724 19944 6730
rect 19892 6666 19944 6672
rect 19708 6452 19760 6458
rect 19708 6394 19760 6400
rect 19616 5364 19668 5370
rect 19616 5306 19668 5312
rect 20536 5160 20588 5166
rect 20536 5102 20588 5108
rect 20548 4826 20576 5102
rect 20536 4820 20588 4826
rect 20536 4762 20588 4768
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 20824 3942 20852 17206
rect 20916 5370 20944 17326
rect 21008 5914 21036 17462
rect 21100 17270 21128 18090
rect 21744 18086 21772 22520
rect 22204 18154 22232 22520
rect 22664 18630 22692 22520
rect 22652 18624 22704 18630
rect 22652 18566 22704 18572
rect 22192 18148 22244 18154
rect 22192 18090 22244 18096
rect 21732 18080 21784 18086
rect 21732 18022 21784 18028
rect 21088 17264 21140 17270
rect 21088 17206 21140 17212
rect 20996 5908 21048 5914
rect 20996 5850 21048 5856
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 20812 3936 20864 3942
rect 20812 3878 20864 3884
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 2686 232 2742 241
rect 2686 167 2742 176
rect 5722 0 5778 480
rect 17222 0 17278 480
<< via2 >>
rect 3790 22616 3846 22672
rect 1858 21120 1914 21176
rect 1582 16632 1638 16688
rect 1766 16088 1822 16144
rect 1582 13096 1638 13152
rect 1950 18128 2006 18184
rect 2134 19760 2190 19816
rect 2778 18264 2834 18320
rect 2778 17856 2834 17912
rect 1950 14048 2006 14104
rect 2042 12588 2044 12608
rect 2044 12588 2096 12608
rect 2096 12588 2098 12608
rect 2042 12552 2098 12588
rect 2042 11600 2098 11656
rect 3238 18536 3294 18592
rect 3330 18148 3386 18184
rect 3330 18128 3332 18148
rect 3332 18128 3384 18148
rect 3384 18128 3386 18148
rect 2226 6568 2282 6624
rect 3330 13640 3386 13696
rect 3514 21528 3570 21584
rect 3790 20032 3846 20088
rect 3514 17040 3570 17096
rect 3514 14612 3570 14648
rect 3514 14592 3516 14612
rect 3516 14592 3568 14612
rect 3568 14592 3570 14612
rect 4066 22072 4122 22128
rect 3974 20596 4030 20632
rect 3974 20576 3976 20596
rect 3976 20576 4028 20596
rect 4028 20576 4030 20596
rect 3974 19624 4030 19680
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 4250 19080 4306 19136
rect 4526 18844 4528 18864
rect 4528 18844 4580 18864
rect 4580 18844 4582 18864
rect 4526 18808 4582 18844
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 4066 17720 4122 17776
rect 3974 17584 4030 17640
rect 4710 17992 4766 18048
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 4066 15544 4122 15600
rect 3882 15136 3938 15192
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 5538 19252 5540 19272
rect 5540 19252 5592 19272
rect 5592 19252 5594 19272
rect 5538 19216 5594 19252
rect 5998 19216 6054 19272
rect 5630 17856 5686 17912
rect 4066 12144 4122 12200
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 4066 11056 4122 11112
rect 3698 9560 3754 9616
rect 3514 8608 3570 8664
rect 4066 10104 4122 10160
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 4894 10784 4950 10840
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 4066 9152 4122 9208
rect 6918 19760 6974 19816
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 7286 17992 7342 18048
rect 7194 17720 7250 17776
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 8298 18808 8354 18864
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 3974 8084 4030 8120
rect 3974 8064 3976 8084
rect 3976 8064 4028 8084
rect 4028 8064 4030 8084
rect 4066 7656 4122 7712
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 3238 4664 3294 4720
rect 3514 3168 3570 3224
rect 3054 1672 3110 1728
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4066 6160 4122 6216
rect 3974 5616 4030 5672
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 4066 5072 4122 5128
rect 6090 7112 6146 7168
rect 4066 4120 4122 4176
rect 4066 3576 4122 3632
rect 4066 2644 4122 2680
rect 4066 2624 4068 2644
rect 4068 2624 4120 2644
rect 4120 2624 4122 2644
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 9954 19760 10010 19816
rect 10782 18264 10838 18320
rect 11150 18264 11206 18320
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 8666 10784 8722 10840
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 9586 10684 9588 10704
rect 9588 10684 9640 10704
rect 9640 10684 9642 10704
rect 9586 10648 9642 10684
rect 10322 11736 10378 11792
rect 10506 11212 10562 11248
rect 10506 11192 10508 11212
rect 10508 11192 10560 11212
rect 10560 11192 10562 11212
rect 9678 9152 9734 9208
rect 10506 9152 10562 9208
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 4158 2080 4214 2136
rect 3882 1128 3938 1184
rect 3422 584 3478 640
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 12806 19760 12862 19816
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 10966 11056 11022 11112
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11518 11348 11574 11384
rect 11518 11328 11520 11348
rect 11520 11328 11572 11348
rect 11572 11328 11574 11348
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11610 9172 11666 9208
rect 11610 9152 11612 9172
rect 11612 9152 11664 9172
rect 11664 9152 11666 9172
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 12162 9052 12164 9072
rect 12164 9052 12216 9072
rect 12216 9052 12218 9072
rect 12162 9016 12218 9052
rect 13266 11736 13322 11792
rect 13082 11092 13084 11112
rect 13084 11092 13136 11112
rect 13136 11092 13138 11112
rect 13082 11056 13138 11092
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 14462 11328 14518 11384
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 15290 11192 15346 11248
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 18050 18148 18106 18184
rect 18050 18128 18052 18148
rect 18052 18128 18104 18148
rect 18104 18128 18106 18148
rect 17958 11464 18014 11520
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 17866 9036 17922 9072
rect 17866 9016 17868 9036
rect 17868 9016 17920 9036
rect 17920 9016 17922 9036
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 2686 176 2742 232
<< metal3 >>
rect 0 22674 480 22704
rect 3785 22674 3851 22677
rect 0 22672 3851 22674
rect 0 22616 3790 22672
rect 3846 22616 3851 22672
rect 0 22614 3851 22616
rect 0 22584 480 22614
rect 3785 22611 3851 22614
rect 0 22130 480 22160
rect 4061 22130 4127 22133
rect 0 22128 4127 22130
rect 0 22072 4066 22128
rect 4122 22072 4127 22128
rect 0 22070 4127 22072
rect 0 22040 480 22070
rect 4061 22067 4127 22070
rect 0 21586 480 21616
rect 3509 21586 3575 21589
rect 0 21584 3575 21586
rect 0 21528 3514 21584
rect 3570 21528 3575 21584
rect 0 21526 3575 21528
rect 0 21496 480 21526
rect 3509 21523 3575 21526
rect 0 21178 480 21208
rect 1853 21178 1919 21181
rect 0 21176 1919 21178
rect 0 21120 1858 21176
rect 1914 21120 1919 21176
rect 0 21118 1919 21120
rect 0 21088 480 21118
rect 1853 21115 1919 21118
rect 4409 20704 4729 20705
rect 0 20634 480 20664
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 20639 18590 20640
rect 3969 20634 4035 20637
rect 0 20632 4035 20634
rect 0 20576 3974 20632
rect 4030 20576 4035 20632
rect 0 20574 4035 20576
rect 0 20544 480 20574
rect 3969 20571 4035 20574
rect 7874 20160 8194 20161
rect 0 20090 480 20120
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 3785 20090 3851 20093
rect 0 20088 3851 20090
rect 0 20032 3790 20088
rect 3846 20032 3851 20088
rect 0 20030 3851 20032
rect 0 20000 480 20030
rect 3785 20027 3851 20030
rect 2129 19818 2195 19821
rect 6913 19818 6979 19821
rect 2129 19816 6979 19818
rect 2129 19760 2134 19816
rect 2190 19760 6918 19816
rect 6974 19760 6979 19816
rect 2129 19758 6979 19760
rect 2129 19755 2195 19758
rect 6913 19755 6979 19758
rect 9949 19818 10015 19821
rect 12801 19818 12867 19821
rect 9949 19816 12867 19818
rect 9949 19760 9954 19816
rect 10010 19760 12806 19816
rect 12862 19760 12867 19816
rect 9949 19758 12867 19760
rect 9949 19755 10015 19758
rect 12801 19755 12867 19758
rect 0 19682 480 19712
rect 3969 19682 4035 19685
rect 0 19680 4035 19682
rect 0 19624 3974 19680
rect 4030 19624 4035 19680
rect 0 19622 4035 19624
rect 0 19592 480 19622
rect 3969 19619 4035 19622
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 5533 19274 5599 19277
rect 5993 19274 6059 19277
rect 5533 19272 6059 19274
rect 5533 19216 5538 19272
rect 5594 19216 5998 19272
rect 6054 19216 6059 19272
rect 5533 19214 6059 19216
rect 5533 19211 5599 19214
rect 5993 19211 6059 19214
rect 0 19138 480 19168
rect 4245 19138 4311 19141
rect 0 19136 4311 19138
rect 0 19080 4250 19136
rect 4306 19080 4311 19136
rect 0 19078 4311 19080
rect 0 19048 480 19078
rect 4245 19075 4311 19078
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 4521 18866 4587 18869
rect 8293 18866 8359 18869
rect 4521 18864 8359 18866
rect 4521 18808 4526 18864
rect 4582 18808 8298 18864
rect 8354 18808 8359 18864
rect 4521 18806 8359 18808
rect 4521 18803 4587 18806
rect 8293 18803 8359 18806
rect 0 18594 480 18624
rect 3233 18594 3299 18597
rect 0 18592 3299 18594
rect 0 18536 3238 18592
rect 3294 18536 3299 18592
rect 0 18534 3299 18536
rect 0 18504 480 18534
rect 3233 18531 3299 18534
rect 4409 18528 4729 18529
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 18463 18590 18464
rect 2773 18322 2839 18325
rect 10777 18322 10843 18325
rect 11145 18322 11211 18325
rect 2773 18320 11211 18322
rect 2773 18264 2778 18320
rect 2834 18264 10782 18320
rect 10838 18264 11150 18320
rect 11206 18264 11211 18320
rect 2773 18262 11211 18264
rect 2773 18259 2839 18262
rect 10777 18259 10843 18262
rect 11145 18259 11211 18262
rect 0 18186 480 18216
rect 1945 18186 2011 18189
rect 0 18184 2011 18186
rect 0 18128 1950 18184
rect 2006 18128 2011 18184
rect 0 18126 2011 18128
rect 0 18096 480 18126
rect 1945 18123 2011 18126
rect 3325 18186 3391 18189
rect 18045 18186 18111 18189
rect 3325 18184 18111 18186
rect 3325 18128 3330 18184
rect 3386 18128 18050 18184
rect 18106 18128 18111 18184
rect 3325 18126 18111 18128
rect 3325 18123 3391 18126
rect 18045 18123 18111 18126
rect 4705 18050 4771 18053
rect 7281 18050 7347 18053
rect 4705 18048 7347 18050
rect 4705 17992 4710 18048
rect 4766 17992 7286 18048
rect 7342 17992 7347 18048
rect 4705 17990 7347 17992
rect 4705 17987 4771 17990
rect 7281 17987 7347 17990
rect 7874 17984 8194 17985
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 17919 15125 17920
rect 2773 17914 2839 17917
rect 5625 17914 5691 17917
rect 2773 17912 5691 17914
rect 2773 17856 2778 17912
rect 2834 17856 5630 17912
rect 5686 17856 5691 17912
rect 2773 17854 5691 17856
rect 2773 17851 2839 17854
rect 5625 17851 5691 17854
rect 4061 17778 4127 17781
rect 7189 17778 7255 17781
rect 4061 17776 7255 17778
rect 4061 17720 4066 17776
rect 4122 17720 7194 17776
rect 7250 17720 7255 17776
rect 4061 17718 7255 17720
rect 4061 17715 4127 17718
rect 7189 17715 7255 17718
rect 0 17642 480 17672
rect 3969 17642 4035 17645
rect 0 17640 4035 17642
rect 0 17584 3974 17640
rect 4030 17584 4035 17640
rect 0 17582 4035 17584
rect 0 17552 480 17582
rect 3969 17579 4035 17582
rect 4409 17440 4729 17441
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 17375 18590 17376
rect 0 17098 480 17128
rect 3509 17098 3575 17101
rect 0 17096 3575 17098
rect 0 17040 3514 17096
rect 3570 17040 3575 17096
rect 0 17038 3575 17040
rect 0 17008 480 17038
rect 3509 17035 3575 17038
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 0 16690 480 16720
rect 1577 16690 1643 16693
rect 0 16688 1643 16690
rect 0 16632 1582 16688
rect 1638 16632 1643 16688
rect 0 16630 1643 16632
rect 0 16600 480 16630
rect 1577 16627 1643 16630
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 0 16146 480 16176
rect 1761 16146 1827 16149
rect 0 16144 1827 16146
rect 0 16088 1766 16144
rect 1822 16088 1827 16144
rect 0 16086 1827 16088
rect 0 16056 480 16086
rect 1761 16083 1827 16086
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 0 15602 480 15632
rect 4061 15602 4127 15605
rect 0 15600 4127 15602
rect 0 15544 4066 15600
rect 4122 15544 4127 15600
rect 0 15542 4127 15544
rect 0 15512 480 15542
rect 4061 15539 4127 15542
rect 4409 15264 4729 15265
rect 0 15194 480 15224
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 15199 18590 15200
rect 3877 15194 3943 15197
rect 0 15192 3943 15194
rect 0 15136 3882 15192
rect 3938 15136 3943 15192
rect 0 15134 3943 15136
rect 0 15104 480 15134
rect 3877 15131 3943 15134
rect 7874 14720 8194 14721
rect 0 14650 480 14680
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 3509 14650 3575 14653
rect 0 14648 3575 14650
rect 0 14592 3514 14648
rect 3570 14592 3575 14648
rect 0 14590 3575 14592
rect 0 14560 480 14590
rect 3509 14587 3575 14590
rect 4409 14176 4729 14177
rect 0 14106 480 14136
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 14111 18590 14112
rect 1945 14106 2011 14109
rect 0 14104 2011 14106
rect 0 14048 1950 14104
rect 2006 14048 2011 14104
rect 0 14046 2011 14048
rect 0 14016 480 14046
rect 1945 14043 2011 14046
rect 0 13698 480 13728
rect 3325 13698 3391 13701
rect 0 13696 3391 13698
rect 0 13640 3330 13696
rect 3386 13640 3391 13696
rect 0 13638 3391 13640
rect 0 13608 480 13638
rect 3325 13635 3391 13638
rect 7874 13632 8194 13633
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 0 13154 480 13184
rect 1577 13154 1643 13157
rect 0 13152 1643 13154
rect 0 13096 1582 13152
rect 1638 13096 1643 13152
rect 0 13094 1643 13096
rect 0 13064 480 13094
rect 1577 13091 1643 13094
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 0 12610 480 12640
rect 2037 12610 2103 12613
rect 0 12608 2103 12610
rect 0 12552 2042 12608
rect 2098 12552 2103 12608
rect 0 12550 2103 12552
rect 0 12520 480 12550
rect 2037 12547 2103 12550
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 12479 15125 12480
rect 0 12202 480 12232
rect 4061 12202 4127 12205
rect 0 12200 4127 12202
rect 0 12144 4066 12200
rect 4122 12144 4127 12200
rect 0 12142 4127 12144
rect 0 12112 480 12142
rect 4061 12139 4127 12142
rect 4409 12000 4729 12001
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 11935 18590 11936
rect 10317 11794 10383 11797
rect 13261 11794 13327 11797
rect 10317 11792 13327 11794
rect 10317 11736 10322 11792
rect 10378 11736 13266 11792
rect 13322 11736 13327 11792
rect 10317 11734 13327 11736
rect 10317 11731 10383 11734
rect 13261 11731 13327 11734
rect 0 11658 480 11688
rect 2037 11658 2103 11661
rect 0 11656 2103 11658
rect 0 11600 2042 11656
rect 2098 11600 2103 11656
rect 0 11598 2103 11600
rect 0 11568 480 11598
rect 2037 11595 2103 11598
rect 17953 11522 18019 11525
rect 22520 11522 23000 11552
rect 17953 11520 23000 11522
rect 17953 11464 17958 11520
rect 18014 11464 23000 11520
rect 17953 11462 23000 11464
rect 17953 11459 18019 11462
rect 7874 11456 8194 11457
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 22520 11432 23000 11462
rect 14805 11391 15125 11392
rect 11513 11386 11579 11389
rect 14457 11386 14523 11389
rect 11513 11384 14523 11386
rect 11513 11328 11518 11384
rect 11574 11328 14462 11384
rect 14518 11328 14523 11384
rect 11513 11326 14523 11328
rect 11513 11323 11579 11326
rect 14457 11323 14523 11326
rect 10501 11250 10567 11253
rect 15285 11250 15351 11253
rect 10501 11248 15351 11250
rect 10501 11192 10506 11248
rect 10562 11192 15290 11248
rect 15346 11192 15351 11248
rect 10501 11190 15351 11192
rect 10501 11187 10567 11190
rect 15285 11187 15351 11190
rect 0 11114 480 11144
rect 4061 11114 4127 11117
rect 0 11112 4127 11114
rect 0 11056 4066 11112
rect 4122 11056 4127 11112
rect 0 11054 4127 11056
rect 0 11024 480 11054
rect 4061 11051 4127 11054
rect 10961 11114 11027 11117
rect 13077 11114 13143 11117
rect 10961 11112 13143 11114
rect 10961 11056 10966 11112
rect 11022 11056 13082 11112
rect 13138 11056 13143 11112
rect 10961 11054 13143 11056
rect 10961 11051 11027 11054
rect 13077 11051 13143 11054
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 10847 18590 10848
rect 4889 10842 4955 10845
rect 8661 10842 8727 10845
rect 4889 10840 8727 10842
rect 4889 10784 4894 10840
rect 4950 10784 8666 10840
rect 8722 10784 8727 10840
rect 4889 10782 8727 10784
rect 4889 10779 4955 10782
rect 8661 10779 8727 10782
rect 0 10706 480 10736
rect 9581 10706 9647 10709
rect 0 10704 9647 10706
rect 0 10648 9586 10704
rect 9642 10648 9647 10704
rect 0 10646 9647 10648
rect 0 10616 480 10646
rect 9581 10643 9647 10646
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 10303 15125 10304
rect 0 10162 480 10192
rect 4061 10162 4127 10165
rect 0 10160 4127 10162
rect 0 10104 4066 10160
rect 4122 10104 4127 10160
rect 0 10102 4127 10104
rect 0 10072 480 10102
rect 4061 10099 4127 10102
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 0 9618 480 9648
rect 3693 9618 3759 9621
rect 0 9616 3759 9618
rect 0 9560 3698 9616
rect 3754 9560 3759 9616
rect 0 9558 3759 9560
rect 0 9528 480 9558
rect 3693 9555 3759 9558
rect 7874 9280 8194 9281
rect 0 9210 480 9240
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 9215 15125 9216
rect 4061 9210 4127 9213
rect 0 9208 4127 9210
rect 0 9152 4066 9208
rect 4122 9152 4127 9208
rect 0 9150 4127 9152
rect 0 9120 480 9150
rect 4061 9147 4127 9150
rect 9673 9210 9739 9213
rect 10501 9210 10567 9213
rect 11605 9210 11671 9213
rect 9673 9208 11671 9210
rect 9673 9152 9678 9208
rect 9734 9152 10506 9208
rect 10562 9152 11610 9208
rect 11666 9152 11671 9208
rect 9673 9150 11671 9152
rect 9673 9147 9739 9150
rect 10501 9147 10567 9150
rect 11605 9147 11671 9150
rect 12157 9074 12223 9077
rect 17861 9074 17927 9077
rect 12157 9072 17927 9074
rect 12157 9016 12162 9072
rect 12218 9016 17866 9072
rect 17922 9016 17927 9072
rect 12157 9014 17927 9016
rect 12157 9011 12223 9014
rect 17861 9011 17927 9014
rect 4409 8736 4729 8737
rect 0 8666 480 8696
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 3509 8666 3575 8669
rect 0 8664 3575 8666
rect 0 8608 3514 8664
rect 3570 8608 3575 8664
rect 0 8606 3575 8608
rect 0 8576 480 8606
rect 3509 8603 3575 8606
rect 7874 8192 8194 8193
rect 0 8122 480 8152
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 3969 8122 4035 8125
rect 0 8120 4035 8122
rect 0 8064 3974 8120
rect 4030 8064 4035 8120
rect 0 8062 4035 8064
rect 0 8032 480 8062
rect 3969 8059 4035 8062
rect 0 7714 480 7744
rect 4061 7714 4127 7717
rect 0 7712 4127 7714
rect 0 7656 4066 7712
rect 4122 7656 4127 7712
rect 0 7654 4127 7656
rect 0 7624 480 7654
rect 4061 7651 4127 7654
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 7583 18590 7584
rect 0 7170 480 7200
rect 6085 7170 6151 7173
rect 0 7168 6151 7170
rect 0 7112 6090 7168
rect 6146 7112 6151 7168
rect 0 7110 6151 7112
rect 0 7080 480 7110
rect 6085 7107 6151 7110
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 7039 15125 7040
rect 0 6626 480 6656
rect 2221 6626 2287 6629
rect 0 6624 2287 6626
rect 0 6568 2226 6624
rect 2282 6568 2287 6624
rect 0 6566 2287 6568
rect 0 6536 480 6566
rect 2221 6563 2287 6566
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 6495 18590 6496
rect 0 6218 480 6248
rect 4061 6218 4127 6221
rect 0 6216 4127 6218
rect 0 6160 4066 6216
rect 4122 6160 4127 6216
rect 0 6158 4127 6160
rect 0 6128 480 6158
rect 4061 6155 4127 6158
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 5951 15125 5952
rect 0 5674 480 5704
rect 3969 5674 4035 5677
rect 0 5672 4035 5674
rect 0 5616 3974 5672
rect 4030 5616 4035 5672
rect 0 5614 4035 5616
rect 0 5584 480 5614
rect 3969 5611 4035 5614
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 0 5130 480 5160
rect 4061 5130 4127 5133
rect 0 5128 4127 5130
rect 0 5072 4066 5128
rect 4122 5072 4127 5128
rect 0 5070 4127 5072
rect 0 5040 480 5070
rect 4061 5067 4127 5070
rect 7874 4928 8194 4929
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 0 4722 480 4752
rect 3233 4722 3299 4725
rect 0 4720 3299 4722
rect 0 4664 3238 4720
rect 3294 4664 3299 4720
rect 0 4662 3299 4664
rect 0 4632 480 4662
rect 3233 4659 3299 4662
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 4319 18590 4320
rect 0 4178 480 4208
rect 4061 4178 4127 4181
rect 0 4176 4127 4178
rect 0 4120 4066 4176
rect 4122 4120 4127 4176
rect 0 4118 4127 4120
rect 0 4088 480 4118
rect 4061 4115 4127 4118
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 3775 15125 3776
rect 0 3634 480 3664
rect 4061 3634 4127 3637
rect 0 3632 4127 3634
rect 0 3576 4066 3632
rect 4122 3576 4127 3632
rect 0 3574 4127 3576
rect 0 3544 480 3574
rect 4061 3571 4127 3574
rect 4409 3296 4729 3297
rect 0 3226 480 3256
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 3231 18590 3232
rect 3509 3226 3575 3229
rect 0 3224 3575 3226
rect 0 3168 3514 3224
rect 3570 3168 3575 3224
rect 0 3166 3575 3168
rect 0 3136 480 3166
rect 3509 3163 3575 3166
rect 7874 2752 8194 2753
rect 0 2682 480 2712
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 4061 2682 4127 2685
rect 0 2680 4127 2682
rect 0 2624 4066 2680
rect 4122 2624 4127 2680
rect 0 2622 4127 2624
rect 0 2592 480 2622
rect 4061 2619 4127 2622
rect 4409 2208 4729 2209
rect 0 2138 480 2168
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 4153 2138 4219 2141
rect 0 2136 4219 2138
rect 0 2080 4158 2136
rect 4214 2080 4219 2136
rect 0 2078 4219 2080
rect 0 2048 480 2078
rect 4153 2075 4219 2078
rect 0 1730 480 1760
rect 3049 1730 3115 1733
rect 0 1728 3115 1730
rect 0 1672 3054 1728
rect 3110 1672 3115 1728
rect 0 1670 3115 1672
rect 0 1640 480 1670
rect 3049 1667 3115 1670
rect 0 1186 480 1216
rect 3877 1186 3943 1189
rect 0 1184 3943 1186
rect 0 1128 3882 1184
rect 3938 1128 3943 1184
rect 0 1126 3943 1128
rect 0 1096 480 1126
rect 3877 1123 3943 1126
rect 0 642 480 672
rect 3417 642 3483 645
rect 0 640 3483 642
rect 0 584 3422 640
rect 3478 584 3483 640
rect 0 582 3483 584
rect 0 552 480 582
rect 3417 579 3483 582
rect 0 234 480 264
rect 2681 234 2747 237
rect 0 232 2747 234
rect 0 176 2686 232
rect 2742 176 2747 232
rect 0 174 2747 176
rect 0 144 480 174
rect 2681 171 2747 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 8736 4729 9760
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7874 19072 8195 20096
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7874 9280 8195 10304
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7874 8192 8195 9216
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7874 4928 8195 5952
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 20704 18590 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 18270 19616 18590 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 18528 18590 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 17440 18590 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 18270 16352 18590 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 15264 18590 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 14176 18590 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 18270 13088 18590 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 12000 18590 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 10912 18590 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 9824 18590 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 8736 18590 9760
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 7648 18590 8672
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 18270 6560 18590 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 5472 18590 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 4384 18590 5408
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 18270 3296 18590 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 2208 18590 3232
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2128 18590 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1604681595
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1604681595
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604681595
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1604681595
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1604681595
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1604681595
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1604681595
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1604681595
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1604681595
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1604681595
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1604681595
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1604681595
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1604681595
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1604681595
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1604681595
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1604681595
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1604681595
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1604681595
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_222 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 21528 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_220
timestamp 1604681595
transform 1 0 21344 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604681595
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1604681595
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1604681595
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1604681595
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1604681595
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1604681595
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1604681595
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1604681595
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1604681595
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1604681595
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1604681595
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1604681595
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1604681595
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_215
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604681595
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1604681595
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1604681595
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1604681595
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1604681595
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1604681595
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1604681595
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1604681595
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_208
timestamp 1604681595
transform 1 0 20240 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _80_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 20516 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_215
timestamp 1604681595
transform 1 0 20884 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1604681595
transform 1 0 1748 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_11
timestamp 1604681595
transform 1 0 2116 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4876 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_23
timestamp 1604681595
transform 1 0 3220 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_40
timestamp 1604681595
transform 1 0 4784 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_50
timestamp 1604681595
transform 1 0 5704 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_62
timestamp 1604681595
transform 1 0 6808 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_74
timestamp 1604681595
transform 1 0 7912 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_86
timestamp 1604681595
transform 1 0 9016 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1604681595
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1604681595
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1604681595
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1604681595
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1604681595
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1604681595
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1604681595
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1604681595
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2024 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_9
timestamp 1604681595
transform 1 0 1932 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_16
timestamp 1604681595
transform 1 0 2576 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3680 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _47_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_44
timestamp 1604681595
transform 1 0 5152 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_56
timestamp 1604681595
transform 1 0 6256 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_60
timestamp 1604681595
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8004 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_5_65
timestamp 1604681595
transform 1 0 7084 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_73
timestamp 1604681595
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10212 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_91
timestamp 1604681595
transform 1 0 9476 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_108
timestamp 1604681595
transform 1 0 11040 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1604681595
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1604681595
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1604681595
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1604681595
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1604681595
transform 1 0 19412 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_196
timestamp 1604681595
transform 1 0 19136 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_203
timestamp 1604681595
transform 1 0 19780 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1604681595
transform 1 0 20516 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_215
timestamp 1604681595
transform 1 0 20884 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 2392 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_11
timestamp 1604681595
transform 1 0 2116 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_11
timestamp 1604681595
transform 1 0 2116 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4600 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_23
timestamp 1604681595
transform 1 0 3220 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_30
timestamp 1604681595
transform 1 0 3864 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_60
timestamp 1604681595
transform 1 0 6624 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_47
timestamp 1604681595
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_71
timestamp 1604681595
transform 1 0 7636 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_83
timestamp 1604681595
transform 1 0 8740 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_78
timestamp 1604681595
transform 1 0 8280 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _56_
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9200 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10672 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1604681595
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1604681595
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_96
timestamp 1604681595
transform 1 0 9936 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_86
timestamp 1604681595
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_104
timestamp 1604681595
transform 1 0 10672 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_113
timestamp 1604681595
transform 1 0 11500 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_125
timestamp 1604681595
transform 1 0 12604 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_116
timestamp 1604681595
transform 1 0 11776 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_137
timestamp 1604681595
transform 1 0 13708 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1604681595
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1604681595
transform 1 0 14812 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1604681595
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1604681595
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1604681595
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1604681595
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1604681595
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1604681595
transform 1 0 19688 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1604681595
transform 1 0 19504 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1604681595
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_206
timestamp 1604681595
transform 1 0 20056 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_196
timestamp 1604681595
transform 1 0 19136 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_204
timestamp 1604681595
transform 1 0 19872 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_215
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_216
timestamp 1604681595
transform 1 0 20976 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_222
timestamp 1604681595
transform 1 0 21528 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l1_in_0_
timestamp 1604681595
transform 1 0 1840 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_7
timestamp 1604681595
transform 1 0 1748 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_17
timestamp 1604681595
transform 1 0 2668 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4508 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1604681595
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_36
timestamp 1604681595
transform 1 0 4416 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_46
timestamp 1604681595
transform 1 0 5336 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_58
timestamp 1604681595
transform 1 0 6440 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_62
timestamp 1604681595
transform 1 0 6808 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6900 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_8_79
timestamp 1604681595
transform 1 0 8372 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10488 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1604681595
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_101
timestamp 1604681595
transform 1 0 10396 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_118
timestamp 1604681595
transform 1 0 11960 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_130
timestamp 1604681595
transform 1 0 13064 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_142
timestamp 1604681595
transform 1 0 14168 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_150
timestamp 1604681595
transform 1 0 14904 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1604681595
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1604681595
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1604681595
transform 1 0 18952 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_190
timestamp 1604681595
transform 1 0 18584 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_198
timestamp 1604681595
transform 1 0 19320 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_210
timestamp 1604681595
transform 1 0 20424 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1656 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 3864 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_9_22
timestamp 1604681595
transform 1 0 3128 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_46
timestamp 1604681595
transform 1 0 5336 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_58
timestamp 1604681595
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_78
timestamp 1604681595
transform 1 0 8280 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9844 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_9_90
timestamp 1604681595
transform 1 0 9384 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_94
timestamp 1604681595
transform 1 0 9752 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_104
timestamp 1604681595
transform 1 0 10672 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12604 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_116
timestamp 1604681595
transform 1 0 11776 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_134
timestamp 1604681595
transform 1 0 13432 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_146
timestamp 1604681595
transform 1 0 14536 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_158
timestamp 1604681595
transform 1 0 15640 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_170
timestamp 1604681595
transform 1 0 16744 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1604681595
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1604681595
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1604681595
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_220
timestamp 1604681595
transform 1 0 21344 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2208 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_11
timestamp 1604681595
transform 1 0 2116 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_21
timestamp 1604681595
transform 1 0 3036 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1604681595
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_40
timestamp 1604681595
transform 1 0 4784 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4968 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_10_58
timestamp 1604681595
transform 1 0 6440 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1604681595
transform 1 0 7176 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_75
timestamp 1604681595
transform 1 0 8004 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_87
timestamp 1604681595
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1604681595
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_102
timestamp 1604681595
transform 1 0 10488 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12512 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11224 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_116
timestamp 1604681595
transform 1 0 11776 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_140
timestamp 1604681595
transform 1 0 13984 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1604681595
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_157
timestamp 1604681595
transform 1 0 15548 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17756 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_169
timestamp 1604681595
transform 1 0 16652 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_187
timestamp 1604681595
transform 1 0 18308 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_199
timestamp 1604681595
transform 1 0 19412 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_211
timestamp 1604681595
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2024 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_9
timestamp 1604681595
transform 1 0 1932 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_16
timestamp 1604681595
transform 1 0 2576 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3680 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_37
timestamp 1604681595
transform 1 0 4508 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1604681595
transform 1 0 5244 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_48
timestamp 1604681595
transform 1 0 5520 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1604681595
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 8648 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7084 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_74
timestamp 1604681595
transform 1 0 7912 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_91
timestamp 1604681595
transform 1 0 9476 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_103
timestamp 1604681595
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_114
timestamp 1604681595
transform 1 0 11592 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_139
timestamp 1604681595
transform 1 0 13892 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 14628 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_11_163
timestamp 1604681595
transform 1 0 16100 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_175
timestamp 1604681595
transform 1 0 17204 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1604681595
transform 1 0 19320 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_190
timestamp 1604681595
transform 1 0 18584 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_202
timestamp 1604681595
transform 1 0 19688 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_214
timestamp 1604681595
transform 1 0 20792 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_222
timestamp 1604681595
transform 1 0 21528 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1604681595
transform 1 0 2852 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604681595
transform 1 0 1748 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_11
timestamp 1604681595
transform 1 0 2116 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4508 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_22
timestamp 1604681595
transform 1 0 3128 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_30
timestamp 1604681595
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_36
timestamp 1604681595
transform 1 0 4416 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6072 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_46
timestamp 1604681595
transform 1 0 5336 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_57
timestamp 1604681595
transform 1 0 6348 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1604681595
transform 1 0 8556 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6900 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_12_72
timestamp 1604681595
transform 1 0 7728 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_80
timestamp 1604681595
transform 1 0 8464 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_84
timestamp 1604681595
transform 1 0 8832 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12604 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 11868 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_109
timestamp 1604681595
transform 1 0 11132 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_120
timestamp 1604681595
transform 1 0 12144 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_124
timestamp 1604681595
transform 1 0 12512 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1604681595
transform 1 0 14168 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_134
timestamp 1604681595
transform 1 0 13432 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_145
timestamp 1604681595
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_160
timestamp 1604681595
transform 1 0 15824 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16560 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17848 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_174
timestamp 1604681595
transform 1 0 17112 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_188
timestamp 1604681595
transform 1 0 18400 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_200
timestamp 1604681595
transform 1 0 19504 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1604681595
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1748 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_19
timestamp 1604681595
transform 1 0 2852 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 3588 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_23
timestamp 1604681595
transform 1 0 3220 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_40
timestamp 1604681595
transform 1 0 4784 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4968 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_43
timestamp 1604681595
transform 1 0 5060 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_55
timestamp 1604681595
transform 1 0 6164 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_58
timestamp 1604681595
transform 1 0 6440 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8556 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 7176 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_13_71
timestamp 1604681595
transform 1 0 7636 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_79
timestamp 1604681595
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_75
timestamp 1604681595
transform 1 0 8004 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_97
timestamp 1604681595
transform 1 0 10028 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_87
timestamp 1604681595
transform 1 0 9108 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1604681595
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_102
timestamp 1604681595
transform 1 0 10488 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 11224 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_114
timestamp 1604681595
transform 1 0 11592 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_119
timestamp 1604681595
transform 1 0 12052 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13156 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_131
timestamp 1604681595
transform 1 0 13156 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_135
timestamp 1604681595
transform 1 0 13524 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_145
timestamp 1604681595
transform 1 0 14444 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15732 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15824 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_147
timestamp 1604681595
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _87_
timestamp 1604681595
transform 1 0 18216 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17388 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_175
timestamp 1604681595
transform 1 0 17204 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_169
timestamp 1604681595
transform 1 0 16652 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_183
timestamp 1604681595
transform 1 0 17940 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_190
timestamp 1604681595
transform 1 0 18584 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_202
timestamp 1604681595
transform 1 0 19688 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_195
timestamp 1604681595
transform 1 0 19044 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_207
timestamp 1604681595
transform 1 0 20148 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_214
timestamp 1604681595
transform 1 0 20792 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_222
timestamp 1604681595
transform 1 0 21528 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1604681595
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 1564 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_14
timestamp 1604681595
transform 1 0 2392 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1604681595
transform 1 0 3312 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4876 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_22
timestamp 1604681595
transform 1 0 3128 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_33
timestamp 1604681595
transform 1 0 4140 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_50
timestamp 1604681595
transform 1 0 5704 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_78
timestamp 1604681595
transform 1 0 8280 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10028 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_15_89
timestamp 1604681595
transform 1 0 9292 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_113
timestamp 1604681595
transform 1 0 11500 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1604681595
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13340 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_131
timestamp 1604681595
transform 1 0 13156 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_142
timestamp 1604681595
transform 1 0 14168 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 14904 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_15_166
timestamp 1604681595
transform 1 0 16376 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_178
timestamp 1604681595
transform 1 0 17480 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1604681595
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_187
timestamp 1604681595
transform 1 0 18308 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_199
timestamp 1604681595
transform 1 0 19412 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_211
timestamp 1604681595
transform 1 0 20516 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_6
timestamp 1604681595
transform 1 0 1656 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_23
timestamp 1604681595
transform 1 0 3220 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_41
timestamp 1604681595
transform 1 0 4876 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5612 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_58
timestamp 1604681595
transform 1 0 6440 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7176 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_16_82
timestamp 1604681595
transform 1 0 8648 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10396 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1604681595
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12604 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_117
timestamp 1604681595
transform 1 0 11868 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 14168 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_134
timestamp 1604681595
transform 1 0 13432 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_145
timestamp 1604681595
transform 1 0 14444 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16100 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_162
timestamp 1604681595
transform 1 0 16008 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18308 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_179
timestamp 1604681595
transform 1 0 17572 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_193
timestamp 1604681595
transform 1 0 18860 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_205
timestamp 1604681595
transform 1 0 19964 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1604681595
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1604681595
transform 1 0 2944 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_11
timestamp 1604681595
transform 1 0 2116 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_19
timestamp 1604681595
transform 1 0 2852 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4508 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_17_29
timestamp 1604681595
transform 1 0 3772 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_53
timestamp 1604681595
transform 1 0 5980 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8464 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_17_71
timestamp 1604681595
transform 1 0 7636 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_79
timestamp 1604681595
transform 1 0 8372 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10672 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_96
timestamp 1604681595
transform 1 0 9936 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_113
timestamp 1604681595
transform 1 0 11500 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1604681595
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_139
timestamp 1604681595
transform 1 0 13892 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 14628 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16192 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_156
timestamp 1604681595
transform 1 0 15456 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_173
timestamp 1604681595
transform 1 0 17020 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1604681595
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1604681595
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1604681595
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_220
timestamp 1604681595
transform 1 0 21344 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1656 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_22
timestamp 1604681595
transform 1 0 3128 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1604681595
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_41
timestamp 1604681595
transform 1 0 4876 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1604681595
transform 1 0 5612 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 6624 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_52
timestamp 1604681595
transform 1 0 5888 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1604681595
transform 1 0 8280 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8556 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_69
timestamp 1604681595
transform 1 0 7452 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_77
timestamp 1604681595
transform 1 0 8188 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1604681595
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_102
timestamp 1604681595
transform 1 0 10488 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 11224 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_119
timestamp 1604681595
transform 1 0 12052 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12788 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 14352 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_136
timestamp 1604681595
transform 1 0 13616 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_147
timestamp 1604681595
transform 1 0 14628 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 17480 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_170
timestamp 1604681595
transform 1 0 16744 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_184
timestamp 1604681595
transform 1 0 18032 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_196
timestamp 1604681595
transform 1 0 19136 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_208
timestamp 1604681595
transform 1 0 20240 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 1564 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_14
timestamp 1604681595
transform 1 0 2392 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_6
timestamp 1604681595
transform 1 0 1656 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 3128 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4784 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_38
timestamp 1604681595
transform 1 0 4600 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_23
timestamp 1604681595
transform 1 0 3220 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 5336 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1604681595
transform 1 0 6440 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_50
timestamp 1604681595
transform 1 0 5704 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_56
timestamp 1604681595
transform 1 0 6256 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1604681595
transform 1 0 8556 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6992 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 6992 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8740 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_8  FILLER_19_73
timestamp 1604681595
transform 1 0 7820 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_81
timestamp 1604681595
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_73
timestamp 1604681595
transform 1 0 7820 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10580 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_84
timestamp 1604681595
transform 1 0 8832 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_102
timestamp 1604681595
transform 1 0 10488 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11776 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 11224 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_112
timestamp 1604681595
transform 1 0 11408 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1604681595
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_113
timestamp 1604681595
transform 1 0 11500 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1604681595
transform 1 0 14168 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13524 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_19_126
timestamp 1604681595
transform 1 0 12696 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_134
timestamp 1604681595
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_132
timestamp 1604681595
transform 1 0 13248 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_140
timestamp 1604681595
transform 1 0 13984 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_145
timestamp 1604681595
transform 1 0 14444 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15732 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_151
timestamp 1604681595
transform 1 0 14996 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_160
timestamp 1604681595
transform 1 0 15824 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_168
timestamp 1604681595
transform 1 0 16560 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_180
timestamp 1604681595
transform 1 0 17664 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_172
timestamp 1604681595
transform 1 0 16928 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_184
timestamp 1604681595
transform 1 0 18032 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1604681595
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1604681595
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_196
timestamp 1604681595
transform 1 0 19136 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_208
timestamp 1604681595
transform 1 0 20240 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_220
timestamp 1604681595
transform 1 0 21344 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 1840 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1604681595
transform 1 0 1748 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4324 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 4048 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_24
timestamp 1604681595
transform 1 0 3312 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_71
timestamp 1604681595
transform 1 0 7636 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_83
timestamp 1604681595
transform 1 0 8740 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9200 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_87
timestamp 1604681595
transform 1 0 9108 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_104
timestamp 1604681595
transform 1 0 10672 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_116
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_132
timestamp 1604681595
transform 1 0 13248 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_144
timestamp 1604681595
transform 1 0 14352 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16008 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14720 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_154
timestamp 1604681595
transform 1 0 15272 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_168
timestamp 1604681595
transform 1 0 16560 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_180
timestamp 1604681595
transform 1 0 17664 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1604681595
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1604681595
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_220
timestamp 1604681595
transform 1 0 21344 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _52_
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_6
timestamp 1604681595
transform 1 0 1656 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_23
timestamp 1604681595
transform 1 0 3220 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_36
timestamp 1604681595
transform 1 0 4416 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6440 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_22_48
timestamp 1604681595
transform 1 0 5520 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_56
timestamp 1604681595
transform 1 0 6256 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8280 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_67
timestamp 1604681595
transform 1 0 7268 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_75
timestamp 1604681595
transform 1 0 8004 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10672 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_84
timestamp 1604681595
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_96
timestamp 1604681595
transform 1 0 9936 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_120
timestamp 1604681595
transform 1 0 12144 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13432 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_132
timestamp 1604681595
transform 1 0 13248 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_140
timestamp 1604681595
transform 1 0 13984 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1604681595
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_160
timestamp 1604681595
transform 1 0 15824 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _94_
timestamp 1604681595
transform 1 0 16560 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_172
timestamp 1604681595
transform 1 0 16928 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_184
timestamp 1604681595
transform 1 0 18032 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_196
timestamp 1604681595
transform 1 0 19136 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_208
timestamp 1604681595
transform 1 0 20240 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 1748 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_11
timestamp 1604681595
transform 1 0 2116 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_19
timestamp 1604681595
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4600 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3036 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_30
timestamp 1604681595
transform 1 0 3864 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _51_
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_47
timestamp 1604681595
transform 1 0 5428 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_58
timestamp 1604681595
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7820 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_23_65
timestamp 1604681595
transform 1 0 7084 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_89
timestamp 1604681595
transform 1 0 9292 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_101
timestamp 1604681595
transform 1 0 10396 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_114
timestamp 1604681595
transform 1 0 11592 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_139
timestamp 1604681595
transform 1 0 13892 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 14628 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_23_163
timestamp 1604681595
transform 1 0 16100 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _59_
timestamp 1604681595
transform 1 0 16836 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_174
timestamp 1604681595
transform 1 0 17112 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1604681595
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1604681595
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1604681595
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_220
timestamp 1604681595
transform 1 0 21344 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2208 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_11
timestamp 1604681595
transform 1 0 2116 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_18
timestamp 1604681595
transform 1 0 2760 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4876 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_30
timestamp 1604681595
transform 1 0 3864 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_40
timestamp 1604681595
transform 1 0 4784 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_57
timestamp 1604681595
transform 1 0 6348 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7084 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_81
timestamp 1604681595
transform 1 0 8556 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_89
timestamp 1604681595
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_102
timestamp 1604681595
transform 1 0 10488 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11592 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 11316 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_110
timestamp 1604681595
transform 1 0 11224 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_123
timestamp 1604681595
transform 1 0 12420 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13156 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_24_140
timestamp 1604681595
transform 1 0 13984 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _93_
timestamp 1604681595
transform 1 0 15456 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_152
timestamp 1604681595
transform 1 0 15088 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_160
timestamp 1604681595
transform 1 0 15824 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_172
timestamp 1604681595
transform 1 0 16928 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_184
timestamp 1604681595
transform 1 0 18032 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_196
timestamp 1604681595
transform 1 0 19136 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_208
timestamp 1604681595
transform 1 0 20240 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2116 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_17
timestamp 1604681595
transform 1 0 2668 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 3772 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_45
timestamp 1604681595
transform 1 0 5244 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1604681595
transform 1 0 6348 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 8464 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_25_71
timestamp 1604681595
transform 1 0 7636 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_79
timestamp 1604681595
transform 1 0 8372 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_96
timestamp 1604681595
transform 1 0 9936 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_104
timestamp 1604681595
transform 1 0 10672 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_114
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13708 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_25_129
timestamp 1604681595
transform 1 0 12972 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _58_
timestamp 1604681595
transform 1 0 15916 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_153
timestamp 1604681595
transform 1 0 15180 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_164
timestamp 1604681595
transform 1 0 16192 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_176
timestamp 1604681595
transform 1 0 17296 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1604681595
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1604681595
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1604681595
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_220
timestamp 1604681595
transform 1 0 21344 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2116 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2116 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_17
timestamp 1604681595
transform 1 0 2668 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_17
timestamp 1604681595
transform 1 0 2668 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 3956 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1604681595
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_41
timestamp 1604681595
transform 1 0 4876 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_29
timestamp 1604681595
transform 1 0 3772 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 5612 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604681595
transform 1 0 6808 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 6164 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_53
timestamp 1604681595
transform 1 0 5980 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_61
timestamp 1604681595
transform 1 0 6716 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 1604681595
transform 1 0 5428 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_58
timestamp 1604681595
transform 1 0 6440 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 8372 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_71
timestamp 1604681595
transform 1 0 7636 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_83
timestamp 1604681595
transform 1 0 8740 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_78
timestamp 1604681595
transform 1 0 8280 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 9016 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1604681595
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_99
timestamp 1604681595
transform 1 0 10212 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_102
timestamp 1604681595
transform 1 0 10488 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604681595
transform 1 0 11224 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11224 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 10948 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_114
timestamp 1604681595
transform 1 0 11592 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 14076 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_26_126
timestamp 1604681595
transform 1 0 12696 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_134
timestamp 1604681595
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_145
timestamp 1604681595
transform 1 0 14444 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_132
timestamp 1604681595
transform 1 0 13248 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_140
timestamp 1604681595
transform 1 0 13984 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604681595
transform 1 0 16284 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_163
timestamp 1604681595
transform 1 0 16100 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_157
timestamp 1604681595
transform 1 0 15548 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_175
timestamp 1604681595
transform 1 0 17204 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_187
timestamp 1604681595
transform 1 0 18308 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_168
timestamp 1604681595
transform 1 0 16560 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_180
timestamp 1604681595
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_199
timestamp 1604681595
transform 1 0 19412 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1604681595
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1604681595
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_211
timestamp 1604681595
transform 1 0 20516 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_220
timestamp 1604681595
transform 1 0 21344 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2208 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_11
timestamp 1604681595
transform 1 0 2116 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_18
timestamp 1604681595
transform 1 0 2760 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_30
timestamp 1604681595
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 6808 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_28_48
timestamp 1604681595
transform 1 0 5520 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_60
timestamp 1604681595
transform 1 0 6624 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_78
timestamp 1604681595
transform 1 0 8280 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1604681595
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_102
timestamp 1604681595
transform 1 0 10488 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11500 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 11224 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13708 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_129
timestamp 1604681595
transform 1 0 12972 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_143
timestamp 1604681595
transform 1 0 14260 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1604681595
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_160
timestamp 1604681595
transform 1 0 15824 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _50_
timestamp 1604681595
transform 1 0 16560 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_171
timestamp 1604681595
transform 1 0 16836 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_183
timestamp 1604681595
transform 1 0 17940 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_195
timestamp 1604681595
transform 1 0 19044 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_207
timestamp 1604681595
transform 1 0 20148 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1604681595
transform 1 0 20700 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2944 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1604681595
transform 1 0 2760 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_11
timestamp 1604681595
transform 1 0 2116 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_17
timestamp 1604681595
transform 1 0 2668 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4508 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_29
timestamp 1604681595
transform 1 0 3772 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_46
timestamp 1604681595
transform 1 0 5336 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_58
timestamp 1604681595
transform 1 0 6440 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8556 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_29_71
timestamp 1604681595
transform 1 0 7636 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_79
timestamp 1604681595
transform 1 0 8372 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_90
timestamp 1604681595
transform 1 0 9384 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_102
timestamp 1604681595
transform 1 0 10488 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 12512 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_114
timestamp 1604681595
transform 1 0 11592 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 14260 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_29_133
timestamp 1604681595
transform 1 0 13340 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_141
timestamp 1604681595
transform 1 0 14076 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_159
timestamp 1604681595
transform 1 0 15732 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _49_
timestamp 1604681595
transform 1 0 16468 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _57_
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1604681595
transform 1 0 18308 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_170
timestamp 1604681595
transform 1 0 16744 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_182
timestamp 1604681595
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_189
timestamp 1604681595
transform 1 0 18492 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_201
timestamp 1604681595
transform 1 0 19596 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_213
timestamp 1604681595
transform 1 0 20700 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1604681595
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _53_
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_6
timestamp 1604681595
transform 1 0 1656 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_23
timestamp 1604681595
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_38
timestamp 1604681595
transform 1 0 4600 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5428 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_30_46
timestamp 1604681595
transform 1 0 5336 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1604681595
transform 1 0 7636 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_30_63
timestamp 1604681595
transform 1 0 6900 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1604681595
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _48_
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 10672 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_96
timestamp 1604681595
transform 1 0 9936 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_120
timestamp 1604681595
transform 1 0 12144 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 12880 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_30_137
timestamp 1604681595
transform 1 0 13708 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _92_
timestamp 1604681595
transform 1 0 16376 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _97_
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_149
timestamp 1604681595
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_158
timestamp 1604681595
transform 1 0 15640 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _90_
timestamp 1604681595
transform 1 0 17480 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_170
timestamp 1604681595
transform 1 0 16744 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_182
timestamp 1604681595
transform 1 0 17848 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_194
timestamp 1604681595
transform 1 0 18952 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_206
timestamp 1604681595
transform 1 0 20056 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 2852 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_11
timestamp 1604681595
transform 1 0 2116 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_35
timestamp 1604681595
transform 1 0 4324 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5152 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_43
timestamp 1604681595
transform 1 0 5060 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_53
timestamp 1604681595
transform 1 0 5980 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 7728 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_70
timestamp 1604681595
transform 1 0 7544 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10028 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_31_88
timestamp 1604681595
transform 1 0 9200 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_96
timestamp 1604681595
transform 1 0 9936 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_106
timestamp 1604681595
transform 1 0 10856 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_118
timestamp 1604681595
transform 1 0 11960 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 13156 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 15364 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_31_147
timestamp 1604681595
transform 1 0 14628 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _91_
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1604681595
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _55_
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_188
timestamp 1604681595
transform 1 0 18400 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_199
timestamp 1604681595
transform 1 0 19412 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_211
timestamp 1604681595
transform 1 0 20516 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_7
timestamp 1604681595
transform 1 0 1748 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_21
timestamp 1604681595
transform 1 0 3036 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1604681595
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_36
timestamp 1604681595
transform 1 0 4416 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5244 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_32_44
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_61
timestamp 1604681595
transform 1 0 6716 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7636 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_32_69
timestamp 1604681595
transform 1 0 7452 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1604681595
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 11868 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_32_109
timestamp 1604681595
transform 1 0 11132 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 14076 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_133
timestamp 1604681595
transform 1 0 13340 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_145
timestamp 1604681595
transform 1 0 14444 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _98_
timestamp 1604681595
transform 1 0 16376 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_158
timestamp 1604681595
transform 1 0 15640 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _95_
timestamp 1604681595
transform 1 0 17480 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_170
timestamp 1604681595
transform 1 0 16744 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_182
timestamp 1604681595
transform 1 0 17848 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _54_
timestamp 1604681595
transform 1 0 19688 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _89_
timestamp 1604681595
transform 1 0 18584 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_194
timestamp 1604681595
transform 1 0 18952 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_205
timestamp 1604681595
transform 1 0 19964 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1604681595
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2116 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_17
timestamp 1604681595
transform 1 0 2668 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 4048 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 3956 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_29
timestamp 1604681595
transform 1 0 3772 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_36
timestamp 1604681595
transform 1 0 4416 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5244 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_44
timestamp 1604681595
transform 1 0 5152 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_54
timestamp 1604681595
transform 1 0 6072 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 6900 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8372 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_67
timestamp 1604681595
transform 1 0 7268 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10212 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9660 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_85
timestamp 1604681595
transform 1 0 8924 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_94
timestamp 1604681595
transform 1 0 9752 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_98
timestamp 1604681595
transform 1 0 10120 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 12604 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 12512 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_108
timestamp 1604681595
transform 1 0 11040 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_120
timestamp 1604681595
transform 1 0 12144 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 13708 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_129
timestamp 1604681595
transform 1 0 12972 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_141
timestamp 1604681595
transform 1 0 14076 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _99_
timestamp 1604681595
transform 1 0 15456 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 15364 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_153
timestamp 1604681595
transform 1 0 15180 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_160
timestamp 1604681595
transform 1 0 15824 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _88_
timestamp 1604681595
transform 1 0 18308 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _96_
timestamp 1604681595
transform 1 0 16560 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 18216 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_172
timestamp 1604681595
transform 1 0 16928 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_184
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_191
timestamp 1604681595
transform 1 0 18676 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_203
timestamp 1604681595
transform 1 0 19780 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 21896 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 21068 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_215
timestamp 1604681595
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_218
timestamp 1604681595
transform 1 0 21160 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_222
timestamp 1604681595
transform 1 0 21528 0 1 20128
box -38 -48 130 592
<< labels >>
rlabel metal3 s 22520 11432 23000 11552 6 ccff_head
port 0 nsew default input
rlabel metal2 s 17222 0 17278 480 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 0 3136 480 3256 6 chanx_left_in[0]
port 2 nsew default input
rlabel metal3 s 0 8032 480 8152 6 chanx_left_in[10]
port 3 nsew default input
rlabel metal3 s 0 8576 480 8696 6 chanx_left_in[11]
port 4 nsew default input
rlabel metal3 s 0 9120 480 9240 6 chanx_left_in[12]
port 5 nsew default input
rlabel metal3 s 0 9528 480 9648 6 chanx_left_in[13]
port 6 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[14]
port 7 nsew default input
rlabel metal3 s 0 10616 480 10736 6 chanx_left_in[15]
port 8 nsew default input
rlabel metal3 s 0 11024 480 11144 6 chanx_left_in[16]
port 9 nsew default input
rlabel metal3 s 0 11568 480 11688 6 chanx_left_in[17]
port 10 nsew default input
rlabel metal3 s 0 12112 480 12232 6 chanx_left_in[18]
port 11 nsew default input
rlabel metal3 s 0 12520 480 12640 6 chanx_left_in[19]
port 12 nsew default input
rlabel metal3 s 0 3544 480 3664 6 chanx_left_in[1]
port 13 nsew default input
rlabel metal3 s 0 4088 480 4208 6 chanx_left_in[2]
port 14 nsew default input
rlabel metal3 s 0 4632 480 4752 6 chanx_left_in[3]
port 15 nsew default input
rlabel metal3 s 0 5040 480 5160 6 chanx_left_in[4]
port 16 nsew default input
rlabel metal3 s 0 5584 480 5704 6 chanx_left_in[5]
port 17 nsew default input
rlabel metal3 s 0 6128 480 6248 6 chanx_left_in[6]
port 18 nsew default input
rlabel metal3 s 0 6536 480 6656 6 chanx_left_in[7]
port 19 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[8]
port 20 nsew default input
rlabel metal3 s 0 7624 480 7744 6 chanx_left_in[9]
port 21 nsew default input
rlabel metal3 s 0 13064 480 13184 6 chanx_left_out[0]
port 22 nsew default tristate
rlabel metal3 s 0 18096 480 18216 6 chanx_left_out[10]
port 23 nsew default tristate
rlabel metal3 s 0 18504 480 18624 6 chanx_left_out[11]
port 24 nsew default tristate
rlabel metal3 s 0 19048 480 19168 6 chanx_left_out[12]
port 25 nsew default tristate
rlabel metal3 s 0 19592 480 19712 6 chanx_left_out[13]
port 26 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 chanx_left_out[14]
port 27 nsew default tristate
rlabel metal3 s 0 20544 480 20664 6 chanx_left_out[15]
port 28 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[16]
port 29 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[17]
port 30 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[18]
port 31 nsew default tristate
rlabel metal3 s 0 22584 480 22704 6 chanx_left_out[19]
port 32 nsew default tristate
rlabel metal3 s 0 13608 480 13728 6 chanx_left_out[1]
port 33 nsew default tristate
rlabel metal3 s 0 14016 480 14136 6 chanx_left_out[2]
port 34 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[3]
port 35 nsew default tristate
rlabel metal3 s 0 15104 480 15224 6 chanx_left_out[4]
port 36 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[5]
port 37 nsew default tristate
rlabel metal3 s 0 16056 480 16176 6 chanx_left_out[6]
port 38 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 chanx_left_out[7]
port 39 nsew default tristate
rlabel metal3 s 0 17008 480 17128 6 chanx_left_out[8]
port 40 nsew default tristate
rlabel metal3 s 0 17552 480 17672 6 chanx_left_out[9]
port 41 nsew default tristate
rlabel metal2 s 3882 22520 3938 23000 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 8574 22520 8630 23000 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 9034 22520 9090 23000 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 9586 22520 9642 23000 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 10046 22520 10102 23000 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 10506 22520 10562 23000 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 10966 22520 11022 23000 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 11426 22520 11482 23000 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 11886 22520 11942 23000 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 12346 22520 12402 23000 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 12806 22520 12862 23000 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 4342 22520 4398 23000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 4894 22520 4950 23000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 5354 22520 5410 23000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 5814 22520 5870 23000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 6274 22520 6330 23000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 6734 22520 6790 23000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 7194 22520 7250 23000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 7654 22520 7710 23000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 8114 22520 8170 23000 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 13266 22520 13322 23000 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 17958 22520 18014 23000 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 18418 22520 18474 23000 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 18970 22520 19026 23000 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 19430 22520 19486 23000 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 19890 22520 19946 23000 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 20350 22520 20406 23000 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 20810 22520 20866 23000 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 21270 22520 21326 23000 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 21730 22520 21786 23000 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 22190 22520 22246 23000 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 13726 22520 13782 23000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 14278 22520 14334 23000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 14738 22520 14794 23000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 15198 22520 15254 23000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 15658 22520 15714 23000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 16118 22520 16174 23000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 16578 22520 16634 23000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 17038 22520 17094 23000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 17498 22520 17554 23000 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 left_bottom_grid_pin_11_
port 82 nsew default input
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_1_
port 83 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_3_
port 84 nsew default input
rlabel metal3 s 0 1096 480 1216 6 left_bottom_grid_pin_5_
port 85 nsew default input
rlabel metal3 s 0 1640 480 1760 6 left_bottom_grid_pin_7_
port 86 nsew default input
rlabel metal3 s 0 2048 480 2168 6 left_bottom_grid_pin_9_
port 87 nsew default input
rlabel metal2 s 5722 0 5778 480 6 prog_clk
port 88 nsew default input
rlabel metal2 s 202 22520 258 23000 6 top_left_grid_pin_42_
port 89 nsew default input
rlabel metal2 s 662 22520 718 23000 6 top_left_grid_pin_43_
port 90 nsew default input
rlabel metal2 s 1122 22520 1178 23000 6 top_left_grid_pin_44_
port 91 nsew default input
rlabel metal2 s 1582 22520 1638 23000 6 top_left_grid_pin_45_
port 92 nsew default input
rlabel metal2 s 2042 22520 2098 23000 6 top_left_grid_pin_46_
port 93 nsew default input
rlabel metal2 s 2502 22520 2558 23000 6 top_left_grid_pin_47_
port 94 nsew default input
rlabel metal2 s 2962 22520 3018 23000 6 top_left_grid_pin_48_
port 95 nsew default input
rlabel metal2 s 3422 22520 3478 23000 6 top_left_grid_pin_49_
port 96 nsew default input
rlabel metal2 s 22650 22520 22706 23000 6 top_right_grid_pin_1_
port 97 nsew default input
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 98 nsew default input
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 99 nsew default input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
