VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_1__1_
  CLASS BLOCK ;
  FOREIGN sb_1__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 140.000 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 2.400 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 2.400 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 2.400 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 2.400 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 2.400 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 2.400 ;
    END
  END address[5]
  PIN address[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 2.400 ;
    END
  END address[6]
  PIN bottom_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 2.400 ;
    END
  END bottom_left_grid_pin_13_
  PIN bottom_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 2.400 ;
    END
  END bottom_right_grid_pin_11_
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 2.400 10.840 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 2.400 17.640 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 2.400 24.440 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 2.400 31.920 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 2.400 38.720 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 2.400 45.520 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 2.400 53.000 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 2.400 59.800 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 2.400 66.600 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 2.400 80.880 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 2.400 87.680 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 2.400 94.480 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 2.400 101.960 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 2.400 108.760 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 2.400 115.560 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 2.400 123.040 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 2.400 129.840 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 2.400 136.640 ;
    END
  END chanx_left_out[8]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 10.240 140.000 10.840 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 17.040 140.000 17.640 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 23.840 140.000 24.440 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 31.320 140.000 31.920 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 38.120 140.000 38.720 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 44.920 140.000 45.520 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 52.400 140.000 53.000 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 59.200 140.000 59.800 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 66.000 140.000 66.600 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 80.280 140.000 80.880 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 87.080 140.000 87.680 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 93.880 140.000 94.480 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 101.360 140.000 101.960 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 108.160 140.000 108.760 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 114.960 140.000 115.560 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 122.440 140.000 123.040 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 129.240 140.000 129.840 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 137.600 136.040 140.000 136.640 ;
    END
  END chanx_right_out[8]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 2.400 ;
    END
  END chany_bottom_out[8]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.310 137.600 3.590 140.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 137.600 10.490 140.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 137.600 17.390 140.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 137.600 24.290 140.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.910 137.600 31.190 140.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.270 137.600 38.550 140.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.170 137.600 45.450 140.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.070 137.600 52.350 140.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 137.600 59.250 140.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.130 137.600 80.410 140.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.030 137.600 87.310 140.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.930 137.600 94.210 140.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.830 137.600 101.110 140.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.190 137.600 108.470 140.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.090 137.600 115.370 140.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.990 137.600 122.270 140.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 128.890 137.600 129.170 140.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.790 137.600 136.070 140.000 ;
    END
  END chany_top_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 2.400 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 2.400 ;
    END
  END enable
  PIN left_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 2.400 74.080 ;
    END
  END left_bottom_grid_pin_12_
  PIN left_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 2.400 4.040 ;
    END
  END left_top_grid_pin_10_
  PIN right_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 73.480 140.000 74.080 ;
    END
  END right_bottom_grid_pin_12_
  PIN right_top_grid_pin_10_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 137.600 3.440 140.000 4.040 ;
    END
  END right_top_grid_pin_10_
  PIN top_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.870 137.600 66.150 140.000 ;
    END
  END top_left_grid_pin_13_
  PIN top_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.230 137.600 73.510 140.000 ;
    END
  END top_right_grid_pin_11_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 28.055 10.640 29.655 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 51.385 10.640 52.985 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 4.745 10.795 134.320 127.925 ;
      LAYER met1 ;
        RECT 0.530 0.380 138.850 137.660 ;
      LAYER met2 ;
        RECT 0.550 137.320 3.030 137.770 ;
        RECT 3.870 137.320 9.930 137.770 ;
        RECT 10.770 137.320 16.830 137.770 ;
        RECT 17.670 137.320 23.730 137.770 ;
        RECT 24.570 137.320 30.630 137.770 ;
        RECT 31.470 137.320 37.990 137.770 ;
        RECT 38.830 137.320 44.890 137.770 ;
        RECT 45.730 137.320 51.790 137.770 ;
        RECT 52.630 137.320 58.690 137.770 ;
        RECT 59.530 137.320 65.590 137.770 ;
        RECT 66.430 137.320 72.950 137.770 ;
        RECT 73.790 137.320 79.850 137.770 ;
        RECT 80.690 137.320 86.750 137.770 ;
        RECT 87.590 137.320 93.650 137.770 ;
        RECT 94.490 137.320 100.550 137.770 ;
        RECT 101.390 137.320 107.910 137.770 ;
        RECT 108.750 137.320 114.810 137.770 ;
        RECT 115.650 137.320 121.710 137.770 ;
        RECT 122.550 137.320 128.610 137.770 ;
        RECT 129.450 137.320 135.510 137.770 ;
        RECT 136.350 137.320 138.830 137.770 ;
        RECT 0.550 2.680 138.830 137.320 ;
        RECT 0.550 0.155 2.110 2.680 ;
        RECT 2.950 0.155 6.710 2.680 ;
        RECT 7.550 0.155 11.310 2.680 ;
        RECT 12.150 0.155 16.370 2.680 ;
        RECT 17.210 0.155 20.970 2.680 ;
        RECT 21.810 0.155 26.030 2.680 ;
        RECT 26.870 0.155 30.630 2.680 ;
        RECT 31.470 0.155 35.690 2.680 ;
        RECT 36.530 0.155 40.290 2.680 ;
        RECT 41.130 0.155 45.350 2.680 ;
        RECT 46.190 0.155 49.950 2.680 ;
        RECT 50.790 0.155 55.010 2.680 ;
        RECT 55.850 0.155 59.610 2.680 ;
        RECT 60.450 0.155 64.670 2.680 ;
        RECT 65.510 0.155 69.270 2.680 ;
        RECT 70.110 0.155 74.330 2.680 ;
        RECT 75.170 0.155 78.930 2.680 ;
        RECT 79.770 0.155 83.990 2.680 ;
        RECT 84.830 0.155 88.590 2.680 ;
        RECT 89.430 0.155 93.650 2.680 ;
        RECT 94.490 0.155 98.250 2.680 ;
        RECT 99.090 0.155 103.310 2.680 ;
        RECT 104.150 0.155 107.910 2.680 ;
        RECT 108.750 0.155 112.970 2.680 ;
        RECT 113.810 0.155 117.570 2.680 ;
        RECT 118.410 0.155 122.630 2.680 ;
        RECT 123.470 0.155 127.230 2.680 ;
        RECT 128.070 0.155 132.290 2.680 ;
        RECT 133.130 0.155 136.890 2.680 ;
        RECT 137.730 0.155 138.830 2.680 ;
      LAYER met3 ;
        RECT 2.800 135.640 137.200 136.040 ;
        RECT 0.270 130.240 138.650 135.640 ;
        RECT 2.800 128.840 137.200 130.240 ;
        RECT 0.270 123.440 138.650 128.840 ;
        RECT 2.800 122.040 137.200 123.440 ;
        RECT 0.270 115.960 138.650 122.040 ;
        RECT 2.800 114.560 137.200 115.960 ;
        RECT 0.270 109.160 138.650 114.560 ;
        RECT 2.800 107.760 137.200 109.160 ;
        RECT 0.270 102.360 138.650 107.760 ;
        RECT 2.800 100.960 137.200 102.360 ;
        RECT 0.270 94.880 138.650 100.960 ;
        RECT 2.800 93.480 137.200 94.880 ;
        RECT 0.270 88.080 138.650 93.480 ;
        RECT 2.800 86.680 137.200 88.080 ;
        RECT 0.270 81.280 138.650 86.680 ;
        RECT 2.800 79.880 137.200 81.280 ;
        RECT 0.270 74.480 138.650 79.880 ;
        RECT 2.800 73.080 137.200 74.480 ;
        RECT 0.270 67.000 138.650 73.080 ;
        RECT 2.800 65.600 137.200 67.000 ;
        RECT 0.270 60.200 138.650 65.600 ;
        RECT 2.800 58.800 137.200 60.200 ;
        RECT 0.270 53.400 138.650 58.800 ;
        RECT 2.800 52.000 137.200 53.400 ;
        RECT 0.270 45.920 138.650 52.000 ;
        RECT 2.800 44.520 137.200 45.920 ;
        RECT 0.270 39.120 138.650 44.520 ;
        RECT 2.800 37.720 137.200 39.120 ;
        RECT 0.270 32.320 138.650 37.720 ;
        RECT 2.800 30.920 137.200 32.320 ;
        RECT 0.270 24.840 138.650 30.920 ;
        RECT 2.800 23.440 137.200 24.840 ;
        RECT 0.270 18.040 138.650 23.440 ;
        RECT 2.800 16.640 137.200 18.040 ;
        RECT 0.270 11.240 138.650 16.640 ;
        RECT 2.800 9.840 137.200 11.240 ;
        RECT 0.270 4.440 138.650 9.840 ;
        RECT 2.800 3.040 137.200 4.440 ;
        RECT 0.270 0.175 138.650 3.040 ;
      LAYER met4 ;
        RECT 0.295 10.375 27.655 128.080 ;
        RECT 30.055 10.375 50.985 128.080 ;
        RECT 53.385 10.375 138.625 128.080 ;
  END
END sb_1__1_
END LIBRARY

