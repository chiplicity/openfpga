magic
tech EFS8A
magscale 1 2
timestamp 1603801476
<< locali >>
rect 9781 12223 9815 12393
rect 10057 11067 10091 11169
rect 12081 3927 12115 4233
<< viali >>
rect 13864 25313 13898 25347
rect 13967 25109 14001 25143
rect 16681 24769 16715 24803
rect 10676 24701 10710 24735
rect 13921 24701 13955 24735
rect 14473 24701 14507 24735
rect 15025 24701 15059 24735
rect 15577 24701 15611 24735
rect 16196 24701 16230 24735
rect 13829 24633 13863 24667
rect 10747 24565 10781 24599
rect 11161 24565 11195 24599
rect 14105 24565 14139 24599
rect 15209 24565 15243 24599
rect 16267 24565 16301 24599
rect 10149 24361 10183 24395
rect 11897 24361 11931 24395
rect 13001 24361 13035 24395
rect 14197 24361 14231 24395
rect 17049 24361 17083 24395
rect 15485 24293 15519 24327
rect 9965 24225 9999 24259
rect 11713 24225 11747 24259
rect 12817 24225 12851 24259
rect 14013 24225 14047 24259
rect 16865 24225 16899 24259
rect 18312 24225 18346 24259
rect 15393 24157 15427 24191
rect 16037 24157 16071 24191
rect 16405 24089 16439 24123
rect 12633 24021 12667 24055
rect 18383 24021 18417 24055
rect 3617 23817 3651 23851
rect 7941 23817 7975 23851
rect 9137 23817 9171 23851
rect 10701 23817 10735 23851
rect 15393 23817 15427 23851
rect 18245 23817 18279 23851
rect 20821 23817 20855 23851
rect 24547 23817 24581 23851
rect 24961 23817 24995 23851
rect 16313 23749 16347 23783
rect 18613 23749 18647 23783
rect 1869 23681 1903 23715
rect 12265 23681 12299 23715
rect 14197 23681 14231 23715
rect 14473 23681 14507 23715
rect 15761 23681 15795 23715
rect 19303 23681 19337 23715
rect 1444 23613 1478 23647
rect 1547 23613 1581 23647
rect 3132 23613 3166 23647
rect 7456 23613 7490 23647
rect 8652 23613 8686 23647
rect 10149 23613 10183 23647
rect 11412 23613 11446 23647
rect 12725 23613 12759 23647
rect 13001 23613 13035 23647
rect 17877 23613 17911 23647
rect 18061 23613 18095 23647
rect 19216 23613 19250 23647
rect 20336 23613 20370 23647
rect 24476 23613 24510 23647
rect 13277 23545 13311 23579
rect 14013 23545 14047 23579
rect 14289 23545 14323 23579
rect 15853 23545 15887 23579
rect 3203 23477 3237 23511
rect 7527 23477 7561 23511
rect 8723 23477 8757 23511
rect 9965 23477 9999 23511
rect 10333 23477 10367 23511
rect 11483 23477 11517 23511
rect 11897 23477 11931 23511
rect 13553 23477 13587 23511
rect 16865 23477 16899 23511
rect 19625 23477 19659 23511
rect 20407 23477 20441 23511
rect 13829 23273 13863 23307
rect 14197 23273 14231 23307
rect 15117 23273 15151 23307
rect 17003 23273 17037 23307
rect 9873 23205 9907 23239
rect 11161 23205 11195 23239
rect 11345 23205 11379 23239
rect 11437 23205 11471 23239
rect 13001 23205 13035 23239
rect 13553 23205 13587 23239
rect 14657 23205 14691 23239
rect 15485 23205 15519 23239
rect 18797 23205 18831 23239
rect 16900 23137 16934 23171
rect 20980 23137 21014 23171
rect 24660 23137 24694 23171
rect 9781 23069 9815 23103
rect 10425 23069 10459 23103
rect 11621 23069 11655 23103
rect 12909 23069 12943 23103
rect 15393 23069 15427 23103
rect 18705 23069 18739 23103
rect 15945 23001 15979 23035
rect 19257 23001 19291 23035
rect 21051 23001 21085 23035
rect 12633 22933 12667 22967
rect 16313 22933 16347 22967
rect 24731 22933 24765 22967
rect 10057 22729 10091 22763
rect 12265 22729 12299 22763
rect 14565 22729 14599 22763
rect 14933 22729 14967 22763
rect 16405 22729 16439 22763
rect 17141 22729 17175 22763
rect 17877 22729 17911 22763
rect 19809 22729 19843 22763
rect 20177 22729 20211 22763
rect 21005 22729 21039 22763
rect 24685 22729 24719 22763
rect 15301 22661 15335 22695
rect 16037 22661 16071 22695
rect 16773 22661 16807 22695
rect 10517 22593 10551 22627
rect 13461 22593 13495 22627
rect 13645 22593 13679 22627
rect 15485 22593 15519 22627
rect 18797 22593 18831 22627
rect 19257 22593 19291 22627
rect 10609 22525 10643 22559
rect 12516 22525 12550 22559
rect 12909 22525 12943 22559
rect 20304 22525 20338 22559
rect 10950 22457 10984 22491
rect 11805 22457 11839 22491
rect 13966 22457 14000 22491
rect 15577 22457 15611 22491
rect 18889 22457 18923 22491
rect 20407 22457 20441 22491
rect 9781 22389 9815 22423
rect 11529 22389 11563 22423
rect 12587 22389 12621 22423
rect 18521 22389 18555 22423
rect 12909 22185 12943 22219
rect 18061 22185 18095 22219
rect 11253 22117 11287 22151
rect 11345 22117 11379 22151
rect 13737 22117 13771 22151
rect 16221 22117 16255 22151
rect 17503 22117 17537 22151
rect 18797 22117 18831 22151
rect 19073 22117 19107 22151
rect 14289 22049 14323 22083
rect 15485 22049 15519 22083
rect 16037 22049 16071 22083
rect 11897 21981 11931 22015
rect 13645 21981 13679 22015
rect 17141 21981 17175 22015
rect 18981 21981 19015 22015
rect 19441 21981 19475 22015
rect 8493 21845 8527 21879
rect 10609 21845 10643 21879
rect 14565 21845 14599 21879
rect 16497 21845 16531 21879
rect 10885 21641 10919 21675
rect 11529 21641 11563 21675
rect 12817 21641 12851 21675
rect 13829 21641 13863 21675
rect 19625 21641 19659 21675
rect 9137 21505 9171 21539
rect 11253 21505 11287 21539
rect 13047 21505 13081 21539
rect 14013 21505 14047 21539
rect 14381 21505 14415 21539
rect 16681 21505 16715 21539
rect 17509 21505 17543 21539
rect 18521 21505 18555 21539
rect 19349 21505 19383 21539
rect 19993 21505 20027 21539
rect 8401 21437 8435 21471
rect 8953 21437 8987 21471
rect 9965 21437 9999 21471
rect 12960 21437 12994 21471
rect 15761 21437 15795 21471
rect 15945 21437 15979 21471
rect 16497 21437 16531 21471
rect 9873 21369 9907 21403
rect 10327 21369 10361 21403
rect 14105 21369 14139 21403
rect 15117 21369 15151 21403
rect 18705 21369 18739 21403
rect 18797 21369 18831 21403
rect 8309 21301 8343 21335
rect 13461 21301 13495 21335
rect 15393 21301 15427 21335
rect 17141 21301 17175 21335
rect 11345 21097 11379 21131
rect 14381 21097 14415 21131
rect 18337 21097 18371 21131
rect 19349 21097 19383 21131
rect 10787 21029 10821 21063
rect 13506 21029 13540 21063
rect 16818 21029 16852 21063
rect 18061 21029 18095 21063
rect 8309 20961 8343 20995
rect 8585 20961 8619 20995
rect 12208 20961 12242 20995
rect 14105 20961 14139 20995
rect 15552 20961 15586 20995
rect 16497 20961 16531 20995
rect 17417 20961 17451 20995
rect 18521 20961 18555 20995
rect 18705 20961 18739 20995
rect 8769 20893 8803 20927
rect 10425 20893 10459 20927
rect 13185 20893 13219 20927
rect 9965 20757 9999 20791
rect 12311 20757 12345 20791
rect 15623 20757 15657 20791
rect 16313 20757 16347 20791
rect 8493 20553 8527 20587
rect 10425 20553 10459 20587
rect 11529 20553 11563 20587
rect 12173 20553 12207 20587
rect 14289 20553 14323 20587
rect 19073 20553 19107 20587
rect 9597 20417 9631 20451
rect 11069 20417 11103 20451
rect 16221 20417 16255 20451
rect 17785 20417 17819 20451
rect 8953 20349 8987 20383
rect 9413 20349 9447 20383
rect 13369 20349 13403 20383
rect 14565 20349 14599 20383
rect 15244 20349 15278 20383
rect 15669 20349 15703 20383
rect 17141 20349 17175 20383
rect 19660 20349 19694 20383
rect 20085 20349 20119 20383
rect 10609 20281 10643 20315
rect 10701 20281 10735 20315
rect 13690 20281 13724 20315
rect 16583 20281 16617 20315
rect 18153 20281 18187 20315
rect 18245 20281 18279 20315
rect 18797 20281 18831 20315
rect 8125 20213 8159 20247
rect 8769 20213 8803 20247
rect 10057 20213 10091 20247
rect 12909 20213 12943 20247
rect 13185 20213 13219 20247
rect 15347 20213 15381 20247
rect 16129 20213 16163 20247
rect 17417 20213 17451 20247
rect 19763 20213 19797 20247
rect 13185 20009 13219 20043
rect 16037 20009 16071 20043
rect 17233 20009 17267 20043
rect 10609 19941 10643 19975
rect 12817 19941 12851 19975
rect 13829 19941 13863 19975
rect 16313 19941 16347 19975
rect 17601 19941 17635 19975
rect 17785 19941 17819 19975
rect 17877 19941 17911 19975
rect 19349 19941 19383 19975
rect 19441 19941 19475 19975
rect 8620 19873 8654 19907
rect 12081 19873 12115 19907
rect 12633 19873 12667 19907
rect 7573 19805 7607 19839
rect 9137 19805 9171 19839
rect 10517 19805 10551 19839
rect 11161 19805 11195 19839
rect 13737 19805 13771 19839
rect 16221 19805 16255 19839
rect 18429 19805 18463 19839
rect 19625 19805 19659 19839
rect 8723 19737 8757 19771
rect 9873 19737 9907 19771
rect 14289 19737 14323 19771
rect 16773 19737 16807 19771
rect 9413 19669 9447 19703
rect 10241 19669 10275 19703
rect 14749 19669 14783 19703
rect 18797 19669 18831 19703
rect 8171 19465 8205 19499
rect 10057 19465 10091 19499
rect 14013 19465 14047 19499
rect 16957 19465 16991 19499
rect 17509 19465 17543 19499
rect 19257 19465 19291 19499
rect 19625 19465 19659 19499
rect 8585 19329 8619 19363
rect 9137 19329 9171 19363
rect 13185 19329 13219 19363
rect 14381 19329 14415 19363
rect 14841 19329 14875 19363
rect 16221 19329 16255 19363
rect 7941 19261 7975 19295
rect 8068 19261 8102 19295
rect 10425 19261 10459 19295
rect 12725 19261 12759 19295
rect 13093 19261 13127 19295
rect 13645 19261 13679 19295
rect 19860 19261 19894 19295
rect 20269 19261 20303 19295
rect 20821 19261 20855 19295
rect 9229 19193 9263 19227
rect 9781 19193 9815 19227
rect 10701 19193 10735 19227
rect 10793 19193 10827 19227
rect 11345 19193 11379 19227
rect 11805 19193 11839 19227
rect 14473 19193 14507 19227
rect 15761 19193 15795 19227
rect 15945 19193 15979 19227
rect 16037 19193 16071 19227
rect 17877 19193 17911 19227
rect 18337 19193 18371 19227
rect 18429 19193 18463 19227
rect 18981 19193 19015 19227
rect 19947 19193 19981 19227
rect 12081 19125 12115 19159
rect 15393 19125 15427 19159
rect 8723 18921 8757 18955
rect 11161 18921 11195 18955
rect 13277 18921 13311 18955
rect 14381 18921 14415 18955
rect 14657 18921 14691 18955
rect 16405 18921 16439 18955
rect 16773 18921 16807 18955
rect 17877 18921 17911 18955
rect 9505 18853 9539 18887
rect 10333 18853 10367 18887
rect 11897 18853 11931 18887
rect 13782 18853 13816 18887
rect 17278 18853 17312 18887
rect 18337 18853 18371 18887
rect 18889 18853 18923 18887
rect 7640 18785 7674 18819
rect 8620 18785 8654 18819
rect 15393 18785 15427 18819
rect 15945 18785 15979 18819
rect 10241 18717 10275 18751
rect 10885 18717 10919 18751
rect 11805 18717 11839 18751
rect 12081 18717 12115 18751
rect 13461 18717 13495 18751
rect 16129 18717 16163 18751
rect 16957 18717 16991 18751
rect 18797 18717 18831 18751
rect 19349 18649 19383 18683
rect 7711 18581 7745 18615
rect 9137 18581 9171 18615
rect 9965 18581 9999 18615
rect 12725 18581 12759 18615
rect 7849 18377 7883 18411
rect 10057 18377 10091 18411
rect 11529 18377 11563 18411
rect 11897 18377 11931 18411
rect 17325 18377 17359 18411
rect 19073 18377 19107 18411
rect 19441 18377 19475 18411
rect 9781 18241 9815 18275
rect 10609 18241 10643 18275
rect 12173 18241 12207 18275
rect 13461 18241 13495 18275
rect 14381 18241 14415 18275
rect 14841 18241 14875 18275
rect 16221 18241 16255 18275
rect 18153 18241 18187 18275
rect 18797 18241 18831 18275
rect 1460 18173 1494 18207
rect 1547 18173 1581 18207
rect 7056 18173 7090 18207
rect 7481 18173 7515 18207
rect 8068 18173 8102 18207
rect 8493 18173 8527 18207
rect 9321 18173 9355 18207
rect 9597 18173 9631 18207
rect 13001 18173 13035 18207
rect 13185 18173 13219 18207
rect 19660 18173 19694 18207
rect 20085 18173 20119 18207
rect 8171 18105 8205 18139
rect 10930 18105 10964 18139
rect 14473 18105 14507 18139
rect 15945 18105 15979 18139
rect 16037 18105 16071 18139
rect 18245 18105 18279 18139
rect 1961 18037 1995 18071
rect 7159 18037 7193 18071
rect 8861 18037 8895 18071
rect 10517 18037 10551 18071
rect 13737 18037 13771 18071
rect 14197 18037 14231 18071
rect 15393 18037 15427 18071
rect 16957 18037 16991 18071
rect 17785 18037 17819 18071
rect 19763 18037 19797 18071
rect 9137 17833 9171 17867
rect 9965 17833 9999 17867
rect 12817 17833 12851 17867
rect 13369 17833 13403 17867
rect 14381 17833 14415 17867
rect 14657 17833 14691 17867
rect 15439 17833 15473 17867
rect 16589 17833 16623 17867
rect 17693 17833 17727 17867
rect 18153 17833 18187 17867
rect 18521 17833 18555 17867
rect 7389 17765 7423 17799
rect 7573 17765 7607 17799
rect 7665 17765 7699 17799
rect 11161 17765 11195 17799
rect 11253 17765 11287 17799
rect 11805 17765 11839 17799
rect 13782 17765 13816 17799
rect 17094 17765 17128 17799
rect 1476 17697 1510 17731
rect 2513 17697 2547 17731
rect 5457 17697 5491 17731
rect 6536 17697 6570 17731
rect 10092 17697 10126 17731
rect 15336 17697 15370 17731
rect 8033 17629 8067 17663
rect 12081 17629 12115 17663
rect 13461 17629 13495 17663
rect 16773 17629 16807 17663
rect 15853 17561 15887 17595
rect 1547 17493 1581 17527
rect 2697 17493 2731 17527
rect 5641 17493 5675 17527
rect 6607 17493 6641 17527
rect 10195 17493 10229 17527
rect 10701 17493 10735 17527
rect 16313 17493 16347 17527
rect 1685 17289 1719 17323
rect 2697 17289 2731 17323
rect 6285 17289 6319 17323
rect 11529 17289 11563 17323
rect 11805 17289 11839 17323
rect 12633 17289 12667 17323
rect 14473 17289 14507 17323
rect 8033 17221 8067 17255
rect 2881 17153 2915 17187
rect 3157 17153 3191 17187
rect 5549 17153 5583 17187
rect 7297 17153 7331 17187
rect 8953 17153 8987 17187
rect 10609 17153 10643 17187
rect 14749 17153 14783 17187
rect 15301 17153 15335 17187
rect 18429 17153 18463 17187
rect 5784 17085 5818 17119
rect 8493 17085 8527 17119
rect 8861 17085 8895 17119
rect 9045 17085 9079 17119
rect 12265 17085 12299 17119
rect 12449 17085 12483 17119
rect 13553 17085 13587 17119
rect 16221 17085 16255 17119
rect 2973 17017 3007 17051
rect 5871 17017 5905 17051
rect 7481 17017 7515 17051
rect 7573 17017 7607 17051
rect 10517 17017 10551 17051
rect 10971 17017 11005 17051
rect 13894 17017 13928 17051
rect 16583 17017 16617 17051
rect 17417 17017 17451 17051
rect 18153 17017 18187 17051
rect 18245 17017 18279 17051
rect 1777 16949 1811 16983
rect 2237 16949 2271 16983
rect 6653 16949 6687 16983
rect 10057 16949 10091 16983
rect 13093 16949 13127 16983
rect 13461 16949 13495 16983
rect 16129 16949 16163 16983
rect 17141 16949 17175 16983
rect 17877 16949 17911 16983
rect 3065 16745 3099 16779
rect 7849 16745 7883 16779
rect 11805 16745 11839 16779
rect 12633 16745 12667 16779
rect 17463 16745 17497 16779
rect 18153 16745 18187 16779
rect 2145 16677 2179 16711
rect 2237 16677 2271 16711
rect 4261 16677 4295 16711
rect 7250 16677 7284 16711
rect 8125 16677 8159 16711
rect 10930 16677 10964 16711
rect 13645 16677 13679 16711
rect 13921 16677 13955 16711
rect 16497 16677 16531 16711
rect 16773 16677 16807 16711
rect 18475 16677 18509 16711
rect 6929 16609 6963 16643
rect 11529 16609 11563 16643
rect 13185 16609 13219 16643
rect 13369 16609 13403 16643
rect 14381 16609 14415 16643
rect 15761 16609 15795 16643
rect 16221 16609 16255 16643
rect 17360 16609 17394 16643
rect 18372 16609 18406 16643
rect 4169 16541 4203 16575
rect 4445 16541 4479 16575
rect 5917 16541 5951 16575
rect 10609 16541 10643 16575
rect 2697 16473 2731 16507
rect 5089 16405 5123 16439
rect 1685 16201 1719 16235
rect 4169 16201 4203 16235
rect 5365 16201 5399 16235
rect 8033 16201 8067 16235
rect 10425 16201 10459 16235
rect 18889 16201 18923 16235
rect 11161 16133 11195 16167
rect 12265 16133 12299 16167
rect 1915 16065 1949 16099
rect 3157 16065 3191 16099
rect 4445 16065 4479 16099
rect 4721 16065 4755 16099
rect 7021 16065 7055 16099
rect 10609 16065 10643 16099
rect 11529 16065 11563 16099
rect 13369 16065 13403 16099
rect 14289 16065 14323 16099
rect 14565 16065 14599 16099
rect 16313 16065 16347 16099
rect 17325 16065 17359 16099
rect 1812 15997 1846 16031
rect 2237 15997 2271 16031
rect 8677 15997 8711 16031
rect 8861 15997 8895 16031
rect 12725 15997 12759 16031
rect 13093 15997 13127 16031
rect 15761 15997 15795 16031
rect 16221 15997 16255 16031
rect 16773 15997 16807 16031
rect 18096 15997 18130 16031
rect 18521 15997 18555 16031
rect 19140 15997 19174 16031
rect 19533 15997 19567 16031
rect 2881 15929 2915 15963
rect 2973 15929 3007 15963
rect 4537 15929 4571 15963
rect 6285 15929 6319 15963
rect 7113 15929 7147 15963
rect 7665 15929 7699 15963
rect 9505 15929 9539 15963
rect 10057 15929 10091 15963
rect 10701 15929 10735 15963
rect 14381 15929 14415 15963
rect 2697 15861 2731 15895
rect 6561 15861 6595 15895
rect 13645 15861 13679 15895
rect 14013 15861 14047 15895
rect 15301 15861 15335 15895
rect 15669 15861 15703 15895
rect 18199 15861 18233 15895
rect 19211 15861 19245 15895
rect 2145 15657 2179 15691
rect 3525 15657 3559 15691
rect 5089 15657 5123 15691
rect 10701 15657 10735 15691
rect 11345 15657 11379 15691
rect 13001 15657 13035 15691
rect 15761 15657 15795 15691
rect 2513 15589 2547 15623
rect 2605 15589 2639 15623
rect 3157 15589 3191 15623
rect 4077 15589 4111 15623
rect 6469 15589 6503 15623
rect 6561 15589 6595 15623
rect 7941 15589 7975 15623
rect 9873 15589 9907 15623
rect 13829 15589 13863 15623
rect 14381 15589 14415 15623
rect 16583 15589 16617 15623
rect 18153 15589 18187 15623
rect 1444 15521 1478 15555
rect 4169 15521 4203 15555
rect 7481 15521 7515 15555
rect 8033 15521 8067 15555
rect 11253 15521 11287 15555
rect 11805 15521 11839 15555
rect 17141 15521 17175 15555
rect 9781 15453 9815 15487
rect 10057 15453 10091 15487
rect 13737 15453 13771 15487
rect 16221 15453 16255 15487
rect 18061 15453 18095 15487
rect 18337 15453 18371 15487
rect 7021 15385 7055 15419
rect 1547 15317 1581 15351
rect 7849 15317 7883 15351
rect 13369 15317 13403 15351
rect 2053 15113 2087 15147
rect 4169 15113 4203 15147
rect 6285 15113 6319 15147
rect 7757 15113 7791 15147
rect 9505 15113 9539 15147
rect 9781 15113 9815 15147
rect 11805 15113 11839 15147
rect 13277 15113 13311 15147
rect 14657 15113 14691 15147
rect 15301 15113 15335 15147
rect 17509 15113 17543 15147
rect 19073 15113 19107 15147
rect 3801 15045 3835 15079
rect 10149 15045 10183 15079
rect 12909 15045 12943 15079
rect 14289 15045 14323 15079
rect 6561 14977 6595 15011
rect 6837 14977 6871 15011
rect 10701 14977 10735 15011
rect 18153 14977 18187 15011
rect 1568 14909 1602 14943
rect 2421 14909 2455 14943
rect 2881 14909 2915 14943
rect 8125 14909 8159 14943
rect 8585 14909 8619 14943
rect 13369 14909 13403 14943
rect 15117 14909 15151 14943
rect 16221 14909 16255 14943
rect 3202 14841 3236 14875
rect 5273 14841 5307 14875
rect 5365 14841 5399 14875
rect 5917 14841 5951 14875
rect 7158 14841 7192 14875
rect 8401 14841 8435 14875
rect 8906 14841 8940 14875
rect 10425 14841 10459 14875
rect 10517 14841 10551 14875
rect 13690 14841 13724 14875
rect 15761 14841 15795 14875
rect 16129 14841 16163 14875
rect 16583 14841 16617 14875
rect 18245 14841 18279 14875
rect 18797 14841 18831 14875
rect 1639 14773 1673 14807
rect 2789 14773 2823 14807
rect 4629 14773 4663 14807
rect 5089 14773 5123 14807
rect 11345 14773 11379 14807
rect 14933 14773 14967 14807
rect 17141 14773 17175 14807
rect 17785 14773 17819 14807
rect 19625 14773 19659 14807
rect 2053 14569 2087 14603
rect 2513 14569 2547 14603
rect 3433 14569 3467 14603
rect 6561 14569 6595 14603
rect 7849 14569 7883 14603
rect 9413 14569 9447 14603
rect 10701 14569 10735 14603
rect 16405 14569 16439 14603
rect 18521 14569 18555 14603
rect 18797 14569 18831 14603
rect 2881 14501 2915 14535
rect 5733 14501 5767 14535
rect 8125 14501 8159 14535
rect 8217 14501 8251 14535
rect 9873 14501 9907 14535
rect 13363 14501 13397 14535
rect 15485 14501 15519 14535
rect 17325 14501 17359 14535
rect 1552 14433 1586 14467
rect 4537 14433 4571 14467
rect 11713 14433 11747 14467
rect 11897 14433 11931 14467
rect 17877 14433 17911 14467
rect 18705 14433 18739 14467
rect 19257 14433 19291 14467
rect 1639 14365 1673 14399
rect 2973 14365 3007 14399
rect 5641 14365 5675 14399
rect 6009 14365 6043 14399
rect 8401 14365 8435 14399
rect 9781 14365 9815 14399
rect 10057 14365 10091 14399
rect 12173 14365 12207 14399
rect 13001 14365 13035 14399
rect 15393 14365 15427 14399
rect 16037 14365 16071 14399
rect 17233 14365 17267 14399
rect 4721 14229 4755 14263
rect 5089 14229 5123 14263
rect 5457 14229 5491 14263
rect 6929 14229 6963 14263
rect 7297 14229 7331 14263
rect 9045 14229 9079 14263
rect 12541 14229 12575 14263
rect 13921 14229 13955 14263
rect 14197 14229 14231 14263
rect 16681 14229 16715 14263
rect 18245 14229 18279 14263
rect 3893 14025 3927 14059
rect 5917 14025 5951 14059
rect 8493 14025 8527 14059
rect 10241 14025 10275 14059
rect 13461 14025 13495 14059
rect 14013 14025 14047 14059
rect 17785 14025 17819 14059
rect 19073 14025 19107 14059
rect 19441 14025 19475 14059
rect 1593 13957 1627 13991
rect 6285 13957 6319 13991
rect 7113 13957 7147 13991
rect 10609 13957 10643 13991
rect 15393 13957 15427 13991
rect 17417 13957 17451 13991
rect 8677 13889 8711 13923
rect 11345 13889 11379 13923
rect 13185 13889 13219 13923
rect 14197 13889 14231 13923
rect 15761 13889 15795 13923
rect 16313 13889 16347 13923
rect 17141 13889 17175 13923
rect 18153 13889 18187 13923
rect 18429 13889 18463 13923
rect 19763 13889 19797 13923
rect 1409 13821 1443 13855
rect 2053 13821 2087 13855
rect 2513 13821 2547 13855
rect 2973 13821 3007 13855
rect 4537 13821 4571 13855
rect 4997 13821 5031 13855
rect 6929 13821 6963 13855
rect 8125 13821 8159 13855
rect 10793 13821 10827 13855
rect 11253 13821 11287 13855
rect 12265 13821 12299 13855
rect 12725 13821 12759 13855
rect 12909 13821 12943 13855
rect 14841 13821 14875 13855
rect 19660 13821 19694 13855
rect 20085 13821 20119 13855
rect 3294 13753 3328 13787
rect 4813 13753 4847 13787
rect 5318 13753 5352 13787
rect 8998 13753 9032 13787
rect 14289 13753 14323 13787
rect 16497 13753 16531 13787
rect 16589 13753 16623 13787
rect 18245 13753 18279 13787
rect 2881 13685 2915 13719
rect 6653 13685 6687 13719
rect 9597 13685 9631 13719
rect 9965 13685 9999 13719
rect 11897 13685 11931 13719
rect 5733 13481 5767 13515
rect 8493 13481 8527 13515
rect 9965 13481 9999 13515
rect 10885 13481 10919 13515
rect 13001 13481 13035 13515
rect 15117 13481 15151 13515
rect 16221 13481 16255 13515
rect 17417 13481 17451 13515
rect 18153 13481 18187 13515
rect 19947 13481 19981 13515
rect 2605 13413 2639 13447
rect 4261 13413 4295 13447
rect 8217 13413 8251 13447
rect 13553 13413 13587 13447
rect 14381 13413 14415 13447
rect 16859 13413 16893 13447
rect 18429 13413 18463 13447
rect 5917 13345 5951 13379
rect 6193 13345 6227 13379
rect 6653 13345 6687 13379
rect 7021 13345 7055 13379
rect 8401 13345 8435 13379
rect 10333 13345 10367 13379
rect 11713 13345 11747 13379
rect 13645 13345 13679 13379
rect 14197 13345 14231 13379
rect 15301 13345 15335 13379
rect 16497 13345 16531 13379
rect 19844 13345 19878 13379
rect 1409 13277 1443 13311
rect 2513 13277 2547 13311
rect 4169 13277 4203 13311
rect 4445 13277 4479 13311
rect 5549 13277 5583 13311
rect 11437 13277 11471 13311
rect 12357 13277 12391 13311
rect 18337 13277 18371 13311
rect 18797 13277 18831 13311
rect 3065 13209 3099 13243
rect 15853 13209 15887 13243
rect 1869 13141 1903 13175
rect 2237 13141 2271 13175
rect 3525 13141 3559 13175
rect 7389 13141 7423 13175
rect 7849 13141 7883 13175
rect 9229 13141 9263 13175
rect 15485 13141 15519 13175
rect 17785 13141 17819 13175
rect 2053 12937 2087 12971
rect 3893 12937 3927 12971
rect 4261 12937 4295 12971
rect 4905 12937 4939 12971
rect 8677 12937 8711 12971
rect 9045 12937 9079 12971
rect 11713 12937 11747 12971
rect 13645 12937 13679 12971
rect 17141 12937 17175 12971
rect 19441 12937 19475 12971
rect 20085 12937 20119 12971
rect 11253 12869 11287 12903
rect 19073 12869 19107 12903
rect 19809 12869 19843 12903
rect 10885 12801 10919 12835
rect 14565 12801 14599 12835
rect 16129 12801 16163 12835
rect 18153 12801 18187 12835
rect 18797 12801 18831 12835
rect 1409 12733 1443 12767
rect 2973 12733 3007 12767
rect 4629 12733 4663 12767
rect 4721 12733 4755 12767
rect 5733 12733 5767 12767
rect 6837 12733 6871 12767
rect 7389 12733 7423 12767
rect 7849 12733 7883 12767
rect 8033 12733 8067 12767
rect 9413 12733 9447 12767
rect 9873 12733 9907 12767
rect 10149 12733 10183 12767
rect 10333 12733 10367 12767
rect 12265 12733 12299 12767
rect 13093 12733 13127 12767
rect 14197 12733 14231 12767
rect 14933 12733 14967 12767
rect 15301 12733 15335 12767
rect 15669 12733 15703 12767
rect 15945 12733 15979 12767
rect 16957 12733 16991 12767
rect 17417 12733 17451 12767
rect 19625 12733 19659 12767
rect 20453 12733 20487 12767
rect 2789 12665 2823 12699
rect 3294 12665 3328 12699
rect 6285 12665 6319 12699
rect 6653 12665 6687 12699
rect 14013 12665 14047 12699
rect 17877 12665 17911 12699
rect 18245 12665 18279 12699
rect 1593 12597 1627 12631
rect 2513 12597 2547 12631
rect 5181 12597 5215 12631
rect 5641 12597 5675 12631
rect 5917 12597 5951 12631
rect 7113 12597 7147 12631
rect 9413 12597 9447 12631
rect 12725 12597 12759 12631
rect 16589 12597 16623 12631
rect 1547 12393 1581 12427
rect 2881 12393 2915 12427
rect 3893 12393 3927 12427
rect 4353 12393 4387 12427
rect 4583 12393 4617 12427
rect 5595 12393 5629 12427
rect 5917 12393 5951 12427
rect 7665 12393 7699 12427
rect 9781 12393 9815 12427
rect 10885 12393 10919 12427
rect 12725 12393 12759 12427
rect 13093 12393 13127 12427
rect 14381 12393 14415 12427
rect 15577 12393 15611 12427
rect 16589 12393 16623 12427
rect 17693 12393 17727 12427
rect 1476 12257 1510 12291
rect 3065 12257 3099 12291
rect 4512 12257 4546 12291
rect 5524 12257 5558 12291
rect 6469 12257 6503 12291
rect 6929 12257 6963 12291
rect 7481 12257 7515 12291
rect 7665 12257 7699 12291
rect 9137 12257 9171 12291
rect 14013 12325 14047 12359
rect 17094 12325 17128 12359
rect 18705 12325 18739 12359
rect 9873 12257 9907 12291
rect 10149 12257 10183 12291
rect 11713 12257 11747 12291
rect 11989 12257 12023 12291
rect 13277 12257 13311 12291
rect 13369 12257 13403 12291
rect 13553 12257 13587 12291
rect 15117 12257 15151 12291
rect 15301 12257 15335 12291
rect 15485 12257 15519 12291
rect 4905 12189 4939 12223
rect 6377 12189 6411 12223
rect 8585 12189 8619 12223
rect 9781 12189 9815 12223
rect 9965 12189 9999 12223
rect 10333 12189 10367 12223
rect 11621 12189 11655 12223
rect 12173 12189 12207 12223
rect 16773 12189 16807 12223
rect 18613 12189 18647 12223
rect 1961 12121 1995 12155
rect 11805 12121 11839 12155
rect 19165 12121 19199 12155
rect 2237 12053 2271 12087
rect 3525 12053 3559 12087
rect 8309 12053 8343 12087
rect 16129 12053 16163 12087
rect 18153 12053 18187 12087
rect 1593 11849 1627 11883
rect 5549 11849 5583 11883
rect 7297 11849 7331 11883
rect 7665 11849 7699 11883
rect 9873 11849 9907 11883
rect 13553 11849 13587 11883
rect 19073 11849 19107 11883
rect 19441 11849 19475 11883
rect 19809 11849 19843 11883
rect 4537 11781 4571 11815
rect 5917 11781 5951 11815
rect 12541 11781 12575 11815
rect 2053 11713 2087 11747
rect 2605 11713 2639 11747
rect 6561 11713 6595 11747
rect 8033 11713 8067 11747
rect 16313 11713 16347 11747
rect 17877 11713 17911 11747
rect 18153 11713 18187 11747
rect 1409 11645 1443 11679
rect 3065 11645 3099 11679
rect 3433 11645 3467 11679
rect 3893 11645 3927 11679
rect 4077 11645 4111 11679
rect 4537 11645 4571 11679
rect 4997 11645 5031 11679
rect 5733 11645 5767 11679
rect 7113 11645 7147 11679
rect 8309 11645 8343 11679
rect 8585 11645 8619 11679
rect 9137 11645 9171 11679
rect 9505 11645 9539 11679
rect 10333 11645 10367 11679
rect 10977 11645 11011 11679
rect 12449 11645 12483 11679
rect 12725 11645 12759 11679
rect 13921 11645 13955 11679
rect 14657 11645 14691 11679
rect 15669 11645 15703 11679
rect 16037 11645 16071 11679
rect 17141 11645 17175 11679
rect 18061 11645 18095 11679
rect 18337 11645 18371 11679
rect 19625 11645 19659 11679
rect 20085 11645 20119 11679
rect 12173 11577 12207 11611
rect 14749 11577 14783 11611
rect 18797 11577 18831 11611
rect 6285 11509 6319 11543
rect 8401 11509 8435 11543
rect 10701 11509 10735 11543
rect 11805 11509 11839 11543
rect 12909 11509 12943 11543
rect 15393 11509 15427 11543
rect 16773 11509 16807 11543
rect 2881 11305 2915 11339
rect 3893 11305 3927 11339
rect 5365 11305 5399 11339
rect 5825 11305 5859 11339
rect 9413 11305 9447 11339
rect 9965 11305 9999 11339
rect 12173 11305 12207 11339
rect 12725 11305 12759 11339
rect 13277 11305 13311 11339
rect 17325 11305 17359 11339
rect 19441 11305 19475 11339
rect 7849 11237 7883 11271
rect 14381 11237 14415 11271
rect 16037 11237 16071 11271
rect 1961 11169 1995 11203
rect 2237 11169 2271 11203
rect 2697 11169 2731 11203
rect 2881 11169 2915 11203
rect 4537 11169 4571 11203
rect 5825 11169 5859 11203
rect 6193 11169 6227 11203
rect 6377 11169 6411 11203
rect 6929 11169 6963 11203
rect 8493 11169 8527 11203
rect 10057 11169 10091 11203
rect 10149 11169 10183 11203
rect 10425 11169 10459 11203
rect 11713 11169 11747 11203
rect 11989 11169 12023 11203
rect 13645 11169 13679 11203
rect 13921 11169 13955 11203
rect 15301 11169 15335 11203
rect 15577 11169 15611 11203
rect 16865 11169 16899 11203
rect 17141 11169 17175 11203
rect 18061 11169 18095 11203
rect 18981 11169 19015 11203
rect 10241 11101 10275 11135
rect 10885 11101 10919 11135
rect 13737 11101 13771 11135
rect 18429 11101 18463 11135
rect 3525 11033 3559 11067
rect 4261 11033 4295 11067
rect 4721 11033 4755 11067
rect 5089 11033 5123 11067
rect 10057 11033 10091 11067
rect 11805 11033 11839 11067
rect 15393 11033 15427 11067
rect 16957 11033 16991 11067
rect 7665 10965 7699 10999
rect 8953 10965 8987 10999
rect 11529 10965 11563 10999
rect 14841 10965 14875 10999
rect 16497 10965 16531 10999
rect 5273 10761 5307 10795
rect 6285 10761 6319 10795
rect 6653 10761 6687 10795
rect 7113 10761 7147 10795
rect 9413 10761 9447 10795
rect 9781 10761 9815 10795
rect 10977 10761 11011 10795
rect 11437 10761 11471 10795
rect 11805 10761 11839 10795
rect 12081 10761 12115 10795
rect 14013 10761 14047 10795
rect 14657 10761 14691 10795
rect 16221 10761 16255 10795
rect 19349 10761 19383 10795
rect 15945 10693 15979 10727
rect 13185 10625 13219 10659
rect 13737 10625 13771 10659
rect 17877 10625 17911 10659
rect 2053 10557 2087 10591
rect 2973 10557 3007 10591
rect 3341 10557 3375 10591
rect 3801 10557 3835 10591
rect 4077 10557 4111 10591
rect 4261 10557 4295 10591
rect 4813 10557 4847 10591
rect 5733 10557 5767 10591
rect 7849 10557 7883 10591
rect 8217 10557 8251 10591
rect 8585 10557 8619 10591
rect 8769 10557 8803 10591
rect 9965 10557 9999 10591
rect 13001 10557 13035 10591
rect 15025 10557 15059 10591
rect 15301 10557 15335 10591
rect 16405 10557 16439 10591
rect 16865 10557 16899 10591
rect 18061 10557 18095 10591
rect 18245 10557 18279 10591
rect 19433 10557 19467 10591
rect 1409 10489 1443 10523
rect 5641 10489 5675 10523
rect 7481 10489 7515 10523
rect 9045 10489 9079 10523
rect 9873 10489 9907 10523
rect 15577 10489 15611 10523
rect 17509 10489 17543 10523
rect 19901 10489 19935 10523
rect 2513 10421 2547 10455
rect 3157 10421 3191 10455
rect 5917 10421 5951 10455
rect 16681 10421 16715 10455
rect 18337 10421 18371 10455
rect 18981 10421 19015 10455
rect 19625 10421 19659 10455
rect 1777 10217 1811 10251
rect 3065 10217 3099 10251
rect 3433 10217 3467 10251
rect 3801 10217 3835 10251
rect 4629 10217 4663 10251
rect 5457 10217 5491 10251
rect 6101 10217 6135 10251
rect 7941 10217 7975 10251
rect 8769 10217 8803 10251
rect 11069 10217 11103 10251
rect 12909 10217 12943 10251
rect 13829 10217 13863 10251
rect 15117 10217 15151 10251
rect 18061 10217 18095 10251
rect 18613 10217 18647 10251
rect 2507 10149 2541 10183
rect 9873 10149 9907 10183
rect 10701 10149 10735 10183
rect 11437 10149 11471 10183
rect 4997 10081 5031 10115
rect 6285 10081 6319 10115
rect 6745 10081 6779 10115
rect 7021 10081 7055 10115
rect 7389 10081 7423 10115
rect 8585 10081 8619 10115
rect 13093 10081 13127 10115
rect 13369 10081 13403 10115
rect 15301 10081 15335 10115
rect 15577 10081 15611 10115
rect 16037 10081 16071 10115
rect 16865 10081 16899 10115
rect 17141 10081 17175 10115
rect 17601 10081 17635 10115
rect 18429 10081 18463 10115
rect 19441 10081 19475 10115
rect 2145 10013 2179 10047
rect 9781 10013 9815 10047
rect 10149 10013 10183 10047
rect 11345 10013 11379 10047
rect 11989 10013 12023 10047
rect 15393 10013 15427 10047
rect 16957 10013 16991 10047
rect 16497 9945 16531 9979
rect 18889 9945 18923 9979
rect 19625 9945 19659 9979
rect 5181 9877 5215 9911
rect 5917 9877 5951 9911
rect 8309 9877 8343 9911
rect 9045 9877 9079 9911
rect 9413 9877 9447 9911
rect 12541 9877 12575 9911
rect 14749 9877 14783 9911
rect 5549 9673 5583 9707
rect 6285 9673 6319 9707
rect 6653 9673 6687 9707
rect 10057 9673 10091 9707
rect 10333 9673 10367 9707
rect 10885 9673 10919 9707
rect 13553 9673 13587 9707
rect 17693 9673 17727 9707
rect 19073 9673 19107 9707
rect 19441 9673 19475 9707
rect 3065 9605 3099 9639
rect 8677 9605 8711 9639
rect 17049 9605 17083 9639
rect 17417 9605 17451 9639
rect 19763 9605 19797 9639
rect 20177 9605 20211 9639
rect 1685 9537 1719 9571
rect 2329 9537 2363 9571
rect 9137 9537 9171 9571
rect 11529 9537 11563 9571
rect 12541 9537 12575 9571
rect 13829 9537 13863 9571
rect 15117 9537 15151 9571
rect 18153 9537 18187 9571
rect 3433 9469 3467 9503
rect 3893 9469 3927 9503
rect 4169 9469 4203 9503
rect 4537 9469 4571 9503
rect 5181 9469 5215 9503
rect 5733 9469 5767 9503
rect 7113 9469 7147 9503
rect 7297 9469 7331 9503
rect 7849 9469 7883 9503
rect 8033 9469 8067 9503
rect 11161 9469 11195 9503
rect 14289 9469 14323 9503
rect 15025 9469 15059 9503
rect 16129 9469 16163 9503
rect 16405 9469 16439 9503
rect 19692 9469 19726 9503
rect 1777 9401 1811 9435
rect 9045 9401 9079 9435
rect 9458 9401 9492 9435
rect 10977 9401 11011 9435
rect 11805 9401 11839 9435
rect 12265 9401 12299 9435
rect 12633 9401 12667 9435
rect 13185 9401 13219 9435
rect 15853 9401 15887 9435
rect 18245 9401 18279 9435
rect 18797 9401 18831 9435
rect 2605 9333 2639 9367
rect 4537 9333 4571 9367
rect 5917 9333 5951 9367
rect 8033 9333 8067 9367
rect 15485 9333 15519 9367
rect 16221 9333 16255 9367
rect 3157 9129 3191 9163
rect 3525 9129 3559 9163
rect 4353 9129 4387 9163
rect 8677 9129 8711 9163
rect 8953 9129 8987 9163
rect 9321 9129 9355 9163
rect 11345 9129 11379 9163
rect 12633 9129 12667 9163
rect 15485 9129 15519 9163
rect 15853 9129 15887 9163
rect 16129 9129 16163 9163
rect 17969 9129 18003 9163
rect 1593 9061 1627 9095
rect 2145 9061 2179 9095
rect 2513 9061 2547 9095
rect 9873 9061 9907 9095
rect 12034 9061 12068 9095
rect 16675 9061 16709 9095
rect 18245 9061 18279 9095
rect 18797 9061 18831 9095
rect 2973 8993 3007 9027
rect 4077 8993 4111 9027
rect 4537 8993 4571 9027
rect 4997 8993 5031 9027
rect 5273 8993 5307 9027
rect 6377 8993 6411 9027
rect 6837 8993 6871 9027
rect 7205 8993 7239 9027
rect 7573 8993 7607 9027
rect 11713 8993 11747 9027
rect 13737 8993 13771 9027
rect 13921 8993 13955 9027
rect 15301 8993 15335 9027
rect 16313 8993 16347 9027
rect 19625 8993 19659 9027
rect 1501 8925 1535 8959
rect 9781 8925 9815 8959
rect 10149 8925 10183 8959
rect 13001 8925 13035 8959
rect 13369 8925 13403 8959
rect 14013 8925 14047 8959
rect 18153 8925 18187 8959
rect 3801 8857 3835 8891
rect 6009 8857 6043 8891
rect 7757 8857 7791 8891
rect 2881 8789 2915 8823
rect 8125 8789 8159 8823
rect 14565 8789 14599 8823
rect 15025 8789 15059 8823
rect 17233 8789 17267 8823
rect 19809 8789 19843 8823
rect 1593 8585 1627 8619
rect 1961 8585 1995 8619
rect 2881 8585 2915 8619
rect 3249 8585 3283 8619
rect 3525 8585 3559 8619
rect 5457 8585 5491 8619
rect 6101 8585 6135 8619
rect 6377 8585 6411 8619
rect 8769 8585 8803 8619
rect 9873 8585 9907 8619
rect 11529 8585 11563 8619
rect 13553 8585 13587 8619
rect 15209 8585 15243 8619
rect 17785 8585 17819 8619
rect 19165 8585 19199 8619
rect 16589 8517 16623 8551
rect 9137 8449 9171 8483
rect 10609 8449 10643 8483
rect 12265 8449 12299 8483
rect 15669 8449 15703 8483
rect 18153 8449 18187 8483
rect 19441 8449 19475 8483
rect 1409 8381 1443 8415
rect 2697 8381 2731 8415
rect 3709 8381 3743 8415
rect 4261 8381 4295 8415
rect 4721 8381 4755 8415
rect 4905 8381 4939 8415
rect 7021 8381 7055 8415
rect 7481 8381 7515 8415
rect 7849 8381 7883 8415
rect 8309 8381 8343 8415
rect 10425 8381 10459 8415
rect 12725 8381 12759 8415
rect 13001 8381 13035 8415
rect 14013 8381 14047 8415
rect 14105 8381 14139 8415
rect 14657 8381 14691 8415
rect 20085 8381 20119 8415
rect 2605 8313 2639 8347
rect 9321 8313 9355 8347
rect 10930 8313 10964 8347
rect 11805 8313 11839 8347
rect 13185 8313 13219 8347
rect 14841 8313 14875 8347
rect 15990 8313 16024 8347
rect 16865 8313 16899 8347
rect 18245 8313 18279 8347
rect 18797 8313 18831 8347
rect 19625 8313 19659 8347
rect 3801 8245 3835 8279
rect 8217 8245 8251 8279
rect 15485 8245 15519 8279
rect 17509 8245 17543 8279
rect 1409 8041 1443 8075
rect 1869 8041 1903 8075
rect 2237 8041 2271 8075
rect 5089 8041 5123 8075
rect 5457 8041 5491 8075
rect 7481 8041 7515 8075
rect 10701 8041 10735 8075
rect 11897 8041 11931 8075
rect 13645 8041 13679 8075
rect 15485 8041 15519 8075
rect 15761 8041 15795 8075
rect 16405 8041 16439 8075
rect 17509 8041 17543 8075
rect 3801 7973 3835 8007
rect 4353 7973 4387 8007
rect 12770 7973 12804 8007
rect 16910 7973 16944 8007
rect 18521 7973 18555 8007
rect 19073 7973 19107 8007
rect 3065 7905 3099 7939
rect 4696 7905 4730 7939
rect 5641 7905 5675 7939
rect 6193 7905 6227 7939
rect 6469 7905 6503 7939
rect 6837 7905 6871 7939
rect 7757 7905 7791 7939
rect 8677 7905 8711 7939
rect 9940 7905 9974 7939
rect 11161 7905 11195 7939
rect 11437 7905 11471 7939
rect 14197 7905 14231 7939
rect 15301 7905 15335 7939
rect 16589 7905 16623 7939
rect 8769 7837 8803 7871
rect 11621 7837 11655 7871
rect 12449 7837 12483 7871
rect 18429 7837 18463 7871
rect 4767 7769 4801 7803
rect 7021 7769 7055 7803
rect 13369 7769 13403 7803
rect 14013 7769 14047 7803
rect 2697 7701 2731 7735
rect 9505 7701 9539 7735
rect 10011 7701 10045 7735
rect 14381 7701 14415 7735
rect 18061 7701 18095 7735
rect 1593 7497 1627 7531
rect 2145 7497 2179 7531
rect 3893 7497 3927 7531
rect 6009 7497 6043 7531
rect 7113 7497 7147 7531
rect 8677 7497 8711 7531
rect 8953 7497 8987 7531
rect 10517 7497 10551 7531
rect 10977 7497 11011 7531
rect 12173 7497 12207 7531
rect 13461 7497 13495 7531
rect 13921 7497 13955 7531
rect 17141 7497 17175 7531
rect 17877 7497 17911 7531
rect 19165 7497 19199 7531
rect 20177 7497 20211 7531
rect 6285 7429 6319 7463
rect 7665 7429 7699 7463
rect 2973 7361 3007 7395
rect 4721 7361 4755 7395
rect 7757 7361 7791 7395
rect 12909 7361 12943 7395
rect 14105 7361 14139 7395
rect 14381 7361 14415 7395
rect 15761 7361 15795 7395
rect 16221 7361 16255 7395
rect 18613 7361 18647 7395
rect 1409 7293 1443 7327
rect 16037 7293 16071 7327
rect 19692 7293 19726 7327
rect 2881 7225 2915 7259
rect 3335 7225 3369 7259
rect 4261 7225 4295 7259
rect 5083 7225 5117 7259
rect 8119 7225 8153 7259
rect 9597 7225 9631 7259
rect 9689 7225 9723 7259
rect 10241 7225 10275 7259
rect 11345 7225 11379 7259
rect 12541 7225 12575 7259
rect 12633 7225 12667 7259
rect 14197 7225 14231 7259
rect 16542 7225 16576 7259
rect 17417 7225 17451 7259
rect 18153 7225 18187 7259
rect 18245 7225 18279 7259
rect 4629 7157 4663 7191
rect 5641 7157 5675 7191
rect 9321 7157 9355 7191
rect 11805 7157 11839 7191
rect 15393 7157 15427 7191
rect 19763 7157 19797 7191
rect 1547 6953 1581 6987
rect 5089 6953 5123 6987
rect 7757 6953 7791 6987
rect 10977 6953 11011 6987
rect 12541 6953 12575 6987
rect 14197 6953 14231 6987
rect 15393 6953 15427 6987
rect 16589 6953 16623 6987
rect 2605 6885 2639 6919
rect 4261 6885 4295 6919
rect 5825 6885 5859 6919
rect 8170 6885 8204 6919
rect 9873 6885 9907 6919
rect 11615 6885 11649 6919
rect 12817 6885 12851 6919
rect 13369 6885 13403 6919
rect 13921 6885 13955 6919
rect 17693 6885 17727 6919
rect 1476 6817 1510 6851
rect 1961 6817 1995 6851
rect 3709 6817 3743 6851
rect 7849 6817 7883 6851
rect 15301 6817 15335 6851
rect 15853 6817 15887 6851
rect 19073 6817 19107 6851
rect 19533 6817 19567 6851
rect 2513 6749 2547 6783
rect 4169 6749 4203 6783
rect 4445 6749 4479 6783
rect 5733 6749 5767 6783
rect 6009 6749 6043 6783
rect 9781 6749 9815 6783
rect 11253 6749 11287 6783
rect 13277 6749 13311 6783
rect 17601 6749 17635 6783
rect 19625 6749 19659 6783
rect 2329 6681 2363 6715
rect 3065 6681 3099 6715
rect 10333 6681 10367 6715
rect 18153 6681 18187 6715
rect 5549 6613 5583 6647
rect 6653 6613 6687 6647
rect 8769 6613 8803 6647
rect 9505 6613 9539 6647
rect 12173 6613 12207 6647
rect 18521 6613 18555 6647
rect 18889 6613 18923 6647
rect 2145 6409 2179 6443
rect 2513 6409 2547 6443
rect 4261 6409 4295 6443
rect 6561 6409 6595 6443
rect 8217 6409 8251 6443
rect 9689 6409 9723 6443
rect 11345 6409 11379 6443
rect 12173 6409 12207 6443
rect 13369 6409 13403 6443
rect 13645 6409 13679 6443
rect 14013 6409 14047 6443
rect 16589 6409 16623 6443
rect 17785 6409 17819 6443
rect 19073 6409 19107 6443
rect 19441 6409 19475 6443
rect 1593 6341 1627 6375
rect 4629 6341 4663 6375
rect 5825 6341 5859 6375
rect 7941 6341 7975 6375
rect 14841 6341 14875 6375
rect 17509 6341 17543 6375
rect 2973 6273 3007 6307
rect 5273 6273 5307 6307
rect 6975 6273 7009 6307
rect 8677 6273 8711 6307
rect 10701 6273 10735 6307
rect 12449 6273 12483 6307
rect 16957 6273 16991 6307
rect 1409 6205 1443 6239
rect 6888 6205 6922 6239
rect 14427 6205 14461 6239
rect 15393 6205 15427 6239
rect 16313 6205 16347 6239
rect 18797 6205 18831 6239
rect 2881 6137 2915 6171
rect 3335 6137 3369 6171
rect 5089 6137 5123 6171
rect 5365 6137 5399 6171
rect 8769 6137 8803 6171
rect 9321 6137 9355 6171
rect 10241 6137 10275 6171
rect 10333 6137 10367 6171
rect 12770 6137 12804 6171
rect 14519 6137 14553 6171
rect 15714 6137 15748 6171
rect 18153 6137 18187 6171
rect 18245 6137 18279 6171
rect 3893 6069 3927 6103
rect 6193 6069 6227 6103
rect 7389 6069 7423 6103
rect 9965 6069 9999 6103
rect 11621 6069 11655 6103
rect 15209 6069 15243 6103
rect 2053 5865 2087 5899
rect 2605 5865 2639 5899
rect 3065 5865 3099 5899
rect 3525 5865 3559 5899
rect 5273 5865 5307 5899
rect 6929 5865 6963 5899
rect 8677 5865 8711 5899
rect 9045 5865 9079 5899
rect 9827 5865 9861 5899
rect 10701 5865 10735 5899
rect 15577 5865 15611 5899
rect 16681 5865 16715 5899
rect 3801 5797 3835 5831
rect 4813 5797 4847 5831
rect 6003 5797 6037 5831
rect 10977 5797 11011 5831
rect 11069 5797 11103 5831
rect 11621 5797 11655 5831
rect 12770 5797 12804 5831
rect 16082 5797 16116 5831
rect 17417 5797 17451 5831
rect 17693 5797 17727 5831
rect 19257 5797 19291 5831
rect 1660 5729 1694 5763
rect 4721 5729 4755 5763
rect 5641 5729 5675 5763
rect 7849 5729 7883 5763
rect 9756 5729 9790 5763
rect 10149 5729 10183 5763
rect 12449 5729 12483 5763
rect 14232 5729 14266 5763
rect 15761 5729 15795 5763
rect 7389 5661 7423 5695
rect 17601 5661 17635 5695
rect 18245 5661 18279 5695
rect 19165 5661 19199 5695
rect 19441 5661 19475 5695
rect 1731 5593 1765 5627
rect 2421 5593 2455 5627
rect 14335 5593 14369 5627
rect 6561 5525 6595 5559
rect 9413 5525 9447 5559
rect 13369 5525 13403 5559
rect 18521 5525 18555 5559
rect 4445 5321 4479 5355
rect 10333 5321 10367 5355
rect 11897 5321 11931 5355
rect 15485 5321 15519 5355
rect 15853 5321 15887 5355
rect 17601 5321 17635 5355
rect 19165 5321 19199 5355
rect 19441 5321 19475 5355
rect 12265 5253 12299 5287
rect 17049 5253 17083 5287
rect 2697 5185 2731 5219
rect 3157 5185 3191 5219
rect 6285 5185 6319 5219
rect 6837 5185 6871 5219
rect 9321 5185 9355 5219
rect 11529 5185 11563 5219
rect 13093 5185 13127 5219
rect 14197 5185 14231 5219
rect 14473 5185 14507 5219
rect 16497 5185 16531 5219
rect 18153 5185 18187 5219
rect 18613 5185 18647 5219
rect 1409 5117 1443 5151
rect 5089 5117 5123 5151
rect 5825 5117 5859 5151
rect 6653 5117 6687 5151
rect 8493 5117 8527 5151
rect 8677 5117 8711 5151
rect 10701 5117 10735 5151
rect 10977 5117 11011 5151
rect 11345 5117 11379 5151
rect 3065 5049 3099 5083
rect 3519 5049 3553 5083
rect 5917 5049 5951 5083
rect 7199 5049 7233 5083
rect 12633 5049 12667 5083
rect 12725 5049 12759 5083
rect 14289 5049 14323 5083
rect 16313 5049 16347 5083
rect 16589 5049 16623 5083
rect 18245 5049 18279 5083
rect 1593 4981 1627 5015
rect 2053 4981 2087 5015
rect 4077 4981 4111 5015
rect 7757 4981 7791 5015
rect 8033 4981 8067 5015
rect 9781 4981 9815 5015
rect 13645 4981 13679 5015
rect 13921 4981 13955 5015
rect 2237 4777 2271 4811
rect 5641 4777 5675 4811
rect 10885 4777 10919 4811
rect 12633 4777 12667 4811
rect 14105 4777 14139 4811
rect 16497 4777 16531 4811
rect 17693 4777 17727 4811
rect 18061 4777 18095 4811
rect 18383 4777 18417 4811
rect 19395 4777 19429 4811
rect 21419 4777 21453 4811
rect 6101 4709 6135 4743
rect 7665 4709 7699 4743
rect 11345 4709 11379 4743
rect 12909 4709 12943 4743
rect 16865 4709 16899 4743
rect 17417 4709 17451 4743
rect 1476 4641 1510 4675
rect 3065 4641 3099 4675
rect 10057 4641 10091 4675
rect 15336 4641 15370 4675
rect 18312 4641 18346 4675
rect 19324 4641 19358 4675
rect 21348 4641 21382 4675
rect 4905 4573 4939 4607
rect 6009 4573 6043 4607
rect 6653 4573 6687 4607
rect 7573 4573 7607 4607
rect 7849 4573 7883 4607
rect 11253 4573 11287 4607
rect 11621 4573 11655 4607
rect 12817 4573 12851 4607
rect 13093 4573 13127 4607
rect 14473 4573 14507 4607
rect 16773 4573 16807 4607
rect 1547 4505 1581 4539
rect 4629 4505 4663 4539
rect 7389 4505 7423 4539
rect 15439 4505 15473 4539
rect 1961 4437 1995 4471
rect 2881 4437 2915 4471
rect 7021 4437 7055 4471
rect 10241 4437 10275 4471
rect 2513 4233 2547 4267
rect 2881 4233 2915 4267
rect 6009 4233 6043 4267
rect 6285 4233 6319 4267
rect 7849 4233 7883 4267
rect 10149 4233 10183 4267
rect 11253 4233 11287 4267
rect 12081 4233 12115 4267
rect 12173 4233 12207 4267
rect 13829 4233 13863 4267
rect 14565 4233 14599 4267
rect 15669 4233 15703 4267
rect 16773 4233 16807 4267
rect 2053 4165 2087 4199
rect 11483 4165 11517 4199
rect 4445 4097 4479 4131
rect 4721 4097 4755 4131
rect 4997 4097 5031 4131
rect 6929 4097 6963 4131
rect 9735 4097 9769 4131
rect 10885 4097 10919 4131
rect 1409 4029 1443 4063
rect 8652 4029 8686 4063
rect 9643 4029 9677 4063
rect 11380 4029 11414 4063
rect 11805 4029 11839 4063
rect 3157 3961 3191 3995
rect 3249 3961 3283 3995
rect 3801 3961 3835 3995
rect 4813 3961 4847 3995
rect 7021 3961 7055 3995
rect 7573 3961 7607 3995
rect 13093 4165 13127 4199
rect 13461 4097 13495 4131
rect 16221 4097 16255 4131
rect 17141 4097 17175 4131
rect 14749 4029 14783 4063
rect 15117 4029 15151 4063
rect 16380 4029 16414 4063
rect 12541 3961 12575 3995
rect 12633 3961 12667 3995
rect 1593 3893 1627 3927
rect 8217 3893 8251 3927
rect 8723 3893 8757 3927
rect 9137 3893 9171 3927
rect 10517 3893 10551 3927
rect 12081 3893 12115 3927
rect 14933 3893 14967 3927
rect 16451 3893 16485 3927
rect 18337 3893 18371 3927
rect 19349 3893 19383 3927
rect 21373 3893 21407 3927
rect 1685 3689 1719 3723
rect 5779 3689 5813 3723
rect 8723 3689 8757 3723
rect 10103 3689 10137 3723
rect 11575 3689 11609 3723
rect 12541 3689 12575 3723
rect 14749 3689 14783 3723
rect 15439 3689 15473 3723
rect 2506 3621 2540 3655
rect 3065 3621 3099 3655
rect 3341 3621 3375 3655
rect 4261 3621 4295 3655
rect 4813 3621 4847 3655
rect 7113 3621 7147 3655
rect 12909 3621 12943 3655
rect 5676 3553 5710 3587
rect 8652 3553 8686 3587
rect 10000 3553 10034 3587
rect 11472 3553 11506 3587
rect 15368 3553 15402 3587
rect 16589 3553 16623 3587
rect 2237 3485 2271 3519
rect 2421 3485 2455 3519
rect 4169 3485 4203 3519
rect 7021 3485 7055 3519
rect 7389 3485 7423 3519
rect 12817 3485 12851 3519
rect 13093 3485 13127 3519
rect 16773 3349 16807 3383
rect 3801 3145 3835 3179
rect 5641 3145 5675 3179
rect 6653 3145 6687 3179
rect 7987 3145 8021 3179
rect 8769 3145 8803 3179
rect 11483 3145 11517 3179
rect 13737 3145 13771 3179
rect 14565 3145 14599 3179
rect 15669 3145 15703 3179
rect 16681 3145 16715 3179
rect 17049 3145 17083 3179
rect 18659 3145 18693 3179
rect 4905 3077 4939 3111
rect 7665 3077 7699 3111
rect 9965 3077 9999 3111
rect 12173 3077 12207 3111
rect 12633 3077 12667 3111
rect 14105 3077 14139 3111
rect 2237 3009 2271 3043
rect 2789 3009 2823 3043
rect 3157 3009 3191 3043
rect 4353 3009 4387 3043
rect 5273 3009 5307 3043
rect 6975 3009 7009 3043
rect 11897 3009 11931 3043
rect 13369 3009 13403 3043
rect 1409 2941 1443 2975
rect 6888 2941 6922 2975
rect 7389 2941 7423 2975
rect 7916 2941 7950 2975
rect 11412 2941 11446 2975
rect 12449 2941 12483 2975
rect 13001 2941 13035 2975
rect 13921 2941 13955 2975
rect 14933 2941 14967 2975
rect 15025 2941 15059 2975
rect 16272 2941 16306 2975
rect 18588 2941 18622 2975
rect 2881 2873 2915 2907
rect 4169 2873 4203 2907
rect 4445 2873 4479 2907
rect 8401 2873 8435 2907
rect 16359 2873 16393 2907
rect 19073 2873 19107 2907
rect 1593 2805 1627 2839
rect 2605 2805 2639 2839
rect 15209 2805 15243 2839
rect 1547 2601 1581 2635
rect 4077 2601 4111 2635
rect 4537 2601 4571 2635
rect 4997 2601 5031 2635
rect 5227 2601 5261 2635
rect 7067 2601 7101 2635
rect 7389 2601 7423 2635
rect 13185 2601 13219 2635
rect 14473 2601 14507 2635
rect 18935 2601 18969 2635
rect 24731 2601 24765 2635
rect 3157 2533 3191 2567
rect 1476 2465 1510 2499
rect 2329 2465 2363 2499
rect 3065 2465 3099 2499
rect 5124 2465 5158 2499
rect 5549 2465 5583 2499
rect 6996 2465 7030 2499
rect 10609 2465 10643 2499
rect 11161 2465 11195 2499
rect 12633 2465 12667 2499
rect 14289 2465 14323 2499
rect 14841 2465 14875 2499
rect 16037 2465 16071 2499
rect 16589 2465 16623 2499
rect 18864 2465 18898 2499
rect 24660 2465 24694 2499
rect 10793 2329 10827 2363
rect 16221 2329 16255 2363
rect 1961 2261 1995 2295
rect 12817 2261 12851 2295
rect 19349 2261 19383 2295
rect 25145 2261 25179 2295
<< metal1 >>
rect 17494 26324 17500 26376
rect 17552 26364 17558 26376
rect 24762 26364 24768 26376
rect 17552 26336 24768 26364
rect 17552 26324 17558 26336
rect 24762 26324 24768 26336
rect 24820 26324 24826 26376
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 13814 25304 13820 25356
rect 13872 25353 13878 25356
rect 13872 25347 13910 25353
rect 13898 25313 13910 25347
rect 13872 25307 13910 25313
rect 13872 25304 13878 25307
rect 13955 25143 14013 25149
rect 13955 25109 13967 25143
rect 14001 25140 14013 25143
rect 14182 25140 14188 25152
rect 14001 25112 14188 25140
rect 14001 25109 14013 25112
rect 13955 25103 14013 25109
rect 14182 25100 14188 25112
rect 14240 25100 14246 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 2958 24828 2964 24880
rect 3016 24868 3022 24880
rect 12526 24868 12532 24880
rect 3016 24840 12532 24868
rect 3016 24828 3022 24840
rect 12526 24828 12532 24840
rect 12584 24828 12590 24880
rect 16666 24800 16672 24812
rect 16627 24772 16672 24800
rect 16666 24760 16672 24772
rect 16724 24760 16730 24812
rect 10664 24735 10722 24741
rect 10664 24701 10676 24735
rect 10710 24732 10722 24735
rect 13909 24735 13967 24741
rect 10710 24704 11192 24732
rect 10710 24701 10722 24704
rect 10664 24695 10722 24701
rect 10686 24556 10692 24608
rect 10744 24605 10750 24608
rect 11164 24605 11192 24704
rect 13909 24701 13921 24735
rect 13955 24732 13967 24735
rect 14274 24732 14280 24744
rect 13955 24704 14280 24732
rect 13955 24701 13967 24704
rect 13909 24695 13967 24701
rect 14274 24692 14280 24704
rect 14332 24732 14338 24744
rect 14461 24735 14519 24741
rect 14461 24732 14473 24735
rect 14332 24704 14473 24732
rect 14332 24692 14338 24704
rect 14461 24701 14473 24704
rect 14507 24701 14519 24735
rect 14461 24695 14519 24701
rect 14734 24692 14740 24744
rect 14792 24732 14798 24744
rect 15013 24735 15071 24741
rect 15013 24732 15025 24735
rect 14792 24704 15025 24732
rect 14792 24692 14798 24704
rect 15013 24701 15025 24704
rect 15059 24732 15071 24735
rect 15565 24735 15623 24741
rect 15565 24732 15577 24735
rect 15059 24704 15577 24732
rect 15059 24701 15071 24704
rect 15013 24695 15071 24701
rect 15565 24701 15577 24704
rect 15611 24701 15623 24735
rect 15565 24695 15623 24701
rect 16184 24735 16242 24741
rect 16184 24701 16196 24735
rect 16230 24732 16242 24735
rect 16684 24732 16712 24760
rect 16230 24704 16712 24732
rect 16230 24701 16242 24704
rect 16184 24695 16242 24701
rect 13814 24664 13820 24676
rect 13727 24636 13820 24664
rect 13814 24624 13820 24636
rect 13872 24664 13878 24676
rect 14752 24664 14780 24692
rect 17034 24664 17040 24676
rect 13872 24636 14780 24664
rect 15212 24636 17040 24664
rect 13872 24624 13878 24636
rect 10744 24599 10793 24605
rect 10744 24565 10747 24599
rect 10781 24565 10793 24599
rect 10744 24559 10793 24565
rect 11149 24599 11207 24605
rect 11149 24565 11161 24599
rect 11195 24596 11207 24599
rect 12066 24596 12072 24608
rect 11195 24568 12072 24596
rect 11195 24565 11207 24568
rect 11149 24559 11207 24565
rect 10744 24556 10750 24559
rect 12066 24556 12072 24568
rect 12124 24556 12130 24608
rect 14090 24596 14096 24608
rect 14051 24568 14096 24596
rect 14090 24556 14096 24568
rect 14148 24556 14154 24608
rect 15212 24605 15240 24636
rect 17034 24624 17040 24636
rect 17092 24624 17098 24676
rect 16298 24605 16304 24608
rect 15197 24599 15255 24605
rect 15197 24565 15209 24599
rect 15243 24565 15255 24599
rect 15197 24559 15255 24565
rect 16255 24599 16304 24605
rect 16255 24565 16267 24599
rect 16301 24565 16304 24599
rect 16255 24559 16304 24565
rect 16298 24556 16304 24559
rect 16356 24556 16362 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 10134 24392 10140 24404
rect 10095 24364 10140 24392
rect 10134 24352 10140 24364
rect 10192 24352 10198 24404
rect 11885 24395 11943 24401
rect 11885 24361 11897 24395
rect 11931 24392 11943 24395
rect 12894 24392 12900 24404
rect 11931 24364 12900 24392
rect 11931 24361 11943 24364
rect 11885 24355 11943 24361
rect 12894 24352 12900 24364
rect 12952 24352 12958 24404
rect 12989 24395 13047 24401
rect 12989 24361 13001 24395
rect 13035 24392 13047 24395
rect 13722 24392 13728 24404
rect 13035 24364 13728 24392
rect 13035 24361 13047 24364
rect 12989 24355 13047 24361
rect 13722 24352 13728 24364
rect 13780 24352 13786 24404
rect 14185 24395 14243 24401
rect 14185 24361 14197 24395
rect 14231 24392 14243 24395
rect 14826 24392 14832 24404
rect 14231 24364 14832 24392
rect 14231 24361 14243 24364
rect 14185 24355 14243 24361
rect 14826 24352 14832 24364
rect 14884 24352 14890 24404
rect 17037 24395 17095 24401
rect 17037 24361 17049 24395
rect 17083 24392 17095 24395
rect 17862 24392 17868 24404
rect 17083 24364 17868 24392
rect 17083 24361 17095 24364
rect 17037 24355 17095 24361
rect 17862 24352 17868 24364
rect 17920 24352 17926 24404
rect 13906 24284 13912 24336
rect 13964 24324 13970 24336
rect 14274 24324 14280 24336
rect 13964 24296 14280 24324
rect 13964 24284 13970 24296
rect 14274 24284 14280 24296
rect 14332 24284 14338 24336
rect 15470 24324 15476 24336
rect 15431 24296 15476 24324
rect 15470 24284 15476 24296
rect 15528 24284 15534 24336
rect 9950 24256 9956 24268
rect 9911 24228 9956 24256
rect 9950 24216 9956 24228
rect 10008 24216 10014 24268
rect 11698 24256 11704 24268
rect 11659 24228 11704 24256
rect 11698 24216 11704 24228
rect 11756 24216 11762 24268
rect 12805 24259 12863 24265
rect 12805 24225 12817 24259
rect 12851 24256 12863 24259
rect 13538 24256 13544 24268
rect 12851 24228 13544 24256
rect 12851 24225 12863 24228
rect 12805 24219 12863 24225
rect 13538 24216 13544 24228
rect 13596 24216 13602 24268
rect 14001 24259 14059 24265
rect 14001 24225 14013 24259
rect 14047 24256 14059 24259
rect 14642 24256 14648 24268
rect 14047 24228 14648 24256
rect 14047 24225 14059 24228
rect 14001 24219 14059 24225
rect 14642 24216 14648 24228
rect 14700 24216 14706 24268
rect 16574 24216 16580 24268
rect 16632 24256 16638 24268
rect 18322 24265 18328 24268
rect 16853 24259 16911 24265
rect 16853 24256 16865 24259
rect 16632 24228 16865 24256
rect 16632 24216 16638 24228
rect 16853 24225 16865 24228
rect 16899 24225 16911 24259
rect 16853 24219 16911 24225
rect 18300 24259 18328 24265
rect 18300 24225 18312 24259
rect 18300 24219 18328 24225
rect 18322 24216 18328 24219
rect 18380 24216 18386 24268
rect 15381 24191 15439 24197
rect 15381 24157 15393 24191
rect 15427 24188 15439 24191
rect 16022 24188 16028 24200
rect 15427 24160 15884 24188
rect 15983 24160 16028 24188
rect 15427 24157 15439 24160
rect 15381 24151 15439 24157
rect 15286 24080 15292 24132
rect 15344 24120 15350 24132
rect 15396 24120 15424 24151
rect 15344 24092 15424 24120
rect 15344 24080 15350 24092
rect 12618 24052 12624 24064
rect 12579 24024 12624 24052
rect 12618 24012 12624 24024
rect 12676 24012 12682 24064
rect 15856 24052 15884 24160
rect 16022 24148 16028 24160
rect 16080 24148 16086 24200
rect 16390 24120 16396 24132
rect 16351 24092 16396 24120
rect 16390 24080 16396 24092
rect 16448 24080 16454 24132
rect 18371 24055 18429 24061
rect 18371 24052 18383 24055
rect 15856 24024 18383 24052
rect 18371 24021 18383 24024
rect 18417 24021 18429 24055
rect 18371 24015 18429 24021
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 3605 23851 3663 23857
rect 3605 23817 3617 23851
rect 3651 23848 3663 23851
rect 4614 23848 4620 23860
rect 3651 23820 4620 23848
rect 3651 23817 3663 23820
rect 3605 23811 3663 23817
rect 1857 23715 1915 23721
rect 1857 23712 1869 23715
rect 1412 23684 1869 23712
rect 474 23604 480 23656
rect 532 23644 538 23656
rect 1412 23653 1440 23684
rect 1857 23681 1869 23684
rect 1903 23681 1915 23715
rect 1857 23675 1915 23681
rect 1412 23647 1490 23653
rect 1412 23644 1444 23647
rect 532 23616 1444 23644
rect 532 23604 538 23616
rect 1432 23613 1444 23616
rect 1478 23613 1490 23647
rect 1432 23607 1490 23613
rect 1535 23647 1593 23653
rect 1535 23613 1547 23647
rect 1581 23644 1593 23647
rect 2682 23644 2688 23656
rect 1581 23616 2688 23644
rect 1581 23613 1593 23616
rect 1535 23607 1593 23613
rect 2682 23604 2688 23616
rect 2740 23604 2746 23656
rect 3120 23647 3178 23653
rect 3120 23613 3132 23647
rect 3166 23644 3178 23647
rect 3620 23644 3648 23811
rect 4614 23808 4620 23820
rect 4672 23808 4678 23860
rect 7929 23851 7987 23857
rect 7929 23817 7941 23851
rect 7975 23848 7987 23851
rect 8754 23848 8760 23860
rect 7975 23820 8760 23848
rect 7975 23817 7987 23820
rect 7929 23811 7987 23817
rect 3166 23616 3648 23644
rect 7444 23647 7502 23653
rect 3166 23613 3178 23616
rect 3120 23607 3178 23613
rect 7444 23613 7456 23647
rect 7490 23644 7502 23647
rect 7944 23644 7972 23811
rect 8754 23808 8760 23820
rect 8812 23808 8818 23860
rect 9125 23851 9183 23857
rect 9125 23817 9137 23851
rect 9171 23848 9183 23851
rect 9582 23848 9588 23860
rect 9171 23820 9588 23848
rect 9171 23817 9183 23820
rect 9125 23811 9183 23817
rect 7490 23616 7972 23644
rect 8640 23647 8698 23653
rect 7490 23613 7502 23616
rect 7444 23607 7502 23613
rect 8640 23613 8652 23647
rect 8686 23644 8698 23647
rect 9140 23644 9168 23811
rect 9582 23808 9588 23820
rect 9640 23808 9646 23860
rect 10686 23848 10692 23860
rect 10647 23820 10692 23848
rect 10686 23808 10692 23820
rect 10744 23808 10750 23860
rect 15381 23851 15439 23857
rect 15381 23817 15393 23851
rect 15427 23848 15439 23851
rect 15470 23848 15476 23860
rect 15427 23820 15476 23848
rect 15427 23817 15439 23820
rect 15381 23811 15439 23817
rect 15470 23808 15476 23820
rect 15528 23808 15534 23860
rect 18233 23851 18291 23857
rect 18233 23817 18245 23851
rect 18279 23848 18291 23851
rect 19058 23848 19064 23860
rect 18279 23820 19064 23848
rect 18279 23817 18291 23820
rect 18233 23811 18291 23817
rect 19058 23808 19064 23820
rect 19116 23808 19122 23860
rect 20809 23851 20867 23857
rect 20809 23817 20821 23851
rect 20855 23848 20867 23851
rect 22186 23848 22192 23860
rect 20855 23820 22192 23848
rect 20855 23817 20867 23820
rect 20809 23811 20867 23817
rect 8686 23616 9168 23644
rect 10137 23647 10195 23653
rect 8686 23613 8698 23616
rect 8640 23607 8698 23613
rect 10137 23613 10149 23647
rect 10183 23644 10195 23647
rect 10704 23644 10732 23808
rect 16022 23740 16028 23792
rect 16080 23780 16086 23792
rect 16301 23783 16359 23789
rect 16301 23780 16313 23783
rect 16080 23752 16313 23780
rect 16080 23740 16086 23752
rect 16301 23749 16313 23752
rect 16347 23749 16359 23783
rect 16301 23743 16359 23749
rect 18322 23740 18328 23792
rect 18380 23780 18386 23792
rect 18601 23783 18659 23789
rect 18601 23780 18613 23783
rect 18380 23752 18613 23780
rect 18380 23740 18386 23752
rect 18601 23749 18613 23752
rect 18647 23749 18659 23783
rect 18601 23743 18659 23749
rect 12250 23712 12256 23724
rect 12211 23684 12256 23712
rect 12250 23672 12256 23684
rect 12308 23672 12314 23724
rect 14182 23712 14188 23724
rect 14143 23684 14188 23712
rect 14182 23672 14188 23684
rect 14240 23672 14246 23724
rect 14274 23672 14280 23724
rect 14332 23712 14338 23724
rect 14461 23715 14519 23721
rect 14461 23712 14473 23715
rect 14332 23684 14473 23712
rect 14332 23672 14338 23684
rect 14461 23681 14473 23684
rect 14507 23681 14519 23715
rect 14461 23675 14519 23681
rect 15749 23715 15807 23721
rect 15749 23681 15761 23715
rect 15795 23712 15807 23715
rect 16390 23712 16396 23724
rect 15795 23684 16396 23712
rect 15795 23681 15807 23684
rect 15749 23675 15807 23681
rect 16390 23672 16396 23684
rect 16448 23672 16454 23724
rect 19291 23715 19349 23721
rect 19291 23712 19303 23715
rect 18064 23684 19303 23712
rect 10183 23616 10732 23644
rect 11400 23647 11458 23653
rect 10183 23613 10195 23616
rect 10137 23607 10195 23613
rect 11400 23613 11412 23647
rect 11446 23644 11458 23647
rect 12268 23644 12296 23672
rect 12710 23644 12716 23656
rect 11446 23616 12296 23644
rect 12671 23616 12716 23644
rect 11446 23613 11458 23616
rect 11400 23607 11458 23613
rect 12710 23604 12716 23616
rect 12768 23604 12774 23656
rect 18064 23653 18092 23684
rect 19291 23681 19303 23684
rect 19337 23681 19349 23715
rect 19291 23675 19349 23681
rect 12989 23647 13047 23653
rect 12989 23613 13001 23647
rect 13035 23613 13047 23647
rect 12989 23607 13047 23613
rect 17865 23647 17923 23653
rect 17865 23613 17877 23647
rect 17911 23644 17923 23647
rect 18049 23647 18107 23653
rect 18049 23644 18061 23647
rect 17911 23616 18061 23644
rect 17911 23613 17923 23616
rect 17865 23607 17923 23613
rect 18049 23613 18061 23616
rect 18095 23613 18107 23647
rect 18049 23607 18107 23613
rect 19204 23647 19262 23653
rect 19204 23613 19216 23647
rect 19250 23644 19262 23647
rect 20324 23647 20382 23653
rect 19250 23616 19472 23644
rect 19250 23613 19262 23616
rect 19204 23607 19262 23613
rect 12618 23536 12624 23588
rect 12676 23576 12682 23588
rect 13004 23576 13032 23607
rect 13262 23576 13268 23588
rect 12676 23548 13032 23576
rect 13223 23548 13268 23576
rect 12676 23536 12682 23548
rect 13262 23536 13268 23548
rect 13320 23536 13326 23588
rect 14001 23579 14059 23585
rect 14001 23545 14013 23579
rect 14047 23576 14059 23579
rect 14277 23579 14335 23585
rect 14277 23576 14289 23579
rect 14047 23548 14289 23576
rect 14047 23545 14059 23548
rect 14001 23539 14059 23545
rect 14108 23520 14136 23548
rect 14277 23545 14289 23548
rect 14323 23576 14335 23579
rect 15010 23576 15016 23588
rect 14323 23548 15016 23576
rect 14323 23545 14335 23548
rect 14277 23539 14335 23545
rect 15010 23536 15016 23548
rect 15068 23536 15074 23588
rect 15838 23536 15844 23588
rect 15896 23576 15902 23588
rect 15896 23548 15941 23576
rect 15896 23536 15902 23548
rect 19444 23520 19472 23616
rect 20324 23613 20336 23647
rect 20370 23644 20382 23647
rect 20824 23644 20852 23811
rect 22186 23808 22192 23820
rect 22244 23808 22250 23860
rect 23474 23808 23480 23860
rect 23532 23848 23538 23860
rect 24535 23851 24593 23857
rect 24535 23848 24547 23851
rect 23532 23820 24547 23848
rect 23532 23808 23538 23820
rect 24535 23817 24547 23820
rect 24581 23817 24593 23851
rect 24535 23811 24593 23817
rect 24949 23851 25007 23857
rect 24949 23817 24961 23851
rect 24995 23848 25007 23851
rect 26142 23848 26148 23860
rect 24995 23820 26148 23848
rect 24995 23817 25007 23820
rect 24949 23811 25007 23817
rect 20370 23616 20852 23644
rect 24464 23647 24522 23653
rect 20370 23613 20382 23616
rect 20324 23607 20382 23613
rect 24464 23613 24476 23647
rect 24510 23644 24522 23647
rect 24964 23644 24992 23811
rect 26142 23808 26148 23820
rect 26200 23808 26206 23860
rect 24510 23616 24992 23644
rect 24510 23613 24522 23616
rect 24464 23607 24522 23613
rect 2866 23468 2872 23520
rect 2924 23508 2930 23520
rect 7558 23517 7564 23520
rect 3191 23511 3249 23517
rect 3191 23508 3203 23511
rect 2924 23480 3203 23508
rect 2924 23468 2930 23480
rect 3191 23477 3203 23480
rect 3237 23477 3249 23511
rect 3191 23471 3249 23477
rect 7515 23511 7564 23517
rect 7515 23477 7527 23511
rect 7561 23477 7564 23511
rect 7515 23471 7564 23477
rect 7558 23468 7564 23471
rect 7616 23468 7622 23520
rect 8711 23511 8769 23517
rect 8711 23477 8723 23511
rect 8757 23508 8769 23511
rect 8846 23508 8852 23520
rect 8757 23480 8852 23508
rect 8757 23477 8769 23480
rect 8711 23471 8769 23477
rect 8846 23468 8852 23480
rect 8904 23468 8910 23520
rect 9950 23508 9956 23520
rect 9911 23480 9956 23508
rect 9950 23468 9956 23480
rect 10008 23468 10014 23520
rect 10321 23511 10379 23517
rect 10321 23477 10333 23511
rect 10367 23508 10379 23511
rect 10778 23508 10784 23520
rect 10367 23480 10784 23508
rect 10367 23477 10379 23480
rect 10321 23471 10379 23477
rect 10778 23468 10784 23480
rect 10836 23468 10842 23520
rect 11330 23468 11336 23520
rect 11388 23508 11394 23520
rect 11471 23511 11529 23517
rect 11471 23508 11483 23511
rect 11388 23480 11483 23508
rect 11388 23468 11394 23480
rect 11471 23477 11483 23480
rect 11517 23477 11529 23511
rect 11471 23471 11529 23477
rect 11698 23468 11704 23520
rect 11756 23508 11762 23520
rect 11885 23511 11943 23517
rect 11885 23508 11897 23511
rect 11756 23480 11897 23508
rect 11756 23468 11762 23480
rect 11885 23477 11897 23480
rect 11931 23508 11943 23511
rect 12434 23508 12440 23520
rect 11931 23480 12440 23508
rect 11931 23477 11943 23480
rect 11885 23471 11943 23477
rect 12434 23468 12440 23480
rect 12492 23468 12498 23520
rect 13538 23508 13544 23520
rect 13499 23480 13544 23508
rect 13538 23468 13544 23480
rect 13596 23468 13602 23520
rect 14090 23468 14096 23520
rect 14148 23468 14154 23520
rect 16574 23468 16580 23520
rect 16632 23508 16638 23520
rect 16853 23511 16911 23517
rect 16853 23508 16865 23511
rect 16632 23480 16865 23508
rect 16632 23468 16638 23480
rect 16853 23477 16865 23480
rect 16899 23477 16911 23511
rect 16853 23471 16911 23477
rect 19426 23468 19432 23520
rect 19484 23508 19490 23520
rect 19613 23511 19671 23517
rect 19613 23508 19625 23511
rect 19484 23480 19625 23508
rect 19484 23468 19490 23480
rect 19613 23477 19625 23480
rect 19659 23477 19671 23511
rect 19613 23471 19671 23477
rect 19978 23468 19984 23520
rect 20036 23508 20042 23520
rect 20395 23511 20453 23517
rect 20395 23508 20407 23511
rect 20036 23480 20407 23508
rect 20036 23468 20042 23480
rect 20395 23477 20407 23480
rect 20441 23477 20453 23511
rect 20395 23471 20453 23477
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 12728 23276 13124 23304
rect 9858 23236 9864 23248
rect 9819 23208 9864 23236
rect 9858 23196 9864 23208
rect 9916 23196 9922 23248
rect 11149 23239 11207 23245
rect 11149 23205 11161 23239
rect 11195 23236 11207 23239
rect 11330 23236 11336 23248
rect 11195 23208 11336 23236
rect 11195 23205 11207 23208
rect 11149 23199 11207 23205
rect 11330 23196 11336 23208
rect 11388 23196 11394 23248
rect 11422 23196 11428 23248
rect 11480 23236 11486 23248
rect 11480 23208 11525 23236
rect 11480 23196 11486 23208
rect 9766 23100 9772 23112
rect 9727 23072 9772 23100
rect 9766 23060 9772 23072
rect 9824 23060 9830 23112
rect 10413 23103 10471 23109
rect 10413 23069 10425 23103
rect 10459 23100 10471 23103
rect 11609 23103 11667 23109
rect 11609 23100 11621 23103
rect 10459 23072 11621 23100
rect 10459 23069 10471 23072
rect 10413 23063 10471 23069
rect 11256 23044 11284 23072
rect 11609 23069 11621 23072
rect 11655 23100 11667 23103
rect 12728 23100 12756 23276
rect 12986 23236 12992 23248
rect 12947 23208 12992 23236
rect 12986 23196 12992 23208
rect 13044 23196 13050 23248
rect 13096 23236 13124 23276
rect 13262 23264 13268 23316
rect 13320 23304 13326 23316
rect 13630 23304 13636 23316
rect 13320 23276 13636 23304
rect 13320 23264 13326 23276
rect 13630 23264 13636 23276
rect 13688 23304 13694 23316
rect 13817 23307 13875 23313
rect 13817 23304 13829 23307
rect 13688 23276 13829 23304
rect 13688 23264 13694 23276
rect 13817 23273 13829 23276
rect 13863 23273 13875 23307
rect 14182 23304 14188 23316
rect 14143 23276 14188 23304
rect 13817 23267 13875 23273
rect 14182 23264 14188 23276
rect 14240 23264 14246 23316
rect 15102 23304 15108 23316
rect 15063 23276 15108 23304
rect 15102 23264 15108 23276
rect 15160 23264 15166 23316
rect 16991 23307 17049 23313
rect 16991 23304 17003 23307
rect 15304 23276 17003 23304
rect 13541 23239 13599 23245
rect 13541 23236 13553 23239
rect 13096 23208 13553 23236
rect 13541 23205 13553 23208
rect 13587 23205 13599 23239
rect 14642 23236 14648 23248
rect 14555 23208 14648 23236
rect 13541 23199 13599 23205
rect 14642 23196 14648 23208
rect 14700 23236 14706 23248
rect 15304 23236 15332 23276
rect 16991 23273 17003 23276
rect 17037 23273 17049 23307
rect 16991 23267 17049 23273
rect 15470 23236 15476 23248
rect 14700 23208 15332 23236
rect 15431 23208 15476 23236
rect 14700 23196 14706 23208
rect 15470 23196 15476 23208
rect 15528 23196 15534 23248
rect 18506 23196 18512 23248
rect 18564 23236 18570 23248
rect 18785 23239 18843 23245
rect 18785 23236 18797 23239
rect 18564 23208 18797 23236
rect 18564 23196 18570 23208
rect 18785 23205 18797 23208
rect 18831 23205 18843 23239
rect 18785 23199 18843 23205
rect 16888 23171 16946 23177
rect 16888 23168 16900 23171
rect 16224 23140 16900 23168
rect 12894 23100 12900 23112
rect 11655 23072 12756 23100
rect 12855 23072 12900 23100
rect 11655 23069 11667 23072
rect 11609 23063 11667 23069
rect 12894 23060 12900 23072
rect 12952 23060 12958 23112
rect 15381 23103 15439 23109
rect 15381 23069 15393 23103
rect 15427 23100 15439 23103
rect 16022 23100 16028 23112
rect 15427 23072 16028 23100
rect 15427 23069 15439 23072
rect 15381 23063 15439 23069
rect 16022 23060 16028 23072
rect 16080 23060 16086 23112
rect 11238 22992 11244 23044
rect 11296 22992 11302 23044
rect 14826 22992 14832 23044
rect 14884 23032 14890 23044
rect 15933 23035 15991 23041
rect 15933 23032 15945 23035
rect 14884 23004 15945 23032
rect 14884 22992 14890 23004
rect 15933 23001 15945 23004
rect 15979 23032 15991 23035
rect 16224 23032 16252 23140
rect 16888 23137 16900 23140
rect 16934 23168 16946 23171
rect 17126 23168 17132 23180
rect 16934 23140 17132 23168
rect 16934 23137 16946 23140
rect 16888 23131 16946 23137
rect 17126 23128 17132 23140
rect 17184 23128 17190 23180
rect 20968 23171 21026 23177
rect 20968 23137 20980 23171
rect 21014 23168 21026 23171
rect 21174 23168 21180 23180
rect 21014 23140 21180 23168
rect 21014 23137 21026 23140
rect 20968 23131 21026 23137
rect 21174 23128 21180 23140
rect 21232 23128 21238 23180
rect 24670 23177 24676 23180
rect 24648 23171 24676 23177
rect 24648 23137 24660 23171
rect 24648 23131 24676 23137
rect 24670 23128 24676 23131
rect 24728 23128 24734 23180
rect 17862 23060 17868 23112
rect 17920 23100 17926 23112
rect 18693 23103 18751 23109
rect 18693 23100 18705 23103
rect 17920 23072 18705 23100
rect 17920 23060 17926 23072
rect 18693 23069 18705 23072
rect 18739 23100 18751 23103
rect 18739 23072 20760 23100
rect 18739 23069 18751 23072
rect 18693 23063 18751 23069
rect 19242 23032 19248 23044
rect 15979 23004 16252 23032
rect 19203 23004 19248 23032
rect 15979 23001 15991 23004
rect 15933 22995 15991 23001
rect 19242 22992 19248 23004
rect 19300 22992 19306 23044
rect 20732 23032 20760 23072
rect 21039 23035 21097 23041
rect 21039 23032 21051 23035
rect 20732 23004 21051 23032
rect 21039 23001 21051 23004
rect 21085 23001 21097 23035
rect 21039 22995 21097 23001
rect 12621 22967 12679 22973
rect 12621 22933 12633 22967
rect 12667 22964 12679 22967
rect 12710 22964 12716 22976
rect 12667 22936 12716 22964
rect 12667 22933 12679 22936
rect 12621 22927 12679 22933
rect 12710 22924 12716 22936
rect 12768 22964 12774 22976
rect 13078 22964 13084 22976
rect 12768 22936 13084 22964
rect 12768 22924 12774 22936
rect 13078 22924 13084 22936
rect 13136 22924 13142 22976
rect 15838 22924 15844 22976
rect 15896 22964 15902 22976
rect 16301 22967 16359 22973
rect 16301 22964 16313 22967
rect 15896 22936 16313 22964
rect 15896 22924 15902 22936
rect 16301 22933 16313 22936
rect 16347 22933 16359 22967
rect 16301 22927 16359 22933
rect 23474 22924 23480 22976
rect 23532 22964 23538 22976
rect 24719 22967 24777 22973
rect 24719 22964 24731 22967
rect 23532 22936 24731 22964
rect 23532 22924 23538 22936
rect 24719 22933 24731 22936
rect 24765 22933 24777 22967
rect 24719 22927 24777 22933
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 9766 22720 9772 22772
rect 9824 22760 9830 22772
rect 10045 22763 10103 22769
rect 10045 22760 10057 22763
rect 9824 22732 10057 22760
rect 9824 22720 9830 22732
rect 10045 22729 10057 22732
rect 10091 22729 10103 22763
rect 10045 22723 10103 22729
rect 12253 22763 12311 22769
rect 12253 22729 12265 22763
rect 12299 22760 12311 22763
rect 12894 22760 12900 22772
rect 12299 22732 12900 22760
rect 12299 22729 12311 22732
rect 12253 22723 12311 22729
rect 12894 22720 12900 22732
rect 12952 22720 12958 22772
rect 14553 22763 14611 22769
rect 14553 22729 14565 22763
rect 14599 22760 14611 22763
rect 14921 22763 14979 22769
rect 14921 22760 14933 22763
rect 14599 22732 14933 22760
rect 14599 22729 14611 22732
rect 14553 22723 14611 22729
rect 14921 22729 14933 22732
rect 14967 22760 14979 22763
rect 15470 22760 15476 22772
rect 14967 22732 15476 22760
rect 14967 22729 14979 22732
rect 14921 22723 14979 22729
rect 15470 22720 15476 22732
rect 15528 22720 15534 22772
rect 16298 22760 16304 22772
rect 15856 22732 16304 22760
rect 12526 22652 12532 22704
rect 12584 22692 12590 22704
rect 12710 22692 12716 22704
rect 12584 22664 12716 22692
rect 12584 22652 12590 22664
rect 12710 22652 12716 22664
rect 12768 22652 12774 22704
rect 15286 22692 15292 22704
rect 15247 22664 15292 22692
rect 15286 22652 15292 22664
rect 15344 22652 15350 22704
rect 10505 22627 10563 22633
rect 10505 22593 10517 22627
rect 10551 22624 10563 22627
rect 10870 22624 10876 22636
rect 10551 22596 10876 22624
rect 10551 22593 10563 22596
rect 10505 22587 10563 22593
rect 10870 22584 10876 22596
rect 10928 22624 10934 22636
rect 13449 22627 13507 22633
rect 13449 22624 13461 22627
rect 10928 22596 13461 22624
rect 10928 22584 10934 22596
rect 10597 22559 10655 22565
rect 10597 22525 10609 22559
rect 10643 22556 10655 22559
rect 10686 22556 10692 22568
rect 10643 22528 10692 22556
rect 10643 22525 10655 22528
rect 10597 22519 10655 22525
rect 10686 22516 10692 22528
rect 10744 22516 10750 22568
rect 10980 22497 11008 22596
rect 13449 22593 13461 22596
rect 13495 22593 13507 22627
rect 13630 22624 13636 22636
rect 13591 22596 13636 22624
rect 13449 22587 13507 22593
rect 12526 22565 12532 22568
rect 12504 22559 12532 22565
rect 12504 22525 12516 22559
rect 12584 22556 12590 22568
rect 12897 22559 12955 22565
rect 12897 22556 12909 22559
rect 12584 22528 12909 22556
rect 12504 22519 12532 22525
rect 12526 22516 12532 22519
rect 12584 22516 12590 22528
rect 12897 22525 12909 22528
rect 12943 22525 12955 22559
rect 12897 22519 12955 22525
rect 10938 22491 11008 22497
rect 10938 22457 10950 22491
rect 10984 22460 11008 22491
rect 10984 22457 10996 22460
rect 10938 22451 10996 22457
rect 11146 22448 11152 22500
rect 11204 22488 11210 22500
rect 11422 22488 11428 22500
rect 11204 22460 11428 22488
rect 11204 22448 11210 22460
rect 11422 22448 11428 22460
rect 11480 22488 11486 22500
rect 11793 22491 11851 22497
rect 11793 22488 11805 22491
rect 11480 22460 11805 22488
rect 11480 22448 11486 22460
rect 11793 22457 11805 22460
rect 11839 22457 11851 22491
rect 13464 22488 13492 22587
rect 13630 22584 13636 22596
rect 13688 22584 13694 22636
rect 15473 22627 15531 22633
rect 15473 22593 15485 22627
rect 15519 22624 15531 22627
rect 15856 22624 15884 22732
rect 16298 22720 16304 22732
rect 16356 22760 16362 22772
rect 16393 22763 16451 22769
rect 16393 22760 16405 22763
rect 16356 22732 16405 22760
rect 16356 22720 16362 22732
rect 16393 22729 16405 22732
rect 16439 22729 16451 22763
rect 17126 22760 17132 22772
rect 17087 22732 17132 22760
rect 16393 22723 16451 22729
rect 17126 22720 17132 22732
rect 17184 22720 17190 22772
rect 17862 22760 17868 22772
rect 17823 22732 17868 22760
rect 17862 22720 17868 22732
rect 17920 22720 17926 22772
rect 19794 22760 19800 22772
rect 19755 22732 19800 22760
rect 19794 22720 19800 22732
rect 19852 22720 19858 22772
rect 20162 22760 20168 22772
rect 20123 22732 20168 22760
rect 20162 22720 20168 22732
rect 20220 22720 20226 22772
rect 20993 22763 21051 22769
rect 20993 22729 21005 22763
rect 21039 22760 21051 22763
rect 21174 22760 21180 22772
rect 21039 22732 21180 22760
rect 21039 22729 21051 22732
rect 20993 22723 21051 22729
rect 21174 22720 21180 22732
rect 21232 22720 21238 22772
rect 24670 22760 24676 22772
rect 24631 22732 24676 22760
rect 24670 22720 24676 22732
rect 24728 22720 24734 22772
rect 16022 22692 16028 22704
rect 15983 22664 16028 22692
rect 16022 22652 16028 22664
rect 16080 22692 16086 22704
rect 16761 22695 16819 22701
rect 16761 22692 16773 22695
rect 16080 22664 16773 22692
rect 16080 22652 16086 22664
rect 16761 22661 16773 22664
rect 16807 22661 16819 22695
rect 19812 22692 19840 22720
rect 16761 22655 16819 22661
rect 18800 22664 19840 22692
rect 18800 22633 18828 22664
rect 15519 22596 15884 22624
rect 18785 22627 18843 22633
rect 15519 22593 15531 22596
rect 15473 22587 15531 22593
rect 18785 22593 18797 22627
rect 18831 22593 18843 22627
rect 19242 22624 19248 22636
rect 19203 22596 19248 22624
rect 18785 22587 18843 22593
rect 19242 22584 19248 22596
rect 19300 22584 19306 22636
rect 20162 22516 20168 22568
rect 20220 22556 20226 22568
rect 20292 22559 20350 22565
rect 20292 22556 20304 22559
rect 20220 22528 20304 22556
rect 20220 22516 20226 22528
rect 20292 22525 20304 22528
rect 20338 22525 20350 22559
rect 20292 22519 20350 22525
rect 13630 22488 13636 22500
rect 13464 22460 13636 22488
rect 11793 22451 11851 22457
rect 13630 22448 13636 22460
rect 13688 22488 13694 22500
rect 13954 22491 14012 22497
rect 13954 22488 13966 22491
rect 13688 22460 13966 22488
rect 13688 22448 13694 22460
rect 13954 22457 13966 22460
rect 14000 22457 14012 22491
rect 13954 22451 14012 22457
rect 15286 22448 15292 22500
rect 15344 22488 15350 22500
rect 15565 22491 15623 22497
rect 15565 22488 15577 22491
rect 15344 22460 15577 22488
rect 15344 22448 15350 22460
rect 15565 22457 15577 22460
rect 15611 22457 15623 22491
rect 15565 22451 15623 22457
rect 18874 22448 18880 22500
rect 18932 22488 18938 22500
rect 20395 22491 20453 22497
rect 20395 22488 20407 22491
rect 18932 22460 18977 22488
rect 19352 22460 20407 22488
rect 18932 22448 18938 22460
rect 19352 22432 19380 22460
rect 20395 22457 20407 22460
rect 20441 22457 20453 22491
rect 20395 22451 20453 22457
rect 9769 22423 9827 22429
rect 9769 22389 9781 22423
rect 9815 22420 9827 22423
rect 9858 22420 9864 22432
rect 9815 22392 9864 22420
rect 9815 22389 9827 22392
rect 9769 22383 9827 22389
rect 9858 22380 9864 22392
rect 9916 22380 9922 22432
rect 11514 22420 11520 22432
rect 11475 22392 11520 22420
rect 11514 22380 11520 22392
rect 11572 22380 11578 22432
rect 12575 22423 12633 22429
rect 12575 22389 12587 22423
rect 12621 22420 12633 22423
rect 12710 22420 12716 22432
rect 12621 22392 12716 22420
rect 12621 22389 12633 22392
rect 12575 22383 12633 22389
rect 12710 22380 12716 22392
rect 12768 22380 12774 22432
rect 18046 22380 18052 22432
rect 18104 22420 18110 22432
rect 18506 22420 18512 22432
rect 18104 22392 18512 22420
rect 18104 22380 18110 22392
rect 18506 22380 18512 22392
rect 18564 22380 18570 22432
rect 19334 22380 19340 22432
rect 19392 22380 19398 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 12897 22219 12955 22225
rect 12897 22185 12909 22219
rect 12943 22216 12955 22219
rect 12986 22216 12992 22228
rect 12943 22188 12992 22216
rect 12943 22185 12955 22188
rect 12897 22179 12955 22185
rect 12986 22176 12992 22188
rect 13044 22176 13050 22228
rect 18049 22219 18107 22225
rect 18049 22185 18061 22219
rect 18095 22216 18107 22219
rect 18095 22188 19104 22216
rect 18095 22185 18107 22188
rect 18049 22179 18107 22185
rect 19076 22160 19104 22188
rect 11238 22148 11244 22160
rect 11199 22120 11244 22148
rect 11238 22108 11244 22120
rect 11296 22108 11302 22160
rect 11333 22151 11391 22157
rect 11333 22117 11345 22151
rect 11379 22148 11391 22151
rect 11514 22148 11520 22160
rect 11379 22120 11520 22148
rect 11379 22117 11391 22120
rect 11333 22111 11391 22117
rect 11514 22108 11520 22120
rect 11572 22108 11578 22160
rect 13722 22148 13728 22160
rect 13683 22120 13728 22148
rect 13722 22108 13728 22120
rect 13780 22108 13786 22160
rect 16206 22148 16212 22160
rect 16167 22120 16212 22148
rect 16206 22108 16212 22120
rect 16264 22108 16270 22160
rect 17494 22157 17500 22160
rect 17491 22148 17500 22157
rect 17455 22120 17500 22148
rect 17491 22111 17500 22120
rect 17494 22108 17500 22111
rect 17552 22108 17558 22160
rect 18782 22148 18788 22160
rect 18743 22120 18788 22148
rect 18782 22108 18788 22120
rect 18840 22108 18846 22160
rect 19058 22148 19064 22160
rect 18971 22120 19064 22148
rect 19058 22108 19064 22120
rect 19116 22108 19122 22160
rect 14274 22040 14280 22092
rect 14332 22080 14338 22092
rect 14332 22052 14377 22080
rect 14332 22040 14338 22052
rect 15378 22040 15384 22092
rect 15436 22080 15442 22092
rect 15473 22083 15531 22089
rect 15473 22080 15485 22083
rect 15436 22052 15485 22080
rect 15436 22040 15442 22052
rect 15473 22049 15485 22052
rect 15519 22049 15531 22083
rect 15473 22043 15531 22049
rect 16025 22083 16083 22089
rect 16025 22049 16037 22083
rect 16071 22080 16083 22083
rect 16482 22080 16488 22092
rect 16071 22052 16488 22080
rect 16071 22049 16083 22052
rect 16025 22043 16083 22049
rect 16482 22040 16488 22052
rect 16540 22040 16546 22092
rect 11885 22015 11943 22021
rect 11885 21981 11897 22015
rect 11931 22012 11943 22015
rect 12066 22012 12072 22024
rect 11931 21984 12072 22012
rect 11931 21981 11943 21984
rect 11885 21975 11943 21981
rect 12066 21972 12072 21984
rect 12124 21972 12130 22024
rect 12802 21972 12808 22024
rect 12860 22012 12866 22024
rect 13633 22015 13691 22021
rect 13633 22012 13645 22015
rect 12860 21984 13645 22012
rect 12860 21972 12866 21984
rect 13633 21981 13645 21984
rect 13679 21981 13691 22015
rect 17126 22012 17132 22024
rect 17087 21984 17132 22012
rect 13633 21975 13691 21981
rect 17126 21972 17132 21984
rect 17184 21972 17190 22024
rect 18966 22012 18972 22024
rect 18927 21984 18972 22012
rect 18966 21972 18972 21984
rect 19024 22012 19030 22024
rect 19242 22012 19248 22024
rect 19024 21984 19248 22012
rect 19024 21972 19030 21984
rect 19242 21972 19248 21984
rect 19300 21972 19306 22024
rect 19426 22012 19432 22024
rect 19387 21984 19432 22012
rect 19426 21972 19432 21984
rect 19484 21972 19490 22024
rect 8481 21879 8539 21885
rect 8481 21845 8493 21879
rect 8527 21876 8539 21879
rect 8938 21876 8944 21888
rect 8527 21848 8944 21876
rect 8527 21845 8539 21848
rect 8481 21839 8539 21845
rect 8938 21836 8944 21848
rect 8996 21836 9002 21888
rect 9122 21836 9128 21888
rect 9180 21876 9186 21888
rect 10597 21879 10655 21885
rect 10597 21876 10609 21879
rect 9180 21848 10609 21876
rect 9180 21836 9186 21848
rect 10597 21845 10609 21848
rect 10643 21876 10655 21879
rect 10686 21876 10692 21888
rect 10643 21848 10692 21876
rect 10643 21845 10655 21848
rect 10597 21839 10655 21845
rect 10686 21836 10692 21848
rect 10744 21836 10750 21888
rect 13998 21836 14004 21888
rect 14056 21876 14062 21888
rect 14553 21879 14611 21885
rect 14553 21876 14565 21879
rect 14056 21848 14565 21876
rect 14056 21836 14062 21848
rect 14553 21845 14565 21848
rect 14599 21845 14611 21879
rect 16482 21876 16488 21888
rect 16443 21848 16488 21876
rect 14553 21839 14611 21845
rect 16482 21836 16488 21848
rect 16540 21836 16546 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 9858 21632 9864 21684
rect 9916 21672 9922 21684
rect 10873 21675 10931 21681
rect 10873 21672 10885 21675
rect 9916 21644 10885 21672
rect 9916 21632 9922 21644
rect 10873 21641 10885 21644
rect 10919 21641 10931 21675
rect 10873 21635 10931 21641
rect 11238 21632 11244 21684
rect 11296 21672 11302 21684
rect 11517 21675 11575 21681
rect 11517 21672 11529 21675
rect 11296 21644 11529 21672
rect 11296 21632 11302 21644
rect 11517 21641 11529 21644
rect 11563 21641 11575 21675
rect 12802 21672 12808 21684
rect 12763 21644 12808 21672
rect 11517 21635 11575 21641
rect 12802 21632 12808 21644
rect 12860 21632 12866 21684
rect 13814 21672 13820 21684
rect 13775 21644 13820 21672
rect 13814 21632 13820 21644
rect 13872 21632 13878 21684
rect 19058 21632 19064 21684
rect 19116 21672 19122 21684
rect 19613 21675 19671 21681
rect 19613 21672 19625 21675
rect 19116 21644 19625 21672
rect 19116 21632 19122 21644
rect 19613 21641 19625 21644
rect 19659 21641 19671 21675
rect 19613 21635 19671 21641
rect 9122 21536 9128 21548
rect 9083 21508 9128 21536
rect 9122 21496 9128 21508
rect 9180 21496 9186 21548
rect 11241 21539 11299 21545
rect 11241 21505 11253 21539
rect 11287 21536 11299 21539
rect 11514 21536 11520 21548
rect 11287 21508 11520 21536
rect 11287 21505 11299 21508
rect 11241 21499 11299 21505
rect 11514 21496 11520 21508
rect 11572 21496 11578 21548
rect 13035 21539 13093 21545
rect 13035 21505 13047 21539
rect 13081 21536 13093 21539
rect 13998 21536 14004 21548
rect 13081 21508 14004 21536
rect 13081 21505 13093 21508
rect 13035 21499 13093 21505
rect 13998 21496 14004 21508
rect 14056 21496 14062 21548
rect 14366 21536 14372 21548
rect 14327 21508 14372 21536
rect 14366 21496 14372 21508
rect 14424 21496 14430 21548
rect 16669 21539 16727 21545
rect 16669 21505 16681 21539
rect 16715 21536 16727 21539
rect 17126 21536 17132 21548
rect 16715 21508 17132 21536
rect 16715 21505 16727 21508
rect 16669 21499 16727 21505
rect 17126 21496 17132 21508
rect 17184 21536 17190 21548
rect 17497 21539 17555 21545
rect 17497 21536 17509 21539
rect 17184 21508 17509 21536
rect 17184 21496 17190 21508
rect 17497 21505 17509 21508
rect 17543 21505 17555 21539
rect 17497 21499 17555 21505
rect 17954 21496 17960 21548
rect 18012 21536 18018 21548
rect 18509 21539 18567 21545
rect 18509 21536 18521 21539
rect 18012 21508 18521 21536
rect 18012 21496 18018 21508
rect 18509 21505 18521 21508
rect 18555 21536 18567 21539
rect 18782 21536 18788 21548
rect 18555 21508 18788 21536
rect 18555 21505 18567 21508
rect 18509 21499 18567 21505
rect 18782 21496 18788 21508
rect 18840 21496 18846 21548
rect 18966 21496 18972 21548
rect 19024 21536 19030 21548
rect 19337 21539 19395 21545
rect 19337 21536 19349 21539
rect 19024 21508 19349 21536
rect 19024 21496 19030 21508
rect 19337 21505 19349 21508
rect 19383 21536 19395 21539
rect 19981 21539 20039 21545
rect 19981 21536 19993 21539
rect 19383 21508 19993 21536
rect 19383 21505 19395 21508
rect 19337 21499 19395 21505
rect 19981 21505 19993 21508
rect 20027 21505 20039 21539
rect 19981 21499 20039 21505
rect 8389 21471 8447 21477
rect 8389 21468 8401 21471
rect 8312 21440 8401 21468
rect 8312 21344 8340 21440
rect 8389 21437 8401 21440
rect 8435 21437 8447 21471
rect 8938 21468 8944 21480
rect 8899 21440 8944 21468
rect 8389 21431 8447 21437
rect 8938 21428 8944 21440
rect 8996 21428 9002 21480
rect 9674 21428 9680 21480
rect 9732 21468 9738 21480
rect 9953 21471 10011 21477
rect 9953 21468 9965 21471
rect 9732 21440 9965 21468
rect 9732 21428 9738 21440
rect 9953 21437 9965 21440
rect 9999 21437 10011 21471
rect 12894 21468 12900 21480
rect 12858 21440 12900 21468
rect 9953 21431 10011 21437
rect 12894 21428 12900 21440
rect 12952 21477 12958 21480
rect 12952 21471 13006 21477
rect 12952 21437 12960 21471
rect 12994 21468 13006 21471
rect 15746 21468 15752 21480
rect 12994 21440 13492 21468
rect 15707 21440 15752 21468
rect 12994 21437 13006 21440
rect 12952 21431 13006 21437
rect 12952 21428 12958 21431
rect 9861 21403 9919 21409
rect 9861 21369 9873 21403
rect 9907 21400 9919 21403
rect 10315 21403 10373 21409
rect 10315 21400 10327 21403
rect 9907 21372 10327 21400
rect 9907 21369 9919 21372
rect 9861 21363 9919 21369
rect 10315 21369 10327 21372
rect 10361 21400 10373 21403
rect 10870 21400 10876 21412
rect 10361 21372 10876 21400
rect 10361 21369 10373 21372
rect 10315 21363 10373 21369
rect 10870 21360 10876 21372
rect 10928 21360 10934 21412
rect 13464 21344 13492 21440
rect 15746 21428 15752 21440
rect 15804 21468 15810 21480
rect 15933 21471 15991 21477
rect 15933 21468 15945 21471
rect 15804 21440 15945 21468
rect 15804 21428 15810 21440
rect 15933 21437 15945 21440
rect 15979 21437 15991 21471
rect 16482 21468 16488 21480
rect 16443 21440 16488 21468
rect 15933 21431 15991 21437
rect 16482 21428 16488 21440
rect 16540 21428 16546 21480
rect 14090 21400 14096 21412
rect 14051 21372 14096 21400
rect 14090 21360 14096 21372
rect 14148 21360 14154 21412
rect 15105 21403 15163 21409
rect 15105 21369 15117 21403
rect 15151 21400 15163 21403
rect 16500 21400 16528 21428
rect 15151 21372 16528 21400
rect 18693 21403 18751 21409
rect 15151 21369 15163 21372
rect 15105 21363 15163 21369
rect 18693 21369 18705 21403
rect 18739 21369 18751 21403
rect 18693 21363 18751 21369
rect 8294 21332 8300 21344
rect 8255 21304 8300 21332
rect 8294 21292 8300 21304
rect 8352 21292 8358 21344
rect 13446 21332 13452 21344
rect 13407 21304 13452 21332
rect 13446 21292 13452 21304
rect 13504 21292 13510 21344
rect 15378 21332 15384 21344
rect 15339 21304 15384 21332
rect 15378 21292 15384 21304
rect 15436 21292 15442 21344
rect 16666 21292 16672 21344
rect 16724 21332 16730 21344
rect 17129 21335 17187 21341
rect 17129 21332 17141 21335
rect 16724 21304 17141 21332
rect 16724 21292 16730 21304
rect 17129 21301 17141 21304
rect 17175 21332 17187 21335
rect 17494 21332 17500 21344
rect 17175 21304 17500 21332
rect 17175 21301 17187 21304
rect 17129 21295 17187 21301
rect 17494 21292 17500 21304
rect 17552 21292 17558 21344
rect 18708 21332 18736 21363
rect 18782 21360 18788 21412
rect 18840 21400 18846 21412
rect 18840 21372 18885 21400
rect 18840 21360 18846 21372
rect 19334 21332 19340 21344
rect 18708 21304 19340 21332
rect 19334 21292 19340 21304
rect 19392 21292 19398 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 10962 21088 10968 21140
rect 11020 21128 11026 21140
rect 11333 21131 11391 21137
rect 11333 21128 11345 21131
rect 11020 21100 11345 21128
rect 11020 21088 11026 21100
rect 11333 21097 11345 21100
rect 11379 21128 11391 21131
rect 12986 21128 12992 21140
rect 11379 21100 12992 21128
rect 11379 21097 11391 21100
rect 11333 21091 11391 21097
rect 12986 21088 12992 21100
rect 13044 21088 13050 21140
rect 14090 21088 14096 21140
rect 14148 21128 14154 21140
rect 14369 21131 14427 21137
rect 14369 21128 14381 21131
rect 14148 21100 14381 21128
rect 14148 21088 14154 21100
rect 14369 21097 14381 21100
rect 14415 21097 14427 21131
rect 17218 21128 17224 21140
rect 14369 21091 14427 21097
rect 16500 21100 17224 21128
rect 10775 21063 10833 21069
rect 10775 21029 10787 21063
rect 10821 21060 10833 21063
rect 10870 21060 10876 21072
rect 10821 21032 10876 21060
rect 10821 21029 10833 21032
rect 10775 21023 10833 21029
rect 10870 21020 10876 21032
rect 10928 21020 10934 21072
rect 13078 21020 13084 21072
rect 13136 21060 13142 21072
rect 13494 21063 13552 21069
rect 13494 21060 13506 21063
rect 13136 21032 13506 21060
rect 13136 21020 13142 21032
rect 13494 21029 13506 21032
rect 13540 21060 13552 21063
rect 13630 21060 13636 21072
rect 13540 21032 13636 21060
rect 13540 21029 13552 21032
rect 13494 21023 13552 21029
rect 13630 21020 13636 21032
rect 13688 21020 13694 21072
rect 8294 20992 8300 21004
rect 8255 20964 8300 20992
rect 8294 20952 8300 20964
rect 8352 20952 8358 21004
rect 8570 20992 8576 21004
rect 8531 20964 8576 20992
rect 8570 20952 8576 20964
rect 8628 20952 8634 21004
rect 11882 20952 11888 21004
rect 11940 20992 11946 21004
rect 12196 20995 12254 21001
rect 12196 20992 12208 20995
rect 11940 20964 12208 20992
rect 11940 20952 11946 20964
rect 12196 20961 12208 20964
rect 12242 20961 12254 20995
rect 12196 20955 12254 20961
rect 13814 20952 13820 21004
rect 13872 20992 13878 21004
rect 14093 20995 14151 21001
rect 14093 20992 14105 20995
rect 13872 20964 14105 20992
rect 13872 20952 13878 20964
rect 14093 20961 14105 20964
rect 14139 20961 14151 20995
rect 14093 20955 14151 20961
rect 15540 20995 15598 21001
rect 15540 20961 15552 20995
rect 15586 20992 15598 20995
rect 16114 20992 16120 21004
rect 15586 20964 16120 20992
rect 15586 20961 15598 20964
rect 15540 20955 15598 20961
rect 16114 20952 16120 20964
rect 16172 20952 16178 21004
rect 16500 21001 16528 21100
rect 17218 21088 17224 21100
rect 17276 21128 17282 21140
rect 18325 21131 18383 21137
rect 18325 21128 18337 21131
rect 17276 21100 18337 21128
rect 17276 21088 17282 21100
rect 18325 21097 18337 21100
rect 18371 21097 18383 21131
rect 19334 21128 19340 21140
rect 19295 21100 19340 21128
rect 18325 21091 18383 21097
rect 19334 21088 19340 21100
rect 19392 21088 19398 21140
rect 16666 21020 16672 21072
rect 16724 21060 16730 21072
rect 16806 21063 16864 21069
rect 16806 21060 16818 21063
rect 16724 21032 16818 21060
rect 16724 21020 16730 21032
rect 16806 21029 16818 21032
rect 16852 21029 16864 21063
rect 18046 21060 18052 21072
rect 16806 21023 16864 21029
rect 17420 21032 18052 21060
rect 17420 21001 17448 21032
rect 18046 21020 18052 21032
rect 18104 21020 18110 21072
rect 16485 20995 16543 21001
rect 16485 20961 16497 20995
rect 16531 20961 16543 20995
rect 16485 20955 16543 20961
rect 17405 20995 17463 21001
rect 17405 20961 17417 20995
rect 17451 20961 17463 20995
rect 18506 20992 18512 21004
rect 18467 20964 18512 20992
rect 17405 20955 17463 20961
rect 18506 20952 18512 20964
rect 18564 20952 18570 21004
rect 18693 20995 18751 21001
rect 18693 20961 18705 20995
rect 18739 20961 18751 20995
rect 18693 20955 18751 20961
rect 8757 20927 8815 20933
rect 8757 20893 8769 20927
rect 8803 20924 8815 20927
rect 10413 20927 10471 20933
rect 10413 20924 10425 20927
rect 8803 20896 10425 20924
rect 8803 20893 8815 20896
rect 8757 20887 8815 20893
rect 10413 20893 10425 20896
rect 10459 20924 10471 20927
rect 11054 20924 11060 20936
rect 10459 20896 11060 20924
rect 10459 20893 10471 20896
rect 10413 20887 10471 20893
rect 11054 20884 11060 20896
rect 11112 20884 11118 20936
rect 13170 20924 13176 20936
rect 13131 20896 13176 20924
rect 13170 20884 13176 20896
rect 13228 20884 13234 20936
rect 16132 20924 16160 20952
rect 16574 20924 16580 20936
rect 16132 20896 16580 20924
rect 16574 20884 16580 20896
rect 16632 20884 16638 20936
rect 17770 20884 17776 20936
rect 17828 20924 17834 20936
rect 18708 20924 18736 20955
rect 17828 20896 18736 20924
rect 17828 20884 17834 20896
rect 9674 20748 9680 20800
rect 9732 20788 9738 20800
rect 9953 20791 10011 20797
rect 9953 20788 9965 20791
rect 9732 20760 9965 20788
rect 9732 20748 9738 20760
rect 9953 20757 9965 20760
rect 9999 20757 10011 20791
rect 9953 20751 10011 20757
rect 12299 20791 12357 20797
rect 12299 20757 12311 20791
rect 12345 20788 12357 20791
rect 12434 20788 12440 20800
rect 12345 20760 12440 20788
rect 12345 20757 12357 20760
rect 12299 20751 12357 20757
rect 12434 20748 12440 20760
rect 12492 20748 12498 20800
rect 15611 20791 15669 20797
rect 15611 20757 15623 20791
rect 15657 20788 15669 20791
rect 16022 20788 16028 20800
rect 15657 20760 16028 20788
rect 15657 20757 15669 20760
rect 15611 20751 15669 20757
rect 16022 20748 16028 20760
rect 16080 20748 16086 20800
rect 16301 20791 16359 20797
rect 16301 20757 16313 20791
rect 16347 20788 16359 20791
rect 16666 20788 16672 20800
rect 16347 20760 16672 20788
rect 16347 20757 16359 20760
rect 16301 20751 16359 20757
rect 16666 20748 16672 20760
rect 16724 20748 16730 20800
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 8481 20587 8539 20593
rect 8481 20553 8493 20587
rect 8527 20584 8539 20587
rect 8570 20584 8576 20596
rect 8527 20556 8576 20584
rect 8527 20553 8539 20556
rect 8481 20547 8539 20553
rect 8570 20544 8576 20556
rect 8628 20544 8634 20596
rect 10413 20587 10471 20593
rect 10413 20553 10425 20587
rect 10459 20584 10471 20587
rect 10870 20584 10876 20596
rect 10459 20556 10876 20584
rect 10459 20553 10471 20556
rect 10413 20547 10471 20553
rect 10870 20544 10876 20556
rect 10928 20544 10934 20596
rect 11054 20544 11060 20596
rect 11112 20584 11118 20596
rect 11517 20587 11575 20593
rect 11517 20584 11529 20587
rect 11112 20556 11529 20584
rect 11112 20544 11118 20556
rect 11517 20553 11529 20556
rect 11563 20553 11575 20587
rect 11517 20547 11575 20553
rect 11882 20544 11888 20596
rect 11940 20584 11946 20596
rect 12161 20587 12219 20593
rect 12161 20584 12173 20587
rect 11940 20556 12173 20584
rect 11940 20544 11946 20556
rect 12161 20553 12173 20556
rect 12207 20584 12219 20587
rect 12342 20584 12348 20596
rect 12207 20556 12348 20584
rect 12207 20553 12219 20556
rect 12161 20547 12219 20553
rect 12342 20544 12348 20556
rect 12400 20544 12406 20596
rect 14090 20544 14096 20596
rect 14148 20584 14154 20596
rect 14277 20587 14335 20593
rect 14277 20584 14289 20587
rect 14148 20556 14289 20584
rect 14148 20544 14154 20556
rect 14277 20553 14289 20556
rect 14323 20553 14335 20587
rect 14277 20547 14335 20553
rect 18506 20544 18512 20596
rect 18564 20584 18570 20596
rect 19061 20587 19119 20593
rect 19061 20584 19073 20587
rect 18564 20556 19073 20584
rect 18564 20544 18570 20556
rect 19061 20553 19073 20556
rect 19107 20553 19119 20587
rect 19061 20547 19119 20553
rect 9585 20451 9643 20457
rect 9585 20417 9597 20451
rect 9631 20448 9643 20451
rect 9674 20448 9680 20460
rect 9631 20420 9680 20448
rect 9631 20417 9643 20420
rect 9585 20411 9643 20417
rect 9674 20408 9680 20420
rect 9732 20408 9738 20460
rect 11054 20448 11060 20460
rect 11015 20420 11060 20448
rect 11054 20408 11060 20420
rect 11112 20408 11118 20460
rect 16206 20448 16212 20460
rect 16167 20420 16212 20448
rect 16206 20408 16212 20420
rect 16264 20408 16270 20460
rect 16574 20408 16580 20460
rect 16632 20448 16638 20460
rect 17770 20448 17776 20460
rect 16632 20420 17776 20448
rect 16632 20408 16638 20420
rect 17770 20408 17776 20420
rect 17828 20408 17834 20460
rect 8941 20383 8999 20389
rect 8941 20380 8953 20383
rect 8772 20352 8953 20380
rect 8772 20256 8800 20352
rect 8941 20349 8953 20352
rect 8987 20349 8999 20383
rect 8941 20343 8999 20349
rect 9122 20340 9128 20392
rect 9180 20380 9186 20392
rect 9401 20383 9459 20389
rect 9401 20380 9413 20383
rect 9180 20352 9413 20380
rect 9180 20340 9186 20352
rect 9401 20349 9413 20352
rect 9447 20349 9459 20383
rect 9401 20343 9459 20349
rect 12802 20340 12808 20392
rect 12860 20380 12866 20392
rect 13357 20383 13415 20389
rect 13357 20380 13369 20383
rect 12860 20352 13369 20380
rect 12860 20340 12866 20352
rect 13357 20349 13369 20352
rect 13403 20380 13415 20383
rect 14553 20383 14611 20389
rect 14553 20380 14565 20383
rect 13403 20352 14565 20380
rect 13403 20349 13415 20352
rect 13357 20343 13415 20349
rect 14553 20349 14565 20352
rect 14599 20349 14611 20383
rect 14553 20343 14611 20349
rect 15194 20340 15200 20392
rect 15252 20389 15258 20392
rect 15252 20383 15290 20389
rect 15278 20380 15290 20383
rect 15657 20383 15715 20389
rect 15657 20380 15669 20383
rect 15278 20352 15669 20380
rect 15278 20349 15290 20352
rect 15252 20343 15290 20349
rect 15657 20349 15669 20352
rect 15703 20349 15715 20383
rect 15657 20343 15715 20349
rect 17129 20383 17187 20389
rect 17129 20349 17141 20383
rect 17175 20380 17187 20383
rect 17862 20380 17868 20392
rect 17175 20352 17868 20380
rect 17175 20349 17187 20352
rect 17129 20343 17187 20349
rect 15252 20340 15258 20343
rect 17862 20340 17868 20352
rect 17920 20340 17926 20392
rect 19610 20340 19616 20392
rect 19668 20389 19674 20392
rect 19668 20383 19706 20389
rect 19694 20380 19706 20383
rect 20073 20383 20131 20389
rect 20073 20380 20085 20383
rect 19694 20352 20085 20380
rect 19694 20349 19706 20352
rect 19668 20343 19706 20349
rect 20073 20349 20085 20352
rect 20119 20380 20131 20383
rect 20162 20380 20168 20392
rect 20119 20352 20168 20380
rect 20119 20349 20131 20352
rect 20073 20343 20131 20349
rect 19668 20340 19674 20343
rect 20162 20340 20168 20352
rect 20220 20340 20226 20392
rect 10134 20272 10140 20324
rect 10192 20312 10198 20324
rect 10597 20315 10655 20321
rect 10597 20312 10609 20315
rect 10192 20284 10609 20312
rect 10192 20272 10198 20284
rect 10597 20281 10609 20284
rect 10643 20281 10655 20315
rect 10597 20275 10655 20281
rect 10689 20315 10747 20321
rect 10689 20281 10701 20315
rect 10735 20312 10747 20315
rect 10962 20312 10968 20324
rect 10735 20284 10968 20312
rect 10735 20281 10747 20284
rect 10689 20275 10747 20281
rect 8113 20247 8171 20253
rect 8113 20213 8125 20247
rect 8159 20244 8171 20247
rect 8294 20244 8300 20256
rect 8159 20216 8300 20244
rect 8159 20213 8171 20216
rect 8113 20207 8171 20213
rect 8294 20204 8300 20216
rect 8352 20244 8358 20256
rect 8754 20244 8760 20256
rect 8352 20216 8760 20244
rect 8352 20204 8358 20216
rect 8754 20204 8760 20216
rect 8812 20204 8818 20256
rect 10042 20244 10048 20256
rect 9955 20216 10048 20244
rect 10042 20204 10048 20216
rect 10100 20244 10106 20256
rect 10704 20244 10732 20275
rect 10962 20272 10968 20284
rect 11020 20272 11026 20324
rect 13678 20315 13736 20321
rect 13678 20312 13690 20315
rect 13188 20284 13690 20312
rect 10100 20216 10732 20244
rect 12897 20247 12955 20253
rect 10100 20204 10106 20216
rect 12897 20213 12909 20247
rect 12943 20244 12955 20247
rect 13078 20244 13084 20256
rect 12943 20216 13084 20244
rect 12943 20213 12955 20216
rect 12897 20207 12955 20213
rect 13078 20204 13084 20216
rect 13136 20244 13142 20256
rect 13188 20253 13216 20284
rect 13678 20281 13690 20284
rect 13724 20281 13736 20315
rect 13678 20275 13736 20281
rect 16571 20315 16629 20321
rect 16571 20281 16583 20315
rect 16617 20312 16629 20315
rect 16666 20312 16672 20324
rect 16617 20284 16672 20312
rect 16617 20281 16629 20284
rect 16571 20275 16629 20281
rect 16666 20272 16672 20284
rect 16724 20312 16730 20324
rect 18138 20312 18144 20324
rect 16724 20284 17080 20312
rect 18099 20284 18144 20312
rect 16724 20272 16730 20284
rect 17052 20256 17080 20284
rect 18138 20272 18144 20284
rect 18196 20272 18202 20324
rect 18233 20315 18291 20321
rect 18233 20281 18245 20315
rect 18279 20281 18291 20315
rect 18233 20275 18291 20281
rect 18785 20315 18843 20321
rect 18785 20281 18797 20315
rect 18831 20312 18843 20315
rect 18966 20312 18972 20324
rect 18831 20284 18972 20312
rect 18831 20281 18843 20284
rect 18785 20275 18843 20281
rect 13173 20247 13231 20253
rect 13173 20244 13185 20247
rect 13136 20216 13185 20244
rect 13136 20204 13142 20216
rect 13173 20213 13185 20216
rect 13219 20213 13231 20247
rect 13173 20207 13231 20213
rect 15335 20247 15393 20253
rect 15335 20213 15347 20247
rect 15381 20244 15393 20247
rect 15562 20244 15568 20256
rect 15381 20216 15568 20244
rect 15381 20213 15393 20216
rect 15335 20207 15393 20213
rect 15562 20204 15568 20216
rect 15620 20204 15626 20256
rect 16114 20244 16120 20256
rect 16075 20216 16120 20244
rect 16114 20204 16120 20216
rect 16172 20204 16178 20256
rect 17034 20204 17040 20256
rect 17092 20244 17098 20256
rect 17405 20247 17463 20253
rect 17405 20244 17417 20247
rect 17092 20216 17417 20244
rect 17092 20204 17098 20216
rect 17405 20213 17417 20216
rect 17451 20213 17463 20247
rect 17405 20207 17463 20213
rect 18046 20204 18052 20256
rect 18104 20244 18110 20256
rect 18248 20244 18276 20275
rect 18966 20272 18972 20284
rect 19024 20272 19030 20324
rect 18104 20216 18276 20244
rect 18104 20204 18110 20216
rect 19334 20204 19340 20256
rect 19392 20244 19398 20256
rect 19751 20247 19809 20253
rect 19751 20244 19763 20247
rect 19392 20216 19763 20244
rect 19392 20204 19398 20216
rect 19751 20213 19763 20216
rect 19797 20213 19809 20247
rect 19751 20207 19809 20213
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 13170 20040 13176 20052
rect 13131 20012 13176 20040
rect 13170 20000 13176 20012
rect 13228 20000 13234 20052
rect 16025 20043 16083 20049
rect 16025 20009 16037 20043
rect 16071 20040 16083 20043
rect 16206 20040 16212 20052
rect 16071 20012 16212 20040
rect 16071 20009 16083 20012
rect 16025 20003 16083 20009
rect 16206 20000 16212 20012
rect 16264 20000 16270 20052
rect 17218 20040 17224 20052
rect 17179 20012 17224 20040
rect 17218 20000 17224 20012
rect 17276 20000 17282 20052
rect 18046 20000 18052 20052
rect 18104 20040 18110 20052
rect 19150 20040 19156 20052
rect 18104 20012 19156 20040
rect 18104 20000 18110 20012
rect 19150 20000 19156 20012
rect 19208 20040 19214 20052
rect 19208 20012 19472 20040
rect 19208 20000 19214 20012
rect 10597 19975 10655 19981
rect 10597 19941 10609 19975
rect 10643 19972 10655 19975
rect 10962 19972 10968 19984
rect 10643 19944 10968 19972
rect 10643 19941 10655 19944
rect 10597 19935 10655 19941
rect 10962 19932 10968 19944
rect 11020 19932 11026 19984
rect 12802 19972 12808 19984
rect 12763 19944 12808 19972
rect 12802 19932 12808 19944
rect 12860 19932 12866 19984
rect 13814 19972 13820 19984
rect 13775 19944 13820 19972
rect 13814 19932 13820 19944
rect 13872 19932 13878 19984
rect 16298 19972 16304 19984
rect 16259 19944 16304 19972
rect 16298 19932 16304 19944
rect 16356 19932 16362 19984
rect 17589 19975 17647 19981
rect 17589 19941 17601 19975
rect 17635 19972 17647 19975
rect 17770 19972 17776 19984
rect 17635 19944 17776 19972
rect 17635 19941 17647 19944
rect 17589 19935 17647 19941
rect 17770 19932 17776 19944
rect 17828 19932 17834 19984
rect 17862 19932 17868 19984
rect 17920 19972 17926 19984
rect 19334 19972 19340 19984
rect 17920 19944 17965 19972
rect 19295 19944 19340 19972
rect 17920 19932 17926 19944
rect 19334 19932 19340 19944
rect 19392 19932 19398 19984
rect 19444 19981 19472 20012
rect 19429 19975 19487 19981
rect 19429 19941 19441 19975
rect 19475 19941 19487 19975
rect 19429 19935 19487 19941
rect 8570 19864 8576 19916
rect 8628 19913 8634 19916
rect 8628 19907 8666 19913
rect 8654 19873 8666 19907
rect 8628 19867 8666 19873
rect 8628 19864 8634 19867
rect 11974 19864 11980 19916
rect 12032 19904 12038 19916
rect 12069 19907 12127 19913
rect 12069 19904 12081 19907
rect 12032 19876 12081 19904
rect 12032 19864 12038 19876
rect 12069 19873 12081 19876
rect 12115 19873 12127 19907
rect 12618 19904 12624 19916
rect 12579 19876 12624 19904
rect 12069 19867 12127 19873
rect 12618 19864 12624 19876
rect 12676 19864 12682 19916
rect 7561 19839 7619 19845
rect 7561 19805 7573 19839
rect 7607 19836 7619 19839
rect 8202 19836 8208 19848
rect 7607 19808 8208 19836
rect 7607 19805 7619 19808
rect 7561 19799 7619 19805
rect 8202 19796 8208 19808
rect 8260 19796 8266 19848
rect 9122 19836 9128 19848
rect 9083 19808 9128 19836
rect 9122 19796 9128 19808
rect 9180 19796 9186 19848
rect 10505 19839 10563 19845
rect 10505 19805 10517 19839
rect 10551 19805 10563 19839
rect 10505 19799 10563 19805
rect 11149 19839 11207 19845
rect 11149 19805 11161 19839
rect 11195 19836 11207 19839
rect 11330 19836 11336 19848
rect 11195 19808 11336 19836
rect 11195 19805 11207 19808
rect 11149 19799 11207 19805
rect 8711 19771 8769 19777
rect 8711 19737 8723 19771
rect 8757 19768 8769 19771
rect 9861 19771 9919 19777
rect 9861 19768 9873 19771
rect 8757 19740 9873 19768
rect 8757 19737 8769 19740
rect 8711 19731 8769 19737
rect 9861 19737 9873 19740
rect 9907 19768 9919 19771
rect 10520 19768 10548 19799
rect 11330 19796 11336 19808
rect 11388 19796 11394 19848
rect 12434 19796 12440 19848
rect 12492 19836 12498 19848
rect 13262 19836 13268 19848
rect 12492 19808 13268 19836
rect 12492 19796 12498 19808
rect 13262 19796 13268 19808
rect 13320 19836 13326 19848
rect 13725 19839 13783 19845
rect 13725 19836 13737 19839
rect 13320 19808 13737 19836
rect 13320 19796 13326 19808
rect 13725 19805 13737 19808
rect 13771 19805 13783 19839
rect 13725 19799 13783 19805
rect 16022 19796 16028 19848
rect 16080 19836 16086 19848
rect 16209 19839 16267 19845
rect 16209 19836 16221 19839
rect 16080 19808 16221 19836
rect 16080 19796 16086 19808
rect 16209 19805 16221 19808
rect 16255 19836 16267 19839
rect 16574 19836 16580 19848
rect 16255 19808 16580 19836
rect 16255 19805 16267 19808
rect 16209 19799 16267 19805
rect 16574 19796 16580 19808
rect 16632 19796 16638 19848
rect 18417 19839 18475 19845
rect 18417 19805 18429 19839
rect 18463 19836 18475 19839
rect 18966 19836 18972 19848
rect 18463 19808 18972 19836
rect 18463 19805 18475 19808
rect 18417 19799 18475 19805
rect 18966 19796 18972 19808
rect 19024 19796 19030 19848
rect 19613 19839 19671 19845
rect 19613 19805 19625 19839
rect 19659 19805 19671 19839
rect 19613 19799 19671 19805
rect 9907 19740 10548 19768
rect 14277 19771 14335 19777
rect 9907 19737 9919 19740
rect 9861 19731 9919 19737
rect 14277 19737 14289 19771
rect 14323 19737 14335 19771
rect 14277 19731 14335 19737
rect 16761 19771 16819 19777
rect 16761 19737 16773 19771
rect 16807 19768 16819 19771
rect 18230 19768 18236 19780
rect 16807 19740 18236 19768
rect 16807 19737 16819 19740
rect 16761 19731 16819 19737
rect 9398 19700 9404 19712
rect 9359 19672 9404 19700
rect 9398 19660 9404 19672
rect 9456 19660 9462 19712
rect 10226 19700 10232 19712
rect 10187 19672 10232 19700
rect 10226 19660 10232 19672
rect 10284 19660 10290 19712
rect 14292 19700 14320 19731
rect 18230 19728 18236 19740
rect 18288 19768 18294 19780
rect 19628 19768 19656 19799
rect 18288 19740 19656 19768
rect 18288 19728 18294 19740
rect 14366 19700 14372 19712
rect 14279 19672 14372 19700
rect 14366 19660 14372 19672
rect 14424 19700 14430 19712
rect 14737 19703 14795 19709
rect 14737 19700 14749 19703
rect 14424 19672 14749 19700
rect 14424 19660 14430 19672
rect 14737 19669 14749 19672
rect 14783 19700 14795 19703
rect 16206 19700 16212 19712
rect 14783 19672 16212 19700
rect 14783 19669 14795 19672
rect 14737 19663 14795 19669
rect 16206 19660 16212 19672
rect 16264 19660 16270 19712
rect 18138 19660 18144 19712
rect 18196 19700 18202 19712
rect 18785 19703 18843 19709
rect 18785 19700 18797 19703
rect 18196 19672 18797 19700
rect 18196 19660 18202 19672
rect 18785 19669 18797 19672
rect 18831 19700 18843 19703
rect 19242 19700 19248 19712
rect 18831 19672 19248 19700
rect 18831 19669 18843 19672
rect 18785 19663 18843 19669
rect 19242 19660 19248 19672
rect 19300 19660 19306 19712
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 8110 19456 8116 19508
rect 8168 19505 8174 19508
rect 8168 19499 8217 19505
rect 8168 19465 8171 19499
rect 8205 19465 8217 19499
rect 10042 19496 10048 19508
rect 10003 19468 10048 19496
rect 8168 19459 8217 19465
rect 8168 19456 8174 19459
rect 10042 19456 10048 19468
rect 10100 19456 10106 19508
rect 13814 19456 13820 19508
rect 13872 19496 13878 19508
rect 14001 19499 14059 19505
rect 14001 19496 14013 19499
rect 13872 19468 14013 19496
rect 13872 19456 13878 19468
rect 14001 19465 14013 19468
rect 14047 19465 14059 19499
rect 14001 19459 14059 19465
rect 16298 19456 16304 19508
rect 16356 19496 16362 19508
rect 16945 19499 17003 19505
rect 16945 19496 16957 19499
rect 16356 19468 16957 19496
rect 16356 19456 16362 19468
rect 16945 19465 16957 19468
rect 16991 19496 17003 19499
rect 17497 19499 17555 19505
rect 17497 19496 17509 19499
rect 16991 19468 17509 19496
rect 16991 19465 17003 19468
rect 16945 19459 17003 19465
rect 17497 19465 17509 19468
rect 17543 19496 17555 19499
rect 17862 19496 17868 19508
rect 17543 19468 17868 19496
rect 17543 19465 17555 19468
rect 17497 19459 17555 19465
rect 17862 19456 17868 19468
rect 17920 19456 17926 19508
rect 19150 19456 19156 19508
rect 19208 19496 19214 19508
rect 19245 19499 19303 19505
rect 19245 19496 19257 19499
rect 19208 19468 19257 19496
rect 19208 19456 19214 19468
rect 19245 19465 19257 19468
rect 19291 19465 19303 19499
rect 19610 19496 19616 19508
rect 19571 19468 19616 19496
rect 19245 19459 19303 19465
rect 19610 19456 19616 19468
rect 19668 19456 19674 19508
rect 6638 19388 6644 19440
rect 6696 19428 6702 19440
rect 9214 19428 9220 19440
rect 6696 19400 9220 19428
rect 6696 19388 6702 19400
rect 9214 19388 9220 19400
rect 9272 19388 9278 19440
rect 7742 19320 7748 19372
rect 7800 19360 7806 19372
rect 7834 19360 7840 19372
rect 7800 19332 7840 19360
rect 7800 19320 7806 19332
rect 7834 19320 7840 19332
rect 7892 19320 7898 19372
rect 8570 19360 8576 19372
rect 8531 19332 8576 19360
rect 8570 19320 8576 19332
rect 8628 19320 8634 19372
rect 9125 19363 9183 19369
rect 9125 19329 9137 19363
rect 9171 19360 9183 19363
rect 9398 19360 9404 19372
rect 9171 19332 9404 19360
rect 9171 19329 9183 19332
rect 9125 19323 9183 19329
rect 9398 19320 9404 19332
rect 9456 19320 9462 19372
rect 12250 19320 12256 19372
rect 12308 19360 12314 19372
rect 12526 19360 12532 19372
rect 12308 19332 12532 19360
rect 12308 19320 12314 19332
rect 12526 19320 12532 19332
rect 12584 19320 12590 19372
rect 13170 19360 13176 19372
rect 13131 19332 13176 19360
rect 13170 19320 13176 19332
rect 13228 19320 13234 19372
rect 14366 19360 14372 19372
rect 14327 19332 14372 19360
rect 14366 19320 14372 19332
rect 14424 19320 14430 19372
rect 14826 19360 14832 19372
rect 14787 19332 14832 19360
rect 14826 19320 14832 19332
rect 14884 19320 14890 19372
rect 16206 19360 16212 19372
rect 16167 19332 16212 19360
rect 16206 19320 16212 19332
rect 16264 19320 16270 19372
rect 7926 19292 7932 19304
rect 7887 19264 7932 19292
rect 7926 19252 7932 19264
rect 7984 19292 7990 19304
rect 8056 19295 8114 19301
rect 8056 19292 8068 19295
rect 7984 19264 8068 19292
rect 7984 19252 7990 19264
rect 8056 19261 8068 19264
rect 8102 19292 8114 19295
rect 8938 19292 8944 19304
rect 8102 19264 8944 19292
rect 8102 19261 8114 19264
rect 8056 19255 8114 19261
rect 8938 19252 8944 19264
rect 8996 19252 9002 19304
rect 10410 19292 10416 19304
rect 10371 19264 10416 19292
rect 10410 19252 10416 19264
rect 10468 19252 10474 19304
rect 12710 19292 12716 19304
rect 12671 19264 12716 19292
rect 12710 19252 12716 19264
rect 12768 19292 12774 19304
rect 12894 19292 12900 19304
rect 12768 19264 12900 19292
rect 12768 19252 12774 19264
rect 12894 19252 12900 19264
rect 12952 19252 12958 19304
rect 13081 19295 13139 19301
rect 13081 19261 13093 19295
rect 13127 19292 13139 19295
rect 13633 19295 13691 19301
rect 13633 19292 13645 19295
rect 13127 19264 13645 19292
rect 13127 19261 13139 19264
rect 13081 19255 13139 19261
rect 13633 19261 13645 19264
rect 13679 19261 13691 19295
rect 13633 19255 13691 19261
rect 19848 19295 19906 19301
rect 19848 19261 19860 19295
rect 19894 19292 19906 19295
rect 20254 19292 20260 19304
rect 19894 19264 20260 19292
rect 19894 19261 19906 19264
rect 19848 19255 19906 19261
rect 9217 19227 9275 19233
rect 9217 19193 9229 19227
rect 9263 19193 9275 19227
rect 9217 19187 9275 19193
rect 9769 19227 9827 19233
rect 9769 19193 9781 19227
rect 9815 19224 9827 19227
rect 10428 19224 10456 19252
rect 10689 19227 10747 19233
rect 10689 19224 10701 19227
rect 9815 19196 10364 19224
rect 10428 19196 10701 19224
rect 9815 19193 9827 19196
rect 9769 19187 9827 19193
rect 9232 19156 9260 19187
rect 9858 19156 9864 19168
rect 9232 19128 9864 19156
rect 9858 19116 9864 19128
rect 9916 19116 9922 19168
rect 10336 19156 10364 19196
rect 10689 19193 10701 19196
rect 10735 19193 10747 19227
rect 10689 19187 10747 19193
rect 10781 19227 10839 19233
rect 10781 19193 10793 19227
rect 10827 19224 10839 19227
rect 11146 19224 11152 19236
rect 10827 19196 11152 19224
rect 10827 19193 10839 19196
rect 10781 19187 10839 19193
rect 11146 19184 11152 19196
rect 11204 19184 11210 19236
rect 11330 19224 11336 19236
rect 11291 19196 11336 19224
rect 11330 19184 11336 19196
rect 11388 19184 11394 19236
rect 11793 19227 11851 19233
rect 11793 19193 11805 19227
rect 11839 19224 11851 19227
rect 12158 19224 12164 19236
rect 11839 19196 12164 19224
rect 11839 19193 11851 19196
rect 11793 19187 11851 19193
rect 12158 19184 12164 19196
rect 12216 19224 12222 19236
rect 12526 19224 12532 19236
rect 12216 19196 12532 19224
rect 12216 19184 12222 19196
rect 12526 19184 12532 19196
rect 12584 19224 12590 19236
rect 13096 19224 13124 19255
rect 20254 19252 20260 19264
rect 20312 19252 20318 19304
rect 20806 19292 20812 19304
rect 20767 19264 20812 19292
rect 20806 19252 20812 19264
rect 20864 19252 20870 19304
rect 12584 19196 13124 19224
rect 12584 19184 12590 19196
rect 14458 19184 14464 19236
rect 14516 19224 14522 19236
rect 15749 19227 15807 19233
rect 14516 19196 14561 19224
rect 14516 19184 14522 19196
rect 15749 19193 15761 19227
rect 15795 19224 15807 19227
rect 15930 19224 15936 19236
rect 15795 19196 15936 19224
rect 15795 19193 15807 19196
rect 15749 19187 15807 19193
rect 15930 19184 15936 19196
rect 15988 19184 15994 19236
rect 16025 19227 16083 19233
rect 16025 19193 16037 19227
rect 16071 19193 16083 19227
rect 16025 19187 16083 19193
rect 17865 19227 17923 19233
rect 17865 19193 17877 19227
rect 17911 19224 17923 19227
rect 18322 19224 18328 19236
rect 17911 19196 18328 19224
rect 17911 19193 17923 19196
rect 17865 19187 17923 19193
rect 11054 19156 11060 19168
rect 10336 19128 11060 19156
rect 11054 19116 11060 19128
rect 11112 19116 11118 19168
rect 11974 19116 11980 19168
rect 12032 19156 12038 19168
rect 12069 19159 12127 19165
rect 12069 19156 12081 19159
rect 12032 19128 12081 19156
rect 12032 19116 12038 19128
rect 12069 19125 12081 19128
rect 12115 19125 12127 19159
rect 12069 19119 12127 19125
rect 15381 19159 15439 19165
rect 15381 19125 15393 19159
rect 15427 19156 15439 19159
rect 15838 19156 15844 19168
rect 15427 19128 15844 19156
rect 15427 19125 15439 19128
rect 15381 19119 15439 19125
rect 15838 19116 15844 19128
rect 15896 19156 15902 19168
rect 16040 19156 16068 19187
rect 18322 19184 18328 19196
rect 18380 19184 18386 19236
rect 18414 19184 18420 19236
rect 18472 19224 18478 19236
rect 18690 19224 18696 19236
rect 18472 19196 18696 19224
rect 18472 19184 18478 19196
rect 18690 19184 18696 19196
rect 18748 19184 18754 19236
rect 18966 19224 18972 19236
rect 18927 19196 18972 19224
rect 18966 19184 18972 19196
rect 19024 19184 19030 19236
rect 19334 19184 19340 19236
rect 19392 19224 19398 19236
rect 19935 19227 19993 19233
rect 19935 19224 19947 19227
rect 19392 19196 19947 19224
rect 19392 19184 19398 19196
rect 19935 19193 19947 19196
rect 19981 19193 19993 19227
rect 19935 19187 19993 19193
rect 15896 19128 16068 19156
rect 15896 19116 15902 19128
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 8711 18955 8769 18961
rect 8711 18921 8723 18955
rect 8757 18952 8769 18955
rect 9398 18952 9404 18964
rect 8757 18924 9404 18952
rect 8757 18921 8769 18924
rect 8711 18915 8769 18921
rect 9398 18912 9404 18924
rect 9456 18912 9462 18964
rect 11146 18952 11152 18964
rect 11107 18924 11152 18952
rect 11146 18912 11152 18924
rect 11204 18912 11210 18964
rect 13262 18952 13268 18964
rect 13223 18924 13268 18952
rect 13262 18912 13268 18924
rect 13320 18912 13326 18964
rect 14369 18955 14427 18961
rect 14369 18921 14381 18955
rect 14415 18952 14427 18955
rect 14458 18952 14464 18964
rect 14415 18924 14464 18952
rect 14415 18921 14427 18924
rect 14369 18915 14427 18921
rect 14458 18912 14464 18924
rect 14516 18952 14522 18964
rect 14645 18955 14703 18961
rect 14645 18952 14657 18955
rect 14516 18924 14657 18952
rect 14516 18912 14522 18924
rect 14645 18921 14657 18924
rect 14691 18921 14703 18955
rect 14645 18915 14703 18921
rect 15838 18912 15844 18964
rect 15896 18952 15902 18964
rect 16022 18952 16028 18964
rect 15896 18924 16028 18952
rect 15896 18912 15902 18924
rect 16022 18912 16028 18924
rect 16080 18952 16086 18964
rect 16393 18955 16451 18961
rect 16393 18952 16405 18955
rect 16080 18924 16405 18952
rect 16080 18912 16086 18924
rect 16393 18921 16405 18924
rect 16439 18921 16451 18955
rect 16393 18915 16451 18921
rect 16574 18912 16580 18964
rect 16632 18952 16638 18964
rect 16761 18955 16819 18961
rect 16761 18952 16773 18955
rect 16632 18924 16773 18952
rect 16632 18912 16638 18924
rect 16761 18921 16773 18924
rect 16807 18921 16819 18955
rect 16761 18915 16819 18921
rect 17865 18955 17923 18961
rect 17865 18921 17877 18955
rect 17911 18952 17923 18955
rect 17911 18924 18920 18952
rect 17911 18921 17923 18924
rect 17865 18915 17923 18921
rect 9493 18887 9551 18893
rect 9493 18853 9505 18887
rect 9539 18884 9551 18887
rect 9858 18884 9864 18896
rect 9539 18856 9864 18884
rect 9539 18853 9551 18856
rect 9493 18847 9551 18853
rect 9858 18844 9864 18856
rect 9916 18884 9922 18896
rect 10321 18887 10379 18893
rect 10321 18884 10333 18887
rect 9916 18856 10333 18884
rect 9916 18844 9922 18856
rect 10321 18853 10333 18856
rect 10367 18853 10379 18887
rect 11882 18884 11888 18896
rect 11843 18856 11888 18884
rect 10321 18847 10379 18853
rect 11882 18844 11888 18856
rect 11940 18844 11946 18896
rect 13078 18844 13084 18896
rect 13136 18884 13142 18896
rect 13770 18887 13828 18893
rect 13770 18884 13782 18887
rect 13136 18856 13782 18884
rect 13136 18844 13142 18856
rect 13770 18853 13782 18856
rect 13816 18853 13828 18887
rect 13770 18847 13828 18853
rect 16850 18844 16856 18896
rect 16908 18884 16914 18896
rect 17034 18884 17040 18896
rect 16908 18856 17040 18884
rect 16908 18844 16914 18856
rect 17034 18844 17040 18856
rect 17092 18884 17098 18896
rect 17266 18887 17324 18893
rect 17266 18884 17278 18887
rect 17092 18856 17278 18884
rect 17092 18844 17098 18856
rect 17266 18853 17278 18856
rect 17312 18853 17324 18887
rect 17266 18847 17324 18853
rect 18325 18887 18383 18893
rect 18325 18853 18337 18887
rect 18371 18884 18383 18887
rect 18414 18884 18420 18896
rect 18371 18856 18420 18884
rect 18371 18853 18383 18856
rect 18325 18847 18383 18853
rect 18414 18844 18420 18856
rect 18472 18844 18478 18896
rect 18892 18893 18920 18924
rect 18877 18887 18935 18893
rect 18877 18853 18889 18887
rect 18923 18884 18935 18887
rect 19058 18884 19064 18896
rect 18923 18856 19064 18884
rect 18923 18853 18935 18856
rect 18877 18847 18935 18853
rect 19058 18844 19064 18856
rect 19116 18844 19122 18896
rect 7628 18819 7686 18825
rect 7628 18785 7640 18819
rect 7674 18816 7686 18819
rect 7742 18816 7748 18828
rect 7674 18788 7748 18816
rect 7674 18785 7686 18788
rect 7628 18779 7686 18785
rect 7742 18776 7748 18788
rect 7800 18776 7806 18828
rect 8478 18776 8484 18828
rect 8536 18816 8542 18828
rect 8608 18819 8666 18825
rect 8608 18816 8620 18819
rect 8536 18788 8620 18816
rect 8536 18776 8542 18788
rect 8608 18785 8620 18788
rect 8654 18816 8666 18819
rect 9950 18816 9956 18828
rect 8654 18788 9956 18816
rect 8654 18785 8666 18788
rect 8608 18779 8666 18785
rect 9950 18776 9956 18788
rect 10008 18776 10014 18828
rect 15378 18816 15384 18828
rect 15339 18788 15384 18816
rect 15378 18776 15384 18788
rect 15436 18776 15442 18828
rect 15933 18819 15991 18825
rect 15933 18785 15945 18819
rect 15979 18816 15991 18819
rect 16206 18816 16212 18828
rect 15979 18788 16212 18816
rect 15979 18785 15991 18788
rect 15933 18779 15991 18785
rect 16206 18776 16212 18788
rect 16264 18816 16270 18828
rect 16482 18816 16488 18828
rect 16264 18788 16488 18816
rect 16264 18776 16270 18788
rect 16482 18776 16488 18788
rect 16540 18776 16546 18828
rect 10042 18708 10048 18760
rect 10100 18748 10106 18760
rect 10229 18751 10287 18757
rect 10229 18748 10241 18751
rect 10100 18720 10241 18748
rect 10100 18708 10106 18720
rect 10229 18717 10241 18720
rect 10275 18717 10287 18751
rect 10229 18711 10287 18717
rect 10873 18751 10931 18757
rect 10873 18717 10885 18751
rect 10919 18748 10931 18751
rect 11330 18748 11336 18760
rect 10919 18720 11336 18748
rect 10919 18717 10931 18720
rect 10873 18711 10931 18717
rect 11330 18708 11336 18720
rect 11388 18748 11394 18760
rect 11790 18748 11796 18760
rect 11388 18720 11796 18748
rect 11388 18708 11394 18720
rect 11790 18708 11796 18720
rect 11848 18708 11854 18760
rect 12066 18748 12072 18760
rect 12027 18720 12072 18748
rect 12066 18708 12072 18720
rect 12124 18708 12130 18760
rect 13446 18748 13452 18760
rect 13407 18720 13452 18748
rect 13446 18708 13452 18720
rect 13504 18708 13510 18760
rect 16117 18751 16175 18757
rect 16117 18717 16129 18751
rect 16163 18748 16175 18751
rect 16945 18751 17003 18757
rect 16945 18748 16957 18751
rect 16163 18720 16957 18748
rect 16163 18717 16175 18720
rect 16117 18711 16175 18717
rect 16945 18717 16957 18720
rect 16991 18748 17003 18751
rect 17310 18748 17316 18760
rect 16991 18720 17316 18748
rect 16991 18717 17003 18720
rect 16945 18711 17003 18717
rect 17310 18708 17316 18720
rect 17368 18708 17374 18760
rect 18785 18751 18843 18757
rect 18785 18717 18797 18751
rect 18831 18748 18843 18751
rect 18966 18748 18972 18760
rect 18831 18720 18972 18748
rect 18831 18717 18843 18720
rect 18785 18711 18843 18717
rect 18966 18708 18972 18720
rect 19024 18748 19030 18760
rect 19426 18748 19432 18760
rect 19024 18720 19432 18748
rect 19024 18708 19030 18720
rect 19426 18708 19432 18720
rect 19484 18708 19490 18760
rect 19334 18680 19340 18692
rect 19295 18652 19340 18680
rect 19334 18640 19340 18652
rect 19392 18640 19398 18692
rect 7699 18615 7757 18621
rect 7699 18581 7711 18615
rect 7745 18612 7757 18615
rect 8662 18612 8668 18624
rect 7745 18584 8668 18612
rect 7745 18581 7757 18584
rect 7699 18575 7757 18581
rect 8662 18572 8668 18584
rect 8720 18572 8726 18624
rect 8754 18572 8760 18624
rect 8812 18612 8818 18624
rect 9125 18615 9183 18621
rect 9125 18612 9137 18615
rect 8812 18584 9137 18612
rect 8812 18572 8818 18584
rect 9125 18581 9137 18584
rect 9171 18612 9183 18615
rect 9582 18612 9588 18624
rect 9171 18584 9588 18612
rect 9171 18581 9183 18584
rect 9125 18575 9183 18581
rect 9582 18572 9588 18584
rect 9640 18572 9646 18624
rect 9950 18612 9956 18624
rect 9911 18584 9956 18612
rect 9950 18572 9956 18584
rect 10008 18572 10014 18624
rect 11698 18572 11704 18624
rect 11756 18612 11762 18624
rect 12710 18612 12716 18624
rect 11756 18584 12716 18612
rect 11756 18572 11762 18584
rect 12710 18572 12716 18584
rect 12768 18572 12774 18624
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 7834 18408 7840 18420
rect 7795 18380 7840 18408
rect 7834 18368 7840 18380
rect 7892 18368 7898 18420
rect 9858 18368 9864 18420
rect 9916 18408 9922 18420
rect 10045 18411 10103 18417
rect 10045 18408 10057 18411
rect 9916 18380 10057 18408
rect 9916 18368 9922 18380
rect 10045 18377 10057 18380
rect 10091 18377 10103 18411
rect 10045 18371 10103 18377
rect 11517 18411 11575 18417
rect 11517 18377 11529 18411
rect 11563 18408 11575 18411
rect 11882 18408 11888 18420
rect 11563 18380 11888 18408
rect 11563 18377 11575 18380
rect 11517 18371 11575 18377
rect 11882 18368 11888 18380
rect 11940 18368 11946 18420
rect 17310 18408 17316 18420
rect 17271 18380 17316 18408
rect 17310 18368 17316 18380
rect 17368 18368 17374 18420
rect 19058 18408 19064 18420
rect 19019 18380 19064 18408
rect 19058 18368 19064 18380
rect 19116 18368 19122 18420
rect 19426 18408 19432 18420
rect 19387 18380 19432 18408
rect 19426 18368 19432 18380
rect 19484 18368 19490 18420
rect 14274 18300 14280 18352
rect 14332 18340 14338 18352
rect 14332 18312 14412 18340
rect 14332 18300 14338 18312
rect 9769 18275 9827 18281
rect 9769 18241 9781 18275
rect 9815 18272 9827 18275
rect 9950 18272 9956 18284
rect 9815 18244 9956 18272
rect 9815 18241 9827 18244
rect 9769 18235 9827 18241
rect 9950 18232 9956 18244
rect 10008 18272 10014 18284
rect 10597 18275 10655 18281
rect 10597 18272 10609 18275
rect 10008 18244 10609 18272
rect 10008 18232 10014 18244
rect 10597 18241 10609 18244
rect 10643 18241 10655 18275
rect 12158 18272 12164 18284
rect 12119 18244 12164 18272
rect 10597 18235 10655 18241
rect 12158 18232 12164 18244
rect 12216 18272 12222 18284
rect 12618 18272 12624 18284
rect 12216 18244 12624 18272
rect 12216 18232 12222 18244
rect 12618 18232 12624 18244
rect 12676 18272 12682 18284
rect 13446 18272 13452 18284
rect 12676 18244 13216 18272
rect 13407 18244 13452 18272
rect 12676 18232 12682 18244
rect 1448 18207 1506 18213
rect 1448 18173 1460 18207
rect 1494 18204 1506 18207
rect 1535 18207 1593 18213
rect 1494 18173 1507 18204
rect 1448 18167 1507 18173
rect 1535 18173 1547 18207
rect 1581 18204 1593 18207
rect 1854 18204 1860 18216
rect 1581 18176 1860 18204
rect 1581 18173 1593 18176
rect 1535 18167 1593 18173
rect 1479 18136 1507 18167
rect 1854 18164 1860 18176
rect 1912 18164 1918 18216
rect 7006 18164 7012 18216
rect 7064 18213 7070 18216
rect 7064 18207 7102 18213
rect 7090 18204 7102 18207
rect 7469 18207 7527 18213
rect 7469 18204 7481 18207
rect 7090 18176 7481 18204
rect 7090 18173 7102 18176
rect 7064 18167 7102 18173
rect 7469 18173 7481 18176
rect 7515 18204 7527 18207
rect 8056 18207 8114 18213
rect 8056 18204 8068 18207
rect 7515 18176 8068 18204
rect 7515 18173 7527 18176
rect 7469 18167 7527 18173
rect 8056 18173 8068 18176
rect 8102 18204 8114 18207
rect 8481 18207 8539 18213
rect 8481 18204 8493 18207
rect 8102 18176 8493 18204
rect 8102 18173 8114 18176
rect 8056 18167 8114 18173
rect 8481 18173 8493 18176
rect 8527 18173 8539 18207
rect 9306 18204 9312 18216
rect 9267 18176 9312 18204
rect 8481 18167 8539 18173
rect 7064 18164 7070 18167
rect 9306 18164 9312 18176
rect 9364 18164 9370 18216
rect 9582 18204 9588 18216
rect 9543 18176 9588 18204
rect 9582 18164 9588 18176
rect 9640 18164 9646 18216
rect 12986 18204 12992 18216
rect 12947 18176 12992 18204
rect 12986 18164 12992 18176
rect 13044 18164 13050 18216
rect 13188 18213 13216 18244
rect 13446 18232 13452 18244
rect 13504 18232 13510 18284
rect 14384 18281 14412 18312
rect 14660 18312 16252 18340
rect 14660 18284 14688 18312
rect 14369 18275 14427 18281
rect 14369 18241 14381 18275
rect 14415 18272 14427 18275
rect 14642 18272 14648 18284
rect 14415 18244 14648 18272
rect 14415 18241 14427 18244
rect 14369 18235 14427 18241
rect 14642 18232 14648 18244
rect 14700 18232 14706 18284
rect 14826 18272 14832 18284
rect 14787 18244 14832 18272
rect 14826 18232 14832 18244
rect 14884 18232 14890 18284
rect 16224 18281 16252 18312
rect 16209 18275 16267 18281
rect 16209 18241 16221 18275
rect 16255 18241 16267 18275
rect 16209 18235 16267 18241
rect 18141 18275 18199 18281
rect 18141 18241 18153 18275
rect 18187 18272 18199 18275
rect 18230 18272 18236 18284
rect 18187 18244 18236 18272
rect 18187 18241 18199 18244
rect 18141 18235 18199 18241
rect 18230 18232 18236 18244
rect 18288 18232 18294 18284
rect 18785 18275 18843 18281
rect 18785 18241 18797 18275
rect 18831 18272 18843 18275
rect 19334 18272 19340 18284
rect 18831 18244 19340 18272
rect 18831 18241 18843 18244
rect 18785 18235 18843 18241
rect 19334 18232 19340 18244
rect 19392 18232 19398 18284
rect 13173 18207 13231 18213
rect 13173 18173 13185 18207
rect 13219 18173 13231 18207
rect 13173 18167 13231 18173
rect 19610 18164 19616 18216
rect 19668 18213 19674 18216
rect 19668 18207 19706 18213
rect 19694 18204 19706 18207
rect 20073 18207 20131 18213
rect 20073 18204 20085 18207
rect 19694 18176 20085 18204
rect 19694 18173 19706 18176
rect 19668 18167 19706 18173
rect 20073 18173 20085 18176
rect 20119 18204 20131 18207
rect 20254 18204 20260 18216
rect 20119 18176 20260 18204
rect 20119 18173 20131 18176
rect 20073 18167 20131 18173
rect 19668 18164 19674 18167
rect 20254 18164 20260 18176
rect 20312 18164 20318 18216
rect 8202 18145 8208 18148
rect 8159 18139 8208 18145
rect 1479 18108 1992 18136
rect 1964 18077 1992 18108
rect 8159 18105 8171 18139
rect 8205 18105 8208 18139
rect 8159 18099 8208 18105
rect 8202 18096 8208 18099
rect 8260 18096 8266 18148
rect 10918 18139 10976 18145
rect 10918 18136 10930 18139
rect 10704 18108 10930 18136
rect 10704 18080 10732 18108
rect 10918 18105 10930 18108
rect 10964 18105 10976 18139
rect 10918 18099 10976 18105
rect 14461 18139 14519 18145
rect 14461 18105 14473 18139
rect 14507 18105 14519 18139
rect 15930 18136 15936 18148
rect 15891 18108 15936 18136
rect 14461 18099 14519 18105
rect 1949 18071 2007 18077
rect 1949 18037 1961 18071
rect 1995 18068 2007 18071
rect 2314 18068 2320 18080
rect 1995 18040 2320 18068
rect 1995 18037 2007 18040
rect 1949 18031 2007 18037
rect 2314 18028 2320 18040
rect 2372 18028 2378 18080
rect 7190 18077 7196 18080
rect 7147 18071 7196 18077
rect 7147 18037 7159 18071
rect 7193 18037 7196 18071
rect 7147 18031 7196 18037
rect 7190 18028 7196 18031
rect 7248 18028 7254 18080
rect 8478 18028 8484 18080
rect 8536 18068 8542 18080
rect 8849 18071 8907 18077
rect 8849 18068 8861 18071
rect 8536 18040 8861 18068
rect 8536 18028 8542 18040
rect 8849 18037 8861 18040
rect 8895 18037 8907 18071
rect 8849 18031 8907 18037
rect 10505 18071 10563 18077
rect 10505 18037 10517 18071
rect 10551 18068 10563 18071
rect 10686 18068 10692 18080
rect 10551 18040 10692 18068
rect 10551 18037 10563 18040
rect 10505 18031 10563 18037
rect 10686 18028 10692 18040
rect 10744 18028 10750 18080
rect 13078 18028 13084 18080
rect 13136 18068 13142 18080
rect 13725 18071 13783 18077
rect 13725 18068 13737 18071
rect 13136 18040 13737 18068
rect 13136 18028 13142 18040
rect 13725 18037 13737 18040
rect 13771 18037 13783 18071
rect 13725 18031 13783 18037
rect 14185 18071 14243 18077
rect 14185 18037 14197 18071
rect 14231 18068 14243 18071
rect 14274 18068 14280 18080
rect 14231 18040 14280 18068
rect 14231 18037 14243 18040
rect 14185 18031 14243 18037
rect 14274 18028 14280 18040
rect 14332 18068 14338 18080
rect 14476 18068 14504 18099
rect 15930 18096 15936 18108
rect 15988 18096 15994 18148
rect 16022 18096 16028 18148
rect 16080 18136 16086 18148
rect 18233 18139 18291 18145
rect 16080 18108 16125 18136
rect 16080 18096 16086 18108
rect 18233 18105 18245 18139
rect 18279 18105 18291 18139
rect 18233 18099 18291 18105
rect 15378 18068 15384 18080
rect 14332 18040 14504 18068
rect 15339 18040 15384 18068
rect 14332 18028 14338 18040
rect 15378 18028 15384 18040
rect 15436 18028 15442 18080
rect 16850 18028 16856 18080
rect 16908 18068 16914 18080
rect 16945 18071 17003 18077
rect 16945 18068 16957 18071
rect 16908 18040 16957 18068
rect 16908 18028 16914 18040
rect 16945 18037 16957 18040
rect 16991 18037 17003 18071
rect 17770 18068 17776 18080
rect 17731 18040 17776 18068
rect 16945 18031 17003 18037
rect 17770 18028 17776 18040
rect 17828 18068 17834 18080
rect 18248 18068 18276 18099
rect 17828 18040 18276 18068
rect 19751 18071 19809 18077
rect 17828 18028 17834 18040
rect 19751 18037 19763 18071
rect 19797 18068 19809 18071
rect 19978 18068 19984 18080
rect 19797 18040 19984 18068
rect 19797 18037 19809 18040
rect 19751 18031 19809 18037
rect 19978 18028 19984 18040
rect 20036 18028 20042 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 9125 17867 9183 17873
rect 9125 17833 9137 17867
rect 9171 17864 9183 17867
rect 9306 17864 9312 17876
rect 9171 17836 9312 17864
rect 9171 17833 9183 17836
rect 9125 17827 9183 17833
rect 9306 17824 9312 17836
rect 9364 17824 9370 17876
rect 9953 17867 10011 17873
rect 9953 17833 9965 17867
rect 9999 17864 10011 17867
rect 10042 17864 10048 17876
rect 9999 17836 10048 17864
rect 9999 17833 10011 17836
rect 9953 17827 10011 17833
rect 10042 17824 10048 17836
rect 10100 17824 10106 17876
rect 11054 17824 11060 17876
rect 11112 17864 11118 17876
rect 12805 17867 12863 17873
rect 11112 17836 11192 17864
rect 11112 17824 11118 17836
rect 1670 17796 1676 17808
rect 1479 17768 1676 17796
rect 1479 17737 1507 17768
rect 1670 17756 1676 17768
rect 1728 17796 1734 17808
rect 2682 17796 2688 17808
rect 1728 17768 2688 17796
rect 1728 17756 1734 17768
rect 2682 17756 2688 17768
rect 2740 17756 2746 17808
rect 7377 17799 7435 17805
rect 7377 17765 7389 17799
rect 7423 17796 7435 17799
rect 7558 17796 7564 17808
rect 7423 17768 7564 17796
rect 7423 17765 7435 17768
rect 7377 17759 7435 17765
rect 7558 17756 7564 17768
rect 7616 17756 7622 17808
rect 7653 17799 7711 17805
rect 7653 17765 7665 17799
rect 7699 17796 7711 17799
rect 7834 17796 7840 17808
rect 7699 17768 7840 17796
rect 7699 17765 7711 17768
rect 7653 17759 7711 17765
rect 7834 17756 7840 17768
rect 7892 17756 7898 17808
rect 11164 17805 11192 17836
rect 12805 17833 12817 17867
rect 12851 17864 12863 17867
rect 12986 17864 12992 17876
rect 12851 17836 12992 17864
rect 12851 17833 12863 17836
rect 12805 17827 12863 17833
rect 12986 17824 12992 17836
rect 13044 17824 13050 17876
rect 13357 17867 13415 17873
rect 13357 17833 13369 17867
rect 13403 17864 13415 17867
rect 13446 17864 13452 17876
rect 13403 17836 13452 17864
rect 13403 17833 13415 17836
rect 13357 17827 13415 17833
rect 13446 17824 13452 17836
rect 13504 17824 13510 17876
rect 14274 17824 14280 17876
rect 14332 17864 14338 17876
rect 14369 17867 14427 17873
rect 14369 17864 14381 17867
rect 14332 17836 14381 17864
rect 14332 17824 14338 17836
rect 14369 17833 14381 17836
rect 14415 17833 14427 17867
rect 14642 17864 14648 17876
rect 14603 17836 14648 17864
rect 14369 17827 14427 17833
rect 14642 17824 14648 17836
rect 14700 17824 14706 17876
rect 15427 17867 15485 17873
rect 15427 17833 15439 17867
rect 15473 17864 15485 17867
rect 15930 17864 15936 17876
rect 15473 17836 15936 17864
rect 15473 17833 15485 17836
rect 15427 17827 15485 17833
rect 15930 17824 15936 17836
rect 15988 17864 15994 17876
rect 16577 17867 16635 17873
rect 16577 17864 16589 17867
rect 15988 17836 16589 17864
rect 15988 17824 15994 17836
rect 16577 17833 16589 17836
rect 16623 17833 16635 17867
rect 16577 17827 16635 17833
rect 17681 17867 17739 17873
rect 17681 17833 17693 17867
rect 17727 17864 17739 17867
rect 17770 17864 17776 17876
rect 17727 17836 17776 17864
rect 17727 17833 17739 17836
rect 17681 17827 17739 17833
rect 17770 17824 17776 17836
rect 17828 17824 17834 17876
rect 18141 17867 18199 17873
rect 18141 17833 18153 17867
rect 18187 17864 18199 17867
rect 18230 17864 18236 17876
rect 18187 17836 18236 17864
rect 18187 17833 18199 17836
rect 18141 17827 18199 17833
rect 18230 17824 18236 17836
rect 18288 17824 18294 17876
rect 18322 17824 18328 17876
rect 18380 17864 18386 17876
rect 18509 17867 18567 17873
rect 18509 17864 18521 17867
rect 18380 17836 18521 17864
rect 18380 17824 18386 17836
rect 18509 17833 18521 17836
rect 18555 17833 18567 17867
rect 18509 17827 18567 17833
rect 11149 17799 11207 17805
rect 11149 17765 11161 17799
rect 11195 17765 11207 17799
rect 11149 17759 11207 17765
rect 11241 17799 11299 17805
rect 11241 17765 11253 17799
rect 11287 17796 11299 17799
rect 11514 17796 11520 17808
rect 11287 17768 11520 17796
rect 11287 17765 11299 17768
rect 11241 17759 11299 17765
rect 11514 17756 11520 17768
rect 11572 17756 11578 17808
rect 11793 17799 11851 17805
rect 11793 17765 11805 17799
rect 11839 17796 11851 17799
rect 12066 17796 12072 17808
rect 11839 17768 12072 17796
rect 11839 17765 11851 17768
rect 11793 17759 11851 17765
rect 12066 17756 12072 17768
rect 12124 17756 12130 17808
rect 13078 17756 13084 17808
rect 13136 17796 13142 17808
rect 13770 17799 13828 17805
rect 13770 17796 13782 17799
rect 13136 17768 13782 17796
rect 13136 17756 13142 17768
rect 13770 17765 13782 17768
rect 13816 17765 13828 17799
rect 13770 17759 13828 17765
rect 16850 17756 16856 17808
rect 16908 17796 16914 17808
rect 17082 17799 17140 17805
rect 17082 17796 17094 17799
rect 16908 17768 17094 17796
rect 16908 17756 16914 17768
rect 17082 17765 17094 17768
rect 17128 17765 17140 17799
rect 17082 17759 17140 17765
rect 1464 17731 1522 17737
rect 1464 17697 1476 17731
rect 1510 17697 1522 17731
rect 1464 17691 1522 17697
rect 2222 17688 2228 17740
rect 2280 17728 2286 17740
rect 2501 17731 2559 17737
rect 2501 17728 2513 17731
rect 2280 17700 2513 17728
rect 2280 17688 2286 17700
rect 2501 17697 2513 17700
rect 2547 17697 2559 17731
rect 5442 17728 5448 17740
rect 5403 17700 5448 17728
rect 2501 17691 2559 17697
rect 5442 17688 5448 17700
rect 5500 17688 5506 17740
rect 6546 17737 6552 17740
rect 6524 17731 6552 17737
rect 6524 17728 6536 17731
rect 6459 17700 6536 17728
rect 6524 17697 6536 17700
rect 6604 17728 6610 17740
rect 6730 17728 6736 17740
rect 6604 17700 6736 17728
rect 6524 17691 6552 17697
rect 6546 17688 6552 17691
rect 6604 17688 6610 17700
rect 6730 17688 6736 17700
rect 6788 17688 6794 17740
rect 9950 17688 9956 17740
rect 10008 17728 10014 17740
rect 10080 17731 10138 17737
rect 10080 17728 10092 17731
rect 10008 17700 10092 17728
rect 10008 17688 10014 17700
rect 10080 17697 10092 17700
rect 10126 17697 10138 17731
rect 10080 17691 10138 17697
rect 15286 17688 15292 17740
rect 15344 17737 15350 17740
rect 15344 17731 15382 17737
rect 15370 17697 15382 17731
rect 15344 17691 15382 17697
rect 15344 17688 15350 17691
rect 8018 17660 8024 17672
rect 7979 17632 8024 17660
rect 8018 17620 8024 17632
rect 8076 17620 8082 17672
rect 11790 17620 11796 17672
rect 11848 17660 11854 17672
rect 12069 17663 12127 17669
rect 12069 17660 12081 17663
rect 11848 17632 12081 17660
rect 11848 17620 11854 17632
rect 12069 17629 12081 17632
rect 12115 17629 12127 17663
rect 13446 17660 13452 17672
rect 13407 17632 13452 17660
rect 12069 17623 12127 17629
rect 13446 17620 13452 17632
rect 13504 17620 13510 17672
rect 16758 17660 16764 17672
rect 16719 17632 16764 17660
rect 16758 17620 16764 17632
rect 16816 17620 16822 17672
rect 15841 17595 15899 17601
rect 15841 17561 15853 17595
rect 15887 17592 15899 17595
rect 16206 17592 16212 17604
rect 15887 17564 16212 17592
rect 15887 17561 15899 17564
rect 15841 17555 15899 17561
rect 16206 17552 16212 17564
rect 16264 17552 16270 17604
rect 1535 17527 1593 17533
rect 1535 17493 1547 17527
rect 1581 17524 1593 17527
rect 2130 17524 2136 17536
rect 1581 17496 2136 17524
rect 1581 17493 1593 17496
rect 1535 17487 1593 17493
rect 2130 17484 2136 17496
rect 2188 17484 2194 17536
rect 2682 17524 2688 17536
rect 2643 17496 2688 17524
rect 2682 17484 2688 17496
rect 2740 17484 2746 17536
rect 5629 17527 5687 17533
rect 5629 17493 5641 17527
rect 5675 17524 5687 17527
rect 6178 17524 6184 17536
rect 5675 17496 6184 17524
rect 5675 17493 5687 17496
rect 5629 17487 5687 17493
rect 6178 17484 6184 17496
rect 6236 17484 6242 17536
rect 6362 17484 6368 17536
rect 6420 17524 6426 17536
rect 6595 17527 6653 17533
rect 6595 17524 6607 17527
rect 6420 17496 6607 17524
rect 6420 17484 6426 17496
rect 6595 17493 6607 17496
rect 6641 17493 6653 17527
rect 6595 17487 6653 17493
rect 10134 17484 10140 17536
rect 10192 17533 10198 17536
rect 10192 17527 10241 17533
rect 10192 17493 10195 17527
rect 10229 17493 10241 17527
rect 10192 17487 10241 17493
rect 10689 17527 10747 17533
rect 10689 17493 10701 17527
rect 10735 17524 10747 17527
rect 10962 17524 10968 17536
rect 10735 17496 10968 17524
rect 10735 17493 10747 17496
rect 10689 17487 10747 17493
rect 10192 17484 10198 17487
rect 10962 17484 10968 17496
rect 11020 17484 11026 17536
rect 16298 17524 16304 17536
rect 16259 17496 16304 17524
rect 16298 17484 16304 17496
rect 16356 17484 16362 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1670 17320 1676 17332
rect 1631 17292 1676 17320
rect 1670 17280 1676 17292
rect 1728 17280 1734 17332
rect 2682 17320 2688 17332
rect 2643 17292 2688 17320
rect 2682 17280 2688 17292
rect 2740 17280 2746 17332
rect 6270 17320 6276 17332
rect 6231 17292 6276 17320
rect 6270 17280 6276 17292
rect 6328 17280 6334 17332
rect 11514 17320 11520 17332
rect 11475 17292 11520 17320
rect 11514 17280 11520 17292
rect 11572 17320 11578 17332
rect 11793 17323 11851 17329
rect 11793 17320 11805 17323
rect 11572 17292 11805 17320
rect 11572 17280 11578 17292
rect 11793 17289 11805 17292
rect 11839 17289 11851 17323
rect 12618 17320 12624 17332
rect 12579 17292 12624 17320
rect 11793 17283 11851 17289
rect 12618 17280 12624 17292
rect 12676 17280 12682 17332
rect 14458 17320 14464 17332
rect 14419 17292 14464 17320
rect 14458 17280 14464 17292
rect 14516 17280 14522 17332
rect 8018 17252 8024 17264
rect 7979 17224 8024 17252
rect 8018 17212 8024 17224
rect 8076 17212 8082 17264
rect 2866 17184 2872 17196
rect 2827 17156 2872 17184
rect 2866 17144 2872 17156
rect 2924 17144 2930 17196
rect 3050 17144 3056 17196
rect 3108 17184 3114 17196
rect 3145 17187 3203 17193
rect 3145 17184 3157 17187
rect 3108 17156 3157 17184
rect 3108 17144 3114 17156
rect 3145 17153 3157 17156
rect 3191 17153 3203 17187
rect 3145 17147 3203 17153
rect 5442 17144 5448 17196
rect 5500 17184 5506 17196
rect 5537 17187 5595 17193
rect 5537 17184 5549 17187
rect 5500 17156 5549 17184
rect 5500 17144 5506 17156
rect 5537 17153 5549 17156
rect 5583 17184 5595 17187
rect 6638 17184 6644 17196
rect 5583 17156 6644 17184
rect 5583 17153 5595 17156
rect 5537 17147 5595 17153
rect 6638 17144 6644 17156
rect 6696 17144 6702 17196
rect 7285 17187 7343 17193
rect 7285 17153 7297 17187
rect 7331 17184 7343 17187
rect 7834 17184 7840 17196
rect 7331 17156 7840 17184
rect 7331 17153 7343 17156
rect 7285 17147 7343 17153
rect 7834 17144 7840 17156
rect 7892 17184 7898 17196
rect 8941 17187 8999 17193
rect 8941 17184 8953 17187
rect 7892 17156 8953 17184
rect 7892 17144 7898 17156
rect 8941 17153 8953 17156
rect 8987 17153 8999 17187
rect 8941 17147 8999 17153
rect 10597 17187 10655 17193
rect 10597 17153 10609 17187
rect 10643 17184 10655 17187
rect 10962 17184 10968 17196
rect 10643 17156 10968 17184
rect 10643 17153 10655 17156
rect 10597 17147 10655 17153
rect 10962 17144 10968 17156
rect 11020 17144 11026 17196
rect 13446 17144 13452 17196
rect 13504 17184 13510 17196
rect 14737 17187 14795 17193
rect 14737 17184 14749 17187
rect 13504 17156 14749 17184
rect 13504 17144 13510 17156
rect 14737 17153 14749 17156
rect 14783 17153 14795 17187
rect 15286 17184 15292 17196
rect 15247 17156 15292 17184
rect 14737 17147 14795 17153
rect 15286 17144 15292 17156
rect 15344 17144 15350 17196
rect 18230 17144 18236 17196
rect 18288 17184 18294 17196
rect 18417 17187 18475 17193
rect 18417 17184 18429 17187
rect 18288 17156 18429 17184
rect 18288 17144 18294 17156
rect 18417 17153 18429 17156
rect 18463 17153 18475 17187
rect 18417 17147 18475 17153
rect 5772 17119 5830 17125
rect 5772 17085 5784 17119
rect 5818 17116 5830 17119
rect 6270 17116 6276 17128
rect 5818 17088 6276 17116
rect 5818 17085 5830 17088
rect 5772 17079 5830 17085
rect 6270 17076 6276 17088
rect 6328 17076 6334 17128
rect 8481 17119 8539 17125
rect 8481 17085 8493 17119
rect 8527 17116 8539 17119
rect 8849 17119 8907 17125
rect 8849 17116 8861 17119
rect 8527 17088 8861 17116
rect 8527 17085 8539 17088
rect 8481 17079 8539 17085
rect 8849 17085 8861 17088
rect 8895 17116 8907 17119
rect 9033 17119 9091 17125
rect 9033 17116 9045 17119
rect 8895 17088 9045 17116
rect 8895 17085 8907 17088
rect 8849 17079 8907 17085
rect 9033 17085 9045 17088
rect 9079 17085 9091 17119
rect 9033 17079 9091 17085
rect 12253 17119 12311 17125
rect 12253 17085 12265 17119
rect 12299 17116 12311 17119
rect 12437 17119 12495 17125
rect 12437 17116 12449 17119
rect 12299 17088 12449 17116
rect 12299 17085 12311 17088
rect 12253 17079 12311 17085
rect 12437 17085 12449 17088
rect 12483 17116 12495 17119
rect 13354 17116 13360 17128
rect 12483 17088 13360 17116
rect 12483 17085 12495 17088
rect 12437 17079 12495 17085
rect 2682 17008 2688 17060
rect 2740 17048 2746 17060
rect 2961 17051 3019 17057
rect 2961 17048 2973 17051
rect 2740 17020 2973 17048
rect 2740 17008 2746 17020
rect 2961 17017 2973 17020
rect 3007 17017 3019 17051
rect 2961 17011 3019 17017
rect 5859 17051 5917 17057
rect 5859 17017 5871 17051
rect 5905 17048 5917 17051
rect 7466 17048 7472 17060
rect 5905 17020 7472 17048
rect 5905 17017 5917 17020
rect 5859 17011 5917 17017
rect 1762 16980 1768 16992
rect 1723 16952 1768 16980
rect 1762 16940 1768 16952
rect 1820 16940 1826 16992
rect 2222 16980 2228 16992
rect 2183 16952 2228 16980
rect 2222 16940 2228 16952
rect 2280 16940 2286 16992
rect 2976 16980 3004 17011
rect 7466 17008 7472 17020
rect 7524 17008 7530 17060
rect 7561 17051 7619 17057
rect 7561 17017 7573 17051
rect 7607 17017 7619 17051
rect 7561 17011 7619 17017
rect 4154 16980 4160 16992
rect 2976 16952 4160 16980
rect 4154 16940 4160 16952
rect 4212 16940 4218 16992
rect 6641 16983 6699 16989
rect 6641 16949 6653 16983
rect 6687 16980 6699 16983
rect 6730 16980 6736 16992
rect 6687 16952 6736 16980
rect 6687 16949 6699 16952
rect 6641 16943 6699 16949
rect 6730 16940 6736 16952
rect 6788 16940 6794 16992
rect 7576 16980 7604 17011
rect 7834 16980 7840 16992
rect 7576 16952 7840 16980
rect 7834 16940 7840 16952
rect 7892 16980 7898 16992
rect 8496 16980 8524 17079
rect 13354 17076 13360 17088
rect 13412 17076 13418 17128
rect 13538 17116 13544 17128
rect 13499 17088 13544 17116
rect 13538 17076 13544 17088
rect 13596 17076 13602 17128
rect 16209 17119 16267 17125
rect 16209 17085 16221 17119
rect 16255 17116 16267 17119
rect 16298 17116 16304 17128
rect 16255 17088 16304 17116
rect 16255 17085 16267 17088
rect 16209 17079 16267 17085
rect 16298 17076 16304 17088
rect 16356 17076 16362 17128
rect 10505 17051 10563 17057
rect 10505 17017 10517 17051
rect 10551 17048 10563 17051
rect 10686 17048 10692 17060
rect 10551 17020 10692 17048
rect 10551 17017 10563 17020
rect 10505 17011 10563 17017
rect 10686 17008 10692 17020
rect 10744 17048 10750 17060
rect 10959 17051 11017 17057
rect 10959 17048 10971 17051
rect 10744 17020 10971 17048
rect 10744 17008 10750 17020
rect 10959 17017 10971 17020
rect 11005 17048 11017 17051
rect 13882 17051 13940 17057
rect 11005 17020 13124 17048
rect 11005 17017 11017 17020
rect 10959 17011 11017 17017
rect 13096 16992 13124 17020
rect 13882 17017 13894 17051
rect 13928 17048 13940 17051
rect 16571 17051 16629 17057
rect 13928 17017 13946 17048
rect 13882 17011 13946 17017
rect 16571 17017 16583 17051
rect 16617 17048 16629 17051
rect 17405 17051 17463 17057
rect 17405 17048 17417 17051
rect 16617 17020 16651 17048
rect 16868 17020 17417 17048
rect 16617 17017 16629 17020
rect 16571 17011 16629 17017
rect 7892 16952 8524 16980
rect 7892 16940 7898 16952
rect 9950 16940 9956 16992
rect 10008 16980 10014 16992
rect 10045 16983 10103 16989
rect 10045 16980 10057 16983
rect 10008 16952 10057 16980
rect 10008 16940 10014 16952
rect 10045 16949 10057 16952
rect 10091 16949 10103 16983
rect 13078 16980 13084 16992
rect 12991 16952 13084 16980
rect 10045 16943 10103 16949
rect 13078 16940 13084 16952
rect 13136 16980 13142 16992
rect 13354 16980 13360 16992
rect 13136 16952 13360 16980
rect 13136 16940 13142 16952
rect 13354 16940 13360 16952
rect 13412 16980 13418 16992
rect 13449 16983 13507 16989
rect 13449 16980 13461 16983
rect 13412 16952 13461 16980
rect 13412 16940 13418 16952
rect 13449 16949 13461 16952
rect 13495 16980 13507 16983
rect 13918 16980 13946 17011
rect 16117 16983 16175 16989
rect 16117 16980 16129 16983
rect 13495 16952 16129 16980
rect 13495 16949 13507 16952
rect 13449 16943 13507 16949
rect 16117 16949 16129 16952
rect 16163 16980 16175 16983
rect 16586 16980 16614 17011
rect 16868 16992 16896 17020
rect 17405 17017 17417 17020
rect 17451 17017 17463 17051
rect 18138 17048 18144 17060
rect 18099 17020 18144 17048
rect 17405 17011 17463 17017
rect 18138 17008 18144 17020
rect 18196 17008 18202 17060
rect 18233 17051 18291 17057
rect 18233 17017 18245 17051
rect 18279 17048 18291 17051
rect 18414 17048 18420 17060
rect 18279 17020 18420 17048
rect 18279 17017 18291 17020
rect 18233 17011 18291 17017
rect 16850 16980 16856 16992
rect 16163 16952 16856 16980
rect 16163 16949 16175 16952
rect 16117 16943 16175 16949
rect 16850 16940 16856 16952
rect 16908 16940 16914 16992
rect 17129 16983 17187 16989
rect 17129 16949 17141 16983
rect 17175 16980 17187 16983
rect 17865 16983 17923 16989
rect 17865 16980 17877 16983
rect 17175 16952 17877 16980
rect 17175 16949 17187 16952
rect 17129 16943 17187 16949
rect 17865 16949 17877 16952
rect 17911 16980 17923 16983
rect 18248 16980 18276 17011
rect 18414 17008 18420 17020
rect 18472 17008 18478 17060
rect 17911 16952 18276 16980
rect 17911 16949 17923 16952
rect 17865 16943 17923 16949
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 2866 16736 2872 16788
rect 2924 16776 2930 16788
rect 3053 16779 3111 16785
rect 3053 16776 3065 16779
rect 2924 16748 3065 16776
rect 2924 16736 2930 16748
rect 3053 16745 3065 16748
rect 3099 16745 3111 16779
rect 7834 16776 7840 16788
rect 7795 16748 7840 16776
rect 3053 16739 3111 16745
rect 7834 16736 7840 16748
rect 7892 16736 7898 16788
rect 11054 16736 11060 16788
rect 11112 16776 11118 16788
rect 11793 16779 11851 16785
rect 11793 16776 11805 16779
rect 11112 16748 11805 16776
rect 11112 16736 11118 16748
rect 11793 16745 11805 16748
rect 11839 16745 11851 16779
rect 12618 16776 12624 16788
rect 12579 16748 12624 16776
rect 11793 16739 11851 16745
rect 12618 16736 12624 16748
rect 12676 16736 12682 16788
rect 17451 16779 17509 16785
rect 17451 16745 17463 16779
rect 17497 16776 17509 16779
rect 18138 16776 18144 16788
rect 17497 16748 18144 16776
rect 17497 16745 17509 16748
rect 17451 16739 17509 16745
rect 18138 16736 18144 16748
rect 18196 16736 18202 16788
rect 2130 16708 2136 16720
rect 2091 16680 2136 16708
rect 2130 16668 2136 16680
rect 2188 16668 2194 16720
rect 2222 16668 2228 16720
rect 2280 16708 2286 16720
rect 2280 16680 2325 16708
rect 2280 16668 2286 16680
rect 4154 16668 4160 16720
rect 4212 16708 4218 16720
rect 4249 16711 4307 16717
rect 4249 16708 4261 16711
rect 4212 16680 4261 16708
rect 4212 16668 4218 16680
rect 4249 16677 4261 16680
rect 4295 16677 4307 16711
rect 4249 16671 4307 16677
rect 7006 16668 7012 16720
rect 7064 16708 7070 16720
rect 7238 16711 7296 16717
rect 7238 16708 7250 16711
rect 7064 16680 7250 16708
rect 7064 16668 7070 16680
rect 7238 16677 7250 16680
rect 7284 16677 7296 16711
rect 7238 16671 7296 16677
rect 7466 16668 7472 16720
rect 7524 16708 7530 16720
rect 8113 16711 8171 16717
rect 8113 16708 8125 16711
rect 7524 16680 8125 16708
rect 7524 16668 7530 16680
rect 8113 16677 8125 16680
rect 8159 16677 8171 16711
rect 8113 16671 8171 16677
rect 10686 16668 10692 16720
rect 10744 16708 10750 16720
rect 10918 16711 10976 16717
rect 10918 16708 10930 16711
rect 10744 16680 10930 16708
rect 10744 16668 10750 16680
rect 10918 16677 10930 16680
rect 10964 16677 10976 16711
rect 12636 16708 12664 16736
rect 13078 16708 13084 16720
rect 12636 16680 13084 16708
rect 10918 16671 10976 16677
rect 13078 16668 13084 16680
rect 13136 16708 13142 16720
rect 13136 16680 13400 16708
rect 13136 16668 13142 16680
rect 6914 16640 6920 16652
rect 6875 16612 6920 16640
rect 6914 16600 6920 16612
rect 6972 16600 6978 16652
rect 11146 16640 11152 16652
rect 11072 16612 11152 16640
rect 4157 16575 4215 16581
rect 4157 16541 4169 16575
rect 4203 16572 4215 16575
rect 4246 16572 4252 16584
rect 4203 16544 4252 16572
rect 4203 16541 4215 16544
rect 4157 16535 4215 16541
rect 4246 16532 4252 16544
rect 4304 16532 4310 16584
rect 4338 16532 4344 16584
rect 4396 16572 4402 16584
rect 4433 16575 4491 16581
rect 4433 16572 4445 16575
rect 4396 16544 4445 16572
rect 4396 16532 4402 16544
rect 4433 16541 4445 16544
rect 4479 16541 4491 16575
rect 4433 16535 4491 16541
rect 5905 16575 5963 16581
rect 5905 16541 5917 16575
rect 5951 16572 5963 16575
rect 6454 16572 6460 16584
rect 5951 16544 6460 16572
rect 5951 16541 5963 16544
rect 5905 16535 5963 16541
rect 6454 16532 6460 16544
rect 6512 16532 6518 16584
rect 10597 16575 10655 16581
rect 10597 16541 10609 16575
rect 10643 16572 10655 16575
rect 10686 16572 10692 16584
rect 10643 16544 10692 16572
rect 10643 16541 10655 16544
rect 10597 16535 10655 16541
rect 10686 16532 10692 16544
rect 10744 16532 10750 16584
rect 10870 16532 10876 16584
rect 10928 16572 10934 16584
rect 11072 16572 11100 16612
rect 11146 16600 11152 16612
rect 11204 16640 11210 16652
rect 13372 16649 13400 16680
rect 13538 16668 13544 16720
rect 13596 16708 13602 16720
rect 13633 16711 13691 16717
rect 13633 16708 13645 16711
rect 13596 16680 13645 16708
rect 13596 16668 13602 16680
rect 13633 16677 13645 16680
rect 13679 16708 13691 16711
rect 13909 16711 13967 16717
rect 13909 16708 13921 16711
rect 13679 16680 13921 16708
rect 13679 16677 13691 16680
rect 13633 16671 13691 16677
rect 13909 16677 13921 16680
rect 13955 16677 13967 16711
rect 13909 16671 13967 16677
rect 16485 16711 16543 16717
rect 16485 16677 16497 16711
rect 16531 16708 16543 16711
rect 16758 16708 16764 16720
rect 16531 16680 16764 16708
rect 16531 16677 16543 16680
rect 16485 16671 16543 16677
rect 16758 16668 16764 16680
rect 16816 16668 16822 16720
rect 17954 16668 17960 16720
rect 18012 16708 18018 16720
rect 18463 16711 18521 16717
rect 18463 16708 18475 16711
rect 18012 16680 18475 16708
rect 18012 16668 18018 16680
rect 18463 16677 18475 16680
rect 18509 16677 18521 16711
rect 18463 16671 18521 16677
rect 11517 16643 11575 16649
rect 11517 16640 11529 16643
rect 11204 16612 11529 16640
rect 11204 16600 11210 16612
rect 11517 16609 11529 16612
rect 11563 16609 11575 16643
rect 11517 16603 11575 16609
rect 13173 16643 13231 16649
rect 13173 16609 13185 16643
rect 13219 16609 13231 16643
rect 13173 16603 13231 16609
rect 13357 16643 13415 16649
rect 13357 16609 13369 16643
rect 13403 16609 13415 16643
rect 14366 16640 14372 16652
rect 14327 16612 14372 16640
rect 13357 16603 13415 16609
rect 10928 16544 11100 16572
rect 13188 16572 13216 16603
rect 14366 16600 14372 16612
rect 14424 16600 14430 16652
rect 15654 16600 15660 16652
rect 15712 16640 15718 16652
rect 15749 16643 15807 16649
rect 15749 16640 15761 16643
rect 15712 16612 15761 16640
rect 15712 16600 15718 16612
rect 15749 16609 15761 16612
rect 15795 16609 15807 16643
rect 16206 16640 16212 16652
rect 16167 16612 16212 16640
rect 15749 16603 15807 16609
rect 16206 16600 16212 16612
rect 16264 16600 16270 16652
rect 17310 16600 17316 16652
rect 17368 16649 17374 16652
rect 17368 16643 17406 16649
rect 17394 16609 17406 16643
rect 17368 16603 17406 16609
rect 17368 16600 17374 16603
rect 18322 16600 18328 16652
rect 18380 16649 18386 16652
rect 18380 16643 18418 16649
rect 18406 16609 18418 16643
rect 18380 16603 18418 16609
rect 18380 16600 18386 16603
rect 13630 16572 13636 16584
rect 13188 16544 13636 16572
rect 10928 16532 10934 16544
rect 13630 16532 13636 16544
rect 13688 16532 13694 16584
rect 2685 16507 2743 16513
rect 2685 16473 2697 16507
rect 2731 16504 2743 16507
rect 2866 16504 2872 16516
rect 2731 16476 2872 16504
rect 2731 16473 2743 16476
rect 2685 16467 2743 16473
rect 2866 16464 2872 16476
rect 2924 16464 2930 16516
rect 4430 16396 4436 16448
rect 4488 16436 4494 16448
rect 5077 16439 5135 16445
rect 5077 16436 5089 16439
rect 4488 16408 5089 16436
rect 4488 16396 4494 16408
rect 5077 16405 5089 16408
rect 5123 16405 5135 16439
rect 5077 16399 5135 16405
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 1673 16235 1731 16241
rect 1673 16201 1685 16235
rect 1719 16232 1731 16235
rect 2222 16232 2228 16244
rect 1719 16204 2228 16232
rect 1719 16201 1731 16204
rect 1673 16195 1731 16201
rect 2222 16192 2228 16204
rect 2280 16192 2286 16244
rect 4154 16232 4160 16244
rect 4115 16204 4160 16232
rect 4154 16192 4160 16204
rect 4212 16192 4218 16244
rect 4246 16192 4252 16244
rect 4304 16232 4310 16244
rect 5353 16235 5411 16241
rect 5353 16232 5365 16235
rect 4304 16204 5365 16232
rect 4304 16192 4310 16204
rect 5353 16201 5365 16204
rect 5399 16201 5411 16235
rect 8018 16232 8024 16244
rect 7979 16204 8024 16232
rect 5353 16195 5411 16201
rect 8018 16192 8024 16204
rect 8076 16192 8082 16244
rect 10413 16235 10471 16241
rect 10413 16201 10425 16235
rect 10459 16232 10471 16235
rect 10594 16232 10600 16244
rect 10459 16204 10600 16232
rect 10459 16201 10471 16204
rect 10413 16195 10471 16201
rect 10594 16192 10600 16204
rect 10652 16192 10658 16244
rect 18322 16192 18328 16244
rect 18380 16232 18386 16244
rect 18877 16235 18935 16241
rect 18877 16232 18889 16235
rect 18380 16204 18889 16232
rect 18380 16192 18386 16204
rect 18877 16201 18889 16204
rect 18923 16201 18935 16235
rect 18877 16195 18935 16201
rect 2240 16164 2268 16192
rect 2774 16164 2780 16176
rect 2240 16136 2780 16164
rect 2774 16124 2780 16136
rect 2832 16124 2838 16176
rect 2976 16136 4476 16164
rect 1903 16099 1961 16105
rect 1903 16065 1915 16099
rect 1949 16096 1961 16099
rect 2976 16096 3004 16136
rect 4448 16108 4476 16136
rect 3142 16096 3148 16108
rect 1949 16068 3004 16096
rect 3103 16068 3148 16096
rect 1949 16065 1961 16068
rect 1903 16059 1961 16065
rect 3142 16056 3148 16068
rect 3200 16056 3206 16108
rect 4430 16096 4436 16108
rect 4391 16068 4436 16096
rect 4430 16056 4436 16068
rect 4488 16056 4494 16108
rect 4706 16096 4712 16108
rect 4667 16068 4712 16096
rect 4706 16056 4712 16068
rect 4764 16056 4770 16108
rect 7009 16099 7067 16105
rect 7009 16065 7021 16099
rect 7055 16096 7067 16099
rect 8036 16096 8064 16192
rect 11054 16124 11060 16176
rect 11112 16164 11118 16176
rect 11149 16167 11207 16173
rect 11149 16164 11161 16167
rect 11112 16136 11161 16164
rect 11112 16124 11118 16136
rect 11149 16133 11161 16136
rect 11195 16133 11207 16167
rect 11149 16127 11207 16133
rect 11606 16124 11612 16176
rect 11664 16164 11670 16176
rect 12253 16167 12311 16173
rect 12253 16164 12265 16167
rect 11664 16136 12265 16164
rect 11664 16124 11670 16136
rect 12253 16133 12265 16136
rect 12299 16164 12311 16167
rect 12710 16164 12716 16176
rect 12299 16136 12716 16164
rect 12299 16133 12311 16136
rect 12253 16127 12311 16133
rect 12710 16124 12716 16136
rect 12768 16164 12774 16176
rect 15654 16164 15660 16176
rect 12768 16136 15660 16164
rect 12768 16124 12774 16136
rect 15654 16124 15660 16136
rect 15712 16124 15718 16176
rect 7055 16068 8064 16096
rect 7055 16065 7067 16068
rect 7009 16059 7067 16065
rect 10134 16056 10140 16108
rect 10192 16096 10198 16108
rect 10597 16099 10655 16105
rect 10597 16096 10609 16099
rect 10192 16068 10609 16096
rect 10192 16056 10198 16068
rect 10597 16065 10609 16068
rect 10643 16096 10655 16099
rect 11517 16099 11575 16105
rect 11517 16096 11529 16099
rect 10643 16068 11529 16096
rect 10643 16065 10655 16068
rect 10597 16059 10655 16065
rect 11517 16065 11529 16068
rect 11563 16065 11575 16099
rect 11517 16059 11575 16065
rect 13357 16099 13415 16105
rect 13357 16065 13369 16099
rect 13403 16096 13415 16099
rect 13446 16096 13452 16108
rect 13403 16068 13452 16096
rect 13403 16065 13415 16068
rect 13357 16059 13415 16065
rect 13446 16056 13452 16068
rect 13504 16056 13510 16108
rect 14277 16099 14335 16105
rect 14277 16065 14289 16099
rect 14323 16096 14335 16099
rect 14366 16096 14372 16108
rect 14323 16068 14372 16096
rect 14323 16065 14335 16068
rect 14277 16059 14335 16065
rect 14366 16056 14372 16068
rect 14424 16056 14430 16108
rect 14550 16096 14556 16108
rect 14511 16068 14556 16096
rect 14550 16056 14556 16068
rect 14608 16056 14614 16108
rect 16298 16096 16304 16108
rect 16259 16068 16304 16096
rect 16298 16056 16304 16068
rect 16356 16056 16362 16108
rect 17310 16096 17316 16108
rect 17271 16068 17316 16096
rect 17310 16056 17316 16068
rect 17368 16056 17374 16108
rect 1578 15988 1584 16040
rect 1636 16028 1642 16040
rect 1762 16028 1768 16040
rect 1820 16037 1826 16040
rect 1820 16031 1858 16037
rect 1636 16000 1768 16028
rect 1636 15988 1642 16000
rect 1762 15988 1768 16000
rect 1846 16028 1858 16031
rect 2225 16031 2283 16037
rect 2225 16028 2237 16031
rect 1846 16000 2237 16028
rect 1846 15997 1858 16000
rect 1820 15991 1858 15997
rect 2225 15997 2237 16000
rect 2271 15997 2283 16031
rect 2225 15991 2283 15997
rect 8665 16031 8723 16037
rect 8665 15997 8677 16031
rect 8711 16028 8723 16031
rect 8846 16028 8852 16040
rect 8711 16000 8852 16028
rect 8711 15997 8723 16000
rect 8665 15991 8723 15997
rect 1820 15988 1826 15991
rect 8846 15988 8852 16000
rect 8904 15988 8910 16040
rect 12710 15988 12716 16040
rect 12768 16028 12774 16040
rect 13078 16028 13084 16040
rect 12768 16000 12813 16028
rect 13039 16000 13084 16028
rect 12768 15988 12774 16000
rect 13078 15988 13084 16000
rect 13136 15988 13142 16040
rect 15746 16028 15752 16040
rect 15707 16000 15752 16028
rect 15746 15988 15752 16000
rect 15804 15988 15810 16040
rect 16206 16028 16212 16040
rect 16119 16000 16212 16028
rect 16206 15988 16212 16000
rect 16264 16028 16270 16040
rect 16761 16031 16819 16037
rect 16761 16028 16773 16031
rect 16264 16000 16773 16028
rect 16264 15988 16270 16000
rect 16761 15997 16773 16000
rect 16807 15997 16819 16031
rect 16761 15991 16819 15997
rect 18046 15988 18052 16040
rect 18104 16037 18110 16040
rect 18104 16031 18142 16037
rect 18130 16028 18142 16031
rect 18509 16031 18567 16037
rect 18509 16028 18521 16031
rect 18130 16000 18521 16028
rect 18130 15997 18142 16000
rect 18104 15991 18142 15997
rect 18509 15997 18521 16000
rect 18555 15997 18567 16031
rect 18509 15991 18567 15997
rect 18104 15988 18110 15991
rect 18598 15988 18604 16040
rect 18656 16028 18662 16040
rect 19128 16031 19186 16037
rect 19128 16028 19140 16031
rect 18656 16000 19140 16028
rect 18656 15988 18662 16000
rect 19128 15997 19140 16000
rect 19174 16028 19186 16031
rect 19521 16031 19579 16037
rect 19521 16028 19533 16031
rect 19174 16000 19533 16028
rect 19174 15997 19186 16000
rect 19128 15991 19186 15997
rect 19521 15997 19533 16000
rect 19567 15997 19579 16031
rect 19521 15991 19579 15997
rect 2866 15960 2872 15972
rect 2827 15932 2872 15960
rect 2866 15920 2872 15932
rect 2924 15920 2930 15972
rect 2961 15963 3019 15969
rect 2961 15929 2973 15963
rect 3007 15960 3019 15963
rect 3234 15960 3240 15972
rect 3007 15932 3240 15960
rect 3007 15929 3019 15932
rect 2961 15923 3019 15929
rect 2685 15895 2743 15901
rect 2685 15861 2697 15895
rect 2731 15892 2743 15895
rect 2976 15892 3004 15923
rect 3234 15920 3240 15932
rect 3292 15920 3298 15972
rect 4154 15920 4160 15972
rect 4212 15960 4218 15972
rect 4525 15963 4583 15969
rect 4525 15960 4537 15963
rect 4212 15932 4537 15960
rect 4212 15920 4218 15932
rect 4525 15929 4537 15932
rect 4571 15960 4583 15963
rect 5074 15960 5080 15972
rect 4571 15932 5080 15960
rect 4571 15929 4583 15932
rect 4525 15923 4583 15929
rect 5074 15920 5080 15932
rect 5132 15920 5138 15972
rect 6273 15963 6331 15969
rect 6273 15929 6285 15963
rect 6319 15960 6331 15963
rect 6822 15960 6828 15972
rect 6319 15932 6828 15960
rect 6319 15929 6331 15932
rect 6273 15923 6331 15929
rect 6822 15920 6828 15932
rect 6880 15920 6886 15972
rect 7006 15960 7012 15972
rect 6932 15932 7012 15960
rect 2731 15864 3004 15892
rect 2731 15861 2743 15864
rect 2685 15855 2743 15861
rect 6086 15852 6092 15904
rect 6144 15892 6150 15904
rect 6549 15895 6607 15901
rect 6549 15892 6561 15895
rect 6144 15864 6561 15892
rect 6144 15852 6150 15864
rect 6549 15861 6561 15864
rect 6595 15892 6607 15895
rect 6932 15892 6960 15932
rect 7006 15920 7012 15932
rect 7064 15920 7070 15972
rect 7098 15920 7104 15972
rect 7156 15960 7162 15972
rect 7156 15932 7201 15960
rect 7156 15920 7162 15932
rect 7282 15920 7288 15972
rect 7340 15960 7346 15972
rect 7653 15963 7711 15969
rect 7653 15960 7665 15963
rect 7340 15932 7665 15960
rect 7340 15920 7346 15932
rect 7653 15929 7665 15932
rect 7699 15929 7711 15963
rect 9490 15960 9496 15972
rect 9451 15932 9496 15960
rect 7653 15923 7711 15929
rect 9490 15920 9496 15932
rect 9548 15920 9554 15972
rect 10045 15963 10103 15969
rect 10045 15929 10057 15963
rect 10091 15960 10103 15963
rect 10689 15963 10747 15969
rect 10689 15960 10701 15963
rect 10091 15932 10701 15960
rect 10091 15929 10103 15932
rect 10045 15923 10103 15929
rect 10689 15929 10701 15932
rect 10735 15960 10747 15963
rect 10870 15960 10876 15972
rect 10735 15932 10876 15960
rect 10735 15929 10747 15932
rect 10689 15923 10747 15929
rect 10870 15920 10876 15932
rect 10928 15920 10934 15972
rect 14369 15963 14427 15969
rect 14369 15929 14381 15963
rect 14415 15929 14427 15963
rect 16224 15960 16252 15988
rect 14369 15923 14427 15929
rect 15304 15932 16252 15960
rect 13630 15892 13636 15904
rect 6595 15864 6960 15892
rect 13591 15864 13636 15892
rect 6595 15861 6607 15864
rect 6549 15855 6607 15861
rect 13630 15852 13636 15864
rect 13688 15852 13694 15904
rect 13998 15892 14004 15904
rect 13959 15864 14004 15892
rect 13998 15852 14004 15864
rect 14056 15892 14062 15904
rect 14384 15892 14412 15923
rect 15304 15904 15332 15932
rect 15286 15892 15292 15904
rect 14056 15864 14412 15892
rect 15247 15864 15292 15892
rect 14056 15852 14062 15864
rect 15286 15852 15292 15864
rect 15344 15852 15350 15904
rect 15654 15892 15660 15904
rect 15615 15864 15660 15892
rect 15654 15852 15660 15864
rect 15712 15852 15718 15904
rect 18138 15852 18144 15904
rect 18196 15901 18202 15904
rect 18196 15895 18245 15901
rect 18196 15861 18199 15895
rect 18233 15861 18245 15895
rect 18196 15855 18245 15861
rect 18196 15852 18202 15855
rect 18966 15852 18972 15904
rect 19024 15892 19030 15904
rect 19199 15895 19257 15901
rect 19199 15892 19211 15895
rect 19024 15864 19211 15892
rect 19024 15852 19030 15864
rect 19199 15861 19211 15864
rect 19245 15861 19257 15895
rect 19199 15855 19257 15861
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 2130 15688 2136 15700
rect 2091 15660 2136 15688
rect 2130 15648 2136 15660
rect 2188 15648 2194 15700
rect 2866 15648 2872 15700
rect 2924 15688 2930 15700
rect 3513 15691 3571 15697
rect 3513 15688 3525 15691
rect 2924 15660 3525 15688
rect 2924 15648 2930 15660
rect 3513 15657 3525 15660
rect 3559 15688 3571 15691
rect 4338 15688 4344 15700
rect 3559 15660 4344 15688
rect 3559 15657 3571 15660
rect 3513 15651 3571 15657
rect 4338 15648 4344 15660
rect 4396 15648 4402 15700
rect 5074 15688 5080 15700
rect 5035 15660 5080 15688
rect 5074 15648 5080 15660
rect 5132 15648 5138 15700
rect 10686 15688 10692 15700
rect 10647 15660 10692 15688
rect 10686 15648 10692 15660
rect 10744 15688 10750 15700
rect 11333 15691 11391 15697
rect 11333 15688 11345 15691
rect 10744 15660 11345 15688
rect 10744 15648 10750 15660
rect 11333 15657 11345 15660
rect 11379 15657 11391 15691
rect 11333 15651 11391 15657
rect 12989 15691 13047 15697
rect 12989 15657 13001 15691
rect 13035 15688 13047 15691
rect 13078 15688 13084 15700
rect 13035 15660 13084 15688
rect 13035 15657 13047 15660
rect 12989 15651 13047 15657
rect 13078 15648 13084 15660
rect 13136 15648 13142 15700
rect 15746 15688 15752 15700
rect 15707 15660 15752 15688
rect 15746 15648 15752 15660
rect 15804 15688 15810 15700
rect 16022 15688 16028 15700
rect 15804 15660 16028 15688
rect 15804 15648 15810 15660
rect 16022 15648 16028 15660
rect 16080 15648 16086 15700
rect 2498 15620 2504 15632
rect 2459 15592 2504 15620
rect 2498 15580 2504 15592
rect 2556 15580 2562 15632
rect 2590 15580 2596 15632
rect 2648 15620 2654 15632
rect 3142 15620 3148 15632
rect 2648 15592 2693 15620
rect 3103 15592 3148 15620
rect 2648 15580 2654 15592
rect 3142 15580 3148 15592
rect 3200 15580 3206 15632
rect 3234 15580 3240 15632
rect 3292 15620 3298 15632
rect 4065 15623 4123 15629
rect 4065 15620 4077 15623
rect 3292 15592 4077 15620
rect 3292 15580 3298 15592
rect 4065 15589 4077 15592
rect 4111 15589 4123 15623
rect 6454 15620 6460 15632
rect 6415 15592 6460 15620
rect 4065 15583 4123 15589
rect 6454 15580 6460 15592
rect 6512 15580 6518 15632
rect 6546 15580 6552 15632
rect 6604 15620 6610 15632
rect 7929 15623 7987 15629
rect 7929 15620 7941 15623
rect 6604 15592 7941 15620
rect 6604 15580 6610 15592
rect 7929 15589 7941 15592
rect 7975 15589 7987 15623
rect 7929 15583 7987 15589
rect 9490 15580 9496 15632
rect 9548 15620 9554 15632
rect 9766 15620 9772 15632
rect 9548 15592 9772 15620
rect 9548 15580 9554 15592
rect 9766 15580 9772 15592
rect 9824 15620 9830 15632
rect 9861 15623 9919 15629
rect 9861 15620 9873 15623
rect 9824 15592 9873 15620
rect 9824 15580 9830 15592
rect 9861 15589 9873 15592
rect 9907 15589 9919 15623
rect 13814 15620 13820 15632
rect 13775 15592 13820 15620
rect 9861 15583 9919 15589
rect 13814 15580 13820 15592
rect 13872 15580 13878 15632
rect 14369 15623 14427 15629
rect 14369 15589 14381 15623
rect 14415 15620 14427 15623
rect 14550 15620 14556 15632
rect 14415 15592 14556 15620
rect 14415 15589 14427 15592
rect 14369 15583 14427 15589
rect 14550 15580 14556 15592
rect 14608 15580 14614 15632
rect 16571 15623 16629 15629
rect 16571 15589 16583 15623
rect 16617 15620 16629 15623
rect 16850 15620 16856 15632
rect 16617 15592 16856 15620
rect 16617 15589 16629 15592
rect 16571 15583 16629 15589
rect 16850 15580 16856 15592
rect 16908 15580 16914 15632
rect 17494 15620 17500 15632
rect 17144 15592 17500 15620
rect 1432 15555 1490 15561
rect 1432 15552 1444 15555
rect 1412 15521 1444 15552
rect 1478 15521 1490 15555
rect 4154 15552 4160 15564
rect 4115 15524 4160 15552
rect 1412 15515 1490 15521
rect 1412 15416 1440 15515
rect 4154 15512 4160 15524
rect 4212 15512 4218 15564
rect 7098 15512 7104 15564
rect 7156 15552 7162 15564
rect 7469 15555 7527 15561
rect 7469 15552 7481 15555
rect 7156 15524 7481 15552
rect 7156 15512 7162 15524
rect 7469 15521 7481 15524
rect 7515 15552 7527 15555
rect 7834 15552 7840 15564
rect 7515 15524 7840 15552
rect 7515 15521 7527 15524
rect 7469 15515 7527 15521
rect 7834 15512 7840 15524
rect 7892 15552 7898 15564
rect 8021 15555 8079 15561
rect 8021 15552 8033 15555
rect 7892 15524 8033 15552
rect 7892 15512 7898 15524
rect 8021 15521 8033 15524
rect 8067 15521 8079 15555
rect 11238 15552 11244 15564
rect 11199 15524 11244 15552
rect 8021 15515 8079 15521
rect 11238 15512 11244 15524
rect 11296 15512 11302 15564
rect 11790 15552 11796 15564
rect 11751 15524 11796 15552
rect 11790 15512 11796 15524
rect 11848 15512 11854 15564
rect 17144 15561 17172 15592
rect 17494 15580 17500 15592
rect 17552 15620 17558 15632
rect 18141 15623 18199 15629
rect 18141 15620 18153 15623
rect 17552 15592 18153 15620
rect 17552 15580 17558 15592
rect 18141 15589 18153 15592
rect 18187 15589 18199 15623
rect 18141 15583 18199 15589
rect 17129 15555 17187 15561
rect 17129 15521 17141 15555
rect 17175 15521 17187 15555
rect 17129 15515 17187 15521
rect 8938 15444 8944 15496
rect 8996 15484 9002 15496
rect 9398 15484 9404 15496
rect 8996 15456 9404 15484
rect 8996 15444 9002 15456
rect 9398 15444 9404 15456
rect 9456 15484 9462 15496
rect 9769 15487 9827 15493
rect 9769 15484 9781 15487
rect 9456 15456 9781 15484
rect 9456 15444 9462 15456
rect 9769 15453 9781 15456
rect 9815 15453 9827 15487
rect 10042 15484 10048 15496
rect 10003 15456 10048 15484
rect 9769 15447 9827 15453
rect 10042 15444 10048 15456
rect 10100 15444 10106 15496
rect 13722 15484 13728 15496
rect 13683 15456 13728 15484
rect 13722 15444 13728 15456
rect 13780 15444 13786 15496
rect 16209 15487 16267 15493
rect 16209 15453 16221 15487
rect 16255 15484 16267 15487
rect 16482 15484 16488 15496
rect 16255 15456 16488 15484
rect 16255 15453 16267 15456
rect 16209 15447 16267 15453
rect 16482 15444 16488 15456
rect 16540 15444 16546 15496
rect 18046 15484 18052 15496
rect 18007 15456 18052 15484
rect 18046 15444 18052 15456
rect 18104 15444 18110 15496
rect 18325 15487 18383 15493
rect 18325 15453 18337 15487
rect 18371 15453 18383 15487
rect 18325 15447 18383 15453
rect 2038 15416 2044 15428
rect 1412 15388 2044 15416
rect 2038 15376 2044 15388
rect 2096 15416 2102 15428
rect 3142 15416 3148 15428
rect 2096 15388 3148 15416
rect 2096 15376 2102 15388
rect 3142 15376 3148 15388
rect 3200 15376 3206 15428
rect 7009 15419 7067 15425
rect 7009 15385 7021 15419
rect 7055 15416 7067 15419
rect 7282 15416 7288 15428
rect 7055 15388 7288 15416
rect 7055 15385 7067 15388
rect 7009 15379 7067 15385
rect 7282 15376 7288 15388
rect 7340 15376 7346 15428
rect 17954 15376 17960 15428
rect 18012 15416 18018 15428
rect 18340 15416 18368 15447
rect 18012 15388 18368 15416
rect 18012 15376 18018 15388
rect 1535 15351 1593 15357
rect 1535 15317 1547 15351
rect 1581 15348 1593 15351
rect 2406 15348 2412 15360
rect 1581 15320 2412 15348
rect 1581 15317 1593 15320
rect 1535 15311 1593 15317
rect 2406 15308 2412 15320
rect 2464 15308 2470 15360
rect 7837 15351 7895 15357
rect 7837 15317 7849 15351
rect 7883 15348 7895 15351
rect 8110 15348 8116 15360
rect 7883 15320 8116 15348
rect 7883 15317 7895 15320
rect 7837 15311 7895 15317
rect 8110 15308 8116 15320
rect 8168 15308 8174 15360
rect 13170 15308 13176 15360
rect 13228 15348 13234 15360
rect 13357 15351 13415 15357
rect 13357 15348 13369 15351
rect 13228 15320 13369 15348
rect 13228 15308 13234 15320
rect 13357 15317 13369 15320
rect 13403 15317 13415 15351
rect 13357 15311 13415 15317
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 2041 15147 2099 15153
rect 2041 15113 2053 15147
rect 2087 15144 2099 15147
rect 2590 15144 2596 15156
rect 2087 15116 2596 15144
rect 2087 15113 2099 15116
rect 2041 15107 2099 15113
rect 2590 15104 2596 15116
rect 2648 15144 2654 15156
rect 4154 15144 4160 15156
rect 2648 15116 4160 15144
rect 2648 15104 2654 15116
rect 4154 15104 4160 15116
rect 4212 15104 4218 15156
rect 6273 15147 6331 15153
rect 6273 15113 6285 15147
rect 6319 15144 6331 15147
rect 6546 15144 6552 15156
rect 6319 15116 6552 15144
rect 6319 15113 6331 15116
rect 6273 15107 6331 15113
rect 6546 15104 6552 15116
rect 6604 15104 6610 15156
rect 7745 15147 7803 15153
rect 7745 15113 7757 15147
rect 7791 15144 7803 15147
rect 7834 15144 7840 15156
rect 7791 15116 7840 15144
rect 7791 15113 7803 15116
rect 7745 15107 7803 15113
rect 7834 15104 7840 15116
rect 7892 15104 7898 15156
rect 8846 15104 8852 15156
rect 8904 15144 8910 15156
rect 9493 15147 9551 15153
rect 9493 15144 9505 15147
rect 8904 15116 9505 15144
rect 8904 15104 8910 15116
rect 9493 15113 9505 15116
rect 9539 15113 9551 15147
rect 9766 15144 9772 15156
rect 9727 15116 9772 15144
rect 9493 15107 9551 15113
rect 2774 15036 2780 15088
rect 2832 15076 2838 15088
rect 3789 15079 3847 15085
rect 3789 15076 3801 15079
rect 2832 15048 3801 15076
rect 2832 15036 2838 15048
rect 3789 15045 3801 15048
rect 3835 15076 3847 15079
rect 4062 15076 4068 15088
rect 3835 15048 4068 15076
rect 3835 15045 3847 15048
rect 3789 15039 3847 15045
rect 4062 15036 4068 15048
rect 4120 15036 4126 15088
rect 9508 15076 9536 15107
rect 9766 15104 9772 15116
rect 9824 15104 9830 15156
rect 11790 15144 11796 15156
rect 11751 15116 11796 15144
rect 11790 15104 11796 15116
rect 11848 15104 11854 15156
rect 13265 15147 13323 15153
rect 13265 15113 13277 15147
rect 13311 15144 13323 15147
rect 13354 15144 13360 15156
rect 13311 15116 13360 15144
rect 13311 15113 13323 15116
rect 13265 15107 13323 15113
rect 13354 15104 13360 15116
rect 13412 15104 13418 15156
rect 14642 15144 14648 15156
rect 14603 15116 14648 15144
rect 14642 15104 14648 15116
rect 14700 15104 14706 15156
rect 15286 15144 15292 15156
rect 15247 15116 15292 15144
rect 15286 15104 15292 15116
rect 15344 15104 15350 15156
rect 17494 15144 17500 15156
rect 17455 15116 17500 15144
rect 17494 15104 17500 15116
rect 17552 15104 17558 15156
rect 18046 15104 18052 15156
rect 18104 15144 18110 15156
rect 19061 15147 19119 15153
rect 19061 15144 19073 15147
rect 18104 15116 19073 15144
rect 18104 15104 18110 15116
rect 19061 15113 19073 15116
rect 19107 15113 19119 15147
rect 19061 15107 19119 15113
rect 10137 15079 10195 15085
rect 10137 15076 10149 15079
rect 9508 15048 10149 15076
rect 10137 15045 10149 15048
rect 10183 15076 10195 15079
rect 10502 15076 10508 15088
rect 10183 15048 10508 15076
rect 10183 15045 10195 15048
rect 10137 15039 10195 15045
rect 10502 15036 10508 15048
rect 10560 15036 10566 15088
rect 12897 15079 12955 15085
rect 12897 15045 12909 15079
rect 12943 15076 12955 15079
rect 13814 15076 13820 15088
rect 12943 15048 13820 15076
rect 12943 15045 12955 15048
rect 12897 15039 12955 15045
rect 13814 15036 13820 15048
rect 13872 15076 13878 15088
rect 14277 15079 14335 15085
rect 14277 15076 14289 15079
rect 13872 15048 14289 15076
rect 13872 15036 13878 15048
rect 14277 15045 14289 15048
rect 14323 15076 14335 15079
rect 15470 15076 15476 15088
rect 14323 15048 15476 15076
rect 14323 15045 14335 15048
rect 14277 15039 14335 15045
rect 15470 15036 15476 15048
rect 15528 15036 15534 15088
rect 2958 15008 2964 15020
rect 2148 14980 2964 15008
rect 1556 14943 1614 14949
rect 1556 14909 1568 14943
rect 1602 14940 1614 14943
rect 2148 14940 2176 14980
rect 2958 14968 2964 14980
rect 3016 15008 3022 15020
rect 3970 15008 3976 15020
rect 3016 14980 3976 15008
rect 3016 14968 3022 14980
rect 3970 14968 3976 14980
rect 4028 14968 4034 15020
rect 5258 14968 5264 15020
rect 5316 15008 5322 15020
rect 6086 15008 6092 15020
rect 5316 14980 6092 15008
rect 5316 14968 5322 14980
rect 6086 14968 6092 14980
rect 6144 15008 6150 15020
rect 6549 15011 6607 15017
rect 6549 15008 6561 15011
rect 6144 14980 6561 15008
rect 6144 14968 6150 14980
rect 6549 14977 6561 14980
rect 6595 14977 6607 15011
rect 6549 14971 6607 14977
rect 6825 15011 6883 15017
rect 6825 14977 6837 15011
rect 6871 15008 6883 15011
rect 7098 15008 7104 15020
rect 6871 14980 7104 15008
rect 6871 14977 6883 14980
rect 6825 14971 6883 14977
rect 1602 14912 2176 14940
rect 2409 14943 2467 14949
rect 1602 14909 1614 14912
rect 1556 14903 1614 14909
rect 2409 14909 2421 14943
rect 2455 14940 2467 14943
rect 2869 14943 2927 14949
rect 2869 14940 2881 14943
rect 2455 14912 2881 14940
rect 2455 14909 2467 14912
rect 2409 14903 2467 14909
rect 2869 14909 2881 14912
rect 2915 14940 2927 14943
rect 3050 14940 3056 14952
rect 2915 14912 3056 14940
rect 2915 14909 2927 14912
rect 2869 14903 2927 14909
rect 3050 14900 3056 14912
rect 3108 14900 3114 14952
rect 3190 14875 3248 14881
rect 3190 14872 3202 14875
rect 2884 14844 3202 14872
rect 2884 14816 2912 14844
rect 3190 14841 3202 14844
rect 3236 14841 3248 14875
rect 5261 14875 5319 14881
rect 5261 14872 5273 14875
rect 3190 14835 3248 14841
rect 4632 14844 5273 14872
rect 4632 14816 4660 14844
rect 5261 14841 5273 14844
rect 5307 14841 5319 14875
rect 5261 14835 5319 14841
rect 5350 14832 5356 14884
rect 5408 14872 5414 14884
rect 5905 14875 5963 14881
rect 5408 14844 5453 14872
rect 5408 14832 5414 14844
rect 5905 14841 5917 14875
rect 5951 14872 5963 14875
rect 5994 14872 6000 14884
rect 5951 14844 6000 14872
rect 5951 14841 5963 14844
rect 5905 14835 5963 14841
rect 5994 14832 6000 14844
rect 6052 14832 6058 14884
rect 6564 14872 6592 14971
rect 7098 14968 7104 14980
rect 7156 14968 7162 15020
rect 10042 14968 10048 15020
rect 10100 15008 10106 15020
rect 10689 15011 10747 15017
rect 10689 15008 10701 15011
rect 10100 14980 10701 15008
rect 10100 14968 10106 14980
rect 10689 14977 10701 14980
rect 10735 14977 10747 15011
rect 18138 15008 18144 15020
rect 18099 14980 18144 15008
rect 10689 14971 10747 14977
rect 18138 14968 18144 14980
rect 18196 14968 18202 15020
rect 8113 14943 8171 14949
rect 8113 14909 8125 14943
rect 8159 14940 8171 14943
rect 8573 14943 8631 14949
rect 8573 14940 8585 14943
rect 8159 14912 8585 14940
rect 8159 14909 8171 14912
rect 8113 14903 8171 14909
rect 8573 14909 8585 14912
rect 8619 14940 8631 14943
rect 9582 14940 9588 14952
rect 8619 14912 9588 14940
rect 8619 14909 8631 14912
rect 8573 14903 8631 14909
rect 9582 14900 9588 14912
rect 9640 14900 9646 14952
rect 13170 14900 13176 14952
rect 13228 14940 13234 14952
rect 13357 14943 13415 14949
rect 13357 14940 13369 14943
rect 13228 14912 13369 14940
rect 13228 14900 13234 14912
rect 13357 14909 13369 14912
rect 13403 14909 13415 14943
rect 15105 14943 15163 14949
rect 15105 14940 15117 14943
rect 13357 14903 13415 14909
rect 14936 14912 15117 14940
rect 7146 14875 7204 14881
rect 7146 14872 7158 14875
rect 6564 14844 7158 14872
rect 7146 14841 7158 14844
rect 7192 14872 7204 14875
rect 8389 14875 8447 14881
rect 8389 14872 8401 14875
rect 7192 14844 8401 14872
rect 7192 14841 7204 14844
rect 7146 14835 7204 14841
rect 8389 14841 8401 14844
rect 8435 14872 8447 14875
rect 8478 14872 8484 14884
rect 8435 14844 8484 14872
rect 8435 14841 8447 14844
rect 8389 14835 8447 14841
rect 8478 14832 8484 14844
rect 8536 14872 8542 14884
rect 8894 14875 8952 14881
rect 8894 14872 8906 14875
rect 8536 14844 8906 14872
rect 8536 14832 8542 14844
rect 8894 14841 8906 14844
rect 8940 14841 8952 14875
rect 10410 14872 10416 14884
rect 10371 14844 10416 14872
rect 8894 14835 8952 14841
rect 10410 14832 10416 14844
rect 10468 14832 10474 14884
rect 10502 14832 10508 14884
rect 10560 14872 10566 14884
rect 10560 14844 10605 14872
rect 10560 14832 10566 14844
rect 13446 14832 13452 14884
rect 13504 14872 13510 14884
rect 13678 14875 13736 14881
rect 13678 14872 13690 14875
rect 13504 14844 13690 14872
rect 13504 14832 13510 14844
rect 13678 14841 13690 14844
rect 13724 14841 13736 14875
rect 13678 14835 13736 14841
rect 1394 14764 1400 14816
rect 1452 14804 1458 14816
rect 1627 14807 1685 14813
rect 1627 14804 1639 14807
rect 1452 14776 1639 14804
rect 1452 14764 1458 14776
rect 1627 14773 1639 14776
rect 1673 14804 1685 14807
rect 2682 14804 2688 14816
rect 1673 14776 2688 14804
rect 1673 14773 1685 14776
rect 1627 14767 1685 14773
rect 2682 14764 2688 14776
rect 2740 14764 2746 14816
rect 2777 14807 2835 14813
rect 2777 14773 2789 14807
rect 2823 14804 2835 14807
rect 2866 14804 2872 14816
rect 2823 14776 2872 14804
rect 2823 14773 2835 14776
rect 2777 14767 2835 14773
rect 2866 14764 2872 14776
rect 2924 14764 2930 14816
rect 4614 14804 4620 14816
rect 4575 14776 4620 14804
rect 4614 14764 4620 14776
rect 4672 14764 4678 14816
rect 5077 14807 5135 14813
rect 5077 14773 5089 14807
rect 5123 14804 5135 14807
rect 5368 14804 5396 14832
rect 5123 14776 5396 14804
rect 10428 14804 10456 14832
rect 10686 14804 10692 14816
rect 10428 14776 10692 14804
rect 5123 14773 5135 14776
rect 5077 14767 5135 14773
rect 10686 14764 10692 14776
rect 10744 14764 10750 14816
rect 10778 14764 10784 14816
rect 10836 14804 10842 14816
rect 11238 14804 11244 14816
rect 10836 14776 11244 14804
rect 10836 14764 10842 14776
rect 11238 14764 11244 14776
rect 11296 14804 11302 14816
rect 11333 14807 11391 14813
rect 11333 14804 11345 14807
rect 11296 14776 11345 14804
rect 11296 14764 11302 14776
rect 11333 14773 11345 14776
rect 11379 14773 11391 14807
rect 11333 14767 11391 14773
rect 14826 14764 14832 14816
rect 14884 14804 14890 14816
rect 14936 14813 14964 14912
rect 15105 14909 15117 14912
rect 15151 14909 15163 14943
rect 16206 14940 16212 14952
rect 16167 14912 16212 14940
rect 15105 14903 15163 14909
rect 16206 14900 16212 14912
rect 16264 14900 16270 14952
rect 15749 14875 15807 14881
rect 15749 14841 15761 14875
rect 15795 14872 15807 14875
rect 16117 14875 16175 14881
rect 16117 14872 16129 14875
rect 15795 14844 16129 14872
rect 15795 14841 15807 14844
rect 15749 14835 15807 14841
rect 16117 14841 16129 14844
rect 16163 14872 16175 14875
rect 16571 14875 16629 14881
rect 16571 14872 16583 14875
rect 16163 14844 16583 14872
rect 16163 14841 16175 14844
rect 16117 14835 16175 14841
rect 16571 14841 16583 14844
rect 16617 14872 16629 14875
rect 16850 14872 16856 14884
rect 16617 14844 16856 14872
rect 16617 14841 16629 14844
rect 16571 14835 16629 14841
rect 16850 14832 16856 14844
rect 16908 14832 16914 14884
rect 18233 14875 18291 14881
rect 18233 14872 18245 14875
rect 17788 14844 18245 14872
rect 14921 14807 14979 14813
rect 14921 14804 14933 14807
rect 14884 14776 14933 14804
rect 14884 14764 14890 14776
rect 14921 14773 14933 14776
rect 14967 14773 14979 14807
rect 14921 14767 14979 14773
rect 17129 14807 17187 14813
rect 17129 14773 17141 14807
rect 17175 14804 17187 14807
rect 17310 14804 17316 14816
rect 17175 14776 17316 14804
rect 17175 14773 17187 14776
rect 17129 14767 17187 14773
rect 17310 14764 17316 14776
rect 17368 14804 17374 14816
rect 17788 14813 17816 14844
rect 18233 14841 18245 14844
rect 18279 14841 18291 14875
rect 18782 14872 18788 14884
rect 18743 14844 18788 14872
rect 18233 14835 18291 14841
rect 18782 14832 18788 14844
rect 18840 14832 18846 14884
rect 17773 14807 17831 14813
rect 17773 14804 17785 14807
rect 17368 14776 17785 14804
rect 17368 14764 17374 14776
rect 17773 14773 17785 14776
rect 17819 14773 17831 14807
rect 17773 14767 17831 14773
rect 19334 14764 19340 14816
rect 19392 14804 19398 14816
rect 19613 14807 19671 14813
rect 19613 14804 19625 14807
rect 19392 14776 19625 14804
rect 19392 14764 19398 14776
rect 19613 14773 19625 14776
rect 19659 14773 19671 14807
rect 19613 14767 19671 14773
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 2038 14600 2044 14612
rect 1999 14572 2044 14600
rect 2038 14560 2044 14572
rect 2096 14560 2102 14612
rect 2498 14600 2504 14612
rect 2459 14572 2504 14600
rect 2498 14560 2504 14572
rect 2556 14560 2562 14612
rect 2682 14560 2688 14612
rect 2740 14600 2746 14612
rect 3421 14603 3479 14609
rect 3421 14600 3433 14603
rect 2740 14572 3433 14600
rect 2740 14560 2746 14572
rect 3421 14569 3433 14572
rect 3467 14569 3479 14603
rect 3421 14563 3479 14569
rect 6454 14560 6460 14612
rect 6512 14600 6518 14612
rect 6549 14603 6607 14609
rect 6549 14600 6561 14603
rect 6512 14572 6561 14600
rect 6512 14560 6518 14572
rect 6549 14569 6561 14572
rect 6595 14569 6607 14603
rect 7834 14600 7840 14612
rect 7795 14572 7840 14600
rect 6549 14563 6607 14569
rect 7834 14560 7840 14572
rect 7892 14560 7898 14612
rect 9398 14600 9404 14612
rect 9359 14572 9404 14600
rect 9398 14560 9404 14572
rect 9456 14560 9462 14612
rect 10686 14600 10692 14612
rect 10647 14572 10692 14600
rect 10686 14560 10692 14572
rect 10744 14560 10750 14612
rect 16206 14560 16212 14612
rect 16264 14600 16270 14612
rect 16393 14603 16451 14609
rect 16393 14600 16405 14603
rect 16264 14572 16405 14600
rect 16264 14560 16270 14572
rect 16393 14569 16405 14572
rect 16439 14600 16451 14603
rect 16439 14572 18000 14600
rect 16439 14569 16451 14572
rect 16393 14563 16451 14569
rect 2869 14535 2927 14541
rect 2869 14501 2881 14535
rect 2915 14532 2927 14535
rect 2958 14532 2964 14544
rect 2915 14504 2964 14532
rect 2915 14501 2927 14504
rect 2869 14495 2927 14501
rect 2958 14492 2964 14504
rect 3016 14492 3022 14544
rect 5721 14535 5779 14541
rect 5721 14501 5733 14535
rect 5767 14532 5779 14535
rect 6270 14532 6276 14544
rect 5767 14504 6276 14532
rect 5767 14501 5779 14504
rect 5721 14495 5779 14501
rect 6270 14492 6276 14504
rect 6328 14492 6334 14544
rect 8110 14532 8116 14544
rect 8071 14504 8116 14532
rect 8110 14492 8116 14504
rect 8168 14492 8174 14544
rect 8202 14492 8208 14544
rect 8260 14532 8266 14544
rect 9861 14535 9919 14541
rect 8260 14504 8305 14532
rect 8260 14492 8266 14504
rect 9861 14501 9873 14535
rect 9907 14532 9919 14535
rect 9950 14532 9956 14544
rect 9907 14504 9956 14532
rect 9907 14501 9919 14504
rect 9861 14495 9919 14501
rect 9950 14492 9956 14504
rect 10008 14492 10014 14544
rect 13354 14541 13360 14544
rect 13351 14532 13360 14541
rect 13315 14504 13360 14532
rect 13351 14495 13360 14504
rect 13354 14492 13360 14495
rect 13412 14492 13418 14544
rect 15470 14532 15476 14544
rect 15431 14504 15476 14532
rect 15470 14492 15476 14504
rect 15528 14492 15534 14544
rect 17310 14532 17316 14544
rect 17271 14504 17316 14532
rect 17310 14492 17316 14504
rect 17368 14492 17374 14544
rect 17972 14532 18000 14572
rect 18138 14560 18144 14612
rect 18196 14600 18202 14612
rect 18509 14603 18567 14609
rect 18509 14600 18521 14603
rect 18196 14572 18521 14600
rect 18196 14560 18202 14572
rect 18509 14569 18521 14572
rect 18555 14569 18567 14603
rect 18509 14563 18567 14569
rect 18785 14603 18843 14609
rect 18785 14569 18797 14603
rect 18831 14569 18843 14603
rect 18785 14563 18843 14569
rect 18800 14532 18828 14563
rect 17972 14504 18828 14532
rect 1540 14467 1598 14473
rect 1540 14433 1552 14467
rect 1586 14464 1598 14467
rect 2038 14464 2044 14476
rect 1586 14436 2044 14464
rect 1586 14433 1598 14436
rect 1540 14427 1598 14433
rect 2038 14424 2044 14436
rect 2096 14424 2102 14476
rect 4522 14464 4528 14476
rect 4483 14436 4528 14464
rect 4522 14424 4528 14436
rect 4580 14424 4586 14476
rect 11698 14464 11704 14476
rect 11659 14436 11704 14464
rect 11698 14424 11704 14436
rect 11756 14424 11762 14476
rect 11885 14467 11943 14473
rect 11885 14433 11897 14467
rect 11931 14464 11943 14467
rect 12894 14464 12900 14476
rect 11931 14436 12900 14464
rect 11931 14433 11943 14436
rect 11885 14427 11943 14433
rect 1627 14399 1685 14405
rect 1627 14365 1639 14399
rect 1673 14396 1685 14399
rect 1946 14396 1952 14408
rect 1673 14368 1952 14396
rect 1673 14365 1685 14368
rect 1627 14359 1685 14365
rect 1946 14356 1952 14368
rect 2004 14356 2010 14408
rect 2958 14396 2964 14408
rect 2919 14368 2964 14396
rect 2958 14356 2964 14368
rect 3016 14356 3022 14408
rect 5629 14399 5687 14405
rect 5629 14396 5641 14399
rect 5552 14368 5641 14396
rect 5552 14272 5580 14368
rect 5629 14365 5641 14368
rect 5675 14365 5687 14399
rect 5994 14396 6000 14408
rect 5955 14368 6000 14396
rect 5629 14359 5687 14365
rect 5994 14356 6000 14368
rect 6052 14356 6058 14408
rect 8386 14396 8392 14408
rect 8347 14368 8392 14396
rect 8386 14356 8392 14368
rect 8444 14356 8450 14408
rect 9766 14396 9772 14408
rect 9727 14368 9772 14396
rect 9766 14356 9772 14368
rect 9824 14356 9830 14408
rect 10045 14399 10103 14405
rect 10045 14365 10057 14399
rect 10091 14365 10103 14399
rect 10045 14359 10103 14365
rect 8404 14328 8432 14356
rect 10060 14328 10088 14359
rect 11422 14356 11428 14408
rect 11480 14396 11486 14408
rect 11900 14396 11928 14427
rect 12894 14424 12900 14436
rect 12952 14424 12958 14476
rect 17865 14467 17923 14473
rect 17865 14433 17877 14467
rect 17911 14464 17923 14467
rect 18046 14464 18052 14476
rect 17911 14436 18052 14464
rect 17911 14433 17923 14436
rect 17865 14427 17923 14433
rect 18046 14424 18052 14436
rect 18104 14424 18110 14476
rect 18693 14467 18751 14473
rect 18693 14433 18705 14467
rect 18739 14433 18751 14467
rect 19242 14464 19248 14476
rect 19203 14436 19248 14464
rect 18693 14427 18751 14433
rect 11480 14368 11928 14396
rect 12161 14399 12219 14405
rect 11480 14356 11486 14368
rect 12161 14365 12173 14399
rect 12207 14396 12219 14399
rect 12986 14396 12992 14408
rect 12207 14368 12992 14396
rect 12207 14365 12219 14368
rect 12161 14359 12219 14365
rect 12986 14356 12992 14368
rect 13044 14356 13050 14408
rect 15381 14399 15439 14405
rect 15381 14365 15393 14399
rect 15427 14396 15439 14399
rect 15746 14396 15752 14408
rect 15427 14368 15752 14396
rect 15427 14365 15439 14368
rect 15381 14359 15439 14365
rect 15746 14356 15752 14368
rect 15804 14356 15810 14408
rect 16025 14399 16083 14405
rect 16025 14365 16037 14399
rect 16071 14396 16083 14399
rect 16298 14396 16304 14408
rect 16071 14368 16304 14396
rect 16071 14365 16083 14368
rect 16025 14359 16083 14365
rect 16298 14356 16304 14368
rect 16356 14356 16362 14408
rect 17218 14396 17224 14408
rect 17179 14368 17224 14396
rect 17218 14356 17224 14368
rect 17276 14356 17282 14408
rect 17586 14356 17592 14408
rect 17644 14396 17650 14408
rect 18708 14396 18736 14427
rect 19242 14424 19248 14436
rect 19300 14424 19306 14476
rect 19058 14396 19064 14408
rect 17644 14368 19064 14396
rect 17644 14356 17650 14368
rect 19058 14356 19064 14368
rect 19116 14356 19122 14408
rect 8404 14300 10088 14328
rect 4706 14260 4712 14272
rect 4667 14232 4712 14260
rect 4706 14220 4712 14232
rect 4764 14220 4770 14272
rect 5074 14260 5080 14272
rect 5035 14232 5080 14260
rect 5074 14220 5080 14232
rect 5132 14220 5138 14272
rect 5445 14263 5503 14269
rect 5445 14229 5457 14263
rect 5491 14260 5503 14263
rect 5534 14260 5540 14272
rect 5491 14232 5540 14260
rect 5491 14229 5503 14232
rect 5445 14223 5503 14229
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 6914 14260 6920 14272
rect 6875 14232 6920 14260
rect 6914 14220 6920 14232
rect 6972 14220 6978 14272
rect 7098 14220 7104 14272
rect 7156 14260 7162 14272
rect 7285 14263 7343 14269
rect 7285 14260 7297 14263
rect 7156 14232 7297 14260
rect 7156 14220 7162 14232
rect 7285 14229 7297 14232
rect 7331 14229 7343 14263
rect 9030 14260 9036 14272
rect 8991 14232 9036 14260
rect 7285 14223 7343 14229
rect 9030 14220 9036 14232
rect 9088 14220 9094 14272
rect 12529 14263 12587 14269
rect 12529 14229 12541 14263
rect 12575 14260 12587 14263
rect 12894 14260 12900 14272
rect 12575 14232 12900 14260
rect 12575 14229 12587 14232
rect 12529 14223 12587 14229
rect 12894 14220 12900 14232
rect 12952 14220 12958 14272
rect 13909 14263 13967 14269
rect 13909 14229 13921 14263
rect 13955 14260 13967 14263
rect 13998 14260 14004 14272
rect 13955 14232 14004 14260
rect 13955 14229 13967 14232
rect 13909 14223 13967 14229
rect 13998 14220 14004 14232
rect 14056 14220 14062 14272
rect 14182 14260 14188 14272
rect 14143 14232 14188 14260
rect 14182 14220 14188 14232
rect 14240 14220 14246 14272
rect 16574 14220 16580 14272
rect 16632 14260 16638 14272
rect 16669 14263 16727 14269
rect 16669 14260 16681 14263
rect 16632 14232 16681 14260
rect 16632 14220 16638 14232
rect 16669 14229 16681 14232
rect 16715 14229 16727 14263
rect 16669 14223 16727 14229
rect 18233 14263 18291 14269
rect 18233 14229 18245 14263
rect 18279 14260 18291 14263
rect 18322 14260 18328 14272
rect 18279 14232 18328 14260
rect 18279 14229 18291 14232
rect 18233 14223 18291 14229
rect 18322 14220 18328 14232
rect 18380 14220 18386 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 3881 14059 3939 14065
rect 3881 14025 3893 14059
rect 3927 14056 3939 14059
rect 4154 14056 4160 14068
rect 3927 14028 4160 14056
rect 3927 14025 3939 14028
rect 3881 14019 3939 14025
rect 4154 14016 4160 14028
rect 4212 14016 4218 14068
rect 5350 14016 5356 14068
rect 5408 14056 5414 14068
rect 5905 14059 5963 14065
rect 5905 14056 5917 14059
rect 5408 14028 5917 14056
rect 5408 14016 5414 14028
rect 5905 14025 5917 14028
rect 5951 14056 5963 14059
rect 6914 14056 6920 14068
rect 5951 14028 6920 14056
rect 5951 14025 5963 14028
rect 5905 14019 5963 14025
rect 6914 14016 6920 14028
rect 6972 14016 6978 14068
rect 8478 14056 8484 14068
rect 8439 14028 8484 14056
rect 8478 14016 8484 14028
rect 8536 14016 8542 14068
rect 9766 14016 9772 14068
rect 9824 14056 9830 14068
rect 10229 14059 10287 14065
rect 10229 14056 10241 14059
rect 9824 14028 10241 14056
rect 9824 14016 9830 14028
rect 10229 14025 10241 14028
rect 10275 14025 10287 14059
rect 10229 14019 10287 14025
rect 13354 14016 13360 14068
rect 13412 14056 13418 14068
rect 13449 14059 13507 14065
rect 13449 14056 13461 14059
rect 13412 14028 13461 14056
rect 13412 14016 13418 14028
rect 13449 14025 13461 14028
rect 13495 14025 13507 14059
rect 13998 14056 14004 14068
rect 13959 14028 14004 14056
rect 13449 14019 13507 14025
rect 13998 14016 14004 14028
rect 14056 14016 14062 14068
rect 17310 14016 17316 14068
rect 17368 14056 17374 14068
rect 17773 14059 17831 14065
rect 17773 14056 17785 14059
rect 17368 14028 17785 14056
rect 17368 14016 17374 14028
rect 17773 14025 17785 14028
rect 17819 14025 17831 14059
rect 19058 14056 19064 14068
rect 19019 14028 19064 14056
rect 17773 14019 17831 14025
rect 1578 13988 1584 14000
rect 1539 13960 1584 13988
rect 1578 13948 1584 13960
rect 1636 13948 1642 14000
rect 6270 13988 6276 14000
rect 6183 13960 6276 13988
rect 6270 13948 6276 13960
rect 6328 13988 6334 14000
rect 7101 13991 7159 13997
rect 7101 13988 7113 13991
rect 6328 13960 7113 13988
rect 6328 13948 6334 13960
rect 7101 13957 7113 13960
rect 7147 13957 7159 13991
rect 10594 13988 10600 14000
rect 10555 13960 10600 13988
rect 7101 13951 7159 13957
rect 10594 13948 10600 13960
rect 10652 13948 10658 14000
rect 15381 13991 15439 13997
rect 15381 13957 15393 13991
rect 15427 13988 15439 13991
rect 15470 13988 15476 14000
rect 15427 13960 15476 13988
rect 15427 13957 15439 13960
rect 15381 13951 15439 13957
rect 15470 13948 15476 13960
rect 15528 13988 15534 14000
rect 16758 13988 16764 14000
rect 15528 13960 16764 13988
rect 15528 13948 15534 13960
rect 16758 13948 16764 13960
rect 16816 13948 16822 14000
rect 17218 13948 17224 14000
rect 17276 13988 17282 14000
rect 17405 13991 17463 13997
rect 17405 13988 17417 13991
rect 17276 13960 17417 13988
rect 17276 13948 17282 13960
rect 17405 13957 17417 13960
rect 17451 13957 17463 13991
rect 17405 13951 17463 13957
rect 8662 13920 8668 13932
rect 8575 13892 8668 13920
rect 8662 13880 8668 13892
rect 8720 13920 8726 13932
rect 9030 13920 9036 13932
rect 8720 13892 9036 13920
rect 8720 13880 8726 13892
rect 9030 13880 9036 13892
rect 9088 13880 9094 13932
rect 1394 13852 1400 13864
rect 1355 13824 1400 13852
rect 1394 13812 1400 13824
rect 1452 13812 1458 13864
rect 2038 13852 2044 13864
rect 1999 13824 2044 13852
rect 2038 13812 2044 13824
rect 2096 13812 2102 13864
rect 2501 13855 2559 13861
rect 2501 13821 2513 13855
rect 2547 13852 2559 13855
rect 2961 13855 3019 13861
rect 2961 13852 2973 13855
rect 2547 13824 2973 13852
rect 2547 13821 2559 13824
rect 2501 13815 2559 13821
rect 2961 13821 2973 13824
rect 3007 13852 3019 13855
rect 4062 13852 4068 13864
rect 3007 13824 4068 13852
rect 3007 13821 3019 13824
rect 2961 13815 3019 13821
rect 4062 13812 4068 13824
rect 4120 13812 4126 13864
rect 4522 13852 4528 13864
rect 4483 13824 4528 13852
rect 4522 13812 4528 13824
rect 4580 13812 4586 13864
rect 4985 13855 5043 13861
rect 4985 13821 4997 13855
rect 5031 13852 5043 13855
rect 5074 13852 5080 13864
rect 5031 13824 5080 13852
rect 5031 13821 5043 13824
rect 4985 13815 5043 13821
rect 5074 13812 5080 13824
rect 5132 13852 5138 13864
rect 5132 13824 5488 13852
rect 5132 13812 5138 13824
rect 3282 13787 3340 13793
rect 3282 13784 3294 13787
rect 2884 13756 3294 13784
rect 2884 13728 2912 13756
rect 3282 13753 3294 13756
rect 3328 13784 3340 13787
rect 4801 13787 4859 13793
rect 4801 13784 4813 13787
rect 3328 13756 4813 13784
rect 3328 13753 3340 13756
rect 3282 13747 3340 13753
rect 4801 13753 4813 13756
rect 4847 13784 4859 13787
rect 5258 13784 5264 13796
rect 4847 13756 5264 13784
rect 4847 13753 4859 13756
rect 4801 13747 4859 13753
rect 5258 13744 5264 13756
rect 5316 13793 5322 13796
rect 5316 13787 5364 13793
rect 5316 13753 5318 13787
rect 5352 13753 5364 13787
rect 5460 13784 5488 13824
rect 6914 13812 6920 13864
rect 6972 13852 6978 13864
rect 8113 13855 8171 13861
rect 6972 13824 7017 13852
rect 6972 13812 6978 13824
rect 8113 13821 8125 13855
rect 8159 13852 8171 13855
rect 8202 13852 8208 13864
rect 8159 13824 8208 13852
rect 8159 13821 8171 13824
rect 8113 13815 8171 13821
rect 8202 13812 8208 13824
rect 8260 13852 8266 13864
rect 10612 13852 10640 13948
rect 10962 13880 10968 13932
rect 11020 13920 11026 13932
rect 11333 13923 11391 13929
rect 11333 13920 11345 13923
rect 11020 13892 11345 13920
rect 11020 13880 11026 13892
rect 11333 13889 11345 13892
rect 11379 13889 11391 13923
rect 13170 13920 13176 13932
rect 11333 13883 11391 13889
rect 12728 13892 13032 13920
rect 13131 13892 13176 13920
rect 10778 13852 10784 13864
rect 8260 13824 9628 13852
rect 10612 13824 10784 13852
rect 8260 13812 8266 13824
rect 5718 13784 5724 13796
rect 5460 13756 5724 13784
rect 5316 13747 5364 13753
rect 5316 13744 5322 13747
rect 5718 13744 5724 13756
rect 5776 13744 5782 13796
rect 8478 13744 8484 13796
rect 8536 13784 8542 13796
rect 8986 13787 9044 13793
rect 8986 13784 8998 13787
rect 8536 13756 8998 13784
rect 8536 13744 8542 13756
rect 8986 13753 8998 13756
rect 9032 13753 9044 13787
rect 8986 13747 9044 13753
rect 2866 13716 2872 13728
rect 2827 13688 2872 13716
rect 2866 13676 2872 13688
rect 2924 13676 2930 13728
rect 6641 13719 6699 13725
rect 6641 13685 6653 13719
rect 6687 13716 6699 13719
rect 6822 13716 6828 13728
rect 6687 13688 6828 13716
rect 6687 13685 6699 13688
rect 6641 13679 6699 13685
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 9600 13725 9628 13824
rect 10778 13812 10784 13824
rect 10836 13812 10842 13864
rect 10870 13812 10876 13864
rect 10928 13852 10934 13864
rect 11241 13855 11299 13861
rect 11241 13852 11253 13855
rect 10928 13824 11253 13852
rect 10928 13812 10934 13824
rect 11241 13821 11253 13824
rect 11287 13852 11299 13855
rect 11606 13852 11612 13864
rect 11287 13824 11612 13852
rect 11287 13821 11299 13824
rect 11241 13815 11299 13821
rect 11606 13812 11612 13824
rect 11664 13812 11670 13864
rect 11974 13812 11980 13864
rect 12032 13852 12038 13864
rect 12728 13861 12756 13892
rect 12253 13855 12311 13861
rect 12253 13852 12265 13855
rect 12032 13824 12265 13852
rect 12032 13812 12038 13824
rect 12253 13821 12265 13824
rect 12299 13852 12311 13855
rect 12713 13855 12771 13861
rect 12713 13852 12725 13855
rect 12299 13824 12725 13852
rect 12299 13821 12311 13824
rect 12253 13815 12311 13821
rect 12713 13821 12725 13824
rect 12759 13821 12771 13855
rect 12894 13852 12900 13864
rect 12855 13824 12900 13852
rect 12713 13815 12771 13821
rect 12894 13812 12900 13824
rect 12952 13812 12958 13864
rect 13004 13852 13032 13892
rect 13170 13880 13176 13892
rect 13228 13880 13234 13932
rect 14182 13920 14188 13932
rect 14143 13892 14188 13920
rect 14182 13880 14188 13892
rect 14240 13880 14246 13932
rect 15746 13920 15752 13932
rect 15707 13892 15752 13920
rect 15746 13880 15752 13892
rect 15804 13880 15810 13932
rect 16301 13923 16359 13929
rect 16301 13889 16313 13923
rect 16347 13920 16359 13923
rect 16574 13920 16580 13932
rect 16347 13892 16580 13920
rect 16347 13889 16359 13892
rect 16301 13883 16359 13889
rect 16574 13880 16580 13892
rect 16632 13880 16638 13932
rect 17126 13920 17132 13932
rect 17039 13892 17132 13920
rect 17126 13880 17132 13892
rect 17184 13920 17190 13932
rect 17678 13920 17684 13932
rect 17184 13892 17684 13920
rect 17184 13880 17190 13892
rect 17678 13880 17684 13892
rect 17736 13880 17742 13932
rect 13722 13852 13728 13864
rect 13004 13824 13728 13852
rect 13722 13812 13728 13824
rect 13780 13812 13786 13864
rect 13998 13812 14004 13864
rect 14056 13812 14062 13864
rect 14829 13855 14887 13861
rect 14829 13821 14841 13855
rect 14875 13852 14887 13855
rect 15102 13852 15108 13864
rect 14875 13824 15108 13852
rect 14875 13821 14887 13824
rect 14829 13815 14887 13821
rect 15102 13812 15108 13824
rect 15160 13852 15166 13864
rect 17788 13852 17816 14019
rect 19058 14016 19064 14028
rect 19116 14016 19122 14068
rect 19242 14016 19248 14068
rect 19300 14056 19306 14068
rect 19429 14059 19487 14065
rect 19429 14056 19441 14059
rect 19300 14028 19441 14056
rect 19300 14016 19306 14028
rect 19429 14025 19441 14028
rect 19475 14025 19487 14059
rect 19429 14019 19487 14025
rect 18141 13923 18199 13929
rect 18141 13889 18153 13923
rect 18187 13920 18199 13923
rect 18322 13920 18328 13932
rect 18187 13892 18328 13920
rect 18187 13889 18199 13892
rect 18141 13883 18199 13889
rect 18322 13880 18328 13892
rect 18380 13880 18386 13932
rect 18414 13880 18420 13932
rect 18472 13920 18478 13932
rect 18472 13892 18517 13920
rect 18472 13880 18478 13892
rect 19334 13880 19340 13932
rect 19392 13920 19398 13932
rect 19751 13923 19809 13929
rect 19751 13920 19763 13923
rect 19392 13892 19763 13920
rect 19392 13880 19398 13892
rect 19751 13889 19763 13892
rect 19797 13889 19809 13923
rect 19751 13883 19809 13889
rect 15160 13824 16344 13852
rect 17788 13824 18000 13852
rect 15160 13812 15166 13824
rect 14016 13784 14044 13812
rect 16316 13796 16344 13824
rect 14277 13787 14335 13793
rect 14277 13784 14289 13787
rect 14016 13756 14289 13784
rect 14277 13753 14289 13756
rect 14323 13753 14335 13787
rect 14277 13747 14335 13753
rect 16298 13744 16304 13796
rect 16356 13784 16362 13796
rect 16485 13787 16543 13793
rect 16485 13784 16497 13787
rect 16356 13756 16497 13784
rect 16356 13744 16362 13756
rect 16485 13753 16497 13756
rect 16531 13753 16543 13787
rect 16485 13747 16543 13753
rect 16574 13744 16580 13796
rect 16632 13784 16638 13796
rect 17972 13784 18000 13824
rect 19426 13812 19432 13864
rect 19484 13852 19490 13864
rect 19648 13855 19706 13861
rect 19648 13852 19660 13855
rect 19484 13824 19660 13852
rect 19484 13812 19490 13824
rect 19648 13821 19660 13824
rect 19694 13852 19706 13855
rect 20073 13855 20131 13861
rect 20073 13852 20085 13855
rect 19694 13824 20085 13852
rect 19694 13821 19706 13824
rect 19648 13815 19706 13821
rect 20073 13821 20085 13824
rect 20119 13821 20131 13855
rect 20073 13815 20131 13821
rect 18138 13784 18144 13796
rect 16632 13756 16677 13784
rect 17972 13756 18144 13784
rect 16632 13744 16638 13756
rect 18138 13744 18144 13756
rect 18196 13784 18202 13796
rect 18233 13787 18291 13793
rect 18233 13784 18245 13787
rect 18196 13756 18245 13784
rect 18196 13744 18202 13756
rect 18233 13753 18245 13756
rect 18279 13753 18291 13787
rect 18233 13747 18291 13753
rect 9585 13719 9643 13725
rect 9585 13685 9597 13719
rect 9631 13716 9643 13719
rect 9766 13716 9772 13728
rect 9631 13688 9772 13716
rect 9631 13685 9643 13688
rect 9585 13679 9643 13685
rect 9766 13676 9772 13688
rect 9824 13676 9830 13728
rect 9950 13716 9956 13728
rect 9911 13688 9956 13716
rect 9950 13676 9956 13688
rect 10008 13676 10014 13728
rect 11698 13676 11704 13728
rect 11756 13716 11762 13728
rect 11885 13719 11943 13725
rect 11885 13716 11897 13719
rect 11756 13688 11897 13716
rect 11756 13676 11762 13688
rect 11885 13685 11897 13688
rect 11931 13716 11943 13719
rect 12618 13716 12624 13728
rect 11931 13688 12624 13716
rect 11931 13685 11943 13688
rect 11885 13679 11943 13685
rect 12618 13676 12624 13688
rect 12676 13676 12682 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 5718 13512 5724 13524
rect 5679 13484 5724 13512
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 8478 13512 8484 13524
rect 8439 13484 8484 13512
rect 8478 13472 8484 13484
rect 8536 13472 8542 13524
rect 9950 13512 9956 13524
rect 9911 13484 9956 13512
rect 9950 13472 9956 13484
rect 10008 13472 10014 13524
rect 10870 13512 10876 13524
rect 10831 13484 10876 13512
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 12986 13512 12992 13524
rect 12947 13484 12992 13512
rect 12986 13472 12992 13484
rect 13044 13472 13050 13524
rect 15102 13512 15108 13524
rect 15063 13484 15108 13512
rect 15102 13472 15108 13484
rect 15160 13472 15166 13524
rect 15194 13472 15200 13524
rect 15252 13512 15258 13524
rect 16209 13515 16267 13521
rect 16209 13512 16221 13515
rect 15252 13484 16221 13512
rect 15252 13472 15258 13484
rect 16209 13481 16221 13484
rect 16255 13512 16267 13515
rect 16298 13512 16304 13524
rect 16255 13484 16304 13512
rect 16255 13481 16267 13484
rect 16209 13475 16267 13481
rect 16298 13472 16304 13484
rect 16356 13472 16362 13524
rect 16574 13472 16580 13524
rect 16632 13512 16638 13524
rect 17405 13515 17463 13521
rect 17405 13512 17417 13515
rect 16632 13484 17417 13512
rect 16632 13472 16638 13484
rect 17405 13481 17417 13484
rect 17451 13481 17463 13515
rect 18138 13512 18144 13524
rect 18099 13484 18144 13512
rect 17405 13475 17463 13481
rect 18138 13472 18144 13484
rect 18196 13472 18202 13524
rect 19334 13472 19340 13524
rect 19392 13512 19398 13524
rect 19935 13515 19993 13521
rect 19935 13512 19947 13515
rect 19392 13484 19947 13512
rect 19392 13472 19398 13484
rect 19935 13481 19947 13484
rect 19981 13481 19993 13515
rect 19935 13475 19993 13481
rect 2593 13447 2651 13453
rect 2593 13413 2605 13447
rect 2639 13444 2651 13447
rect 2682 13444 2688 13456
rect 2639 13416 2688 13444
rect 2639 13413 2651 13416
rect 2593 13407 2651 13413
rect 2682 13404 2688 13416
rect 2740 13404 2746 13456
rect 4246 13444 4252 13456
rect 4207 13416 4252 13444
rect 4246 13404 4252 13416
rect 4304 13404 4310 13456
rect 8205 13447 8263 13453
rect 8205 13444 8217 13447
rect 6656 13416 8217 13444
rect 5905 13379 5963 13385
rect 5905 13345 5917 13379
rect 5951 13345 5963 13379
rect 6178 13376 6184 13388
rect 6139 13348 6184 13376
rect 5905 13339 5963 13345
rect 1397 13311 1455 13317
rect 1397 13277 1409 13311
rect 1443 13308 1455 13311
rect 2038 13308 2044 13320
rect 1443 13280 2044 13308
rect 1443 13277 1455 13280
rect 1397 13271 1455 13277
rect 2038 13268 2044 13280
rect 2096 13308 2102 13320
rect 2501 13311 2559 13317
rect 2501 13308 2513 13311
rect 2096 13280 2513 13308
rect 2096 13268 2102 13280
rect 2501 13277 2513 13280
rect 2547 13277 2559 13311
rect 2501 13271 2559 13277
rect 4157 13311 4215 13317
rect 4157 13277 4169 13311
rect 4203 13308 4215 13311
rect 4338 13308 4344 13320
rect 4203 13280 4344 13308
rect 4203 13277 4215 13280
rect 4157 13271 4215 13277
rect 4338 13268 4344 13280
rect 4396 13268 4402 13320
rect 4433 13311 4491 13317
rect 4433 13277 4445 13311
rect 4479 13277 4491 13311
rect 4433 13271 4491 13277
rect 5537 13311 5595 13317
rect 5537 13277 5549 13311
rect 5583 13308 5595 13311
rect 5920 13308 5948 13339
rect 6178 13336 6184 13348
rect 6236 13336 6242 13388
rect 6362 13336 6368 13388
rect 6420 13376 6426 13388
rect 6656 13385 6684 13416
rect 8205 13413 8217 13416
rect 8251 13444 8263 13447
rect 9030 13444 9036 13456
rect 8251 13416 9036 13444
rect 8251 13413 8263 13416
rect 8205 13407 8263 13413
rect 9030 13404 9036 13416
rect 9088 13404 9094 13456
rect 12894 13404 12900 13456
rect 12952 13444 12958 13456
rect 16850 13453 16856 13456
rect 13541 13447 13599 13453
rect 13541 13444 13553 13447
rect 12952 13416 13553 13444
rect 12952 13404 12958 13416
rect 13541 13413 13553 13416
rect 13587 13444 13599 13447
rect 14369 13447 14427 13453
rect 13587 13416 14228 13444
rect 13587 13413 13599 13416
rect 13541 13407 13599 13413
rect 6641 13379 6699 13385
rect 6641 13376 6653 13379
rect 6420 13348 6653 13376
rect 6420 13336 6426 13348
rect 6641 13345 6653 13348
rect 6687 13345 6699 13379
rect 6641 13339 6699 13345
rect 7009 13379 7067 13385
rect 7009 13345 7021 13379
rect 7055 13376 7067 13379
rect 7466 13376 7472 13388
rect 7055 13348 7472 13376
rect 7055 13345 7067 13348
rect 7009 13339 7067 13345
rect 7466 13336 7472 13348
rect 7524 13336 7530 13388
rect 8389 13379 8447 13385
rect 8389 13345 8401 13379
rect 8435 13376 8447 13379
rect 8754 13376 8760 13388
rect 8435 13348 8760 13376
rect 8435 13345 8447 13348
rect 8389 13339 8447 13345
rect 8754 13336 8760 13348
rect 8812 13336 8818 13388
rect 9766 13336 9772 13388
rect 9824 13376 9830 13388
rect 10321 13379 10379 13385
rect 10321 13376 10333 13379
rect 9824 13348 10333 13376
rect 9824 13336 9830 13348
rect 10321 13345 10333 13348
rect 10367 13376 10379 13379
rect 10870 13376 10876 13388
rect 10367 13348 10876 13376
rect 10367 13345 10379 13348
rect 10321 13339 10379 13345
rect 10870 13336 10876 13348
rect 10928 13336 10934 13388
rect 11698 13376 11704 13388
rect 11659 13348 11704 13376
rect 11698 13336 11704 13348
rect 11756 13336 11762 13388
rect 13630 13376 13636 13388
rect 13591 13348 13636 13376
rect 13630 13336 13636 13348
rect 13688 13336 13694 13388
rect 14200 13385 14228 13416
rect 14369 13413 14381 13447
rect 14415 13444 14427 13447
rect 14415 13416 16528 13444
rect 14415 13413 14427 13416
rect 14369 13407 14427 13413
rect 14185 13379 14243 13385
rect 14185 13345 14197 13379
rect 14231 13376 14243 13379
rect 15194 13376 15200 13388
rect 14231 13348 15200 13376
rect 14231 13345 14243 13348
rect 14185 13339 14243 13345
rect 15194 13336 15200 13348
rect 15252 13336 15258 13388
rect 16500 13385 16528 13416
rect 16847 13407 16856 13453
rect 16908 13444 16914 13456
rect 16908 13416 16995 13444
rect 16850 13404 16856 13407
rect 16908 13404 16914 13416
rect 18046 13404 18052 13456
rect 18104 13444 18110 13456
rect 18417 13447 18475 13453
rect 18417 13444 18429 13447
rect 18104 13416 18429 13444
rect 18104 13404 18110 13416
rect 18417 13413 18429 13416
rect 18463 13444 18475 13447
rect 19058 13444 19064 13456
rect 18463 13416 19064 13444
rect 18463 13413 18475 13416
rect 18417 13407 18475 13413
rect 19058 13404 19064 13416
rect 19116 13404 19122 13456
rect 15289 13379 15347 13385
rect 15289 13345 15301 13379
rect 15335 13376 15347 13379
rect 16485 13379 16543 13385
rect 15335 13348 15884 13376
rect 15335 13345 15347 13348
rect 15289 13339 15347 13345
rect 6086 13308 6092 13320
rect 5583 13280 6092 13308
rect 5583 13277 5595 13280
rect 5537 13271 5595 13277
rect 3053 13243 3111 13249
rect 3053 13240 3065 13243
rect 1872 13212 3065 13240
rect 1486 13132 1492 13184
rect 1544 13172 1550 13184
rect 1872 13181 1900 13212
rect 3053 13209 3065 13212
rect 3099 13240 3111 13243
rect 4448 13240 4476 13271
rect 6086 13268 6092 13280
rect 6144 13268 6150 13320
rect 11422 13308 11428 13320
rect 11383 13280 11428 13308
rect 11422 13268 11428 13280
rect 11480 13268 11486 13320
rect 12345 13311 12403 13317
rect 12345 13277 12357 13311
rect 12391 13308 12403 13311
rect 12434 13308 12440 13320
rect 12391 13280 12440 13308
rect 12391 13277 12403 13280
rect 12345 13271 12403 13277
rect 12434 13268 12440 13280
rect 12492 13268 12498 13320
rect 15856 13249 15884 13348
rect 16485 13345 16497 13379
rect 16531 13376 16543 13379
rect 16666 13376 16672 13388
rect 16531 13348 16672 13376
rect 16531 13345 16543 13348
rect 16485 13339 16543 13345
rect 16666 13336 16672 13348
rect 16724 13336 16730 13388
rect 16574 13268 16580 13320
rect 16632 13308 16638 13320
rect 16862 13308 16890 13404
rect 19794 13336 19800 13388
rect 19852 13385 19858 13388
rect 19852 13379 19890 13385
rect 19878 13345 19890 13379
rect 19852 13339 19890 13345
rect 19852 13336 19858 13339
rect 16632 13280 16890 13308
rect 18325 13311 18383 13317
rect 16632 13268 16638 13280
rect 18325 13277 18337 13311
rect 18371 13308 18383 13311
rect 18598 13308 18604 13320
rect 18371 13280 18604 13308
rect 18371 13277 18383 13280
rect 18325 13271 18383 13277
rect 18598 13268 18604 13280
rect 18656 13268 18662 13320
rect 18782 13308 18788 13320
rect 18743 13280 18788 13308
rect 18782 13268 18788 13280
rect 18840 13268 18846 13320
rect 3099 13212 4476 13240
rect 15841 13243 15899 13249
rect 3099 13209 3111 13212
rect 3053 13203 3111 13209
rect 15841 13209 15853 13243
rect 15887 13240 15899 13243
rect 16850 13240 16856 13252
rect 15887 13212 16856 13240
rect 15887 13209 15899 13212
rect 15841 13203 15899 13209
rect 16850 13200 16856 13212
rect 16908 13200 16914 13252
rect 1857 13175 1915 13181
rect 1857 13172 1869 13175
rect 1544 13144 1869 13172
rect 1544 13132 1550 13144
rect 1857 13141 1869 13144
rect 1903 13141 1915 13175
rect 2222 13172 2228 13184
rect 2183 13144 2228 13172
rect 1857 13135 1915 13141
rect 2222 13132 2228 13144
rect 2280 13132 2286 13184
rect 3510 13172 3516 13184
rect 3471 13144 3516 13172
rect 3510 13132 3516 13144
rect 3568 13132 3574 13184
rect 7374 13172 7380 13184
rect 7335 13144 7380 13172
rect 7374 13132 7380 13144
rect 7432 13132 7438 13184
rect 7837 13175 7895 13181
rect 7837 13141 7849 13175
rect 7883 13172 7895 13175
rect 7926 13172 7932 13184
rect 7883 13144 7932 13172
rect 7883 13141 7895 13144
rect 7837 13135 7895 13141
rect 7926 13132 7932 13144
rect 7984 13132 7990 13184
rect 9217 13175 9275 13181
rect 9217 13141 9229 13175
rect 9263 13172 9275 13175
rect 10134 13172 10140 13184
rect 9263 13144 10140 13172
rect 9263 13141 9275 13144
rect 9217 13135 9275 13141
rect 10134 13132 10140 13144
rect 10192 13132 10198 13184
rect 15473 13175 15531 13181
rect 15473 13141 15485 13175
rect 15519 13172 15531 13175
rect 15654 13172 15660 13184
rect 15519 13144 15660 13172
rect 15519 13141 15531 13144
rect 15473 13135 15531 13141
rect 15654 13132 15660 13144
rect 15712 13132 15718 13184
rect 17770 13172 17776 13184
rect 17731 13144 17776 13172
rect 17770 13132 17776 13144
rect 17828 13132 17834 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 2038 12968 2044 12980
rect 1999 12940 2044 12968
rect 2038 12928 2044 12940
rect 2096 12928 2102 12980
rect 3878 12968 3884 12980
rect 3791 12940 3884 12968
rect 3878 12928 3884 12940
rect 3936 12968 3942 12980
rect 4246 12968 4252 12980
rect 3936 12940 4252 12968
rect 3936 12928 3942 12940
rect 4246 12928 4252 12940
rect 4304 12928 4310 12980
rect 4890 12968 4896 12980
rect 4851 12940 4896 12968
rect 4890 12928 4896 12940
rect 4948 12928 4954 12980
rect 8665 12971 8723 12977
rect 8665 12937 8677 12971
rect 8711 12968 8723 12971
rect 8754 12968 8760 12980
rect 8711 12940 8760 12968
rect 8711 12937 8723 12940
rect 8665 12931 8723 12937
rect 8754 12928 8760 12940
rect 8812 12928 8818 12980
rect 9030 12968 9036 12980
rect 8943 12940 9036 12968
rect 9030 12928 9036 12940
rect 9088 12968 9094 12980
rect 9766 12968 9772 12980
rect 9088 12940 9772 12968
rect 9088 12928 9094 12940
rect 9766 12928 9772 12940
rect 9824 12928 9830 12980
rect 11698 12968 11704 12980
rect 11659 12940 11704 12968
rect 11698 12928 11704 12940
rect 11756 12928 11762 12980
rect 13630 12968 13636 12980
rect 13591 12940 13636 12968
rect 13630 12928 13636 12940
rect 13688 12968 13694 12980
rect 14458 12968 14464 12980
rect 13688 12940 14464 12968
rect 13688 12928 13694 12940
rect 14458 12928 14464 12940
rect 14516 12928 14522 12980
rect 16114 12928 16120 12980
rect 16172 12968 16178 12980
rect 17129 12971 17187 12977
rect 17129 12968 17141 12971
rect 16172 12940 17141 12968
rect 16172 12928 16178 12940
rect 17129 12937 17141 12940
rect 17175 12968 17187 12971
rect 17586 12968 17592 12980
rect 17175 12940 17592 12968
rect 17175 12937 17187 12940
rect 17129 12931 17187 12937
rect 17586 12928 17592 12940
rect 17644 12928 17650 12980
rect 18598 12928 18604 12980
rect 18656 12968 18662 12980
rect 19429 12971 19487 12977
rect 19429 12968 19441 12971
rect 18656 12940 19441 12968
rect 18656 12928 18662 12940
rect 19429 12937 19441 12940
rect 19475 12937 19487 12971
rect 19429 12931 19487 12937
rect 19886 12928 19892 12980
rect 19944 12968 19950 12980
rect 20073 12971 20131 12977
rect 20073 12968 20085 12971
rect 19944 12940 20085 12968
rect 19944 12928 19950 12940
rect 20073 12937 20085 12940
rect 20119 12937 20131 12971
rect 20073 12931 20131 12937
rect 5902 12860 5908 12912
rect 5960 12900 5966 12912
rect 6178 12900 6184 12912
rect 5960 12872 6184 12900
rect 5960 12860 5966 12872
rect 6178 12860 6184 12872
rect 6236 12860 6242 12912
rect 11241 12903 11299 12909
rect 11241 12900 11253 12903
rect 9600 12872 11253 12900
rect 1397 12767 1455 12773
rect 1397 12733 1409 12767
rect 1443 12764 1455 12767
rect 1578 12764 1584 12776
rect 1443 12736 1584 12764
rect 1443 12733 1455 12736
rect 1397 12727 1455 12733
rect 1578 12724 1584 12736
rect 1636 12764 1642 12776
rect 2222 12764 2228 12776
rect 1636 12736 2228 12764
rect 1636 12724 1642 12736
rect 2222 12724 2228 12736
rect 2280 12724 2286 12776
rect 2961 12767 3019 12773
rect 2961 12733 2973 12767
rect 3007 12764 3019 12767
rect 3510 12764 3516 12776
rect 3007 12736 3516 12764
rect 3007 12733 3019 12736
rect 2961 12727 3019 12733
rect 3510 12724 3516 12736
rect 3568 12724 3574 12776
rect 4617 12767 4675 12773
rect 4617 12733 4629 12767
rect 4663 12764 4675 12767
rect 4706 12764 4712 12776
rect 4663 12736 4712 12764
rect 4663 12733 4675 12736
rect 4617 12727 4675 12733
rect 4706 12724 4712 12736
rect 4764 12724 4770 12776
rect 5721 12767 5779 12773
rect 5721 12733 5733 12767
rect 5767 12733 5779 12767
rect 5721 12727 5779 12733
rect 2590 12656 2596 12708
rect 2648 12696 2654 12708
rect 2777 12699 2835 12705
rect 2777 12696 2789 12699
rect 2648 12668 2789 12696
rect 2648 12656 2654 12668
rect 2777 12665 2789 12668
rect 2823 12696 2835 12699
rect 2866 12696 2872 12708
rect 2823 12668 2872 12696
rect 2823 12665 2835 12668
rect 2777 12659 2835 12665
rect 2866 12656 2872 12668
rect 2924 12696 2930 12708
rect 3282 12699 3340 12705
rect 3282 12696 3294 12699
rect 2924 12668 3294 12696
rect 2924 12656 2930 12668
rect 3282 12665 3294 12668
rect 3328 12665 3340 12699
rect 5736 12696 5764 12727
rect 6454 12724 6460 12776
rect 6512 12764 6518 12776
rect 6822 12764 6828 12776
rect 6512 12736 6828 12764
rect 6512 12724 6518 12736
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 7374 12764 7380 12776
rect 7335 12736 7380 12764
rect 7374 12724 7380 12736
rect 7432 12764 7438 12776
rect 7558 12764 7564 12776
rect 7432 12736 7564 12764
rect 7432 12724 7438 12736
rect 7558 12724 7564 12736
rect 7616 12724 7622 12776
rect 7837 12767 7895 12773
rect 7837 12733 7849 12767
rect 7883 12764 7895 12767
rect 7926 12764 7932 12776
rect 7883 12736 7932 12764
rect 7883 12733 7895 12736
rect 7837 12727 7895 12733
rect 7926 12724 7932 12736
rect 7984 12724 7990 12776
rect 8021 12767 8079 12773
rect 8021 12733 8033 12767
rect 8067 12733 8079 12767
rect 8021 12727 8079 12733
rect 6270 12696 6276 12708
rect 5736 12668 6276 12696
rect 3282 12659 3340 12665
rect 6270 12656 6276 12668
rect 6328 12656 6334 12708
rect 6546 12656 6552 12708
rect 6604 12696 6610 12708
rect 6641 12699 6699 12705
rect 6641 12696 6653 12699
rect 6604 12668 6653 12696
rect 6604 12656 6610 12668
rect 6641 12665 6653 12668
rect 6687 12696 6699 12699
rect 8036 12696 8064 12727
rect 8938 12724 8944 12776
rect 8996 12764 9002 12776
rect 9401 12767 9459 12773
rect 9401 12764 9413 12767
rect 8996 12736 9413 12764
rect 8996 12724 9002 12736
rect 9401 12733 9413 12736
rect 9447 12764 9459 12767
rect 9600 12764 9628 12872
rect 11241 12869 11253 12872
rect 11287 12869 11299 12903
rect 16482 12900 16488 12912
rect 11241 12863 11299 12869
rect 16132 12872 16488 12900
rect 10873 12835 10931 12841
rect 10873 12832 10885 12835
rect 9876 12804 10885 12832
rect 9876 12776 9904 12804
rect 10873 12801 10885 12804
rect 10919 12801 10931 12835
rect 10873 12795 10931 12801
rect 14553 12835 14611 12841
rect 14553 12801 14565 12835
rect 14599 12832 14611 12835
rect 14826 12832 14832 12844
rect 14599 12804 14832 12832
rect 14599 12801 14611 12804
rect 14553 12795 14611 12801
rect 14826 12792 14832 12804
rect 14884 12792 14890 12844
rect 16132 12841 16160 12872
rect 16482 12860 16488 12872
rect 16540 12860 16546 12912
rect 19058 12900 19064 12912
rect 19019 12872 19064 12900
rect 19058 12860 19064 12872
rect 19116 12860 19122 12912
rect 19794 12900 19800 12912
rect 19755 12872 19800 12900
rect 19794 12860 19800 12872
rect 19852 12860 19858 12912
rect 16117 12835 16175 12841
rect 16117 12801 16129 12835
rect 16163 12801 16175 12835
rect 16117 12795 16175 12801
rect 17770 12792 17776 12844
rect 17828 12832 17834 12844
rect 18141 12835 18199 12841
rect 18141 12832 18153 12835
rect 17828 12804 18153 12832
rect 17828 12792 17834 12804
rect 18141 12801 18153 12804
rect 18187 12832 18199 12835
rect 18506 12832 18512 12844
rect 18187 12804 18512 12832
rect 18187 12801 18199 12804
rect 18141 12795 18199 12801
rect 18506 12792 18512 12804
rect 18564 12792 18570 12844
rect 18782 12832 18788 12844
rect 18743 12804 18788 12832
rect 18782 12792 18788 12804
rect 18840 12792 18846 12844
rect 9447 12736 9628 12764
rect 9447 12733 9459 12736
rect 9401 12727 9459 12733
rect 9674 12724 9680 12776
rect 9732 12724 9738 12776
rect 9858 12764 9864 12776
rect 9771 12736 9864 12764
rect 9858 12724 9864 12736
rect 9916 12724 9922 12776
rect 10134 12764 10140 12776
rect 10095 12736 10140 12764
rect 10134 12724 10140 12736
rect 10192 12724 10198 12776
rect 10321 12767 10379 12773
rect 10321 12764 10333 12767
rect 10244 12736 10333 12764
rect 9692 12696 9720 12724
rect 6687 12668 8064 12696
rect 9416 12668 9720 12696
rect 6687 12665 6699 12668
rect 6641 12659 6699 12665
rect 1394 12588 1400 12640
rect 1452 12628 1458 12640
rect 1581 12631 1639 12637
rect 1581 12628 1593 12631
rect 1452 12600 1593 12628
rect 1452 12588 1458 12600
rect 1581 12597 1593 12600
rect 1627 12597 1639 12631
rect 1581 12591 1639 12597
rect 2501 12631 2559 12637
rect 2501 12597 2513 12631
rect 2547 12628 2559 12631
rect 2682 12628 2688 12640
rect 2547 12600 2688 12628
rect 2547 12597 2559 12600
rect 2501 12591 2559 12597
rect 2682 12588 2688 12600
rect 2740 12588 2746 12640
rect 5166 12628 5172 12640
rect 5127 12600 5172 12628
rect 5166 12588 5172 12600
rect 5224 12588 5230 12640
rect 5629 12631 5687 12637
rect 5629 12597 5641 12631
rect 5675 12628 5687 12631
rect 5905 12631 5963 12637
rect 5905 12628 5917 12631
rect 5675 12600 5917 12628
rect 5675 12597 5687 12600
rect 5629 12591 5687 12597
rect 5905 12597 5917 12600
rect 5951 12628 5963 12631
rect 6362 12628 6368 12640
rect 5951 12600 6368 12628
rect 5951 12597 5963 12600
rect 5905 12591 5963 12597
rect 6362 12588 6368 12600
rect 6420 12588 6426 12640
rect 7098 12628 7104 12640
rect 7059 12600 7104 12628
rect 7098 12588 7104 12600
rect 7156 12588 7162 12640
rect 9416 12637 9444 12668
rect 9401 12631 9459 12637
rect 9401 12597 9413 12631
rect 9447 12597 9459 12631
rect 9401 12591 9459 12597
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 10244 12628 10272 12736
rect 10321 12733 10333 12736
rect 10367 12764 10379 12767
rect 10367 12736 11928 12764
rect 10367 12733 10379 12736
rect 10321 12727 10379 12733
rect 11900 12696 11928 12736
rect 11974 12724 11980 12776
rect 12032 12764 12038 12776
rect 12253 12767 12311 12773
rect 12253 12764 12265 12767
rect 12032 12736 12265 12764
rect 12032 12724 12038 12736
rect 12253 12733 12265 12736
rect 12299 12764 12311 12767
rect 13081 12767 13139 12773
rect 13081 12764 13093 12767
rect 12299 12736 13093 12764
rect 12299 12733 12311 12736
rect 12253 12727 12311 12733
rect 13081 12733 13093 12736
rect 13127 12764 13139 12767
rect 13538 12764 13544 12776
rect 13127 12736 13544 12764
rect 13127 12733 13139 12736
rect 13081 12727 13139 12733
rect 13538 12724 13544 12736
rect 13596 12724 13602 12776
rect 14182 12764 14188 12776
rect 14143 12736 14188 12764
rect 14182 12724 14188 12736
rect 14240 12764 14246 12776
rect 14921 12767 14979 12773
rect 14921 12764 14933 12767
rect 14240 12736 14933 12764
rect 14240 12724 14246 12736
rect 14921 12733 14933 12736
rect 14967 12764 14979 12767
rect 15194 12764 15200 12776
rect 14967 12736 15200 12764
rect 14967 12733 14979 12736
rect 14921 12727 14979 12733
rect 15194 12724 15200 12736
rect 15252 12724 15258 12776
rect 15289 12767 15347 12773
rect 15289 12733 15301 12767
rect 15335 12764 15347 12767
rect 15378 12764 15384 12776
rect 15335 12736 15384 12764
rect 15335 12733 15347 12736
rect 15289 12727 15347 12733
rect 15378 12724 15384 12736
rect 15436 12764 15442 12776
rect 15657 12767 15715 12773
rect 15657 12764 15669 12767
rect 15436 12736 15669 12764
rect 15436 12724 15442 12736
rect 15657 12733 15669 12736
rect 15703 12764 15715 12767
rect 15746 12764 15752 12776
rect 15703 12736 15752 12764
rect 15703 12733 15715 12736
rect 15657 12727 15715 12733
rect 15746 12724 15752 12736
rect 15804 12724 15810 12776
rect 15838 12724 15844 12776
rect 15896 12764 15902 12776
rect 15933 12767 15991 12773
rect 15933 12764 15945 12767
rect 15896 12736 15945 12764
rect 15896 12724 15902 12736
rect 15933 12733 15945 12736
rect 15979 12764 15991 12767
rect 16298 12764 16304 12776
rect 15979 12736 16304 12764
rect 15979 12733 15991 12736
rect 15933 12727 15991 12733
rect 16298 12724 16304 12736
rect 16356 12724 16362 12776
rect 16482 12724 16488 12776
rect 16540 12764 16546 12776
rect 16945 12767 17003 12773
rect 16945 12764 16957 12767
rect 16540 12736 16957 12764
rect 16540 12724 16546 12736
rect 16945 12733 16957 12736
rect 16991 12764 17003 12767
rect 17405 12767 17463 12773
rect 17405 12764 17417 12767
rect 16991 12736 17417 12764
rect 16991 12733 17003 12736
rect 16945 12727 17003 12733
rect 17405 12733 17417 12736
rect 17451 12733 17463 12767
rect 17405 12727 17463 12733
rect 19334 12724 19340 12776
rect 19392 12764 19398 12776
rect 19613 12767 19671 12773
rect 19613 12764 19625 12767
rect 19392 12736 19625 12764
rect 19392 12724 19398 12736
rect 19613 12733 19625 12736
rect 19659 12764 19671 12767
rect 20441 12767 20499 12773
rect 20441 12764 20453 12767
rect 19659 12736 20453 12764
rect 19659 12733 19671 12736
rect 19613 12727 19671 12733
rect 20441 12733 20453 12736
rect 20487 12733 20499 12767
rect 20441 12727 20499 12733
rect 13998 12696 14004 12708
rect 11900 12668 13860 12696
rect 13959 12668 14004 12696
rect 12710 12628 12716 12640
rect 9732 12600 10272 12628
rect 12671 12600 12716 12628
rect 9732 12588 9738 12600
rect 12710 12588 12716 12600
rect 12768 12588 12774 12640
rect 13832 12628 13860 12668
rect 13998 12656 14004 12668
rect 14056 12656 14062 12708
rect 16758 12656 16764 12708
rect 16816 12696 16822 12708
rect 17865 12699 17923 12705
rect 17865 12696 17877 12699
rect 16816 12668 17877 12696
rect 16816 12656 16822 12668
rect 17865 12665 17877 12668
rect 17911 12696 17923 12699
rect 18233 12699 18291 12705
rect 18233 12696 18245 12699
rect 17911 12668 18245 12696
rect 17911 12665 17923 12668
rect 17865 12659 17923 12665
rect 18233 12665 18245 12668
rect 18279 12665 18291 12699
rect 18233 12659 18291 12665
rect 14182 12628 14188 12640
rect 13832 12600 14188 12628
rect 14182 12588 14188 12600
rect 14240 12588 14246 12640
rect 16574 12628 16580 12640
rect 16535 12600 16580 12628
rect 16574 12588 16580 12600
rect 16632 12588 16638 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1578 12433 1584 12436
rect 1535 12427 1584 12433
rect 1535 12393 1547 12427
rect 1581 12393 1584 12427
rect 1535 12387 1584 12393
rect 1578 12384 1584 12387
rect 1636 12384 1642 12436
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 2869 12427 2927 12433
rect 2869 12424 2881 12427
rect 2832 12396 2881 12424
rect 2832 12384 2838 12396
rect 2869 12393 2881 12396
rect 2915 12393 2927 12427
rect 3878 12424 3884 12436
rect 3839 12396 3884 12424
rect 2869 12387 2927 12393
rect 3878 12384 3884 12396
rect 3936 12384 3942 12436
rect 4338 12424 4344 12436
rect 4299 12396 4344 12424
rect 4338 12384 4344 12396
rect 4396 12384 4402 12436
rect 4614 12433 4620 12436
rect 4571 12427 4620 12433
rect 4571 12393 4583 12427
rect 4617 12393 4620 12427
rect 4571 12387 4620 12393
rect 4614 12384 4620 12387
rect 4672 12384 4678 12436
rect 5534 12384 5540 12436
rect 5592 12433 5598 12436
rect 5592 12427 5641 12433
rect 5592 12393 5595 12427
rect 5629 12393 5641 12427
rect 5902 12424 5908 12436
rect 5863 12396 5908 12424
rect 5592 12387 5641 12393
rect 5592 12384 5598 12387
rect 5902 12384 5908 12396
rect 5960 12424 5966 12436
rect 6178 12424 6184 12436
rect 5960 12396 6184 12424
rect 5960 12384 5966 12396
rect 6178 12384 6184 12396
rect 6236 12384 6242 12436
rect 7006 12384 7012 12436
rect 7064 12424 7070 12436
rect 7653 12427 7711 12433
rect 7653 12424 7665 12427
rect 7064 12396 7665 12424
rect 7064 12384 7070 12396
rect 7653 12393 7665 12396
rect 7699 12393 7711 12427
rect 7653 12387 7711 12393
rect 9769 12427 9827 12433
rect 9769 12393 9781 12427
rect 9815 12424 9827 12427
rect 9858 12424 9864 12436
rect 9815 12396 9864 12424
rect 9815 12393 9827 12396
rect 9769 12387 9827 12393
rect 9858 12384 9864 12396
rect 9916 12384 9922 12436
rect 10134 12384 10140 12436
rect 10192 12424 10198 12436
rect 10870 12424 10876 12436
rect 10192 12384 10226 12424
rect 10831 12396 10876 12424
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 12713 12427 12771 12433
rect 12713 12424 12725 12427
rect 12492 12396 12725 12424
rect 12492 12384 12498 12396
rect 12713 12393 12725 12396
rect 12759 12424 12771 12427
rect 13081 12427 13139 12433
rect 13081 12424 13093 12427
rect 12759 12396 13093 12424
rect 12759 12393 12771 12396
rect 12713 12387 12771 12393
rect 13081 12393 13093 12396
rect 13127 12393 13139 12427
rect 14366 12424 14372 12436
rect 13081 12387 13139 12393
rect 14016 12396 14372 12424
rect 1486 12297 1492 12300
rect 1464 12291 1492 12297
rect 1464 12257 1476 12291
rect 1464 12251 1492 12257
rect 1486 12248 1492 12251
rect 1544 12248 1550 12300
rect 3053 12291 3111 12297
rect 3053 12257 3065 12291
rect 3099 12288 3111 12291
rect 3896 12288 3924 12384
rect 7926 12356 7932 12368
rect 7484 12328 7932 12356
rect 3099 12260 3924 12288
rect 4500 12291 4558 12297
rect 3099 12257 3111 12260
rect 3053 12251 3111 12257
rect 4500 12257 4512 12291
rect 4546 12288 4558 12291
rect 5350 12288 5356 12300
rect 4546 12260 5356 12288
rect 4546 12257 4558 12260
rect 4500 12251 4558 12257
rect 5350 12248 5356 12260
rect 5408 12248 5414 12300
rect 5534 12297 5540 12300
rect 5512 12291 5540 12297
rect 5512 12257 5524 12291
rect 5512 12251 5540 12257
rect 5534 12248 5540 12251
rect 5592 12248 5598 12300
rect 6454 12288 6460 12300
rect 5644 12260 6460 12288
rect 4890 12220 4896 12232
rect 4851 12192 4896 12220
rect 4890 12180 4896 12192
rect 4948 12180 4954 12232
rect 1949 12155 2007 12161
rect 1949 12121 1961 12155
rect 1995 12152 2007 12155
rect 2866 12152 2872 12164
rect 1995 12124 2872 12152
rect 1995 12121 2007 12124
rect 1949 12115 2007 12121
rect 2866 12112 2872 12124
rect 2924 12112 2930 12164
rect 5350 12112 5356 12164
rect 5408 12152 5414 12164
rect 5644 12152 5672 12260
rect 6454 12248 6460 12260
rect 6512 12248 6518 12300
rect 6917 12291 6975 12297
rect 6917 12257 6929 12291
rect 6963 12257 6975 12291
rect 6917 12251 6975 12257
rect 6365 12223 6423 12229
rect 6365 12189 6377 12223
rect 6411 12220 6423 12223
rect 6638 12220 6644 12232
rect 6411 12192 6644 12220
rect 6411 12189 6423 12192
rect 6365 12183 6423 12189
rect 6638 12180 6644 12192
rect 6696 12220 6702 12232
rect 6932 12220 6960 12251
rect 7098 12248 7104 12300
rect 7156 12288 7162 12300
rect 7484 12297 7512 12328
rect 7926 12316 7932 12328
rect 7984 12316 7990 12368
rect 9950 12316 9956 12368
rect 10008 12356 10014 12368
rect 10198 12356 10226 12384
rect 13096 12356 13124 12387
rect 14016 12365 14044 12396
rect 14366 12384 14372 12396
rect 14424 12384 14430 12436
rect 15562 12424 15568 12436
rect 15523 12396 15568 12424
rect 15562 12384 15568 12396
rect 15620 12384 15626 12436
rect 16577 12427 16635 12433
rect 16577 12393 16589 12427
rect 16623 12424 16635 12427
rect 16666 12424 16672 12436
rect 16623 12396 16672 12424
rect 16623 12393 16635 12396
rect 16577 12387 16635 12393
rect 16666 12384 16672 12396
rect 16724 12384 16730 12436
rect 17681 12427 17739 12433
rect 17681 12393 17693 12427
rect 17727 12424 17739 12427
rect 17727 12396 18736 12424
rect 17727 12393 17739 12396
rect 17681 12387 17739 12393
rect 14001 12359 14059 12365
rect 10008 12328 12848 12356
rect 13096 12328 13400 12356
rect 10008 12316 10014 12328
rect 7469 12291 7527 12297
rect 7469 12288 7481 12291
rect 7156 12260 7481 12288
rect 7156 12248 7162 12260
rect 7469 12257 7481 12260
rect 7515 12257 7527 12291
rect 7650 12288 7656 12300
rect 7611 12260 7656 12288
rect 7469 12251 7527 12257
rect 7650 12248 7656 12260
rect 7708 12288 7714 12300
rect 9125 12291 9183 12297
rect 9125 12288 9137 12291
rect 7708 12260 9137 12288
rect 7708 12248 7714 12260
rect 9125 12257 9137 12260
rect 9171 12288 9183 12291
rect 9674 12288 9680 12300
rect 9171 12260 9680 12288
rect 9171 12257 9183 12260
rect 9125 12251 9183 12257
rect 9674 12248 9680 12260
rect 9732 12248 9738 12300
rect 9858 12288 9864 12300
rect 9819 12260 9864 12288
rect 9858 12248 9864 12260
rect 9916 12248 9922 12300
rect 10134 12288 10140 12300
rect 10095 12260 10140 12288
rect 10134 12248 10140 12260
rect 10192 12248 10198 12300
rect 11701 12291 11759 12297
rect 11701 12257 11713 12291
rect 11747 12288 11759 12291
rect 11790 12288 11796 12300
rect 11747 12260 11796 12288
rect 11747 12257 11759 12260
rect 11701 12251 11759 12257
rect 11790 12248 11796 12260
rect 11848 12248 11854 12300
rect 11977 12291 12035 12297
rect 11977 12257 11989 12291
rect 12023 12288 12035 12291
rect 12710 12288 12716 12300
rect 12023 12260 12716 12288
rect 12023 12257 12035 12260
rect 11977 12251 12035 12257
rect 7558 12220 7564 12232
rect 6696 12192 7564 12220
rect 6696 12180 6702 12192
rect 7558 12180 7564 12192
rect 7616 12220 7622 12232
rect 8570 12220 8576 12232
rect 7616 12192 8576 12220
rect 7616 12180 7622 12192
rect 8570 12180 8576 12192
rect 8628 12220 8634 12232
rect 9769 12223 9827 12229
rect 9769 12220 9781 12223
rect 8628 12192 9781 12220
rect 8628 12180 8634 12192
rect 9769 12189 9781 12192
rect 9815 12220 9827 12223
rect 9953 12223 10011 12229
rect 9953 12220 9965 12223
rect 9815 12192 9965 12220
rect 9815 12189 9827 12192
rect 9769 12183 9827 12189
rect 9953 12189 9965 12192
rect 9999 12189 10011 12223
rect 10318 12220 10324 12232
rect 10279 12192 10324 12220
rect 9953 12183 10011 12189
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 11609 12223 11667 12229
rect 11609 12189 11621 12223
rect 11655 12220 11667 12223
rect 11992 12220 12020 12251
rect 12710 12248 12716 12260
rect 12768 12248 12774 12300
rect 12158 12220 12164 12232
rect 11655 12192 12020 12220
rect 12119 12192 12164 12220
rect 11655 12189 11667 12192
rect 11609 12183 11667 12189
rect 12158 12180 12164 12192
rect 12216 12180 12222 12232
rect 12820 12220 12848 12328
rect 13170 12248 13176 12300
rect 13228 12288 13234 12300
rect 13372 12297 13400 12328
rect 14001 12325 14013 12359
rect 14047 12325 14059 12359
rect 14001 12319 14059 12325
rect 15194 12316 15200 12368
rect 15252 12356 15258 12368
rect 18708 12365 18736 12396
rect 17082 12359 17140 12365
rect 17082 12356 17094 12359
rect 15252 12328 15516 12356
rect 15252 12316 15258 12328
rect 15488 12300 15516 12328
rect 16684 12328 17094 12356
rect 16684 12300 16712 12328
rect 17082 12325 17094 12328
rect 17128 12325 17140 12359
rect 17082 12319 17140 12325
rect 18693 12359 18751 12365
rect 18693 12325 18705 12359
rect 18739 12356 18751 12359
rect 19058 12356 19064 12368
rect 18739 12328 19064 12356
rect 18739 12325 18751 12328
rect 18693 12319 18751 12325
rect 19058 12316 19064 12328
rect 19116 12316 19122 12368
rect 13265 12291 13323 12297
rect 13265 12288 13277 12291
rect 13228 12260 13277 12288
rect 13228 12248 13234 12260
rect 13265 12257 13277 12260
rect 13311 12257 13323 12291
rect 13265 12251 13323 12257
rect 13357 12291 13415 12297
rect 13357 12257 13369 12291
rect 13403 12257 13415 12291
rect 13538 12288 13544 12300
rect 13499 12260 13544 12288
rect 13357 12251 13415 12257
rect 13538 12248 13544 12260
rect 13596 12248 13602 12300
rect 15105 12291 15163 12297
rect 15105 12257 15117 12291
rect 15151 12288 15163 12291
rect 15289 12291 15347 12297
rect 15289 12288 15301 12291
rect 15151 12260 15301 12288
rect 15151 12257 15163 12260
rect 15105 12251 15163 12257
rect 15289 12257 15301 12260
rect 15335 12257 15347 12291
rect 15470 12288 15476 12300
rect 15431 12260 15476 12288
rect 15289 12251 15347 12257
rect 15120 12220 15148 12251
rect 15470 12248 15476 12260
rect 15528 12248 15534 12300
rect 16666 12248 16672 12300
rect 16724 12248 16730 12300
rect 16758 12220 16764 12232
rect 12820 12192 15148 12220
rect 16719 12192 16764 12220
rect 16758 12180 16764 12192
rect 16816 12180 16822 12232
rect 18601 12223 18659 12229
rect 18601 12189 18613 12223
rect 18647 12220 18659 12223
rect 18782 12220 18788 12232
rect 18647 12192 18788 12220
rect 18647 12189 18659 12192
rect 18601 12183 18659 12189
rect 18782 12180 18788 12192
rect 18840 12220 18846 12232
rect 19426 12220 19432 12232
rect 18840 12192 19432 12220
rect 18840 12180 18846 12192
rect 19426 12180 19432 12192
rect 19484 12180 19490 12232
rect 5408 12124 5672 12152
rect 5408 12112 5414 12124
rect 11698 12112 11704 12164
rect 11756 12152 11762 12164
rect 11793 12155 11851 12161
rect 11793 12152 11805 12155
rect 11756 12124 11805 12152
rect 11756 12112 11762 12124
rect 11793 12121 11805 12124
rect 11839 12152 11851 12155
rect 12066 12152 12072 12164
rect 11839 12124 12072 12152
rect 11839 12121 11851 12124
rect 11793 12115 11851 12121
rect 12066 12112 12072 12124
rect 12124 12112 12130 12164
rect 17126 12112 17132 12164
rect 17184 12152 17190 12164
rect 19153 12155 19211 12161
rect 19153 12152 19165 12155
rect 17184 12124 19165 12152
rect 17184 12112 17190 12124
rect 19153 12121 19165 12124
rect 19199 12121 19211 12155
rect 19153 12115 19211 12121
rect 2038 12044 2044 12096
rect 2096 12084 2102 12096
rect 2225 12087 2283 12093
rect 2225 12084 2237 12087
rect 2096 12056 2237 12084
rect 2096 12044 2102 12056
rect 2225 12053 2237 12056
rect 2271 12053 2283 12087
rect 2225 12047 2283 12053
rect 3513 12087 3571 12093
rect 3513 12053 3525 12087
rect 3559 12084 3571 12087
rect 4062 12084 4068 12096
rect 3559 12056 4068 12084
rect 3559 12053 3571 12056
rect 3513 12047 3571 12053
rect 4062 12044 4068 12056
rect 4120 12044 4126 12096
rect 7282 12044 7288 12096
rect 7340 12084 7346 12096
rect 8297 12087 8355 12093
rect 8297 12084 8309 12087
rect 7340 12056 8309 12084
rect 7340 12044 7346 12056
rect 8297 12053 8309 12056
rect 8343 12084 8355 12087
rect 9122 12084 9128 12096
rect 8343 12056 9128 12084
rect 8343 12053 8355 12056
rect 8297 12047 8355 12053
rect 9122 12044 9128 12056
rect 9180 12044 9186 12096
rect 13538 12044 13544 12096
rect 13596 12084 13602 12096
rect 15286 12084 15292 12096
rect 13596 12056 15292 12084
rect 13596 12044 13602 12056
rect 15286 12044 15292 12056
rect 15344 12044 15350 12096
rect 15654 12044 15660 12096
rect 15712 12084 15718 12096
rect 16117 12087 16175 12093
rect 16117 12084 16129 12087
rect 15712 12056 16129 12084
rect 15712 12044 15718 12056
rect 16117 12053 16129 12056
rect 16163 12053 16175 12087
rect 16117 12047 16175 12053
rect 18141 12087 18199 12093
rect 18141 12053 18153 12087
rect 18187 12084 18199 12087
rect 18230 12084 18236 12096
rect 18187 12056 18236 12084
rect 18187 12053 18199 12056
rect 18141 12047 18199 12053
rect 18230 12044 18236 12056
rect 18288 12044 18294 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1578 11880 1584 11892
rect 1539 11852 1584 11880
rect 1578 11840 1584 11852
rect 1636 11840 1642 11892
rect 5534 11880 5540 11892
rect 5447 11852 5540 11880
rect 5534 11840 5540 11852
rect 5592 11880 5598 11892
rect 6270 11880 6276 11892
rect 5592 11852 6276 11880
rect 5592 11840 5598 11852
rect 6270 11840 6276 11852
rect 6328 11840 6334 11892
rect 7282 11880 7288 11892
rect 7243 11852 7288 11880
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 7650 11880 7656 11892
rect 7611 11852 7656 11880
rect 7650 11840 7656 11852
rect 7708 11840 7714 11892
rect 9858 11880 9864 11892
rect 9819 11852 9864 11880
rect 9858 11840 9864 11852
rect 9916 11840 9922 11892
rect 13538 11880 13544 11892
rect 13499 11852 13544 11880
rect 13538 11840 13544 11852
rect 13596 11840 13602 11892
rect 19058 11880 19064 11892
rect 19019 11852 19064 11880
rect 19058 11840 19064 11852
rect 19116 11840 19122 11892
rect 19334 11840 19340 11892
rect 19392 11880 19398 11892
rect 19429 11883 19487 11889
rect 19429 11880 19441 11883
rect 19392 11852 19441 11880
rect 19392 11840 19398 11852
rect 19429 11849 19441 11852
rect 19475 11849 19487 11883
rect 19794 11880 19800 11892
rect 19755 11852 19800 11880
rect 19429 11843 19487 11849
rect 19794 11840 19800 11852
rect 19852 11840 19858 11892
rect 4154 11772 4160 11824
rect 4212 11812 4218 11824
rect 4525 11815 4583 11821
rect 4525 11812 4537 11815
rect 4212 11784 4537 11812
rect 4212 11772 4218 11784
rect 4525 11781 4537 11784
rect 4571 11781 4583 11815
rect 5902 11812 5908 11824
rect 5815 11784 5908 11812
rect 4525 11775 4583 11781
rect 5902 11772 5908 11784
rect 5960 11812 5966 11824
rect 7926 11812 7932 11824
rect 5960 11784 7932 11812
rect 5960 11772 5966 11784
rect 7926 11772 7932 11784
rect 7984 11772 7990 11824
rect 12434 11772 12440 11824
rect 12492 11812 12498 11824
rect 12529 11815 12587 11821
rect 12529 11812 12541 11815
rect 12492 11784 12541 11812
rect 12492 11772 12498 11784
rect 12529 11781 12541 11784
rect 12575 11781 12587 11815
rect 12529 11775 12587 11781
rect 2041 11747 2099 11753
rect 2041 11713 2053 11747
rect 2087 11744 2099 11747
rect 2222 11744 2228 11756
rect 2087 11716 2228 11744
rect 2087 11713 2099 11716
rect 2041 11707 2099 11713
rect 2222 11704 2228 11716
rect 2280 11744 2286 11756
rect 2593 11747 2651 11753
rect 2593 11744 2605 11747
rect 2280 11716 2605 11744
rect 2280 11704 2286 11716
rect 2593 11713 2605 11716
rect 2639 11744 2651 11747
rect 2639 11716 3924 11744
rect 2639 11713 2651 11716
rect 2593 11707 2651 11713
rect 3896 11688 3924 11716
rect 5166 11704 5172 11756
rect 5224 11744 5230 11756
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 5224 11716 6561 11744
rect 5224 11704 5230 11716
rect 6549 11713 6561 11716
rect 6595 11744 6607 11747
rect 7466 11744 7472 11756
rect 6595 11716 7472 11744
rect 6595 11713 6607 11716
rect 6549 11707 6607 11713
rect 7466 11704 7472 11716
rect 7524 11704 7530 11756
rect 7558 11704 7564 11756
rect 7616 11744 7622 11756
rect 8021 11747 8079 11753
rect 8021 11744 8033 11747
rect 7616 11716 8033 11744
rect 7616 11704 7622 11716
rect 8021 11713 8033 11716
rect 8067 11744 8079 11747
rect 16301 11747 16359 11753
rect 8067 11716 9536 11744
rect 8067 11713 8079 11716
rect 8021 11707 8079 11713
rect 9508 11688 9536 11716
rect 16301 11713 16313 11747
rect 16347 11744 16359 11747
rect 16758 11744 16764 11756
rect 16347 11716 16764 11744
rect 16347 11713 16359 11716
rect 16301 11707 16359 11713
rect 16758 11704 16764 11716
rect 16816 11704 16822 11756
rect 17865 11747 17923 11753
rect 17865 11713 17877 11747
rect 17911 11744 17923 11747
rect 18141 11747 18199 11753
rect 18141 11744 18153 11747
rect 17911 11716 18153 11744
rect 17911 11713 17923 11716
rect 17865 11707 17923 11713
rect 18141 11713 18153 11716
rect 18187 11744 18199 11747
rect 18414 11744 18420 11756
rect 18187 11716 18420 11744
rect 18187 11713 18199 11716
rect 18141 11707 18199 11713
rect 18414 11704 18420 11716
rect 18472 11704 18478 11756
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 1946 11676 1952 11688
rect 1443 11648 1952 11676
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 1946 11636 1952 11648
rect 2004 11636 2010 11688
rect 2130 11636 2136 11688
rect 2188 11676 2194 11688
rect 2406 11676 2412 11688
rect 2188 11648 2412 11676
rect 2188 11636 2194 11648
rect 2406 11636 2412 11648
rect 2464 11636 2470 11688
rect 3053 11679 3111 11685
rect 3053 11645 3065 11679
rect 3099 11676 3111 11679
rect 3418 11676 3424 11688
rect 3099 11648 3424 11676
rect 3099 11645 3111 11648
rect 3053 11639 3111 11645
rect 3418 11636 3424 11648
rect 3476 11636 3482 11688
rect 3878 11676 3884 11688
rect 3839 11648 3884 11676
rect 3878 11636 3884 11648
rect 3936 11636 3942 11688
rect 4062 11676 4068 11688
rect 4023 11648 4068 11676
rect 4062 11636 4068 11648
rect 4120 11636 4126 11688
rect 4522 11676 4528 11688
rect 4483 11648 4528 11676
rect 4522 11636 4528 11648
rect 4580 11636 4586 11688
rect 4985 11679 5043 11685
rect 4985 11645 4997 11679
rect 5031 11676 5043 11679
rect 5442 11676 5448 11688
rect 5031 11648 5448 11676
rect 5031 11645 5043 11648
rect 4985 11639 5043 11645
rect 5442 11636 5448 11648
rect 5500 11636 5506 11688
rect 5721 11679 5779 11685
rect 5721 11645 5733 11679
rect 5767 11676 5779 11679
rect 7101 11679 7159 11685
rect 5767 11648 6316 11676
rect 5767 11645 5779 11648
rect 5721 11639 5779 11645
rect 6288 11552 6316 11648
rect 7101 11645 7113 11679
rect 7147 11676 7159 11679
rect 7650 11676 7656 11688
rect 7147 11648 7656 11676
rect 7147 11645 7159 11648
rect 7101 11639 7159 11645
rect 7650 11636 7656 11648
rect 7708 11636 7714 11688
rect 8294 11676 8300 11688
rect 8255 11648 8300 11676
rect 8294 11636 8300 11648
rect 8352 11636 8358 11688
rect 8570 11676 8576 11688
rect 8531 11648 8576 11676
rect 8570 11636 8576 11648
rect 8628 11636 8634 11688
rect 9122 11676 9128 11688
rect 9035 11648 9128 11676
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 9490 11676 9496 11688
rect 9451 11648 9496 11676
rect 9490 11636 9496 11648
rect 9548 11636 9554 11688
rect 10321 11679 10379 11685
rect 10321 11645 10333 11679
rect 10367 11676 10379 11679
rect 10962 11676 10968 11688
rect 10367 11648 10968 11676
rect 10367 11645 10379 11648
rect 10321 11639 10379 11645
rect 10962 11636 10968 11648
rect 11020 11636 11026 11688
rect 12437 11679 12495 11685
rect 12437 11645 12449 11679
rect 12483 11676 12495 11679
rect 12710 11676 12716 11688
rect 12483 11648 12517 11676
rect 12671 11648 12716 11676
rect 12483 11645 12495 11648
rect 12437 11639 12495 11645
rect 8754 11568 8760 11620
rect 8812 11608 8818 11620
rect 9140 11608 9168 11636
rect 9950 11608 9956 11620
rect 8812 11580 9956 11608
rect 8812 11568 8818 11580
rect 9950 11568 9956 11580
rect 10008 11568 10014 11620
rect 11698 11568 11704 11620
rect 11756 11608 11762 11620
rect 12161 11611 12219 11617
rect 12161 11608 12173 11611
rect 11756 11580 12173 11608
rect 11756 11568 11762 11580
rect 12161 11577 12173 11580
rect 12207 11608 12219 11611
rect 12452 11608 12480 11639
rect 12710 11636 12716 11648
rect 12768 11636 12774 11688
rect 13909 11679 13967 11685
rect 13909 11645 13921 11679
rect 13955 11676 13967 11679
rect 14645 11679 14703 11685
rect 14645 11676 14657 11679
rect 13955 11648 14657 11676
rect 13955 11645 13967 11648
rect 13909 11639 13967 11645
rect 14645 11645 14657 11648
rect 14691 11676 14703 11679
rect 14918 11676 14924 11688
rect 14691 11648 14924 11676
rect 14691 11645 14703 11648
rect 14645 11639 14703 11645
rect 14918 11636 14924 11648
rect 14976 11636 14982 11688
rect 15654 11676 15660 11688
rect 15615 11648 15660 11676
rect 15654 11636 15660 11648
rect 15712 11636 15718 11688
rect 15838 11636 15844 11688
rect 15896 11676 15902 11688
rect 16025 11679 16083 11685
rect 16025 11676 16037 11679
rect 15896 11648 16037 11676
rect 15896 11636 15902 11648
rect 16025 11645 16037 11648
rect 16071 11676 16083 11679
rect 17129 11679 17187 11685
rect 17129 11676 17141 11679
rect 16071 11648 17141 11676
rect 16071 11645 16083 11648
rect 16025 11639 16083 11645
rect 17129 11645 17141 11648
rect 17175 11645 17187 11679
rect 18046 11676 18052 11688
rect 18007 11648 18052 11676
rect 17129 11639 17187 11645
rect 18046 11636 18052 11648
rect 18104 11636 18110 11688
rect 18230 11636 18236 11688
rect 18288 11676 18294 11688
rect 18325 11679 18383 11685
rect 18325 11676 18337 11679
rect 18288 11648 18337 11676
rect 18288 11636 18294 11648
rect 18325 11645 18337 11648
rect 18371 11645 18383 11679
rect 19610 11676 19616 11688
rect 19571 11648 19616 11676
rect 18325 11639 18383 11645
rect 19610 11636 19616 11648
rect 19668 11676 19674 11688
rect 20073 11679 20131 11685
rect 20073 11676 20085 11679
rect 19668 11648 20085 11676
rect 19668 11636 19674 11648
rect 20073 11645 20085 11648
rect 20119 11645 20131 11679
rect 20073 11639 20131 11645
rect 13170 11608 13176 11620
rect 12207 11580 13176 11608
rect 12207 11577 12219 11580
rect 12161 11571 12219 11577
rect 13170 11568 13176 11580
rect 13228 11568 13234 11620
rect 14734 11608 14740 11620
rect 14695 11580 14740 11608
rect 14734 11568 14740 11580
rect 14792 11568 14798 11620
rect 18785 11611 18843 11617
rect 18785 11577 18797 11611
rect 18831 11608 18843 11611
rect 19242 11608 19248 11620
rect 18831 11580 19248 11608
rect 18831 11577 18843 11580
rect 18785 11571 18843 11577
rect 19242 11568 19248 11580
rect 19300 11568 19306 11620
rect 6270 11540 6276 11552
rect 6231 11512 6276 11540
rect 6270 11500 6276 11512
rect 6328 11500 6334 11552
rect 8389 11543 8447 11549
rect 8389 11509 8401 11543
rect 8435 11540 8447 11543
rect 8662 11540 8668 11552
rect 8435 11512 8668 11540
rect 8435 11509 8447 11512
rect 8389 11503 8447 11509
rect 8662 11500 8668 11512
rect 8720 11500 8726 11552
rect 10686 11540 10692 11552
rect 10647 11512 10692 11540
rect 10686 11500 10692 11512
rect 10744 11500 10750 11552
rect 11793 11543 11851 11549
rect 11793 11509 11805 11543
rect 11839 11540 11851 11543
rect 12066 11540 12072 11552
rect 11839 11512 12072 11540
rect 11839 11509 11851 11512
rect 11793 11503 11851 11509
rect 12066 11500 12072 11512
rect 12124 11500 12130 11552
rect 12894 11540 12900 11552
rect 12855 11512 12900 11540
rect 12894 11500 12900 11512
rect 12952 11500 12958 11552
rect 15381 11543 15439 11549
rect 15381 11509 15393 11543
rect 15427 11540 15439 11543
rect 15470 11540 15476 11552
rect 15427 11512 15476 11540
rect 15427 11509 15439 11512
rect 15381 11503 15439 11509
rect 15470 11500 15476 11512
rect 15528 11540 15534 11552
rect 16298 11540 16304 11552
rect 15528 11512 16304 11540
rect 15528 11500 15534 11512
rect 16298 11500 16304 11512
rect 16356 11500 16362 11552
rect 16666 11500 16672 11552
rect 16724 11540 16730 11552
rect 16761 11543 16819 11549
rect 16761 11540 16773 11543
rect 16724 11512 16773 11540
rect 16724 11500 16730 11512
rect 16761 11509 16773 11512
rect 16807 11509 16819 11543
rect 16761 11503 16819 11509
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 2406 11296 2412 11348
rect 2464 11336 2470 11348
rect 2869 11339 2927 11345
rect 2869 11336 2881 11339
rect 2464 11308 2881 11336
rect 2464 11296 2470 11308
rect 2869 11305 2881 11308
rect 2915 11305 2927 11339
rect 2869 11299 2927 11305
rect 3881 11339 3939 11345
rect 3881 11305 3893 11339
rect 3927 11336 3939 11339
rect 4522 11336 4528 11348
rect 3927 11308 4528 11336
rect 3927 11305 3939 11308
rect 3881 11299 3939 11305
rect 4522 11296 4528 11308
rect 4580 11296 4586 11348
rect 5350 11336 5356 11348
rect 5311 11308 5356 11336
rect 5350 11296 5356 11308
rect 5408 11296 5414 11348
rect 5813 11339 5871 11345
rect 5813 11305 5825 11339
rect 5859 11336 5871 11339
rect 5994 11336 6000 11348
rect 5859 11308 6000 11336
rect 5859 11305 5871 11308
rect 5813 11299 5871 11305
rect 5994 11296 6000 11308
rect 6052 11296 6058 11348
rect 8570 11296 8576 11348
rect 8628 11336 8634 11348
rect 9401 11339 9459 11345
rect 9401 11336 9413 11339
rect 8628 11308 9413 11336
rect 8628 11296 8634 11308
rect 9401 11305 9413 11308
rect 9447 11305 9459 11339
rect 9401 11299 9459 11305
rect 9953 11339 10011 11345
rect 9953 11305 9965 11339
rect 9999 11336 10011 11339
rect 10134 11336 10140 11348
rect 9999 11308 10140 11336
rect 9999 11305 10011 11308
rect 9953 11299 10011 11305
rect 3418 11268 3424 11280
rect 1964 11240 3424 11268
rect 1762 11160 1768 11212
rect 1820 11200 1826 11212
rect 1964 11209 1992 11240
rect 3418 11228 3424 11240
rect 3476 11228 3482 11280
rect 5368 11268 5396 11296
rect 7837 11271 7895 11277
rect 7837 11268 7849 11271
rect 5368 11240 7849 11268
rect 1949 11203 2007 11209
rect 1949 11200 1961 11203
rect 1820 11172 1961 11200
rect 1820 11160 1826 11172
rect 1949 11169 1961 11172
rect 1995 11169 2007 11203
rect 2222 11200 2228 11212
rect 2183 11172 2228 11200
rect 1949 11163 2007 11169
rect 2222 11160 2228 11172
rect 2280 11160 2286 11212
rect 2682 11200 2688 11212
rect 2643 11172 2688 11200
rect 2682 11160 2688 11172
rect 2740 11160 2746 11212
rect 2866 11200 2872 11212
rect 2827 11172 2872 11200
rect 2866 11160 2872 11172
rect 2924 11160 2930 11212
rect 4525 11203 4583 11209
rect 4525 11169 4537 11203
rect 4571 11200 4583 11203
rect 4614 11200 4620 11212
rect 4571 11172 4620 11200
rect 4571 11169 4583 11172
rect 4525 11163 4583 11169
rect 4614 11160 4620 11172
rect 4672 11200 4678 11212
rect 5368 11200 5396 11240
rect 7837 11237 7849 11240
rect 7883 11237 7895 11271
rect 7837 11231 7895 11237
rect 4672 11172 5396 11200
rect 5813 11203 5871 11209
rect 4672 11160 4678 11172
rect 5813 11169 5825 11203
rect 5859 11200 5871 11203
rect 5994 11200 6000 11212
rect 5859 11172 6000 11200
rect 5859 11169 5871 11172
rect 5813 11163 5871 11169
rect 5994 11160 6000 11172
rect 6052 11160 6058 11212
rect 6178 11200 6184 11212
rect 6139 11172 6184 11200
rect 6178 11160 6184 11172
rect 6236 11160 6242 11212
rect 6362 11200 6368 11212
rect 6323 11172 6368 11200
rect 6362 11160 6368 11172
rect 6420 11160 6426 11212
rect 6546 11160 6552 11212
rect 6604 11200 6610 11212
rect 6917 11203 6975 11209
rect 6917 11200 6929 11203
rect 6604 11172 6929 11200
rect 6604 11160 6610 11172
rect 6917 11169 6929 11172
rect 6963 11200 6975 11203
rect 7558 11200 7564 11212
rect 6963 11172 7564 11200
rect 6963 11169 6975 11172
rect 6917 11163 6975 11169
rect 7558 11160 7564 11172
rect 7616 11160 7622 11212
rect 7926 11160 7932 11212
rect 7984 11200 7990 11212
rect 8481 11203 8539 11209
rect 8481 11200 8493 11203
rect 7984 11172 8493 11200
rect 7984 11160 7990 11172
rect 8481 11169 8493 11172
rect 8527 11200 8539 11203
rect 9968 11200 9996 11299
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 11054 11296 11060 11348
rect 11112 11336 11118 11348
rect 12161 11339 12219 11345
rect 12161 11336 12173 11339
rect 11112 11308 12173 11336
rect 11112 11296 11118 11308
rect 12161 11305 12173 11308
rect 12207 11305 12219 11339
rect 12710 11336 12716 11348
rect 12671 11308 12716 11336
rect 12161 11299 12219 11305
rect 12710 11296 12716 11308
rect 12768 11296 12774 11348
rect 13170 11296 13176 11348
rect 13228 11336 13234 11348
rect 13265 11339 13323 11345
rect 13265 11336 13277 11339
rect 13228 11308 13277 11336
rect 13228 11296 13234 11308
rect 13265 11305 13277 11308
rect 13311 11305 13323 11339
rect 13265 11299 13323 11305
rect 16850 11296 16856 11348
rect 16908 11336 16914 11348
rect 17313 11339 17371 11345
rect 17313 11336 17325 11339
rect 16908 11308 17325 11336
rect 16908 11296 16914 11308
rect 17313 11305 17325 11308
rect 17359 11305 17371 11339
rect 19426 11336 19432 11348
rect 19387 11308 19432 11336
rect 17313 11299 17371 11305
rect 19426 11296 19432 11308
rect 19484 11296 19490 11348
rect 14366 11268 14372 11280
rect 14327 11240 14372 11268
rect 14366 11228 14372 11240
rect 14424 11228 14430 11280
rect 14826 11268 14832 11280
rect 14568 11240 14832 11268
rect 8527 11172 9996 11200
rect 10045 11203 10103 11209
rect 8527 11169 8539 11172
rect 8481 11163 8539 11169
rect 10045 11169 10057 11203
rect 10091 11200 10103 11203
rect 10137 11203 10195 11209
rect 10137 11200 10149 11203
rect 10091 11172 10149 11200
rect 10091 11169 10103 11172
rect 10045 11163 10103 11169
rect 10137 11169 10149 11172
rect 10183 11169 10195 11203
rect 10137 11163 10195 11169
rect 10413 11203 10471 11209
rect 10413 11169 10425 11203
rect 10459 11200 10471 11203
rect 10962 11200 10968 11212
rect 10459 11172 10968 11200
rect 10459 11169 10471 11172
rect 10413 11163 10471 11169
rect 10962 11160 10968 11172
rect 11020 11160 11026 11212
rect 11698 11200 11704 11212
rect 11532 11172 11704 11200
rect 2884 11132 2912 11160
rect 2884 11104 4108 11132
rect 3513 11067 3571 11073
rect 3513 11033 3525 11067
rect 3559 11064 3571 11067
rect 3878 11064 3884 11076
rect 3559 11036 3884 11064
rect 3559 11033 3571 11036
rect 3513 11027 3571 11033
rect 3878 11024 3884 11036
rect 3936 11024 3942 11076
rect 4080 10996 4108 11104
rect 5350 11092 5356 11144
rect 5408 11132 5414 11144
rect 6196 11132 6224 11160
rect 5408 11104 6224 11132
rect 5408 11092 5414 11104
rect 9674 11092 9680 11144
rect 9732 11132 9738 11144
rect 10229 11135 10287 11141
rect 10229 11132 10241 11135
rect 9732 11104 10241 11132
rect 9732 11092 9738 11104
rect 10229 11101 10241 11104
rect 10275 11132 10287 11135
rect 10686 11132 10692 11144
rect 10275 11104 10692 11132
rect 10275 11101 10287 11104
rect 10229 11095 10287 11101
rect 10686 11092 10692 11104
rect 10744 11092 10750 11144
rect 10870 11132 10876 11144
rect 10831 11104 10876 11132
rect 10870 11092 10876 11104
rect 10928 11092 10934 11144
rect 4246 11064 4252 11076
rect 4207 11036 4252 11064
rect 4246 11024 4252 11036
rect 4304 11024 4310 11076
rect 4709 11067 4767 11073
rect 4709 11033 4721 11067
rect 4755 11064 4767 11067
rect 5077 11067 5135 11073
rect 5077 11064 5089 11067
rect 4755 11036 5089 11064
rect 4755 11033 4767 11036
rect 4709 11027 4767 11033
rect 5077 11033 5089 11036
rect 5123 11064 5135 11067
rect 6086 11064 6092 11076
rect 5123 11036 6092 11064
rect 5123 11033 5135 11036
rect 5077 11027 5135 11033
rect 6086 11024 6092 11036
rect 6144 11024 6150 11076
rect 9950 11024 9956 11076
rect 10008 11064 10014 11076
rect 10045 11067 10103 11073
rect 10045 11064 10057 11067
rect 10008 11036 10057 11064
rect 10008 11024 10014 11036
rect 10045 11033 10057 11036
rect 10091 11033 10103 11067
rect 10045 11027 10103 11033
rect 4154 10996 4160 11008
rect 4080 10968 4160 10996
rect 4154 10956 4160 10968
rect 4212 10956 4218 11008
rect 7006 10956 7012 11008
rect 7064 10996 7070 11008
rect 7653 10999 7711 11005
rect 7653 10996 7665 10999
rect 7064 10968 7665 10996
rect 7064 10956 7070 10968
rect 7653 10965 7665 10968
rect 7699 10996 7711 10999
rect 8662 10996 8668 11008
rect 7699 10968 8668 10996
rect 7699 10965 7711 10968
rect 7653 10959 7711 10965
rect 8662 10956 8668 10968
rect 8720 10956 8726 11008
rect 8938 10996 8944 11008
rect 8899 10968 8944 10996
rect 8938 10956 8944 10968
rect 8996 10956 9002 11008
rect 11422 10956 11428 11008
rect 11480 10996 11486 11008
rect 11532 11005 11560 11172
rect 11698 11160 11704 11172
rect 11756 11160 11762 11212
rect 11974 11200 11980 11212
rect 11935 11172 11980 11200
rect 11974 11160 11980 11172
rect 12032 11160 12038 11212
rect 13630 11200 13636 11212
rect 13591 11172 13636 11200
rect 13630 11160 13636 11172
rect 13688 11160 13694 11212
rect 13909 11203 13967 11209
rect 13909 11169 13921 11203
rect 13955 11200 13967 11203
rect 13998 11200 14004 11212
rect 13955 11172 14004 11200
rect 13955 11169 13967 11172
rect 13909 11163 13967 11169
rect 13998 11160 14004 11172
rect 14056 11200 14062 11212
rect 14568 11200 14596 11240
rect 14826 11228 14832 11240
rect 14884 11228 14890 11280
rect 16025 11271 16083 11277
rect 16025 11237 16037 11271
rect 16071 11268 16083 11271
rect 16482 11268 16488 11280
rect 16071 11240 16488 11268
rect 16071 11237 16083 11240
rect 16025 11231 16083 11237
rect 16482 11228 16488 11240
rect 16540 11228 16546 11280
rect 14056 11172 14596 11200
rect 14056 11160 14062 11172
rect 14642 11160 14648 11212
rect 14700 11200 14706 11212
rect 15289 11203 15347 11209
rect 15289 11200 15301 11203
rect 14700 11172 15301 11200
rect 14700 11160 14706 11172
rect 15289 11169 15301 11172
rect 15335 11169 15347 11203
rect 15289 11163 15347 11169
rect 15378 11160 15384 11212
rect 15436 11200 15442 11212
rect 15565 11203 15623 11209
rect 15565 11200 15577 11203
rect 15436 11172 15577 11200
rect 15436 11160 15442 11172
rect 15565 11169 15577 11172
rect 15611 11169 15623 11203
rect 16850 11200 16856 11212
rect 16811 11172 16856 11200
rect 15565 11163 15623 11169
rect 13725 11135 13783 11141
rect 13725 11101 13737 11135
rect 13771 11132 13783 11135
rect 13814 11132 13820 11144
rect 13771 11104 13820 11132
rect 13771 11101 13783 11104
rect 13725 11095 13783 11101
rect 13814 11092 13820 11104
rect 13872 11132 13878 11144
rect 14734 11132 14740 11144
rect 13872 11104 14740 11132
rect 13872 11092 13878 11104
rect 14734 11092 14740 11104
rect 14792 11092 14798 11144
rect 15580 11132 15608 11163
rect 16850 11160 16856 11172
rect 16908 11160 16914 11212
rect 17126 11200 17132 11212
rect 17087 11172 17132 11200
rect 17126 11160 17132 11172
rect 17184 11160 17190 11212
rect 18046 11200 18052 11212
rect 18007 11172 18052 11200
rect 18046 11160 18052 11172
rect 18104 11160 18110 11212
rect 18966 11200 18972 11212
rect 18927 11172 18972 11200
rect 18966 11160 18972 11172
rect 19024 11160 19030 11212
rect 18230 11132 18236 11144
rect 15580 11104 18236 11132
rect 18230 11092 18236 11104
rect 18288 11132 18294 11144
rect 18417 11135 18475 11141
rect 18417 11132 18429 11135
rect 18288 11104 18429 11132
rect 18288 11092 18294 11104
rect 18417 11101 18429 11104
rect 18463 11101 18475 11135
rect 18417 11095 18475 11101
rect 11793 11067 11851 11073
rect 11793 11033 11805 11067
rect 11839 11064 11851 11067
rect 12066 11064 12072 11076
rect 11839 11036 12072 11064
rect 11839 11033 11851 11036
rect 11793 11027 11851 11033
rect 12066 11024 12072 11036
rect 12124 11024 12130 11076
rect 14918 11024 14924 11076
rect 14976 11064 14982 11076
rect 15381 11067 15439 11073
rect 15381 11064 15393 11067
rect 14976 11036 15393 11064
rect 14976 11024 14982 11036
rect 15381 11033 15393 11036
rect 15427 11064 15439 11067
rect 15930 11064 15936 11076
rect 15427 11036 15936 11064
rect 15427 11033 15439 11036
rect 15381 11027 15439 11033
rect 15930 11024 15936 11036
rect 15988 11024 15994 11076
rect 16942 11064 16948 11076
rect 16903 11036 16948 11064
rect 16942 11024 16948 11036
rect 17000 11024 17006 11076
rect 11517 10999 11575 11005
rect 11517 10996 11529 10999
rect 11480 10968 11529 10996
rect 11480 10956 11486 10968
rect 11517 10965 11529 10968
rect 11563 10965 11575 10999
rect 11517 10959 11575 10965
rect 14550 10956 14556 11008
rect 14608 10996 14614 11008
rect 14829 10999 14887 11005
rect 14829 10996 14841 10999
rect 14608 10968 14841 10996
rect 14608 10956 14614 10968
rect 14829 10965 14841 10968
rect 14875 10965 14887 10999
rect 16482 10996 16488 11008
rect 16443 10968 16488 10996
rect 14829 10959 14887 10965
rect 16482 10956 16488 10968
rect 16540 10956 16546 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 3878 10752 3884 10804
rect 3936 10792 3942 10804
rect 5261 10795 5319 10801
rect 5261 10792 5273 10795
rect 3936 10764 5273 10792
rect 3936 10752 3942 10764
rect 5261 10761 5273 10764
rect 5307 10792 5319 10795
rect 5350 10792 5356 10804
rect 5307 10764 5356 10792
rect 5307 10761 5319 10764
rect 5261 10755 5319 10761
rect 5350 10752 5356 10764
rect 5408 10752 5414 10804
rect 6273 10795 6331 10801
rect 6273 10761 6285 10795
rect 6319 10792 6331 10795
rect 6362 10792 6368 10804
rect 6319 10764 6368 10792
rect 6319 10761 6331 10764
rect 6273 10755 6331 10761
rect 6362 10752 6368 10764
rect 6420 10752 6426 10804
rect 6638 10792 6644 10804
rect 6599 10764 6644 10792
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 7098 10792 7104 10804
rect 7059 10764 7104 10792
rect 7098 10752 7104 10764
rect 7156 10752 7162 10804
rect 9401 10795 9459 10801
rect 9401 10761 9413 10795
rect 9447 10792 9459 10795
rect 9582 10792 9588 10804
rect 9447 10764 9588 10792
rect 9447 10761 9459 10764
rect 9401 10755 9459 10761
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 9769 10795 9827 10801
rect 9769 10761 9781 10795
rect 9815 10792 9827 10795
rect 9950 10792 9956 10804
rect 9815 10764 9956 10792
rect 9815 10761 9827 10764
rect 9769 10755 9827 10761
rect 9950 10752 9956 10764
rect 10008 10752 10014 10804
rect 10962 10792 10968 10804
rect 10923 10764 10968 10792
rect 10962 10752 10968 10764
rect 11020 10752 11026 10804
rect 11422 10792 11428 10804
rect 11383 10764 11428 10792
rect 11422 10752 11428 10764
rect 11480 10752 11486 10804
rect 11793 10795 11851 10801
rect 11793 10761 11805 10795
rect 11839 10792 11851 10795
rect 11974 10792 11980 10804
rect 11839 10764 11980 10792
rect 11839 10761 11851 10764
rect 11793 10755 11851 10761
rect 11974 10752 11980 10764
rect 12032 10752 12038 10804
rect 12066 10752 12072 10804
rect 12124 10792 12130 10804
rect 12124 10764 12169 10792
rect 12124 10752 12130 10764
rect 13630 10752 13636 10804
rect 13688 10792 13694 10804
rect 14001 10795 14059 10801
rect 14001 10792 14013 10795
rect 13688 10764 14013 10792
rect 13688 10752 13694 10764
rect 14001 10761 14013 10764
rect 14047 10761 14059 10795
rect 14001 10755 14059 10761
rect 3896 10656 3924 10752
rect 14016 10724 14044 10755
rect 14182 10752 14188 10804
rect 14240 10792 14246 10804
rect 14642 10792 14648 10804
rect 14240 10764 14648 10792
rect 14240 10752 14246 10764
rect 14642 10752 14648 10764
rect 14700 10792 14706 10804
rect 15470 10792 15476 10804
rect 14700 10764 15476 10792
rect 14700 10752 14706 10764
rect 15470 10752 15476 10764
rect 15528 10792 15534 10804
rect 16209 10795 16267 10801
rect 16209 10792 16221 10795
rect 15528 10764 16221 10792
rect 15528 10752 15534 10764
rect 16209 10761 16221 10764
rect 16255 10792 16267 10795
rect 16850 10792 16856 10804
rect 16255 10764 16856 10792
rect 16255 10761 16267 10764
rect 16209 10755 16267 10761
rect 16850 10752 16856 10764
rect 16908 10752 16914 10804
rect 19334 10792 19340 10804
rect 19295 10764 19340 10792
rect 19334 10752 19340 10764
rect 19392 10752 19398 10804
rect 15378 10724 15384 10736
rect 14016 10696 15384 10724
rect 15378 10684 15384 10696
rect 15436 10684 15442 10736
rect 15930 10724 15936 10736
rect 15843 10696 15936 10724
rect 15930 10684 15936 10696
rect 15988 10724 15994 10736
rect 17402 10724 17408 10736
rect 15988 10696 17408 10724
rect 15988 10684 15994 10696
rect 17402 10684 17408 10696
rect 17460 10684 17466 10736
rect 3804 10628 3924 10656
rect 2038 10588 2044 10600
rect 1999 10560 2044 10588
rect 2038 10548 2044 10560
rect 2096 10548 2102 10600
rect 2961 10591 3019 10597
rect 2961 10557 2973 10591
rect 3007 10588 3019 10591
rect 3329 10591 3387 10597
rect 3329 10588 3341 10591
rect 3007 10560 3341 10588
rect 3007 10557 3019 10560
rect 2961 10551 3019 10557
rect 3329 10557 3341 10560
rect 3375 10588 3387 10591
rect 3418 10588 3424 10600
rect 3375 10560 3424 10588
rect 3375 10557 3387 10560
rect 3329 10551 3387 10557
rect 3418 10548 3424 10560
rect 3476 10548 3482 10600
rect 3804 10597 3832 10628
rect 6270 10616 6276 10668
rect 6328 10656 6334 10668
rect 8294 10656 8300 10668
rect 6328 10628 8300 10656
rect 6328 10616 6334 10628
rect 3789 10591 3847 10597
rect 3789 10557 3801 10591
rect 3835 10557 3847 10591
rect 4062 10588 4068 10600
rect 4023 10560 4068 10588
rect 3789 10551 3847 10557
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 4154 10548 4160 10600
rect 4212 10588 4218 10600
rect 4249 10591 4307 10597
rect 4249 10588 4261 10591
rect 4212 10560 4261 10588
rect 4212 10548 4218 10560
rect 4249 10557 4261 10560
rect 4295 10588 4307 10591
rect 4801 10591 4859 10597
rect 4801 10588 4813 10591
rect 4295 10560 4813 10588
rect 4295 10557 4307 10560
rect 4249 10551 4307 10557
rect 4801 10557 4813 10560
rect 4847 10588 4859 10591
rect 5258 10588 5264 10600
rect 4847 10560 5264 10588
rect 4847 10557 4859 10560
rect 4801 10551 4859 10557
rect 5258 10548 5264 10560
rect 5316 10548 5322 10600
rect 5721 10591 5779 10597
rect 5721 10557 5733 10591
rect 5767 10588 5779 10591
rect 6638 10588 6644 10600
rect 5767 10560 6644 10588
rect 5767 10557 5779 10560
rect 5721 10551 5779 10557
rect 6638 10548 6644 10560
rect 6696 10548 6702 10600
rect 7852 10597 7880 10628
rect 8294 10616 8300 10628
rect 8352 10656 8358 10668
rect 8938 10656 8944 10668
rect 8352 10628 8944 10656
rect 8352 10616 8358 10628
rect 8938 10616 8944 10628
rect 8996 10616 9002 10668
rect 13170 10656 13176 10668
rect 13131 10628 13176 10656
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 13725 10659 13783 10665
rect 13725 10625 13737 10659
rect 13771 10656 13783 10659
rect 13998 10656 14004 10668
rect 13771 10628 14004 10656
rect 13771 10625 13783 10628
rect 13725 10619 13783 10625
rect 13998 10616 14004 10628
rect 14056 10616 14062 10668
rect 16298 10616 16304 10668
rect 16356 10656 16362 10668
rect 17865 10659 17923 10665
rect 17865 10656 17877 10659
rect 16356 10628 17877 10656
rect 16356 10616 16362 10628
rect 17865 10625 17877 10628
rect 17911 10656 17923 10659
rect 17911 10628 18276 10656
rect 17911 10625 17923 10628
rect 17865 10619 17923 10625
rect 7837 10591 7895 10597
rect 7837 10557 7849 10591
rect 7883 10557 7895 10591
rect 8202 10588 8208 10600
rect 8163 10560 8208 10588
rect 7837 10551 7895 10557
rect 8202 10548 8208 10560
rect 8260 10548 8266 10600
rect 8573 10591 8631 10597
rect 8573 10557 8585 10591
rect 8619 10588 8631 10591
rect 8662 10588 8668 10600
rect 8619 10560 8668 10588
rect 8619 10557 8631 10560
rect 8573 10551 8631 10557
rect 8662 10548 8668 10560
rect 8720 10548 8726 10600
rect 8757 10591 8815 10597
rect 8757 10557 8769 10591
rect 8803 10557 8815 10591
rect 9950 10588 9956 10600
rect 9911 10560 9956 10588
rect 8757 10551 8815 10557
rect 1397 10523 1455 10529
rect 1397 10489 1409 10523
rect 1443 10520 1455 10523
rect 1486 10520 1492 10532
rect 1443 10492 1492 10520
rect 1443 10489 1455 10492
rect 1397 10483 1455 10489
rect 1486 10480 1492 10492
rect 1544 10480 1550 10532
rect 5629 10523 5687 10529
rect 5629 10489 5641 10523
rect 5675 10520 5687 10523
rect 5994 10520 6000 10532
rect 5675 10492 6000 10520
rect 5675 10489 5687 10492
rect 5629 10483 5687 10489
rect 5994 10480 6000 10492
rect 6052 10520 6058 10532
rect 6546 10520 6552 10532
rect 6052 10492 6552 10520
rect 6052 10480 6058 10492
rect 6546 10480 6552 10492
rect 6604 10480 6610 10532
rect 6730 10480 6736 10532
rect 6788 10520 6794 10532
rect 7469 10523 7527 10529
rect 7469 10520 7481 10523
rect 6788 10492 7481 10520
rect 6788 10480 6794 10492
rect 7469 10489 7481 10492
rect 7515 10520 7527 10523
rect 8220 10520 8248 10548
rect 7515 10492 8248 10520
rect 7515 10489 7527 10492
rect 7469 10483 7527 10489
rect 8294 10480 8300 10532
rect 8352 10520 8358 10532
rect 8772 10520 8800 10551
rect 9950 10548 9956 10560
rect 10008 10548 10014 10600
rect 12986 10588 12992 10600
rect 12947 10560 12992 10588
rect 12986 10548 12992 10560
rect 13044 10548 13050 10600
rect 14550 10548 14556 10600
rect 14608 10588 14614 10600
rect 15010 10588 15016 10600
rect 14608 10560 15016 10588
rect 14608 10548 14614 10560
rect 15010 10548 15016 10560
rect 15068 10548 15074 10600
rect 15289 10591 15347 10597
rect 15289 10557 15301 10591
rect 15335 10557 15347 10591
rect 16390 10588 16396 10600
rect 16351 10560 16396 10588
rect 15289 10551 15347 10557
rect 9030 10520 9036 10532
rect 8352 10492 8800 10520
rect 8991 10492 9036 10520
rect 8352 10480 8358 10492
rect 9030 10480 9036 10492
rect 9088 10480 9094 10532
rect 9858 10520 9864 10532
rect 9819 10492 9864 10520
rect 9858 10480 9864 10492
rect 9916 10480 9922 10532
rect 13722 10480 13728 10532
rect 13780 10520 13786 10532
rect 14568 10520 14596 10548
rect 13780 10492 14596 10520
rect 13780 10480 13786 10492
rect 14734 10480 14740 10532
rect 14792 10520 14798 10532
rect 15304 10520 15332 10551
rect 16390 10548 16396 10560
rect 16448 10548 16454 10600
rect 16482 10548 16488 10600
rect 16540 10588 16546 10600
rect 16853 10591 16911 10597
rect 16853 10588 16865 10591
rect 16540 10560 16865 10588
rect 16540 10548 16546 10560
rect 16853 10557 16865 10560
rect 16899 10557 16911 10591
rect 18046 10588 18052 10600
rect 18007 10560 18052 10588
rect 16853 10551 16911 10557
rect 18046 10548 18052 10560
rect 18104 10548 18110 10600
rect 18248 10597 18276 10628
rect 19334 10616 19340 10668
rect 19392 10656 19398 10668
rect 19392 10628 19472 10656
rect 19392 10616 19398 10628
rect 19444 10597 19472 10628
rect 18233 10591 18291 10597
rect 18233 10557 18245 10591
rect 18279 10557 18291 10591
rect 18233 10551 18291 10557
rect 19421 10591 19479 10597
rect 19421 10557 19433 10591
rect 19467 10557 19479 10591
rect 19421 10551 19479 10557
rect 15562 10520 15568 10532
rect 14792 10492 15332 10520
rect 15523 10492 15568 10520
rect 14792 10480 14798 10492
rect 15562 10480 15568 10492
rect 15620 10480 15626 10532
rect 17126 10480 17132 10532
rect 17184 10520 17190 10532
rect 17497 10523 17555 10529
rect 17497 10520 17509 10523
rect 17184 10492 17509 10520
rect 17184 10480 17190 10492
rect 17497 10489 17509 10492
rect 17543 10520 17555 10523
rect 19444 10520 19472 10551
rect 19889 10523 19947 10529
rect 19889 10520 19901 10523
rect 17543 10492 19012 10520
rect 19444 10492 19901 10520
rect 17543 10489 17555 10492
rect 17497 10483 17555 10489
rect 18984 10464 19012 10492
rect 19889 10489 19901 10492
rect 19935 10489 19947 10523
rect 19889 10483 19947 10489
rect 2501 10455 2559 10461
rect 2501 10421 2513 10455
rect 2547 10452 2559 10455
rect 2682 10452 2688 10464
rect 2547 10424 2688 10452
rect 2547 10421 2559 10424
rect 2501 10415 2559 10421
rect 2682 10412 2688 10424
rect 2740 10452 2746 10464
rect 2958 10452 2964 10464
rect 2740 10424 2964 10452
rect 2740 10412 2746 10424
rect 2958 10412 2964 10424
rect 3016 10412 3022 10464
rect 3050 10412 3056 10464
rect 3108 10452 3114 10464
rect 3145 10455 3203 10461
rect 3145 10452 3157 10455
rect 3108 10424 3157 10452
rect 3108 10412 3114 10424
rect 3145 10421 3157 10424
rect 3191 10421 3203 10455
rect 3145 10415 3203 10421
rect 5534 10412 5540 10464
rect 5592 10452 5598 10464
rect 5905 10455 5963 10461
rect 5905 10452 5917 10455
rect 5592 10424 5917 10452
rect 5592 10412 5598 10424
rect 5905 10421 5917 10424
rect 5951 10452 5963 10455
rect 7006 10452 7012 10464
rect 5951 10424 7012 10452
rect 5951 10421 5963 10424
rect 5905 10415 5963 10421
rect 7006 10412 7012 10424
rect 7064 10412 7070 10464
rect 16574 10412 16580 10464
rect 16632 10452 16638 10464
rect 16669 10455 16727 10461
rect 16669 10452 16681 10455
rect 16632 10424 16681 10452
rect 16632 10412 16638 10424
rect 16669 10421 16681 10424
rect 16715 10421 16727 10455
rect 16669 10415 16727 10421
rect 18138 10412 18144 10464
rect 18196 10452 18202 10464
rect 18325 10455 18383 10461
rect 18325 10452 18337 10455
rect 18196 10424 18337 10452
rect 18196 10412 18202 10424
rect 18325 10421 18337 10424
rect 18371 10421 18383 10455
rect 18966 10452 18972 10464
rect 18927 10424 18972 10452
rect 18325 10415 18383 10421
rect 18966 10412 18972 10424
rect 19024 10412 19030 10464
rect 19334 10412 19340 10464
rect 19392 10452 19398 10464
rect 19613 10455 19671 10461
rect 19613 10452 19625 10455
rect 19392 10424 19625 10452
rect 19392 10412 19398 10424
rect 19613 10421 19625 10424
rect 19659 10421 19671 10455
rect 19613 10415 19671 10421
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 1762 10248 1768 10260
rect 1723 10220 1768 10248
rect 1762 10208 1768 10220
rect 1820 10208 1826 10260
rect 2038 10208 2044 10260
rect 2096 10248 2102 10260
rect 3053 10251 3111 10257
rect 3053 10248 3065 10251
rect 2096 10220 3065 10248
rect 2096 10208 2102 10220
rect 3053 10217 3065 10220
rect 3099 10217 3111 10251
rect 3418 10248 3424 10260
rect 3379 10220 3424 10248
rect 3053 10211 3111 10217
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 3789 10251 3847 10257
rect 3789 10217 3801 10251
rect 3835 10248 3847 10251
rect 4062 10248 4068 10260
rect 3835 10220 4068 10248
rect 3835 10217 3847 10220
rect 3789 10211 3847 10217
rect 4062 10208 4068 10220
rect 4120 10208 4126 10260
rect 4614 10248 4620 10260
rect 4575 10220 4620 10248
rect 4614 10208 4620 10220
rect 4672 10248 4678 10260
rect 5445 10251 5503 10257
rect 5445 10248 5457 10251
rect 4672 10220 5457 10248
rect 4672 10208 4678 10220
rect 2495 10183 2553 10189
rect 2495 10149 2507 10183
rect 2541 10180 2553 10183
rect 2590 10180 2596 10192
rect 2541 10152 2596 10180
rect 2541 10149 2553 10152
rect 2495 10143 2553 10149
rect 2590 10140 2596 10152
rect 2648 10140 2654 10192
rect 5000 10121 5028 10220
rect 5445 10217 5457 10220
rect 5491 10217 5503 10251
rect 6086 10248 6092 10260
rect 6047 10220 6092 10248
rect 5445 10211 5503 10217
rect 6086 10208 6092 10220
rect 6144 10208 6150 10260
rect 7926 10248 7932 10260
rect 7887 10220 7932 10248
rect 7926 10208 7932 10220
rect 7984 10208 7990 10260
rect 8570 10208 8576 10260
rect 8628 10248 8634 10260
rect 8757 10251 8815 10257
rect 8757 10248 8769 10251
rect 8628 10220 8769 10248
rect 8628 10208 8634 10220
rect 8757 10217 8769 10220
rect 8803 10217 8815 10251
rect 11054 10248 11060 10260
rect 11015 10220 11060 10248
rect 8757 10211 8815 10217
rect 11054 10208 11060 10220
rect 11112 10208 11118 10260
rect 12434 10208 12440 10260
rect 12492 10248 12498 10260
rect 12897 10251 12955 10257
rect 12897 10248 12909 10251
rect 12492 10220 12909 10248
rect 12492 10208 12498 10220
rect 12897 10217 12909 10220
rect 12943 10217 12955 10251
rect 13814 10248 13820 10260
rect 13775 10220 13820 10248
rect 12897 10211 12955 10217
rect 13814 10208 13820 10220
rect 13872 10208 13878 10260
rect 15102 10248 15108 10260
rect 15063 10220 15108 10248
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 18046 10248 18052 10260
rect 18007 10220 18052 10248
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 18598 10248 18604 10260
rect 18559 10220 18604 10248
rect 18598 10208 18604 10220
rect 18656 10208 18662 10260
rect 9861 10183 9919 10189
rect 9861 10149 9873 10183
rect 9907 10180 9919 10183
rect 9950 10180 9956 10192
rect 9907 10152 9956 10180
rect 9907 10149 9919 10152
rect 9861 10143 9919 10149
rect 9950 10140 9956 10152
rect 10008 10180 10014 10192
rect 10689 10183 10747 10189
rect 10689 10180 10701 10183
rect 10008 10152 10701 10180
rect 10008 10140 10014 10152
rect 10689 10149 10701 10152
rect 10735 10149 10747 10183
rect 11422 10180 11428 10192
rect 11383 10152 11428 10180
rect 10689 10143 10747 10149
rect 11422 10140 11428 10152
rect 11480 10140 11486 10192
rect 14826 10140 14832 10192
rect 14884 10180 14890 10192
rect 14884 10152 15608 10180
rect 14884 10140 14890 10152
rect 4985 10115 5043 10121
rect 4985 10081 4997 10115
rect 5031 10081 5043 10115
rect 6270 10112 6276 10124
rect 6231 10084 6276 10112
rect 4985 10075 5043 10081
rect 6270 10072 6276 10084
rect 6328 10072 6334 10124
rect 6730 10112 6736 10124
rect 6691 10084 6736 10112
rect 6730 10072 6736 10084
rect 6788 10072 6794 10124
rect 7006 10112 7012 10124
rect 6967 10084 7012 10112
rect 7006 10072 7012 10084
rect 7064 10072 7070 10124
rect 7377 10115 7435 10121
rect 7377 10081 7389 10115
rect 7423 10112 7435 10115
rect 7926 10112 7932 10124
rect 7423 10084 7932 10112
rect 7423 10081 7435 10084
rect 7377 10075 7435 10081
rect 7926 10072 7932 10084
rect 7984 10072 7990 10124
rect 8573 10115 8631 10121
rect 8573 10081 8585 10115
rect 8619 10112 8631 10115
rect 8662 10112 8668 10124
rect 8619 10084 8668 10112
rect 8619 10081 8631 10084
rect 8573 10075 8631 10081
rect 8662 10072 8668 10084
rect 8720 10112 8726 10124
rect 9582 10112 9588 10124
rect 8720 10084 9588 10112
rect 8720 10072 8726 10084
rect 9582 10072 9588 10084
rect 9640 10072 9646 10124
rect 12618 10072 12624 10124
rect 12676 10112 12682 10124
rect 13081 10115 13139 10121
rect 13081 10112 13093 10115
rect 12676 10084 13093 10112
rect 12676 10072 12682 10084
rect 13081 10081 13093 10084
rect 13127 10081 13139 10115
rect 13081 10075 13139 10081
rect 13357 10115 13415 10121
rect 13357 10081 13369 10115
rect 13403 10112 13415 10115
rect 13630 10112 13636 10124
rect 13403 10084 13636 10112
rect 13403 10081 13415 10084
rect 13357 10075 13415 10081
rect 2130 10044 2136 10056
rect 2091 10016 2136 10044
rect 2130 10004 2136 10016
rect 2188 10004 2194 10056
rect 9769 10047 9827 10053
rect 9769 10044 9781 10047
rect 9416 10016 9781 10044
rect 5169 9911 5227 9917
rect 5169 9877 5181 9911
rect 5215 9908 5227 9911
rect 5350 9908 5356 9920
rect 5215 9880 5356 9908
rect 5215 9877 5227 9880
rect 5169 9871 5227 9877
rect 5350 9868 5356 9880
rect 5408 9868 5414 9920
rect 5905 9911 5963 9917
rect 5905 9877 5917 9911
rect 5951 9908 5963 9911
rect 6178 9908 6184 9920
rect 5951 9880 6184 9908
rect 5951 9877 5963 9880
rect 5905 9871 5963 9877
rect 6178 9868 6184 9880
rect 6236 9868 6242 9920
rect 8294 9908 8300 9920
rect 8255 9880 8300 9908
rect 8294 9868 8300 9880
rect 8352 9868 8358 9920
rect 8938 9868 8944 9920
rect 8996 9908 9002 9920
rect 9033 9911 9091 9917
rect 9033 9908 9045 9911
rect 8996 9880 9045 9908
rect 8996 9868 9002 9880
rect 9033 9877 9045 9880
rect 9079 9877 9091 9911
rect 9033 9871 9091 9877
rect 9122 9868 9128 9920
rect 9180 9908 9186 9920
rect 9416 9917 9444 10016
rect 9769 10013 9781 10016
rect 9815 10013 9827 10047
rect 10134 10044 10140 10056
rect 10095 10016 10140 10044
rect 9769 10007 9827 10013
rect 10134 10004 10140 10016
rect 10192 10004 10198 10056
rect 11054 10004 11060 10056
rect 11112 10044 11118 10056
rect 11333 10047 11391 10053
rect 11333 10044 11345 10047
rect 11112 10016 11345 10044
rect 11112 10004 11118 10016
rect 11333 10013 11345 10016
rect 11379 10013 11391 10047
rect 11333 10007 11391 10013
rect 11977 10047 12035 10053
rect 11977 10013 11989 10047
rect 12023 10044 12035 10047
rect 12526 10044 12532 10056
rect 12023 10016 12532 10044
rect 12023 10013 12035 10016
rect 11977 10007 12035 10013
rect 12526 10004 12532 10016
rect 12584 10004 12590 10056
rect 13096 10044 13124 10075
rect 13630 10072 13636 10084
rect 13688 10072 13694 10124
rect 15286 10112 15292 10124
rect 15247 10084 15292 10112
rect 15286 10072 15292 10084
rect 15344 10072 15350 10124
rect 15580 10121 15608 10152
rect 15565 10115 15623 10121
rect 15565 10081 15577 10115
rect 15611 10112 15623 10115
rect 15654 10112 15660 10124
rect 15611 10084 15660 10112
rect 15611 10081 15623 10084
rect 15565 10075 15623 10081
rect 15654 10072 15660 10084
rect 15712 10072 15718 10124
rect 16022 10112 16028 10124
rect 15983 10084 16028 10112
rect 16022 10072 16028 10084
rect 16080 10072 16086 10124
rect 16850 10112 16856 10124
rect 16811 10084 16856 10112
rect 16850 10072 16856 10084
rect 16908 10072 16914 10124
rect 17126 10112 17132 10124
rect 17087 10084 17132 10112
rect 17126 10072 17132 10084
rect 17184 10072 17190 10124
rect 17589 10115 17647 10121
rect 17589 10081 17601 10115
rect 17635 10112 17647 10115
rect 18414 10112 18420 10124
rect 17635 10084 18420 10112
rect 17635 10081 17647 10084
rect 17589 10075 17647 10081
rect 18414 10072 18420 10084
rect 18472 10072 18478 10124
rect 19426 10112 19432 10124
rect 19387 10084 19432 10112
rect 19426 10072 19432 10084
rect 19484 10072 19490 10124
rect 13538 10044 13544 10056
rect 13096 10016 13544 10044
rect 13538 10004 13544 10016
rect 13596 10004 13602 10056
rect 15381 10047 15439 10053
rect 15381 10013 15393 10047
rect 15427 10044 15439 10047
rect 15838 10044 15844 10056
rect 15427 10016 15844 10044
rect 15427 10013 15439 10016
rect 15381 10007 15439 10013
rect 15838 10004 15844 10016
rect 15896 10044 15902 10056
rect 16945 10047 17003 10053
rect 16945 10044 16957 10047
rect 15896 10016 16957 10044
rect 15896 10004 15902 10016
rect 16945 10013 16957 10016
rect 16991 10044 17003 10047
rect 17402 10044 17408 10056
rect 16991 10016 17408 10044
rect 16991 10013 17003 10016
rect 16945 10007 17003 10013
rect 17402 10004 17408 10016
rect 17460 10004 17466 10056
rect 16390 9936 16396 9988
rect 16448 9976 16454 9988
rect 16485 9979 16543 9985
rect 16485 9976 16497 9979
rect 16448 9948 16497 9976
rect 16448 9936 16454 9948
rect 16485 9945 16497 9948
rect 16531 9976 16543 9979
rect 16758 9976 16764 9988
rect 16531 9948 16764 9976
rect 16531 9945 16543 9948
rect 16485 9939 16543 9945
rect 16758 9936 16764 9948
rect 16816 9936 16822 9988
rect 18230 9936 18236 9988
rect 18288 9976 18294 9988
rect 18877 9979 18935 9985
rect 18877 9976 18889 9979
rect 18288 9948 18889 9976
rect 18288 9936 18294 9948
rect 18877 9945 18889 9948
rect 18923 9945 18935 9979
rect 19610 9976 19616 9988
rect 19571 9948 19616 9976
rect 18877 9939 18935 9945
rect 19610 9936 19616 9948
rect 19668 9936 19674 9988
rect 9401 9911 9459 9917
rect 9401 9908 9413 9911
rect 9180 9880 9413 9908
rect 9180 9868 9186 9880
rect 9401 9877 9413 9880
rect 9447 9877 9459 9911
rect 9401 9871 9459 9877
rect 12529 9911 12587 9917
rect 12529 9877 12541 9911
rect 12575 9908 12587 9911
rect 12986 9908 12992 9920
rect 12575 9880 12992 9908
rect 12575 9877 12587 9880
rect 12529 9871 12587 9877
rect 12986 9868 12992 9880
rect 13044 9868 13050 9920
rect 14734 9908 14740 9920
rect 14695 9880 14740 9908
rect 14734 9868 14740 9880
rect 14792 9868 14798 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 5534 9704 5540 9716
rect 5495 9676 5540 9704
rect 5534 9664 5540 9676
rect 5592 9664 5598 9716
rect 6273 9707 6331 9713
rect 6273 9673 6285 9707
rect 6319 9704 6331 9707
rect 6641 9707 6699 9713
rect 6641 9704 6653 9707
rect 6319 9676 6653 9704
rect 6319 9673 6331 9676
rect 6273 9667 6331 9673
rect 6641 9673 6653 9676
rect 6687 9704 6699 9707
rect 6730 9704 6736 9716
rect 6687 9676 6736 9704
rect 6687 9673 6699 9676
rect 6641 9667 6699 9673
rect 2958 9596 2964 9648
rect 3016 9636 3022 9648
rect 3053 9639 3111 9645
rect 3053 9636 3065 9639
rect 3016 9608 3065 9636
rect 3016 9596 3022 9608
rect 3053 9605 3065 9608
rect 3099 9636 3111 9639
rect 3099 9608 4200 9636
rect 3099 9605 3111 9608
rect 3053 9599 3111 9605
rect 1670 9568 1676 9580
rect 1631 9540 1676 9568
rect 1670 9528 1676 9540
rect 1728 9528 1734 9580
rect 2314 9568 2320 9580
rect 2275 9540 2320 9568
rect 2314 9528 2320 9540
rect 2372 9528 2378 9580
rect 4172 9568 4200 9608
rect 5552 9568 5580 9664
rect 4172 9540 5580 9568
rect 3418 9500 3424 9512
rect 3379 9472 3424 9500
rect 3418 9460 3424 9472
rect 3476 9460 3482 9512
rect 3878 9500 3884 9512
rect 3839 9472 3884 9500
rect 3878 9460 3884 9472
rect 3936 9460 3942 9512
rect 4172 9509 4200 9540
rect 4157 9503 4215 9509
rect 4157 9469 4169 9503
rect 4203 9469 4215 9503
rect 4522 9500 4528 9512
rect 4483 9472 4528 9500
rect 4157 9463 4215 9469
rect 4522 9460 4528 9472
rect 4580 9500 4586 9512
rect 5169 9503 5227 9509
rect 5169 9500 5181 9503
rect 4580 9472 5181 9500
rect 4580 9460 4586 9472
rect 5169 9469 5181 9472
rect 5215 9469 5227 9503
rect 5169 9463 5227 9469
rect 5721 9503 5779 9509
rect 5721 9469 5733 9503
rect 5767 9500 5779 9503
rect 6288 9500 6316 9667
rect 6730 9664 6736 9676
rect 6788 9664 6794 9716
rect 7742 9664 7748 9716
rect 7800 9704 7806 9716
rect 7800 9676 7880 9704
rect 7800 9664 7806 9676
rect 7852 9636 7880 9676
rect 9950 9664 9956 9716
rect 10008 9704 10014 9716
rect 10045 9707 10103 9713
rect 10045 9704 10057 9707
rect 10008 9676 10057 9704
rect 10008 9664 10014 9676
rect 10045 9673 10057 9676
rect 10091 9704 10103 9707
rect 10321 9707 10379 9713
rect 10321 9704 10333 9707
rect 10091 9676 10333 9704
rect 10091 9673 10103 9676
rect 10045 9667 10103 9673
rect 10321 9673 10333 9676
rect 10367 9673 10379 9707
rect 10321 9667 10379 9673
rect 10873 9707 10931 9713
rect 10873 9673 10885 9707
rect 10919 9704 10931 9707
rect 10962 9704 10968 9716
rect 10919 9676 10968 9704
rect 10919 9673 10931 9676
rect 10873 9667 10931 9673
rect 10962 9664 10968 9676
rect 11020 9664 11026 9716
rect 12526 9704 12532 9716
rect 12452 9676 12532 9704
rect 7392 9608 7880 9636
rect 8665 9639 8723 9645
rect 7392 9580 7420 9608
rect 8665 9605 8677 9639
rect 8711 9636 8723 9639
rect 8754 9636 8760 9648
rect 8711 9608 8760 9636
rect 8711 9605 8723 9608
rect 8665 9599 8723 9605
rect 7374 9528 7380 9580
rect 7432 9528 7438 9580
rect 8680 9568 8708 9599
rect 8754 9596 8760 9608
rect 8812 9596 8818 9648
rect 7852 9540 8708 9568
rect 7852 9512 7880 9540
rect 9030 9528 9036 9580
rect 9088 9568 9094 9580
rect 9125 9571 9183 9577
rect 9125 9568 9137 9571
rect 9088 9540 9137 9568
rect 9088 9528 9094 9540
rect 9125 9537 9137 9540
rect 9171 9537 9183 9571
rect 9125 9531 9183 9537
rect 7098 9500 7104 9512
rect 5767 9472 6316 9500
rect 7059 9472 7104 9500
rect 5767 9469 5779 9472
rect 5721 9463 5779 9469
rect 7098 9460 7104 9472
rect 7156 9460 7162 9512
rect 7285 9503 7343 9509
rect 7285 9469 7297 9503
rect 7331 9469 7343 9503
rect 7834 9500 7840 9512
rect 7747 9472 7840 9500
rect 7285 9463 7343 9469
rect 1765 9435 1823 9441
rect 1765 9401 1777 9435
rect 1811 9432 1823 9435
rect 2038 9432 2044 9444
rect 1811 9404 2044 9432
rect 1811 9401 1823 9404
rect 1765 9395 1823 9401
rect 2038 9392 2044 9404
rect 2096 9392 2102 9444
rect 2590 9364 2596 9376
rect 2551 9336 2596 9364
rect 2590 9324 2596 9336
rect 2648 9324 2654 9376
rect 4430 9324 4436 9376
rect 4488 9364 4494 9376
rect 4525 9367 4583 9373
rect 4525 9364 4537 9367
rect 4488 9336 4537 9364
rect 4488 9324 4494 9336
rect 4525 9333 4537 9336
rect 4571 9333 4583 9367
rect 4525 9327 4583 9333
rect 5905 9367 5963 9373
rect 5905 9333 5917 9367
rect 5951 9364 5963 9367
rect 6178 9364 6184 9376
rect 5951 9336 6184 9364
rect 5951 9333 5963 9336
rect 5905 9327 5963 9333
rect 6178 9324 6184 9336
rect 6236 9364 6242 9376
rect 6822 9364 6828 9376
rect 6236 9336 6828 9364
rect 6236 9324 6242 9336
rect 6822 9324 6828 9336
rect 6880 9364 6886 9376
rect 7300 9364 7328 9463
rect 7834 9460 7840 9472
rect 7892 9460 7898 9512
rect 7926 9460 7932 9512
rect 7984 9500 7990 9512
rect 8021 9503 8079 9509
rect 8021 9500 8033 9503
rect 7984 9472 8033 9500
rect 7984 9460 7990 9472
rect 8021 9469 8033 9472
rect 8067 9469 8079 9503
rect 10980 9500 11008 9664
rect 12452 9636 12480 9676
rect 12526 9664 12532 9676
rect 12584 9664 12590 9716
rect 13538 9704 13544 9716
rect 13451 9676 13544 9704
rect 13538 9664 13544 9676
rect 13596 9704 13602 9716
rect 16390 9704 16396 9716
rect 13596 9676 16396 9704
rect 13596 9664 13602 9676
rect 16390 9664 16396 9676
rect 16448 9664 16454 9716
rect 16850 9664 16856 9716
rect 16908 9704 16914 9716
rect 17681 9707 17739 9713
rect 17681 9704 17693 9707
rect 16908 9676 17693 9704
rect 16908 9664 16914 9676
rect 17681 9673 17693 9676
rect 17727 9673 17739 9707
rect 17681 9667 17739 9673
rect 18414 9664 18420 9716
rect 18472 9704 18478 9716
rect 19061 9707 19119 9713
rect 19061 9704 19073 9707
rect 18472 9676 19073 9704
rect 18472 9664 18478 9676
rect 19061 9673 19073 9676
rect 19107 9673 19119 9707
rect 19426 9704 19432 9716
rect 19387 9676 19432 9704
rect 19061 9667 19119 9673
rect 19426 9664 19432 9676
rect 19484 9664 19490 9716
rect 12894 9636 12900 9648
rect 12452 9608 12900 9636
rect 12894 9596 12900 9608
rect 12952 9596 12958 9648
rect 11514 9568 11520 9580
rect 11475 9540 11520 9568
rect 11514 9528 11520 9540
rect 11572 9528 11578 9580
rect 12526 9568 12532 9580
rect 12487 9540 12532 9568
rect 12526 9528 12532 9540
rect 12584 9568 12590 9580
rect 13817 9571 13875 9577
rect 13817 9568 13829 9571
rect 12584 9540 13829 9568
rect 12584 9528 12590 9540
rect 13817 9537 13829 9540
rect 13863 9537 13875 9571
rect 13817 9531 13875 9537
rect 15105 9571 15163 9577
rect 15105 9537 15117 9571
rect 15151 9568 15163 9571
rect 15286 9568 15292 9580
rect 15151 9540 15292 9568
rect 15151 9537 15163 9540
rect 15105 9531 15163 9537
rect 15286 9528 15292 9540
rect 15344 9568 15350 9580
rect 16868 9568 16896 9664
rect 17037 9639 17095 9645
rect 17037 9605 17049 9639
rect 17083 9636 17095 9639
rect 17126 9636 17132 9648
rect 17083 9608 17132 9636
rect 17083 9605 17095 9608
rect 17037 9599 17095 9605
rect 15344 9540 16896 9568
rect 15344 9528 15350 9540
rect 11149 9503 11207 9509
rect 11149 9500 11161 9503
rect 10980 9472 11161 9500
rect 8021 9463 8079 9469
rect 11149 9469 11161 9472
rect 11195 9469 11207 9503
rect 11149 9463 11207 9469
rect 14277 9503 14335 9509
rect 14277 9469 14289 9503
rect 14323 9500 14335 9503
rect 15013 9503 15071 9509
rect 15013 9500 15025 9503
rect 14323 9472 15025 9500
rect 14323 9469 14335 9472
rect 14277 9463 14335 9469
rect 15013 9469 15025 9472
rect 15059 9500 15071 9503
rect 15194 9500 15200 9512
rect 15059 9472 15200 9500
rect 15059 9469 15071 9472
rect 15013 9463 15071 9469
rect 15194 9460 15200 9472
rect 15252 9500 15258 9512
rect 16114 9500 16120 9512
rect 15252 9472 15516 9500
rect 16075 9472 16120 9500
rect 15252 9460 15258 9472
rect 9490 9441 9496 9444
rect 9033 9435 9091 9441
rect 9033 9401 9045 9435
rect 9079 9432 9091 9435
rect 9446 9435 9496 9441
rect 9446 9432 9458 9435
rect 9079 9404 9458 9432
rect 9079 9401 9091 9404
rect 9033 9395 9091 9401
rect 9446 9401 9458 9404
rect 9492 9401 9496 9435
rect 9446 9395 9496 9401
rect 9490 9392 9496 9395
rect 9548 9432 9554 9444
rect 9548 9404 9594 9432
rect 9548 9392 9554 9404
rect 10778 9392 10784 9444
rect 10836 9432 10842 9444
rect 10965 9435 11023 9441
rect 10965 9432 10977 9435
rect 10836 9404 10977 9432
rect 10836 9392 10842 9404
rect 10965 9401 10977 9404
rect 11011 9432 11023 9435
rect 11793 9435 11851 9441
rect 11793 9432 11805 9435
rect 11011 9404 11805 9432
rect 11011 9401 11023 9404
rect 10965 9395 11023 9401
rect 11793 9401 11805 9404
rect 11839 9401 11851 9435
rect 11793 9395 11851 9401
rect 12253 9435 12311 9441
rect 12253 9401 12265 9435
rect 12299 9432 12311 9435
rect 12618 9432 12624 9444
rect 12299 9404 12624 9432
rect 12299 9401 12311 9404
rect 12253 9395 12311 9401
rect 12618 9392 12624 9404
rect 12676 9392 12682 9444
rect 12894 9392 12900 9444
rect 12952 9432 12958 9444
rect 13173 9435 13231 9441
rect 13173 9432 13185 9435
rect 12952 9404 13185 9432
rect 12952 9392 12958 9404
rect 13173 9401 13185 9404
rect 13219 9401 13231 9435
rect 13173 9395 13231 9401
rect 8018 9364 8024 9376
rect 6880 9336 7328 9364
rect 7979 9336 8024 9364
rect 6880 9324 6886 9336
rect 8018 9324 8024 9336
rect 8076 9324 8082 9376
rect 15488 9373 15516 9472
rect 16114 9460 16120 9472
rect 16172 9460 16178 9512
rect 16298 9460 16304 9512
rect 16356 9500 16362 9512
rect 16393 9503 16451 9509
rect 16393 9500 16405 9503
rect 16356 9472 16405 9500
rect 16356 9460 16362 9472
rect 16393 9469 16405 9472
rect 16439 9500 16451 9503
rect 16482 9500 16488 9512
rect 16439 9472 16488 9500
rect 16439 9469 16451 9472
rect 16393 9463 16451 9469
rect 16482 9460 16488 9472
rect 16540 9460 16546 9512
rect 15654 9392 15660 9444
rect 15712 9432 15718 9444
rect 15841 9435 15899 9441
rect 15841 9432 15853 9435
rect 15712 9404 15853 9432
rect 15712 9392 15718 9404
rect 15841 9401 15853 9404
rect 15887 9432 15899 9435
rect 17052 9432 17080 9599
rect 17126 9596 17132 9608
rect 17184 9596 17190 9648
rect 17402 9636 17408 9648
rect 17363 9608 17408 9636
rect 17402 9596 17408 9608
rect 17460 9596 17466 9648
rect 19751 9639 19809 9645
rect 19751 9636 19763 9639
rect 18156 9608 19763 9636
rect 17954 9528 17960 9580
rect 18012 9568 18018 9580
rect 18156 9577 18184 9608
rect 19751 9605 19763 9608
rect 19797 9605 19809 9639
rect 20162 9636 20168 9648
rect 20123 9608 20168 9636
rect 19751 9599 19809 9605
rect 20162 9596 20168 9608
rect 20220 9596 20226 9648
rect 18141 9571 18199 9577
rect 18141 9568 18153 9571
rect 18012 9540 18153 9568
rect 18012 9528 18018 9540
rect 18141 9537 18153 9540
rect 18187 9537 18199 9571
rect 18141 9531 18199 9537
rect 19680 9503 19738 9509
rect 19680 9469 19692 9503
rect 19726 9500 19738 9503
rect 20180 9500 20208 9596
rect 19726 9472 20208 9500
rect 19726 9469 19738 9472
rect 19680 9463 19738 9469
rect 18230 9432 18236 9444
rect 15887 9404 17080 9432
rect 18191 9404 18236 9432
rect 15887 9401 15899 9404
rect 15841 9395 15899 9401
rect 18230 9392 18236 9404
rect 18288 9392 18294 9444
rect 18782 9432 18788 9444
rect 18743 9404 18788 9432
rect 18782 9392 18788 9404
rect 18840 9392 18846 9444
rect 15473 9367 15531 9373
rect 15473 9333 15485 9367
rect 15519 9364 15531 9367
rect 15746 9364 15752 9376
rect 15519 9336 15752 9364
rect 15519 9333 15531 9336
rect 15473 9327 15531 9333
rect 15746 9324 15752 9336
rect 15804 9324 15810 9376
rect 16206 9364 16212 9376
rect 16167 9336 16212 9364
rect 16206 9324 16212 9336
rect 16264 9324 16270 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 2866 9120 2872 9172
rect 2924 9160 2930 9172
rect 3145 9163 3203 9169
rect 3145 9160 3157 9163
rect 2924 9132 3157 9160
rect 2924 9120 2930 9132
rect 3145 9129 3157 9132
rect 3191 9129 3203 9163
rect 3145 9123 3203 9129
rect 3513 9163 3571 9169
rect 3513 9129 3525 9163
rect 3559 9160 3571 9163
rect 3878 9160 3884 9172
rect 3559 9132 3884 9160
rect 3559 9129 3571 9132
rect 3513 9123 3571 9129
rect 3878 9120 3884 9132
rect 3936 9120 3942 9172
rect 4338 9160 4344 9172
rect 4299 9132 4344 9160
rect 4338 9120 4344 9132
rect 4396 9120 4402 9172
rect 8662 9160 8668 9172
rect 8623 9132 8668 9160
rect 8662 9120 8668 9132
rect 8720 9120 8726 9172
rect 8938 9160 8944 9172
rect 8899 9132 8944 9160
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 9030 9120 9036 9172
rect 9088 9160 9094 9172
rect 9309 9163 9367 9169
rect 9309 9160 9321 9163
rect 9088 9132 9321 9160
rect 9088 9120 9094 9132
rect 9309 9129 9321 9132
rect 9355 9129 9367 9163
rect 9309 9123 9367 9129
rect 11333 9163 11391 9169
rect 11333 9129 11345 9163
rect 11379 9160 11391 9163
rect 11422 9160 11428 9172
rect 11379 9132 11428 9160
rect 11379 9129 11391 9132
rect 11333 9123 11391 9129
rect 11422 9120 11428 9132
rect 11480 9120 11486 9172
rect 12618 9160 12624 9172
rect 12579 9132 12624 9160
rect 12618 9120 12624 9132
rect 12676 9120 12682 9172
rect 15378 9120 15384 9172
rect 15436 9160 15442 9172
rect 15473 9163 15531 9169
rect 15473 9160 15485 9163
rect 15436 9132 15485 9160
rect 15436 9120 15442 9132
rect 15473 9129 15485 9132
rect 15519 9129 15531 9163
rect 15838 9160 15844 9172
rect 15799 9132 15844 9160
rect 15473 9123 15531 9129
rect 15838 9120 15844 9132
rect 15896 9120 15902 9172
rect 16114 9160 16120 9172
rect 16075 9132 16120 9160
rect 16114 9120 16120 9132
rect 16172 9120 16178 9172
rect 17954 9160 17960 9172
rect 17915 9132 17960 9160
rect 17954 9120 17960 9132
rect 18012 9120 18018 9172
rect 1486 9052 1492 9104
rect 1544 9092 1550 9104
rect 1581 9095 1639 9101
rect 1581 9092 1593 9095
rect 1544 9064 1593 9092
rect 1544 9052 1550 9064
rect 1581 9061 1593 9064
rect 1627 9092 1639 9095
rect 1762 9092 1768 9104
rect 1627 9064 1768 9092
rect 1627 9061 1639 9064
rect 1581 9055 1639 9061
rect 1762 9052 1768 9064
rect 1820 9052 1826 9104
rect 2133 9095 2191 9101
rect 2133 9061 2145 9095
rect 2179 9092 2191 9095
rect 2314 9092 2320 9104
rect 2179 9064 2320 9092
rect 2179 9061 2191 9064
rect 2133 9055 2191 9061
rect 2314 9052 2320 9064
rect 2372 9052 2378 9104
rect 2501 9095 2559 9101
rect 2501 9061 2513 9095
rect 2547 9092 2559 9095
rect 3694 9092 3700 9104
rect 2547 9064 3700 9092
rect 2547 9061 2559 9064
rect 2501 9055 2559 9061
rect 3694 9052 3700 9064
rect 3752 9092 3758 9104
rect 4246 9092 4252 9104
rect 3752 9064 4252 9092
rect 3752 9052 3758 9064
rect 4246 9052 4252 9064
rect 4304 9092 4310 9104
rect 4304 9064 4568 9092
rect 4304 9052 4310 9064
rect 2961 9027 3019 9033
rect 2961 8993 2973 9027
rect 3007 9024 3019 9027
rect 3510 9024 3516 9036
rect 3007 8996 3516 9024
rect 3007 8993 3019 8996
rect 2961 8987 3019 8993
rect 3510 8984 3516 8996
rect 3568 8984 3574 9036
rect 4062 9024 4068 9036
rect 4023 8996 4068 9024
rect 4062 8984 4068 8996
rect 4120 8984 4126 9036
rect 4540 9033 4568 9064
rect 6454 9052 6460 9104
rect 6512 9092 6518 9104
rect 9858 9092 9864 9104
rect 6512 9064 7236 9092
rect 9819 9064 9864 9092
rect 6512 9052 6518 9064
rect 4525 9027 4583 9033
rect 4525 8993 4537 9027
rect 4571 8993 4583 9027
rect 4982 9024 4988 9036
rect 4943 8996 4988 9024
rect 4525 8987 4583 8993
rect 4982 8984 4988 8996
rect 5040 8984 5046 9036
rect 5258 9024 5264 9036
rect 5219 8996 5264 9024
rect 5258 8984 5264 8996
rect 5316 8984 5322 9036
rect 5350 8984 5356 9036
rect 5408 9024 5414 9036
rect 5994 9024 6000 9036
rect 5408 8996 6000 9024
rect 5408 8984 5414 8996
rect 5994 8984 6000 8996
rect 6052 9024 6058 9036
rect 6365 9027 6423 9033
rect 6365 9024 6377 9027
rect 6052 8996 6377 9024
rect 6052 8984 6058 8996
rect 6365 8993 6377 8996
rect 6411 8993 6423 9027
rect 6822 9024 6828 9036
rect 6783 8996 6828 9024
rect 6365 8987 6423 8993
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 7208 9033 7236 9064
rect 9858 9052 9864 9064
rect 9916 9052 9922 9104
rect 11790 9052 11796 9104
rect 11848 9092 11854 9104
rect 16666 9101 16672 9104
rect 12022 9095 12080 9101
rect 12022 9092 12034 9095
rect 11848 9064 12034 9092
rect 11848 9052 11854 9064
rect 12022 9061 12034 9064
rect 12068 9061 12080 9095
rect 16663 9092 16672 9101
rect 16627 9064 16672 9092
rect 12022 9055 12080 9061
rect 16663 9055 16672 9064
rect 16666 9052 16672 9055
rect 16724 9052 16730 9104
rect 17770 9052 17776 9104
rect 17828 9092 17834 9104
rect 18233 9095 18291 9101
rect 18233 9092 18245 9095
rect 17828 9064 18245 9092
rect 17828 9052 17834 9064
rect 18233 9061 18245 9064
rect 18279 9061 18291 9095
rect 18782 9092 18788 9104
rect 18743 9064 18788 9092
rect 18233 9055 18291 9061
rect 18782 9052 18788 9064
rect 18840 9052 18846 9104
rect 7193 9027 7251 9033
rect 7193 8993 7205 9027
rect 7239 8993 7251 9027
rect 7193 8987 7251 8993
rect 7561 9027 7619 9033
rect 7561 8993 7573 9027
rect 7607 9024 7619 9027
rect 7926 9024 7932 9036
rect 7607 8996 7932 9024
rect 7607 8993 7619 8996
rect 7561 8987 7619 8993
rect 1486 8956 1492 8968
rect 1447 8928 1492 8956
rect 1486 8916 1492 8928
rect 1544 8916 1550 8968
rect 7576 8956 7604 8987
rect 7926 8984 7932 8996
rect 7984 8984 7990 9036
rect 11701 9027 11759 9033
rect 11701 8993 11713 9027
rect 11747 9024 11759 9027
rect 11882 9024 11888 9036
rect 11747 8996 11888 9024
rect 11747 8993 11759 8996
rect 11701 8987 11759 8993
rect 11882 8984 11888 8996
rect 11940 9024 11946 9036
rect 12342 9024 12348 9036
rect 11940 8996 12348 9024
rect 11940 8984 11946 8996
rect 12342 8984 12348 8996
rect 12400 8984 12406 9036
rect 13722 9024 13728 9036
rect 13683 8996 13728 9024
rect 13722 8984 13728 8996
rect 13780 8984 13786 9036
rect 13909 9027 13967 9033
rect 13909 9024 13921 9027
rect 13832 8996 13921 9024
rect 9766 8956 9772 8968
rect 6104 8928 7604 8956
rect 9727 8928 9772 8956
rect 6104 8900 6132 8928
rect 9766 8916 9772 8928
rect 9824 8916 9830 8968
rect 10134 8956 10140 8968
rect 10095 8928 10140 8956
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 12989 8959 13047 8965
rect 12989 8925 13001 8959
rect 13035 8956 13047 8959
rect 13357 8959 13415 8965
rect 13357 8956 13369 8959
rect 13035 8928 13369 8956
rect 13035 8925 13047 8928
rect 12989 8919 13047 8925
rect 13357 8925 13369 8928
rect 13403 8956 13415 8959
rect 13630 8956 13636 8968
rect 13403 8928 13636 8956
rect 13403 8925 13415 8928
rect 13357 8919 13415 8925
rect 13630 8916 13636 8928
rect 13688 8956 13694 8968
rect 13832 8956 13860 8996
rect 13909 8993 13921 8996
rect 13955 9024 13967 9027
rect 14274 9024 14280 9036
rect 13955 8996 14280 9024
rect 13955 8993 13967 8996
rect 13909 8987 13967 8993
rect 14274 8984 14280 8996
rect 14332 8984 14338 9036
rect 15286 9024 15292 9036
rect 15247 8996 15292 9024
rect 15286 8984 15292 8996
rect 15344 8984 15350 9036
rect 16301 9027 16359 9033
rect 16301 8993 16313 9027
rect 16347 9024 16359 9027
rect 16482 9024 16488 9036
rect 16347 8996 16488 9024
rect 16347 8993 16359 8996
rect 16301 8987 16359 8993
rect 16482 8984 16488 8996
rect 16540 8984 16546 9036
rect 19613 9027 19671 9033
rect 19613 8993 19625 9027
rect 19659 9024 19671 9027
rect 20070 9024 20076 9036
rect 19659 8996 20076 9024
rect 19659 8993 19671 8996
rect 19613 8987 19671 8993
rect 20070 8984 20076 8996
rect 20128 8984 20134 9036
rect 13998 8956 14004 8968
rect 13688 8928 13860 8956
rect 13959 8928 14004 8956
rect 13688 8916 13694 8928
rect 13998 8916 14004 8928
rect 14056 8916 14062 8968
rect 18138 8956 18144 8968
rect 18099 8928 18144 8956
rect 18138 8916 18144 8928
rect 18196 8916 18202 8968
rect 3789 8891 3847 8897
rect 3789 8888 3801 8891
rect 2884 8860 3801 8888
rect 2884 8832 2912 8860
rect 3789 8857 3801 8860
rect 3835 8888 3847 8891
rect 4522 8888 4528 8900
rect 3835 8860 4528 8888
rect 3835 8857 3847 8860
rect 3789 8851 3847 8857
rect 4522 8848 4528 8860
rect 4580 8888 4586 8900
rect 4890 8888 4896 8900
rect 4580 8860 4896 8888
rect 4580 8848 4586 8860
rect 4890 8848 4896 8860
rect 4948 8888 4954 8900
rect 5997 8891 6055 8897
rect 5997 8888 6009 8891
rect 4948 8860 6009 8888
rect 4948 8848 4954 8860
rect 5997 8857 6009 8860
rect 6043 8888 6055 8891
rect 6086 8888 6092 8900
rect 6043 8860 6092 8888
rect 6043 8857 6055 8860
rect 5997 8851 6055 8857
rect 6086 8848 6092 8860
rect 6144 8848 6150 8900
rect 7006 8848 7012 8900
rect 7064 8888 7070 8900
rect 7745 8891 7803 8897
rect 7745 8888 7757 8891
rect 7064 8860 7757 8888
rect 7064 8848 7070 8860
rect 7745 8857 7757 8860
rect 7791 8857 7803 8891
rect 7745 8851 7803 8857
rect 2866 8820 2872 8832
rect 2827 8792 2872 8820
rect 2866 8780 2872 8792
rect 2924 8780 2930 8832
rect 7098 8780 7104 8832
rect 7156 8820 7162 8832
rect 8113 8823 8171 8829
rect 8113 8820 8125 8823
rect 7156 8792 8125 8820
rect 7156 8780 7162 8792
rect 8113 8789 8125 8792
rect 8159 8820 8171 8823
rect 8754 8820 8760 8832
rect 8159 8792 8760 8820
rect 8159 8789 8171 8792
rect 8113 8783 8171 8789
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 14553 8823 14611 8829
rect 14553 8789 14565 8823
rect 14599 8820 14611 8823
rect 14734 8820 14740 8832
rect 14599 8792 14740 8820
rect 14599 8789 14611 8792
rect 14553 8783 14611 8789
rect 14734 8780 14740 8792
rect 14792 8820 14798 8832
rect 15013 8823 15071 8829
rect 15013 8820 15025 8823
rect 14792 8792 15025 8820
rect 14792 8780 14798 8792
rect 15013 8789 15025 8792
rect 15059 8820 15071 8823
rect 16298 8820 16304 8832
rect 15059 8792 16304 8820
rect 15059 8789 15071 8792
rect 15013 8783 15071 8789
rect 16298 8780 16304 8792
rect 16356 8780 16362 8832
rect 17221 8823 17279 8829
rect 17221 8789 17233 8823
rect 17267 8820 17279 8823
rect 17770 8820 17776 8832
rect 17267 8792 17776 8820
rect 17267 8789 17279 8792
rect 17221 8783 17279 8789
rect 17770 8780 17776 8792
rect 17828 8780 17834 8832
rect 19794 8820 19800 8832
rect 19755 8792 19800 8820
rect 19794 8780 19800 8792
rect 19852 8780 19858 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1578 8616 1584 8628
rect 1539 8588 1584 8616
rect 1578 8576 1584 8588
rect 1636 8576 1642 8628
rect 1762 8576 1768 8628
rect 1820 8616 1826 8628
rect 1949 8619 2007 8625
rect 1949 8616 1961 8619
rect 1820 8588 1961 8616
rect 1820 8576 1826 8588
rect 1949 8585 1961 8588
rect 1995 8585 2007 8619
rect 2866 8616 2872 8628
rect 2827 8588 2872 8616
rect 1949 8579 2007 8585
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 3234 8616 3240 8628
rect 3195 8588 3240 8616
rect 3234 8576 3240 8588
rect 3292 8576 3298 8628
rect 3510 8616 3516 8628
rect 3471 8588 3516 8616
rect 3510 8576 3516 8588
rect 3568 8576 3574 8628
rect 5258 8576 5264 8628
rect 5316 8616 5322 8628
rect 5445 8619 5503 8625
rect 5445 8616 5457 8619
rect 5316 8588 5457 8616
rect 5316 8576 5322 8588
rect 5445 8585 5457 8588
rect 5491 8585 5503 8619
rect 6086 8616 6092 8628
rect 6047 8588 6092 8616
rect 5445 8579 5503 8585
rect 5460 8548 5488 8579
rect 6086 8576 6092 8588
rect 6144 8576 6150 8628
rect 6362 8616 6368 8628
rect 6323 8588 6368 8616
rect 6362 8576 6368 8588
rect 6420 8576 6426 8628
rect 8754 8616 8760 8628
rect 8715 8588 8760 8616
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 9858 8616 9864 8628
rect 9819 8588 9864 8616
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 11422 8576 11428 8628
rect 11480 8616 11486 8628
rect 11517 8619 11575 8625
rect 11517 8616 11529 8619
rect 11480 8588 11529 8616
rect 11480 8576 11486 8588
rect 11517 8585 11529 8588
rect 11563 8585 11575 8619
rect 11517 8579 11575 8585
rect 13541 8619 13599 8625
rect 13541 8585 13553 8619
rect 13587 8616 13599 8619
rect 13722 8616 13728 8628
rect 13587 8588 13728 8616
rect 13587 8585 13599 8588
rect 13541 8579 13599 8585
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 15197 8619 15255 8625
rect 15197 8585 15209 8619
rect 15243 8616 15255 8619
rect 15286 8616 15292 8628
rect 15243 8588 15292 8616
rect 15243 8585 15255 8588
rect 15197 8579 15255 8585
rect 15286 8576 15292 8588
rect 15344 8576 15350 8628
rect 17770 8616 17776 8628
rect 17731 8588 17776 8616
rect 17770 8576 17776 8588
rect 17828 8576 17834 8628
rect 18138 8576 18144 8628
rect 18196 8616 18202 8628
rect 19153 8619 19211 8625
rect 19153 8616 19165 8619
rect 18196 8588 19165 8616
rect 18196 8576 18202 8588
rect 19153 8585 19165 8588
rect 19199 8616 19211 8619
rect 19978 8616 19984 8628
rect 19199 8588 19984 8616
rect 19199 8585 19211 8588
rect 19153 8579 19211 8585
rect 19978 8576 19984 8588
rect 20036 8576 20042 8628
rect 6270 8548 6276 8560
rect 5460 8520 6276 8548
rect 6270 8508 6276 8520
rect 6328 8508 6334 8560
rect 16577 8551 16635 8557
rect 16577 8517 16589 8551
rect 16623 8548 16635 8551
rect 18230 8548 18236 8560
rect 16623 8520 18236 8548
rect 16623 8517 16635 8520
rect 16577 8511 16635 8517
rect 18230 8508 18236 8520
rect 18288 8548 18294 8560
rect 19242 8548 19248 8560
rect 18288 8520 19248 8548
rect 18288 8508 18294 8520
rect 19242 8508 19248 8520
rect 19300 8508 19306 8560
rect 4982 8480 4988 8492
rect 4724 8452 4988 8480
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 1946 8412 1952 8424
rect 1443 8384 1952 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 1946 8372 1952 8384
rect 2004 8372 2010 8424
rect 2685 8415 2743 8421
rect 2685 8381 2697 8415
rect 2731 8412 2743 8415
rect 3234 8412 3240 8424
rect 2731 8384 3240 8412
rect 2731 8381 2743 8384
rect 2685 8375 2743 8381
rect 3234 8372 3240 8384
rect 3292 8372 3298 8424
rect 3697 8415 3755 8421
rect 3697 8381 3709 8415
rect 3743 8412 3755 8415
rect 4062 8412 4068 8424
rect 3743 8384 4068 8412
rect 3743 8381 3755 8384
rect 3697 8375 3755 8381
rect 2593 8347 2651 8353
rect 2593 8313 2605 8347
rect 2639 8344 2651 8347
rect 3712 8344 3740 8375
rect 4062 8372 4068 8384
rect 4120 8372 4126 8424
rect 4246 8412 4252 8424
rect 4207 8384 4252 8412
rect 4246 8372 4252 8384
rect 4304 8372 4310 8424
rect 4724 8421 4752 8452
rect 4982 8440 4988 8452
rect 5040 8440 5046 8492
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 9125 8483 9183 8489
rect 9125 8480 9137 8483
rect 6880 8452 9137 8480
rect 6880 8440 6886 8452
rect 4709 8415 4767 8421
rect 4709 8381 4721 8415
rect 4755 8381 4767 8415
rect 4890 8412 4896 8424
rect 4851 8384 4896 8412
rect 4709 8375 4767 8381
rect 4890 8372 4896 8384
rect 4948 8372 4954 8424
rect 5994 8372 6000 8424
rect 6052 8412 6058 8424
rect 7009 8415 7067 8421
rect 7009 8412 7021 8415
rect 6052 8384 7021 8412
rect 6052 8372 6058 8384
rect 7009 8381 7021 8384
rect 7055 8412 7067 8415
rect 7098 8412 7104 8424
rect 7055 8384 7104 8412
rect 7055 8381 7067 8384
rect 7009 8375 7067 8381
rect 7098 8372 7104 8384
rect 7156 8372 7162 8424
rect 7484 8421 7512 8452
rect 9125 8449 9137 8452
rect 9171 8449 9183 8483
rect 10594 8480 10600 8492
rect 10555 8452 10600 8480
rect 9125 8443 9183 8449
rect 10594 8440 10600 8452
rect 10652 8440 10658 8492
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8480 12311 8483
rect 12299 8452 14044 8480
rect 12299 8449 12311 8452
rect 12253 8443 12311 8449
rect 7469 8415 7527 8421
rect 7469 8381 7481 8415
rect 7515 8381 7527 8415
rect 7834 8412 7840 8424
rect 7795 8384 7840 8412
rect 7469 8375 7527 8381
rect 7834 8372 7840 8384
rect 7892 8372 7898 8424
rect 8294 8412 8300 8424
rect 8255 8384 8300 8412
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 9490 8372 9496 8424
rect 9548 8412 9554 8424
rect 12728 8421 12756 8452
rect 10413 8415 10471 8421
rect 10413 8412 10425 8415
rect 9548 8384 10425 8412
rect 9548 8372 9554 8384
rect 10413 8381 10425 8384
rect 10459 8381 10471 8415
rect 10413 8375 10471 8381
rect 12713 8415 12771 8421
rect 12713 8381 12725 8415
rect 12759 8381 12771 8415
rect 12713 8375 12771 8381
rect 12989 8415 13047 8421
rect 12989 8381 13001 8415
rect 13035 8412 13047 8415
rect 13630 8412 13636 8424
rect 13035 8384 13636 8412
rect 13035 8381 13047 8384
rect 12989 8375 13047 8381
rect 2639 8316 3740 8344
rect 9309 8347 9367 8353
rect 2639 8313 2651 8316
rect 2593 8307 2651 8313
rect 9309 8313 9321 8347
rect 9355 8344 9367 8347
rect 9398 8344 9404 8356
rect 9355 8316 9404 8344
rect 9355 8313 9367 8316
rect 9309 8307 9367 8313
rect 9398 8304 9404 8316
rect 9456 8304 9462 8356
rect 10428 8344 10456 8375
rect 13630 8372 13636 8384
rect 13688 8372 13694 8424
rect 14016 8421 14044 8452
rect 15562 8440 15568 8492
rect 15620 8480 15626 8492
rect 15657 8483 15715 8489
rect 15657 8480 15669 8483
rect 15620 8452 15669 8480
rect 15620 8440 15626 8452
rect 15657 8449 15669 8452
rect 15703 8449 15715 8483
rect 15657 8443 15715 8449
rect 18141 8483 18199 8489
rect 18141 8449 18153 8483
rect 18187 8480 18199 8483
rect 18782 8480 18788 8492
rect 18187 8452 18788 8480
rect 18187 8449 18199 8452
rect 18141 8443 18199 8449
rect 18782 8440 18788 8452
rect 18840 8480 18846 8492
rect 19429 8483 19487 8489
rect 19429 8480 19441 8483
rect 18840 8452 19441 8480
rect 18840 8440 18846 8452
rect 19429 8449 19441 8452
rect 19475 8449 19487 8483
rect 19429 8443 19487 8449
rect 14001 8415 14059 8421
rect 14001 8381 14013 8415
rect 14047 8412 14059 8415
rect 14090 8412 14096 8424
rect 14047 8384 14096 8412
rect 14047 8381 14059 8384
rect 14001 8375 14059 8381
rect 14090 8372 14096 8384
rect 14148 8372 14154 8424
rect 14645 8415 14703 8421
rect 14645 8381 14657 8415
rect 14691 8412 14703 8415
rect 14734 8412 14740 8424
rect 14691 8384 14740 8412
rect 14691 8381 14703 8384
rect 14645 8375 14703 8381
rect 14734 8372 14740 8384
rect 14792 8372 14798 8424
rect 20070 8412 20076 8424
rect 20031 8384 20076 8412
rect 20070 8372 20076 8384
rect 20128 8372 20134 8424
rect 10918 8347 10976 8353
rect 10918 8344 10930 8347
rect 10428 8316 10930 8344
rect 10918 8313 10930 8316
rect 10964 8344 10976 8347
rect 11790 8344 11796 8356
rect 10964 8316 11796 8344
rect 10964 8313 10976 8316
rect 10918 8307 10976 8313
rect 11790 8304 11796 8316
rect 11848 8304 11854 8356
rect 13170 8344 13176 8356
rect 13131 8316 13176 8344
rect 13170 8304 13176 8316
rect 13228 8304 13234 8356
rect 14826 8344 14832 8356
rect 14787 8316 14832 8344
rect 14826 8304 14832 8316
rect 14884 8304 14890 8356
rect 15978 8347 16036 8353
rect 15978 8344 15990 8347
rect 15488 8316 15990 8344
rect 3786 8276 3792 8288
rect 3747 8248 3792 8276
rect 3786 8236 3792 8248
rect 3844 8236 3850 8288
rect 7834 8236 7840 8288
rect 7892 8276 7898 8288
rect 8205 8279 8263 8285
rect 8205 8276 8217 8279
rect 7892 8248 8217 8276
rect 7892 8236 7898 8248
rect 8205 8245 8217 8248
rect 8251 8245 8263 8279
rect 8205 8239 8263 8245
rect 15286 8236 15292 8288
rect 15344 8276 15350 8288
rect 15488 8285 15516 8316
rect 15978 8313 15990 8316
rect 16024 8344 16036 8347
rect 16666 8344 16672 8356
rect 16024 8316 16672 8344
rect 16024 8313 16036 8316
rect 15978 8307 16036 8313
rect 16666 8304 16672 8316
rect 16724 8344 16730 8356
rect 16853 8347 16911 8353
rect 16853 8344 16865 8347
rect 16724 8316 16865 8344
rect 16724 8304 16730 8316
rect 16853 8313 16865 8316
rect 16899 8313 16911 8347
rect 18233 8347 18291 8353
rect 16853 8307 16911 8313
rect 17512 8316 18092 8344
rect 17512 8288 17540 8316
rect 15473 8279 15531 8285
rect 15473 8276 15485 8279
rect 15344 8248 15485 8276
rect 15344 8236 15350 8248
rect 15473 8245 15485 8248
rect 15519 8245 15531 8279
rect 17494 8276 17500 8288
rect 17455 8248 17500 8276
rect 15473 8239 15531 8245
rect 17494 8236 17500 8248
rect 17552 8236 17558 8288
rect 18064 8276 18092 8316
rect 18233 8313 18245 8347
rect 18279 8313 18291 8347
rect 18233 8307 18291 8313
rect 18248 8276 18276 8307
rect 18598 8304 18604 8356
rect 18656 8344 18662 8356
rect 18785 8347 18843 8353
rect 18785 8344 18797 8347
rect 18656 8316 18797 8344
rect 18656 8304 18662 8316
rect 18785 8313 18797 8316
rect 18831 8313 18843 8347
rect 19613 8347 19671 8353
rect 19613 8344 19625 8347
rect 18785 8307 18843 8313
rect 19260 8316 19625 8344
rect 18064 8248 18276 8276
rect 19150 8236 19156 8288
rect 19208 8276 19214 8288
rect 19260 8276 19288 8316
rect 19613 8313 19625 8316
rect 19659 8313 19671 8347
rect 19613 8307 19671 8313
rect 19208 8248 19288 8276
rect 19208 8236 19214 8248
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1397 8075 1455 8081
rect 1397 8041 1409 8075
rect 1443 8072 1455 8075
rect 1486 8072 1492 8084
rect 1443 8044 1492 8072
rect 1443 8041 1455 8044
rect 1397 8035 1455 8041
rect 1486 8032 1492 8044
rect 1544 8072 1550 8084
rect 1857 8075 1915 8081
rect 1857 8072 1869 8075
rect 1544 8044 1869 8072
rect 1544 8032 1550 8044
rect 1857 8041 1869 8044
rect 1903 8041 1915 8075
rect 1857 8035 1915 8041
rect 2038 8032 2044 8084
rect 2096 8072 2102 8084
rect 2225 8075 2283 8081
rect 2225 8072 2237 8075
rect 2096 8044 2237 8072
rect 2096 8032 2102 8044
rect 2225 8041 2237 8044
rect 2271 8041 2283 8075
rect 2225 8035 2283 8041
rect 4154 8032 4160 8084
rect 4212 8072 4218 8084
rect 5077 8075 5135 8081
rect 5077 8072 5089 8075
rect 4212 8044 5089 8072
rect 4212 8032 4218 8044
rect 5077 8041 5089 8044
rect 5123 8072 5135 8075
rect 5445 8075 5503 8081
rect 5445 8072 5457 8075
rect 5123 8044 5457 8072
rect 5123 8041 5135 8044
rect 5077 8035 5135 8041
rect 5445 8041 5457 8044
rect 5491 8041 5503 8075
rect 5445 8035 5503 8041
rect 7469 8075 7527 8081
rect 7469 8041 7481 8075
rect 7515 8072 7527 8075
rect 7742 8072 7748 8084
rect 7515 8044 7748 8072
rect 7515 8041 7527 8044
rect 7469 8035 7527 8041
rect 3789 8007 3847 8013
rect 3789 7973 3801 8007
rect 3835 8004 3847 8007
rect 4341 8007 4399 8013
rect 4341 8004 4353 8007
rect 3835 7976 4353 8004
rect 3835 7973 3847 7976
rect 3789 7967 3847 7973
rect 4341 7973 4353 7976
rect 4387 8004 4399 8007
rect 4982 8004 4988 8016
rect 4387 7976 4988 8004
rect 4387 7973 4399 7976
rect 4341 7967 4399 7973
rect 4982 7964 4988 7976
rect 5040 7964 5046 8016
rect 3050 7936 3056 7948
rect 3011 7908 3056 7936
rect 3050 7896 3056 7908
rect 3108 7896 3114 7948
rect 4706 7945 4712 7948
rect 4684 7939 4712 7945
rect 4684 7905 4696 7939
rect 4684 7899 4712 7905
rect 4706 7896 4712 7899
rect 4764 7896 4770 7948
rect 5460 7936 5488 8035
rect 7742 8032 7748 8044
rect 7800 8032 7806 8084
rect 10686 8072 10692 8084
rect 10647 8044 10692 8072
rect 10686 8032 10692 8044
rect 10744 8032 10750 8084
rect 11882 8072 11888 8084
rect 11843 8044 11888 8072
rect 11882 8032 11888 8044
rect 11940 8032 11946 8084
rect 13630 8072 13636 8084
rect 13591 8044 13636 8072
rect 13630 8032 13636 8044
rect 13688 8032 13694 8084
rect 15470 8072 15476 8084
rect 15431 8044 15476 8072
rect 15470 8032 15476 8044
rect 15528 8032 15534 8084
rect 15562 8032 15568 8084
rect 15620 8072 15626 8084
rect 15749 8075 15807 8081
rect 15749 8072 15761 8075
rect 15620 8044 15761 8072
rect 15620 8032 15626 8044
rect 15749 8041 15761 8044
rect 15795 8041 15807 8075
rect 15749 8035 15807 8041
rect 16393 8075 16451 8081
rect 16393 8041 16405 8075
rect 16439 8072 16451 8075
rect 16482 8072 16488 8084
rect 16439 8044 16488 8072
rect 16439 8041 16451 8044
rect 16393 8035 16451 8041
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 17494 8072 17500 8084
rect 17455 8044 17500 8072
rect 17494 8032 17500 8044
rect 17552 8032 17558 8084
rect 6270 7964 6276 8016
rect 6328 8004 6334 8016
rect 6328 7976 6868 8004
rect 6328 7964 6334 7976
rect 5629 7939 5687 7945
rect 5629 7936 5641 7939
rect 5460 7908 5641 7936
rect 5629 7905 5641 7908
rect 5675 7936 5687 7939
rect 5994 7936 6000 7948
rect 5675 7908 6000 7936
rect 5675 7905 5687 7908
rect 5629 7899 5687 7905
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 6178 7936 6184 7948
rect 6139 7908 6184 7936
rect 6178 7896 6184 7908
rect 6236 7896 6242 7948
rect 6362 7896 6368 7948
rect 6420 7936 6426 7948
rect 6840 7945 6868 7976
rect 11790 7964 11796 8016
rect 11848 8004 11854 8016
rect 12758 8007 12816 8013
rect 12758 8004 12770 8007
rect 11848 7976 12770 8004
rect 11848 7964 11854 7976
rect 12758 7973 12770 7976
rect 12804 7973 12816 8007
rect 12758 7967 12816 7973
rect 6457 7939 6515 7945
rect 6457 7936 6469 7939
rect 6420 7908 6469 7936
rect 6420 7896 6426 7908
rect 6457 7905 6469 7908
rect 6503 7905 6515 7939
rect 6457 7899 6515 7905
rect 6825 7939 6883 7945
rect 6825 7905 6837 7939
rect 6871 7936 6883 7939
rect 7745 7939 7803 7945
rect 7745 7936 7757 7939
rect 6871 7908 7757 7936
rect 6871 7905 6883 7908
rect 6825 7899 6883 7905
rect 7745 7905 7757 7908
rect 7791 7936 7803 7939
rect 8202 7936 8208 7948
rect 7791 7908 8208 7936
rect 7791 7905 7803 7908
rect 7745 7899 7803 7905
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 8662 7936 8668 7948
rect 8623 7908 8668 7936
rect 8662 7896 8668 7908
rect 8720 7896 8726 7948
rect 9928 7939 9986 7945
rect 9928 7905 9940 7939
rect 9974 7936 9986 7939
rect 10042 7936 10048 7948
rect 9974 7908 10048 7936
rect 9974 7905 9986 7908
rect 9928 7899 9986 7905
rect 10042 7896 10048 7908
rect 10100 7896 10106 7948
rect 11146 7936 11152 7948
rect 11107 7908 11152 7936
rect 11146 7896 11152 7908
rect 11204 7896 11210 7948
rect 11422 7936 11428 7948
rect 11335 7908 11428 7936
rect 11422 7896 11428 7908
rect 11480 7936 11486 7948
rect 13648 7936 13676 8032
rect 16666 7964 16672 8016
rect 16724 8004 16730 8016
rect 16898 8007 16956 8013
rect 16898 8004 16910 8007
rect 16724 7976 16910 8004
rect 16724 7964 16730 7976
rect 16898 7973 16910 7976
rect 16944 7973 16956 8007
rect 16898 7967 16956 7973
rect 17862 7964 17868 8016
rect 17920 8004 17926 8016
rect 18509 8007 18567 8013
rect 18509 8004 18521 8007
rect 17920 7976 18521 8004
rect 17920 7964 17926 7976
rect 18509 7973 18521 7976
rect 18555 7973 18567 8007
rect 18509 7967 18567 7973
rect 18782 7964 18788 8016
rect 18840 8004 18846 8016
rect 19061 8007 19119 8013
rect 19061 8004 19073 8007
rect 18840 7976 19073 8004
rect 18840 7964 18846 7976
rect 19061 7973 19073 7976
rect 19107 7973 19119 8007
rect 19061 7967 19119 7973
rect 14182 7936 14188 7948
rect 11480 7908 13676 7936
rect 14143 7908 14188 7936
rect 11480 7896 11486 7908
rect 14182 7896 14188 7908
rect 14240 7896 14246 7948
rect 15289 7939 15347 7945
rect 15289 7905 15301 7939
rect 15335 7936 15347 7939
rect 15470 7936 15476 7948
rect 15335 7908 15476 7936
rect 15335 7905 15347 7908
rect 15289 7899 15347 7905
rect 15470 7896 15476 7908
rect 15528 7936 15534 7948
rect 15746 7936 15752 7948
rect 15528 7908 15752 7936
rect 15528 7896 15534 7908
rect 15746 7896 15752 7908
rect 15804 7896 15810 7948
rect 16574 7936 16580 7948
rect 16535 7908 16580 7936
rect 16574 7896 16580 7908
rect 16632 7896 16638 7948
rect 4724 7868 4752 7896
rect 8110 7868 8116 7880
rect 4724 7840 8116 7868
rect 8110 7828 8116 7840
rect 8168 7828 8174 7880
rect 8757 7871 8815 7877
rect 8757 7837 8769 7871
rect 8803 7868 8815 7871
rect 9306 7868 9312 7880
rect 8803 7840 9312 7868
rect 8803 7837 8815 7840
rect 8757 7831 8815 7837
rect 9306 7828 9312 7840
rect 9364 7828 9370 7880
rect 11609 7871 11667 7877
rect 11609 7837 11621 7871
rect 11655 7868 11667 7871
rect 12342 7868 12348 7880
rect 11655 7840 12348 7868
rect 11655 7837 11667 7840
rect 11609 7831 11667 7837
rect 12342 7828 12348 7840
rect 12400 7828 12406 7880
rect 12437 7871 12495 7877
rect 12437 7837 12449 7871
rect 12483 7868 12495 7871
rect 13170 7868 13176 7880
rect 12483 7840 13176 7868
rect 12483 7837 12495 7840
rect 12437 7831 12495 7837
rect 13170 7828 13176 7840
rect 13228 7828 13234 7880
rect 18417 7871 18475 7877
rect 18417 7837 18429 7871
rect 18463 7868 18475 7871
rect 19150 7868 19156 7880
rect 18463 7840 19156 7868
rect 18463 7837 18475 7840
rect 18417 7831 18475 7837
rect 19150 7828 19156 7840
rect 19208 7828 19214 7880
rect 4755 7803 4813 7809
rect 4755 7769 4767 7803
rect 4801 7800 4813 7803
rect 5534 7800 5540 7812
rect 4801 7772 5540 7800
rect 4801 7769 4813 7772
rect 4755 7763 4813 7769
rect 5534 7760 5540 7772
rect 5592 7760 5598 7812
rect 6914 7760 6920 7812
rect 6972 7800 6978 7812
rect 7009 7803 7067 7809
rect 7009 7800 7021 7803
rect 6972 7772 7021 7800
rect 6972 7760 6978 7772
rect 7009 7769 7021 7772
rect 7055 7769 7067 7803
rect 7009 7763 7067 7769
rect 13357 7803 13415 7809
rect 13357 7769 13369 7803
rect 13403 7800 13415 7803
rect 14001 7803 14059 7809
rect 14001 7800 14013 7803
rect 13403 7772 14013 7800
rect 13403 7769 13415 7772
rect 13357 7763 13415 7769
rect 14001 7769 14013 7772
rect 14047 7800 14059 7803
rect 14182 7800 14188 7812
rect 14047 7772 14188 7800
rect 14047 7769 14059 7772
rect 14001 7763 14059 7769
rect 14182 7760 14188 7772
rect 14240 7760 14246 7812
rect 2682 7732 2688 7744
rect 2643 7704 2688 7732
rect 2682 7692 2688 7704
rect 2740 7692 2746 7744
rect 9493 7735 9551 7741
rect 9493 7701 9505 7735
rect 9539 7732 9551 7735
rect 9582 7732 9588 7744
rect 9539 7704 9588 7732
rect 9539 7701 9551 7704
rect 9493 7695 9551 7701
rect 9582 7692 9588 7704
rect 9640 7692 9646 7744
rect 9999 7735 10057 7741
rect 9999 7701 10011 7735
rect 10045 7732 10057 7735
rect 10134 7732 10140 7744
rect 10045 7704 10140 7732
rect 10045 7701 10057 7704
rect 9999 7695 10057 7701
rect 10134 7692 10140 7704
rect 10192 7692 10198 7744
rect 14369 7735 14427 7741
rect 14369 7701 14381 7735
rect 14415 7732 14427 7735
rect 14734 7732 14740 7744
rect 14415 7704 14740 7732
rect 14415 7701 14427 7704
rect 14369 7695 14427 7701
rect 14734 7692 14740 7704
rect 14792 7692 14798 7744
rect 17954 7692 17960 7744
rect 18012 7732 18018 7744
rect 18049 7735 18107 7741
rect 18049 7732 18061 7735
rect 18012 7704 18061 7732
rect 18012 7692 18018 7704
rect 18049 7701 18061 7704
rect 18095 7701 18107 7735
rect 18049 7695 18107 7701
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1578 7528 1584 7540
rect 1539 7500 1584 7528
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 2130 7528 2136 7540
rect 2091 7500 2136 7528
rect 2130 7488 2136 7500
rect 2188 7488 2194 7540
rect 2774 7488 2780 7540
rect 2832 7528 2838 7540
rect 3050 7528 3056 7540
rect 2832 7500 3056 7528
rect 2832 7488 2838 7500
rect 3050 7488 3056 7500
rect 3108 7528 3114 7540
rect 3878 7528 3884 7540
rect 3108 7500 3884 7528
rect 3108 7488 3114 7500
rect 3878 7488 3884 7500
rect 3936 7488 3942 7540
rect 5997 7531 6055 7537
rect 5997 7497 6009 7531
rect 6043 7528 6055 7531
rect 6362 7528 6368 7540
rect 6043 7500 6368 7528
rect 6043 7497 6055 7500
rect 5997 7491 6055 7497
rect 6362 7488 6368 7500
rect 6420 7488 6426 7540
rect 7098 7528 7104 7540
rect 7059 7500 7104 7528
rect 7098 7488 7104 7500
rect 7156 7488 7162 7540
rect 8662 7528 8668 7540
rect 8623 7500 8668 7528
rect 8662 7488 8668 7500
rect 8720 7528 8726 7540
rect 8941 7531 8999 7537
rect 8941 7528 8953 7531
rect 8720 7500 8953 7528
rect 8720 7488 8726 7500
rect 8941 7497 8953 7500
rect 8987 7497 8999 7531
rect 8941 7491 8999 7497
rect 10042 7488 10048 7540
rect 10100 7528 10106 7540
rect 10505 7531 10563 7537
rect 10505 7528 10517 7531
rect 10100 7500 10517 7528
rect 10100 7488 10106 7500
rect 10505 7497 10517 7500
rect 10551 7497 10563 7531
rect 10505 7491 10563 7497
rect 10965 7531 11023 7537
rect 10965 7497 10977 7531
rect 11011 7528 11023 7531
rect 11146 7528 11152 7540
rect 11011 7500 11152 7528
rect 11011 7497 11023 7500
rect 10965 7491 11023 7497
rect 11146 7488 11152 7500
rect 11204 7488 11210 7540
rect 11790 7488 11796 7540
rect 11848 7528 11854 7540
rect 12161 7531 12219 7537
rect 12161 7528 12173 7531
rect 11848 7500 12173 7528
rect 11848 7488 11854 7500
rect 12161 7497 12173 7500
rect 12207 7497 12219 7531
rect 12161 7491 12219 7497
rect 13170 7488 13176 7540
rect 13228 7528 13234 7540
rect 13449 7531 13507 7537
rect 13449 7528 13461 7531
rect 13228 7500 13461 7528
rect 13228 7488 13234 7500
rect 13449 7497 13461 7500
rect 13495 7497 13507 7531
rect 13449 7491 13507 7497
rect 13909 7531 13967 7537
rect 13909 7497 13921 7531
rect 13955 7528 13967 7531
rect 14090 7528 14096 7540
rect 13955 7500 14096 7528
rect 13955 7497 13967 7500
rect 13909 7491 13967 7497
rect 14090 7488 14096 7500
rect 14148 7488 14154 7540
rect 17129 7531 17187 7537
rect 17129 7497 17141 7531
rect 17175 7528 17187 7531
rect 17678 7528 17684 7540
rect 17175 7500 17684 7528
rect 17175 7497 17187 7500
rect 17129 7491 17187 7497
rect 17678 7488 17684 7500
rect 17736 7528 17742 7540
rect 17862 7528 17868 7540
rect 17736 7500 17868 7528
rect 17736 7488 17742 7500
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 18230 7488 18236 7540
rect 18288 7528 18294 7540
rect 18506 7528 18512 7540
rect 18288 7500 18512 7528
rect 18288 7488 18294 7500
rect 18506 7488 18512 7500
rect 18564 7488 18570 7540
rect 19150 7528 19156 7540
rect 19111 7500 19156 7528
rect 19150 7488 19156 7500
rect 19208 7488 19214 7540
rect 20165 7531 20223 7537
rect 20165 7497 20177 7531
rect 20211 7528 20223 7531
rect 20254 7528 20260 7540
rect 20211 7500 20260 7528
rect 20211 7497 20223 7500
rect 20165 7491 20223 7497
rect 6270 7460 6276 7472
rect 6231 7432 6276 7460
rect 6270 7420 6276 7432
rect 6328 7420 6334 7472
rect 7653 7463 7711 7469
rect 7653 7429 7665 7463
rect 7699 7460 7711 7463
rect 9490 7460 9496 7472
rect 7699 7432 9496 7460
rect 7699 7429 7711 7432
rect 7653 7423 7711 7429
rect 2314 7352 2320 7404
rect 2372 7392 2378 7404
rect 2961 7395 3019 7401
rect 2961 7392 2973 7395
rect 2372 7364 2973 7392
rect 2372 7352 2378 7364
rect 2961 7361 2973 7364
rect 3007 7392 3019 7395
rect 3786 7392 3792 7404
rect 3007 7364 3792 7392
rect 3007 7361 3019 7364
rect 2961 7355 3019 7361
rect 3786 7352 3792 7364
rect 3844 7352 3850 7404
rect 4338 7352 4344 7404
rect 4396 7392 4402 7404
rect 4709 7395 4767 7401
rect 4709 7392 4721 7395
rect 4396 7364 4721 7392
rect 4396 7352 4402 7364
rect 4709 7361 4721 7364
rect 4755 7392 4767 7395
rect 5074 7392 5080 7404
rect 4755 7364 5080 7392
rect 4755 7361 4767 7364
rect 4709 7355 4767 7361
rect 5074 7352 5080 7364
rect 5132 7352 5138 7404
rect 7745 7395 7803 7401
rect 7745 7361 7757 7395
rect 7791 7392 7803 7395
rect 8018 7392 8024 7404
rect 7791 7364 8024 7392
rect 7791 7361 7803 7364
rect 7745 7355 7803 7361
rect 8018 7352 8024 7364
rect 8076 7352 8082 7404
rect 1394 7324 1400 7336
rect 1355 7296 1400 7324
rect 1394 7284 1400 7296
rect 1452 7284 1458 7336
rect 8128 7268 8156 7432
rect 9490 7420 9496 7432
rect 9548 7420 9554 7472
rect 12894 7392 12900 7404
rect 12855 7364 12900 7392
rect 12894 7352 12900 7364
rect 12952 7392 12958 7404
rect 14090 7392 14096 7404
rect 12952 7364 14096 7392
rect 12952 7352 12958 7364
rect 14090 7352 14096 7364
rect 14148 7352 14154 7404
rect 14366 7392 14372 7404
rect 14327 7364 14372 7392
rect 14366 7352 14372 7364
rect 14424 7352 14430 7404
rect 15749 7395 15807 7401
rect 15749 7361 15761 7395
rect 15795 7392 15807 7395
rect 16206 7392 16212 7404
rect 15795 7364 16212 7392
rect 15795 7361 15807 7364
rect 15749 7355 15807 7361
rect 16206 7352 16212 7364
rect 16264 7352 16270 7404
rect 18598 7392 18604 7404
rect 18559 7364 18604 7392
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 8938 7284 8944 7336
rect 8996 7324 9002 7336
rect 9214 7324 9220 7336
rect 8996 7296 9220 7324
rect 8996 7284 9002 7296
rect 9214 7284 9220 7296
rect 9272 7284 9278 7336
rect 15286 7284 15292 7336
rect 15344 7324 15350 7336
rect 16025 7327 16083 7333
rect 16025 7324 16037 7327
rect 15344 7296 16037 7324
rect 15344 7284 15350 7296
rect 16025 7293 16037 7296
rect 16071 7293 16083 7327
rect 16025 7287 16083 7293
rect 19680 7327 19738 7333
rect 19680 7293 19692 7327
rect 19726 7324 19738 7327
rect 20180 7324 20208 7491
rect 20254 7488 20260 7500
rect 20312 7488 20318 7540
rect 19726 7296 20208 7324
rect 19726 7293 19738 7296
rect 19680 7287 19738 7293
rect 2590 7216 2596 7268
rect 2648 7256 2654 7268
rect 2869 7259 2927 7265
rect 2869 7256 2881 7259
rect 2648 7228 2881 7256
rect 2648 7216 2654 7228
rect 2869 7225 2881 7228
rect 2915 7256 2927 7259
rect 3323 7259 3381 7265
rect 3323 7256 3335 7259
rect 2915 7228 3335 7256
rect 2915 7225 2927 7228
rect 2869 7219 2927 7225
rect 3323 7225 3335 7228
rect 3369 7256 3381 7259
rect 4249 7259 4307 7265
rect 4249 7256 4261 7259
rect 3369 7228 4261 7256
rect 3369 7225 3381 7228
rect 3323 7219 3381 7225
rect 4249 7225 4261 7228
rect 4295 7256 4307 7259
rect 5071 7259 5129 7265
rect 5071 7256 5083 7259
rect 4295 7228 5083 7256
rect 4295 7225 4307 7228
rect 4249 7219 4307 7225
rect 5071 7225 5083 7228
rect 5117 7256 5129 7259
rect 6270 7256 6276 7268
rect 5117 7228 6276 7256
rect 5117 7225 5129 7228
rect 5071 7219 5129 7225
rect 6270 7216 6276 7228
rect 6328 7216 6334 7268
rect 8110 7265 8116 7268
rect 8107 7256 8116 7265
rect 8023 7228 8116 7256
rect 8107 7219 8116 7228
rect 8110 7216 8116 7219
rect 8168 7216 8174 7268
rect 9585 7259 9643 7265
rect 9585 7225 9597 7259
rect 9631 7225 9643 7259
rect 9585 7219 9643 7225
rect 4617 7191 4675 7197
rect 4617 7157 4629 7191
rect 4663 7188 4675 7191
rect 4706 7188 4712 7200
rect 4663 7160 4712 7188
rect 4663 7157 4675 7160
rect 4617 7151 4675 7157
rect 4706 7148 4712 7160
rect 4764 7188 4770 7200
rect 5350 7188 5356 7200
rect 4764 7160 5356 7188
rect 4764 7148 4770 7160
rect 5350 7148 5356 7160
rect 5408 7148 5414 7200
rect 5442 7148 5448 7200
rect 5500 7188 5506 7200
rect 5629 7191 5687 7197
rect 5629 7188 5641 7191
rect 5500 7160 5641 7188
rect 5500 7148 5506 7160
rect 5629 7157 5641 7160
rect 5675 7157 5687 7191
rect 5629 7151 5687 7157
rect 9214 7148 9220 7200
rect 9272 7188 9278 7200
rect 9309 7191 9367 7197
rect 9309 7188 9321 7191
rect 9272 7160 9321 7188
rect 9272 7148 9278 7160
rect 9309 7157 9321 7160
rect 9355 7157 9367 7191
rect 9309 7151 9367 7157
rect 9490 7148 9496 7200
rect 9548 7188 9554 7200
rect 9600 7188 9628 7219
rect 9674 7216 9680 7268
rect 9732 7256 9738 7268
rect 10229 7259 10287 7265
rect 9732 7228 9777 7256
rect 9732 7216 9738 7228
rect 10229 7225 10241 7259
rect 10275 7256 10287 7259
rect 10686 7256 10692 7268
rect 10275 7228 10692 7256
rect 10275 7225 10287 7228
rect 10229 7219 10287 7225
rect 10686 7216 10692 7228
rect 10744 7216 10750 7268
rect 11333 7259 11391 7265
rect 11333 7225 11345 7259
rect 11379 7256 11391 7259
rect 12526 7256 12532 7268
rect 11379 7228 12532 7256
rect 11379 7225 11391 7228
rect 11333 7219 11391 7225
rect 12526 7216 12532 7228
rect 12584 7216 12590 7268
rect 12621 7259 12679 7265
rect 12621 7225 12633 7259
rect 12667 7225 12679 7259
rect 12621 7219 12679 7225
rect 11790 7188 11796 7200
rect 9548 7160 9628 7188
rect 11751 7160 11796 7188
rect 9548 7148 9554 7160
rect 11790 7148 11796 7160
rect 11848 7148 11854 7200
rect 12250 7148 12256 7200
rect 12308 7188 12314 7200
rect 12636 7188 12664 7219
rect 14182 7216 14188 7268
rect 14240 7256 14246 7268
rect 16040 7256 16068 7287
rect 16530 7259 16588 7265
rect 16530 7256 16542 7259
rect 14240 7228 14285 7256
rect 16040 7228 16542 7256
rect 14240 7216 14246 7228
rect 16530 7225 16542 7228
rect 16576 7256 16588 7259
rect 17405 7259 17463 7265
rect 17405 7256 17417 7259
rect 16576 7228 17417 7256
rect 16576 7225 16588 7228
rect 16530 7219 16588 7225
rect 17405 7225 17417 7228
rect 17451 7225 17463 7259
rect 18138 7256 18144 7268
rect 18099 7228 18144 7256
rect 17405 7219 17463 7225
rect 18138 7216 18144 7228
rect 18196 7216 18202 7268
rect 18233 7259 18291 7265
rect 18233 7225 18245 7259
rect 18279 7225 18291 7259
rect 18233 7219 18291 7225
rect 12308 7160 12664 7188
rect 15381 7191 15439 7197
rect 12308 7148 12314 7160
rect 15381 7157 15393 7191
rect 15427 7188 15439 7191
rect 15470 7188 15476 7200
rect 15427 7160 15476 7188
rect 15427 7157 15439 7160
rect 15381 7151 15439 7157
rect 15470 7148 15476 7160
rect 15528 7148 15534 7200
rect 17954 7148 17960 7200
rect 18012 7188 18018 7200
rect 18248 7188 18276 7219
rect 18012 7160 18276 7188
rect 18012 7148 18018 7160
rect 19334 7148 19340 7200
rect 19392 7188 19398 7200
rect 19751 7191 19809 7197
rect 19751 7188 19763 7191
rect 19392 7160 19763 7188
rect 19392 7148 19398 7160
rect 19751 7157 19763 7160
rect 19797 7157 19809 7191
rect 19751 7151 19809 7157
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 1394 6944 1400 6996
rect 1452 6984 1458 6996
rect 1535 6987 1593 6993
rect 1535 6984 1547 6987
rect 1452 6956 1547 6984
rect 1452 6944 1458 6956
rect 1535 6953 1547 6956
rect 1581 6984 1593 6987
rect 2498 6984 2504 6996
rect 1581 6956 2504 6984
rect 1581 6953 1593 6956
rect 1535 6947 1593 6953
rect 2498 6944 2504 6956
rect 2556 6944 2562 6996
rect 5074 6984 5080 6996
rect 5035 6956 5080 6984
rect 5074 6944 5080 6956
rect 5132 6944 5138 6996
rect 7745 6987 7803 6993
rect 7745 6953 7757 6987
rect 7791 6984 7803 6987
rect 8018 6984 8024 6996
rect 7791 6956 8024 6984
rect 7791 6953 7803 6956
rect 7745 6947 7803 6953
rect 8018 6944 8024 6956
rect 8076 6944 8082 6996
rect 9214 6944 9220 6996
rect 9272 6984 9278 6996
rect 9674 6984 9680 6996
rect 9272 6956 9680 6984
rect 9272 6944 9278 6956
rect 9674 6944 9680 6956
rect 9732 6944 9738 6996
rect 10965 6987 11023 6993
rect 10965 6953 10977 6987
rect 11011 6984 11023 6987
rect 11422 6984 11428 6996
rect 11011 6956 11428 6984
rect 11011 6953 11023 6956
rect 10965 6947 11023 6953
rect 11422 6944 11428 6956
rect 11480 6944 11486 6996
rect 12526 6984 12532 6996
rect 12487 6956 12532 6984
rect 12526 6944 12532 6956
rect 12584 6944 12590 6996
rect 14090 6944 14096 6996
rect 14148 6984 14154 6996
rect 14185 6987 14243 6993
rect 14185 6984 14197 6987
rect 14148 6956 14197 6984
rect 14148 6944 14154 6956
rect 14185 6953 14197 6956
rect 14231 6953 14243 6987
rect 15378 6984 15384 6996
rect 15339 6956 15384 6984
rect 14185 6947 14243 6953
rect 15378 6944 15384 6956
rect 15436 6944 15442 6996
rect 16574 6984 16580 6996
rect 16535 6956 16580 6984
rect 16574 6944 16580 6956
rect 16632 6944 16638 6996
rect 2593 6919 2651 6925
rect 2593 6885 2605 6919
rect 2639 6916 2651 6919
rect 2682 6916 2688 6928
rect 2639 6888 2688 6916
rect 2639 6885 2651 6888
rect 2593 6879 2651 6885
rect 2682 6876 2688 6888
rect 2740 6876 2746 6928
rect 3878 6876 3884 6928
rect 3936 6916 3942 6928
rect 4246 6916 4252 6928
rect 3936 6888 4252 6916
rect 3936 6876 3942 6888
rect 4246 6876 4252 6888
rect 4304 6876 4310 6928
rect 5813 6919 5871 6925
rect 5813 6885 5825 6919
rect 5859 6916 5871 6919
rect 6086 6916 6092 6928
rect 5859 6888 6092 6916
rect 5859 6885 5871 6888
rect 5813 6879 5871 6885
rect 6086 6876 6092 6888
rect 6144 6876 6150 6928
rect 8110 6876 8116 6928
rect 8168 6925 8174 6928
rect 8168 6919 8216 6925
rect 8168 6885 8170 6919
rect 8204 6885 8216 6919
rect 8168 6879 8216 6885
rect 8168 6876 8174 6879
rect 9306 6876 9312 6928
rect 9364 6916 9370 6928
rect 9858 6916 9864 6928
rect 9364 6888 9864 6916
rect 9364 6876 9370 6888
rect 9858 6876 9864 6888
rect 9916 6876 9922 6928
rect 11603 6919 11661 6925
rect 11603 6885 11615 6919
rect 11649 6916 11661 6919
rect 11698 6916 11704 6928
rect 11649 6888 11704 6916
rect 11649 6885 11661 6888
rect 11603 6879 11661 6885
rect 11698 6876 11704 6888
rect 11756 6876 11762 6928
rect 12342 6876 12348 6928
rect 12400 6916 12406 6928
rect 12805 6919 12863 6925
rect 12805 6916 12817 6919
rect 12400 6888 12817 6916
rect 12400 6876 12406 6888
rect 12805 6885 12817 6888
rect 12851 6885 12863 6919
rect 13354 6916 13360 6928
rect 13315 6888 13360 6916
rect 12805 6879 12863 6885
rect 13354 6876 13360 6888
rect 13412 6876 13418 6928
rect 13909 6919 13967 6925
rect 13909 6885 13921 6919
rect 13955 6916 13967 6919
rect 14366 6916 14372 6928
rect 13955 6888 14372 6916
rect 13955 6885 13967 6888
rect 13909 6879 13967 6885
rect 14366 6876 14372 6888
rect 14424 6876 14430 6928
rect 17678 6916 17684 6928
rect 17639 6888 17684 6916
rect 17678 6876 17684 6888
rect 17736 6876 17742 6928
rect 1464 6851 1522 6857
rect 1464 6817 1476 6851
rect 1510 6817 1522 6851
rect 1464 6811 1522 6817
rect 1949 6851 2007 6857
rect 1949 6817 1961 6851
rect 1995 6848 2007 6851
rect 2314 6848 2320 6860
rect 1995 6820 2320 6848
rect 1995 6817 2007 6820
rect 1949 6811 2007 6817
rect 1479 6712 1507 6811
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 3694 6848 3700 6860
rect 3655 6820 3700 6848
rect 3694 6808 3700 6820
rect 3752 6808 3758 6860
rect 7834 6848 7840 6860
rect 7795 6820 7840 6848
rect 7834 6808 7840 6820
rect 7892 6808 7898 6860
rect 14642 6808 14648 6860
rect 14700 6848 14706 6860
rect 15289 6851 15347 6857
rect 15289 6848 15301 6851
rect 14700 6820 15301 6848
rect 14700 6808 14706 6820
rect 15289 6817 15301 6820
rect 15335 6848 15347 6851
rect 15562 6848 15568 6860
rect 15335 6820 15568 6848
rect 15335 6817 15347 6820
rect 15289 6811 15347 6817
rect 15562 6808 15568 6820
rect 15620 6808 15626 6860
rect 15841 6851 15899 6857
rect 15841 6817 15853 6851
rect 15887 6848 15899 6851
rect 16390 6848 16396 6860
rect 15887 6820 16396 6848
rect 15887 6817 15899 6820
rect 15841 6811 15899 6817
rect 16390 6808 16396 6820
rect 16448 6808 16454 6860
rect 19058 6848 19064 6860
rect 19019 6820 19064 6848
rect 19058 6808 19064 6820
rect 19116 6808 19122 6860
rect 19426 6808 19432 6860
rect 19484 6848 19490 6860
rect 19521 6851 19579 6857
rect 19521 6848 19533 6851
rect 19484 6820 19533 6848
rect 19484 6808 19490 6820
rect 19521 6817 19533 6820
rect 19567 6817 19579 6851
rect 19521 6811 19579 6817
rect 2130 6740 2136 6792
rect 2188 6780 2194 6792
rect 2501 6783 2559 6789
rect 2501 6780 2513 6783
rect 2188 6752 2513 6780
rect 2188 6740 2194 6752
rect 2501 6749 2513 6752
rect 2547 6749 2559 6783
rect 4154 6780 4160 6792
rect 4115 6752 4160 6780
rect 2501 6743 2559 6749
rect 4154 6740 4160 6752
rect 4212 6740 4218 6792
rect 4433 6783 4491 6789
rect 4433 6749 4445 6783
rect 4479 6749 4491 6783
rect 4433 6743 4491 6749
rect 2317 6715 2375 6721
rect 1479 6684 2084 6712
rect 2056 6644 2084 6684
rect 2317 6681 2329 6715
rect 2363 6712 2375 6715
rect 2682 6712 2688 6724
rect 2363 6684 2688 6712
rect 2363 6681 2375 6684
rect 2317 6675 2375 6681
rect 2682 6672 2688 6684
rect 2740 6672 2746 6724
rect 3053 6715 3111 6721
rect 3053 6681 3065 6715
rect 3099 6712 3111 6715
rect 3510 6712 3516 6724
rect 3099 6684 3516 6712
rect 3099 6681 3111 6684
rect 3053 6675 3111 6681
rect 3068 6644 3096 6675
rect 3510 6672 3516 6684
rect 3568 6712 3574 6724
rect 4448 6712 4476 6743
rect 5534 6740 5540 6792
rect 5592 6780 5598 6792
rect 5721 6783 5779 6789
rect 5721 6780 5733 6783
rect 5592 6752 5733 6780
rect 5592 6740 5598 6752
rect 5721 6749 5733 6752
rect 5767 6749 5779 6783
rect 5994 6780 6000 6792
rect 5955 6752 6000 6780
rect 5721 6743 5779 6749
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 9398 6740 9404 6792
rect 9456 6780 9462 6792
rect 9769 6783 9827 6789
rect 9769 6780 9781 6783
rect 9456 6752 9781 6780
rect 9456 6740 9462 6752
rect 9769 6749 9781 6752
rect 9815 6780 9827 6783
rect 10042 6780 10048 6792
rect 9815 6752 10048 6780
rect 9815 6749 9827 6752
rect 9769 6743 9827 6749
rect 10042 6740 10048 6752
rect 10100 6740 10106 6792
rect 11241 6783 11299 6789
rect 11241 6749 11253 6783
rect 11287 6780 11299 6783
rect 11514 6780 11520 6792
rect 11287 6752 11520 6780
rect 11287 6749 11299 6752
rect 11241 6743 11299 6749
rect 11514 6740 11520 6752
rect 11572 6740 11578 6792
rect 11606 6740 11612 6792
rect 11664 6780 11670 6792
rect 13265 6783 13323 6789
rect 13265 6780 13277 6783
rect 11664 6752 13277 6780
rect 11664 6740 11670 6752
rect 13265 6749 13277 6752
rect 13311 6780 13323 6783
rect 13998 6780 14004 6792
rect 13311 6752 14004 6780
rect 13311 6749 13323 6752
rect 13265 6743 13323 6749
rect 13998 6740 14004 6752
rect 14056 6740 14062 6792
rect 17586 6780 17592 6792
rect 17547 6752 17592 6780
rect 17586 6740 17592 6752
rect 17644 6740 17650 6792
rect 19610 6780 19616 6792
rect 19571 6752 19616 6780
rect 19610 6740 19616 6752
rect 19668 6740 19674 6792
rect 3568 6684 4476 6712
rect 3568 6672 3574 6684
rect 9306 6672 9312 6724
rect 9364 6712 9370 6724
rect 10321 6715 10379 6721
rect 10321 6712 10333 6715
rect 9364 6684 10333 6712
rect 9364 6672 9370 6684
rect 10321 6681 10333 6684
rect 10367 6681 10379 6715
rect 18138 6712 18144 6724
rect 18051 6684 18144 6712
rect 10321 6675 10379 6681
rect 18138 6672 18144 6684
rect 18196 6712 18202 6724
rect 18196 6684 18920 6712
rect 18196 6672 18202 6684
rect 18892 6656 18920 6684
rect 2056 6616 3096 6644
rect 3694 6604 3700 6656
rect 3752 6644 3758 6656
rect 5537 6647 5595 6653
rect 5537 6644 5549 6647
rect 3752 6616 5549 6644
rect 3752 6604 3758 6616
rect 5537 6613 5549 6616
rect 5583 6644 5595 6647
rect 6178 6644 6184 6656
rect 5583 6616 6184 6644
rect 5583 6613 5595 6616
rect 5537 6607 5595 6613
rect 6178 6604 6184 6616
rect 6236 6644 6242 6656
rect 6641 6647 6699 6653
rect 6641 6644 6653 6647
rect 6236 6616 6653 6644
rect 6236 6604 6242 6616
rect 6641 6613 6653 6616
rect 6687 6613 6699 6647
rect 6641 6607 6699 6613
rect 8662 6604 8668 6656
rect 8720 6644 8726 6656
rect 8757 6647 8815 6653
rect 8757 6644 8769 6647
rect 8720 6616 8769 6644
rect 8720 6604 8726 6616
rect 8757 6613 8769 6616
rect 8803 6644 8815 6647
rect 9214 6644 9220 6656
rect 8803 6616 9220 6644
rect 8803 6613 8815 6616
rect 8757 6607 8815 6613
rect 9214 6604 9220 6616
rect 9272 6604 9278 6656
rect 9490 6644 9496 6656
rect 9451 6616 9496 6644
rect 9490 6604 9496 6616
rect 9548 6604 9554 6656
rect 11054 6604 11060 6656
rect 11112 6644 11118 6656
rect 11790 6644 11796 6656
rect 11112 6616 11796 6644
rect 11112 6604 11118 6616
rect 11790 6604 11796 6616
rect 11848 6644 11854 6656
rect 12161 6647 12219 6653
rect 12161 6644 12173 6647
rect 11848 6616 12173 6644
rect 11848 6604 11854 6616
rect 12161 6613 12173 6616
rect 12207 6644 12219 6647
rect 12250 6644 12256 6656
rect 12207 6616 12256 6644
rect 12207 6613 12219 6616
rect 12161 6607 12219 6613
rect 12250 6604 12256 6616
rect 12308 6604 12314 6656
rect 18046 6604 18052 6656
rect 18104 6644 18110 6656
rect 18509 6647 18567 6653
rect 18509 6644 18521 6647
rect 18104 6616 18521 6644
rect 18104 6604 18110 6616
rect 18509 6613 18521 6616
rect 18555 6613 18567 6647
rect 18874 6644 18880 6656
rect 18835 6616 18880 6644
rect 18509 6607 18567 6613
rect 18874 6604 18880 6616
rect 18932 6604 18938 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 2130 6440 2136 6452
rect 2091 6412 2136 6440
rect 2130 6400 2136 6412
rect 2188 6400 2194 6452
rect 2501 6443 2559 6449
rect 2501 6409 2513 6443
rect 2547 6440 2559 6443
rect 2590 6440 2596 6452
rect 2547 6412 2596 6440
rect 2547 6409 2559 6412
rect 2501 6403 2559 6409
rect 2590 6400 2596 6412
rect 2648 6400 2654 6452
rect 4246 6440 4252 6452
rect 4207 6412 4252 6440
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 5534 6400 5540 6452
rect 5592 6440 5598 6452
rect 6549 6443 6607 6449
rect 6549 6440 6561 6443
rect 5592 6412 6561 6440
rect 5592 6400 5598 6412
rect 6549 6409 6561 6412
rect 6595 6409 6607 6443
rect 6549 6403 6607 6409
rect 7834 6400 7840 6452
rect 7892 6440 7898 6452
rect 8205 6443 8263 6449
rect 8205 6440 8217 6443
rect 7892 6412 8217 6440
rect 7892 6400 7898 6412
rect 8205 6409 8217 6412
rect 8251 6409 8263 6443
rect 8205 6403 8263 6409
rect 9677 6443 9735 6449
rect 9677 6409 9689 6443
rect 9723 6440 9735 6443
rect 9858 6440 9864 6452
rect 9723 6412 9864 6440
rect 9723 6409 9735 6412
rect 9677 6403 9735 6409
rect 9858 6400 9864 6412
rect 9916 6400 9922 6452
rect 11333 6443 11391 6449
rect 11333 6409 11345 6443
rect 11379 6440 11391 6443
rect 11698 6440 11704 6452
rect 11379 6412 11704 6440
rect 11379 6409 11391 6412
rect 11333 6403 11391 6409
rect 11698 6400 11704 6412
rect 11756 6440 11762 6452
rect 12161 6443 12219 6449
rect 12161 6440 12173 6443
rect 11756 6412 12173 6440
rect 11756 6400 11762 6412
rect 12161 6409 12173 6412
rect 12207 6409 12219 6443
rect 13354 6440 13360 6452
rect 13315 6412 13360 6440
rect 12161 6403 12219 6409
rect 1578 6372 1584 6384
rect 1539 6344 1584 6372
rect 1578 6332 1584 6344
rect 1636 6332 1642 6384
rect 4154 6332 4160 6384
rect 4212 6372 4218 6384
rect 4617 6375 4675 6381
rect 4617 6372 4629 6375
rect 4212 6344 4629 6372
rect 4212 6332 4218 6344
rect 4617 6341 4629 6344
rect 4663 6372 4675 6375
rect 5813 6375 5871 6381
rect 5813 6372 5825 6375
rect 4663 6344 5825 6372
rect 4663 6341 4675 6344
rect 4617 6335 4675 6341
rect 5813 6341 5825 6344
rect 5859 6372 5871 6375
rect 5994 6372 6000 6384
rect 5859 6344 6000 6372
rect 5859 6341 5871 6344
rect 5813 6335 5871 6341
rect 5994 6332 6000 6344
rect 6052 6332 6058 6384
rect 7929 6375 7987 6381
rect 7929 6341 7941 6375
rect 7975 6372 7987 6375
rect 8110 6372 8116 6384
rect 7975 6344 8116 6372
rect 7975 6341 7987 6344
rect 7929 6335 7987 6341
rect 8110 6332 8116 6344
rect 8168 6332 8174 6384
rect 2958 6304 2964 6316
rect 2919 6276 2964 6304
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 5258 6304 5264 6316
rect 5171 6276 5264 6304
rect 5258 6264 5264 6276
rect 5316 6304 5322 6316
rect 6963 6307 7021 6313
rect 6963 6304 6975 6307
rect 5316 6276 6975 6304
rect 5316 6264 5322 6276
rect 6963 6273 6975 6276
rect 7009 6273 7021 6307
rect 6963 6267 7021 6273
rect 8665 6307 8723 6313
rect 8665 6273 8677 6307
rect 8711 6304 8723 6307
rect 9030 6304 9036 6316
rect 8711 6276 9036 6304
rect 8711 6273 8723 6276
rect 8665 6267 8723 6273
rect 9030 6264 9036 6276
rect 9088 6304 9094 6316
rect 10686 6304 10692 6316
rect 9088 6276 10692 6304
rect 9088 6264 9094 6276
rect 10686 6264 10692 6276
rect 10744 6264 10750 6316
rect 1394 6236 1400 6248
rect 1355 6208 1400 6236
rect 1394 6196 1400 6208
rect 1452 6196 1458 6248
rect 6876 6239 6934 6245
rect 6876 6205 6888 6239
rect 6922 6236 6934 6239
rect 6922 6208 7420 6236
rect 6922 6205 6934 6208
rect 6876 6199 6934 6205
rect 3326 6177 3332 6180
rect 2869 6171 2927 6177
rect 2869 6137 2881 6171
rect 2915 6168 2927 6171
rect 3323 6168 3332 6177
rect 2915 6140 3332 6168
rect 2915 6137 2927 6140
rect 2869 6131 2927 6137
rect 3323 6131 3332 6140
rect 3326 6128 3332 6131
rect 3384 6128 3390 6180
rect 4706 6128 4712 6180
rect 4764 6168 4770 6180
rect 5077 6171 5135 6177
rect 5077 6168 5089 6171
rect 4764 6140 5089 6168
rect 4764 6128 4770 6140
rect 5077 6137 5089 6140
rect 5123 6168 5135 6171
rect 5353 6171 5411 6177
rect 5353 6168 5365 6171
rect 5123 6140 5365 6168
rect 5123 6137 5135 6140
rect 5077 6131 5135 6137
rect 5353 6137 5365 6140
rect 5399 6168 5411 6171
rect 5442 6168 5448 6180
rect 5399 6140 5448 6168
rect 5399 6137 5411 6140
rect 5353 6131 5411 6137
rect 5442 6128 5448 6140
rect 5500 6128 5506 6180
rect 7392 6112 7420 6208
rect 8754 6128 8760 6180
rect 8812 6168 8818 6180
rect 9306 6168 9312 6180
rect 8812 6140 8857 6168
rect 9267 6140 9312 6168
rect 8812 6128 8818 6140
rect 9306 6128 9312 6140
rect 9364 6128 9370 6180
rect 9858 6128 9864 6180
rect 9916 6168 9922 6180
rect 10229 6171 10287 6177
rect 10229 6168 10241 6171
rect 9916 6140 10241 6168
rect 9916 6128 9922 6140
rect 10229 6137 10241 6140
rect 10275 6137 10287 6171
rect 10229 6131 10287 6137
rect 10321 6171 10379 6177
rect 10321 6137 10333 6171
rect 10367 6137 10379 6171
rect 12176 6168 12204 6403
rect 13354 6400 13360 6412
rect 13412 6440 13418 6452
rect 13633 6443 13691 6449
rect 13633 6440 13645 6443
rect 13412 6412 13645 6440
rect 13412 6400 13418 6412
rect 13633 6409 13645 6412
rect 13679 6409 13691 6443
rect 13998 6440 14004 6452
rect 13959 6412 14004 6440
rect 13633 6403 13691 6409
rect 13998 6400 14004 6412
rect 14056 6400 14062 6452
rect 16390 6400 16396 6452
rect 16448 6440 16454 6452
rect 16577 6443 16635 6449
rect 16577 6440 16589 6443
rect 16448 6412 16589 6440
rect 16448 6400 16454 6412
rect 16577 6409 16589 6412
rect 16623 6409 16635 6443
rect 17770 6440 17776 6452
rect 17731 6412 17776 6440
rect 16577 6403 16635 6409
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 19058 6440 19064 6452
rect 19019 6412 19064 6440
rect 19058 6400 19064 6412
rect 19116 6400 19122 6452
rect 19426 6440 19432 6452
rect 19387 6412 19432 6440
rect 19426 6400 19432 6412
rect 19484 6400 19490 6452
rect 14550 6372 14556 6384
rect 14419 6344 14556 6372
rect 12342 6264 12348 6316
rect 12400 6304 12406 6316
rect 12437 6307 12495 6313
rect 12437 6304 12449 6307
rect 12400 6276 12449 6304
rect 12400 6264 12406 6276
rect 12437 6273 12449 6276
rect 12483 6273 12495 6307
rect 12437 6267 12495 6273
rect 14419 6245 14447 6344
rect 14550 6332 14556 6344
rect 14608 6372 14614 6384
rect 14826 6372 14832 6384
rect 14608 6344 14832 6372
rect 14608 6332 14614 6344
rect 14826 6332 14832 6344
rect 14884 6332 14890 6384
rect 17497 6375 17555 6381
rect 17497 6341 17509 6375
rect 17543 6372 17555 6375
rect 17678 6372 17684 6384
rect 17543 6344 17684 6372
rect 17543 6341 17555 6344
rect 17497 6335 17555 6341
rect 17678 6332 17684 6344
rect 17736 6372 17742 6384
rect 17954 6372 17960 6384
rect 17736 6344 17960 6372
rect 17736 6332 17742 6344
rect 17954 6332 17960 6344
rect 18012 6332 18018 6384
rect 16945 6307 17003 6313
rect 16945 6304 16957 6307
rect 15396 6276 16957 6304
rect 14415 6239 14473 6245
rect 14415 6205 14427 6239
rect 14461 6205 14473 6239
rect 14415 6199 14473 6205
rect 14826 6196 14832 6248
rect 14884 6236 14890 6248
rect 15396 6245 15424 6276
rect 16945 6273 16957 6276
rect 16991 6273 17003 6307
rect 16945 6267 17003 6273
rect 15381 6239 15439 6245
rect 15381 6236 15393 6239
rect 14884 6208 15393 6236
rect 14884 6196 14890 6208
rect 15381 6205 15393 6208
rect 15427 6205 15439 6239
rect 15381 6199 15439 6205
rect 16301 6239 16359 6245
rect 16301 6205 16313 6239
rect 16347 6236 16359 6239
rect 16574 6236 16580 6248
rect 16347 6208 16580 6236
rect 16347 6205 16359 6208
rect 16301 6199 16359 6205
rect 16574 6196 16580 6208
rect 16632 6196 16638 6248
rect 18785 6239 18843 6245
rect 18785 6205 18797 6239
rect 18831 6236 18843 6239
rect 18874 6236 18880 6248
rect 18831 6208 18880 6236
rect 18831 6205 18843 6208
rect 18785 6199 18843 6205
rect 18874 6196 18880 6208
rect 18932 6236 18938 6248
rect 19426 6236 19432 6248
rect 18932 6208 19432 6236
rect 18932 6196 18938 6208
rect 19426 6196 19432 6208
rect 19484 6196 19490 6248
rect 12710 6168 12716 6180
rect 12176 6140 12716 6168
rect 10321 6131 10379 6137
rect 3878 6100 3884 6112
rect 3839 6072 3884 6100
rect 3878 6060 3884 6072
rect 3936 6060 3942 6112
rect 5810 6060 5816 6112
rect 5868 6100 5874 6112
rect 6086 6100 6092 6112
rect 5868 6072 6092 6100
rect 5868 6060 5874 6072
rect 6086 6060 6092 6072
rect 6144 6100 6150 6112
rect 6181 6103 6239 6109
rect 6181 6100 6193 6103
rect 6144 6072 6193 6100
rect 6144 6060 6150 6072
rect 6181 6069 6193 6072
rect 6227 6069 6239 6103
rect 7374 6100 7380 6112
rect 7335 6072 7380 6100
rect 6181 6063 6239 6069
rect 7374 6060 7380 6072
rect 7432 6060 7438 6112
rect 9674 6060 9680 6112
rect 9732 6100 9738 6112
rect 9953 6103 10011 6109
rect 9953 6100 9965 6103
rect 9732 6072 9965 6100
rect 9732 6060 9738 6072
rect 9953 6069 9965 6072
rect 9999 6100 10011 6103
rect 10336 6100 10364 6131
rect 12710 6128 12716 6140
rect 12768 6177 12774 6180
rect 12768 6171 12816 6177
rect 12768 6137 12770 6171
rect 12804 6137 12816 6171
rect 12768 6131 12816 6137
rect 14507 6171 14565 6177
rect 14507 6137 14519 6171
rect 14553 6168 14565 6171
rect 15286 6168 15292 6180
rect 14553 6140 15292 6168
rect 14553 6137 14565 6140
rect 14507 6131 14565 6137
rect 12768 6128 12801 6131
rect 15286 6128 15292 6140
rect 15344 6128 15350 6180
rect 15702 6171 15760 6177
rect 15702 6168 15714 6171
rect 15396 6140 15714 6168
rect 9999 6072 10364 6100
rect 9999 6069 10011 6072
rect 9953 6063 10011 6069
rect 11514 6060 11520 6112
rect 11572 6100 11578 6112
rect 11609 6103 11667 6109
rect 11609 6100 11621 6103
rect 11572 6072 11621 6100
rect 11572 6060 11578 6072
rect 11609 6069 11621 6072
rect 11655 6069 11667 6103
rect 12773 6100 12801 6128
rect 15194 6100 15200 6112
rect 12773 6072 15200 6100
rect 11609 6063 11667 6069
rect 15194 6060 15200 6072
rect 15252 6100 15258 6112
rect 15396 6100 15424 6140
rect 15702 6137 15714 6140
rect 15748 6168 15760 6171
rect 15838 6168 15844 6180
rect 15748 6140 15844 6168
rect 15748 6137 15760 6140
rect 15702 6131 15760 6137
rect 15838 6128 15844 6140
rect 15896 6128 15902 6180
rect 18138 6168 18144 6180
rect 18099 6140 18144 6168
rect 18138 6128 18144 6140
rect 18196 6128 18202 6180
rect 18233 6171 18291 6177
rect 18233 6137 18245 6171
rect 18279 6137 18291 6171
rect 18233 6131 18291 6137
rect 15252 6072 15424 6100
rect 15252 6060 15258 6072
rect 17770 6060 17776 6112
rect 17828 6100 17834 6112
rect 18248 6100 18276 6131
rect 17828 6072 18276 6100
rect 17828 6060 17834 6072
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 2038 5896 2044 5908
rect 1999 5868 2044 5896
rect 2038 5856 2044 5868
rect 2096 5856 2102 5908
rect 2130 5856 2136 5908
rect 2188 5896 2194 5908
rect 2593 5899 2651 5905
rect 2593 5896 2605 5899
rect 2188 5868 2605 5896
rect 2188 5856 2194 5868
rect 2593 5865 2605 5868
rect 2639 5865 2651 5899
rect 2593 5859 2651 5865
rect 2958 5856 2964 5908
rect 3016 5896 3022 5908
rect 3053 5899 3111 5905
rect 3053 5896 3065 5899
rect 3016 5868 3065 5896
rect 3016 5856 3022 5868
rect 3053 5865 3065 5868
rect 3099 5865 3111 5899
rect 3510 5896 3516 5908
rect 3471 5868 3516 5896
rect 3053 5859 3111 5865
rect 3510 5856 3516 5868
rect 3568 5856 3574 5908
rect 5258 5896 5264 5908
rect 5219 5868 5264 5896
rect 5258 5856 5264 5868
rect 5316 5856 5322 5908
rect 6914 5896 6920 5908
rect 6875 5868 6920 5896
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 8665 5899 8723 5905
rect 8665 5865 8677 5899
rect 8711 5896 8723 5899
rect 8754 5896 8760 5908
rect 8711 5868 8760 5896
rect 8711 5865 8723 5868
rect 8665 5859 8723 5865
rect 8754 5856 8760 5868
rect 8812 5856 8818 5908
rect 9030 5896 9036 5908
rect 8991 5868 9036 5896
rect 9030 5856 9036 5868
rect 9088 5856 9094 5908
rect 9490 5856 9496 5908
rect 9548 5896 9554 5908
rect 9815 5899 9873 5905
rect 9815 5896 9827 5899
rect 9548 5868 9827 5896
rect 9548 5856 9554 5868
rect 9815 5865 9827 5868
rect 9861 5865 9873 5899
rect 9815 5859 9873 5865
rect 10134 5856 10140 5908
rect 10192 5896 10198 5908
rect 10689 5899 10747 5905
rect 10689 5896 10701 5899
rect 10192 5868 10701 5896
rect 10192 5856 10198 5868
rect 10689 5865 10701 5868
rect 10735 5896 10747 5899
rect 15562 5896 15568 5908
rect 10735 5868 11008 5896
rect 15523 5868 15568 5896
rect 10735 5865 10747 5868
rect 10689 5859 10747 5865
rect 2498 5788 2504 5840
rect 2556 5828 2562 5840
rect 3789 5831 3847 5837
rect 3789 5828 3801 5831
rect 2556 5800 3801 5828
rect 2556 5788 2562 5800
rect 3789 5797 3801 5800
rect 3835 5797 3847 5831
rect 3789 5791 3847 5797
rect 4801 5831 4859 5837
rect 4801 5797 4813 5831
rect 4847 5828 4859 5831
rect 5810 5828 5816 5840
rect 4847 5800 5816 5828
rect 4847 5797 4859 5800
rect 4801 5791 4859 5797
rect 5810 5788 5816 5800
rect 5868 5788 5874 5840
rect 5991 5831 6049 5837
rect 5991 5797 6003 5831
rect 6037 5828 6049 5831
rect 6270 5828 6276 5840
rect 6037 5800 6276 5828
rect 6037 5797 6049 5800
rect 5991 5791 6049 5797
rect 6270 5788 6276 5800
rect 6328 5788 6334 5840
rect 10980 5837 11008 5868
rect 15562 5856 15568 5868
rect 15620 5856 15626 5908
rect 16669 5899 16727 5905
rect 16669 5865 16681 5899
rect 16715 5896 16727 5899
rect 17862 5896 17868 5908
rect 16715 5868 17868 5896
rect 16715 5865 16727 5868
rect 16669 5859 16727 5865
rect 17862 5856 17868 5868
rect 17920 5856 17926 5908
rect 10965 5831 11023 5837
rect 10965 5797 10977 5831
rect 11011 5797 11023 5831
rect 10965 5791 11023 5797
rect 11054 5788 11060 5840
rect 11112 5828 11118 5840
rect 11606 5828 11612 5840
rect 11112 5800 11157 5828
rect 11567 5800 11612 5828
rect 11112 5788 11118 5800
rect 11606 5788 11612 5800
rect 11664 5788 11670 5840
rect 12710 5788 12716 5840
rect 12768 5837 12774 5840
rect 12768 5831 12816 5837
rect 12768 5797 12770 5831
rect 12804 5797 12816 5831
rect 12768 5791 12816 5797
rect 12768 5788 12774 5791
rect 15838 5788 15844 5840
rect 15896 5828 15902 5840
rect 16070 5831 16128 5837
rect 16070 5828 16082 5831
rect 15896 5800 16082 5828
rect 15896 5788 15902 5800
rect 16070 5797 16082 5800
rect 16116 5797 16128 5831
rect 16070 5791 16128 5797
rect 17405 5831 17463 5837
rect 17405 5797 17417 5831
rect 17451 5828 17463 5831
rect 17586 5828 17592 5840
rect 17451 5800 17592 5828
rect 17451 5797 17463 5800
rect 17405 5791 17463 5797
rect 17586 5788 17592 5800
rect 17644 5788 17650 5840
rect 17681 5831 17739 5837
rect 17681 5797 17693 5831
rect 17727 5828 17739 5831
rect 17770 5828 17776 5840
rect 17727 5800 17776 5828
rect 17727 5797 17739 5800
rect 17681 5791 17739 5797
rect 17770 5788 17776 5800
rect 17828 5788 17834 5840
rect 19242 5828 19248 5840
rect 19203 5800 19248 5828
rect 19242 5788 19248 5800
rect 19300 5788 19306 5840
rect 1670 5769 1676 5772
rect 1648 5763 1676 5769
rect 1648 5729 1660 5763
rect 1648 5723 1676 5729
rect 1670 5720 1676 5723
rect 1728 5720 1734 5772
rect 4706 5760 4712 5772
rect 4667 5732 4712 5760
rect 4706 5720 4712 5732
rect 4764 5720 4770 5772
rect 5534 5720 5540 5772
rect 5592 5760 5598 5772
rect 5629 5763 5687 5769
rect 5629 5760 5641 5763
rect 5592 5732 5641 5760
rect 5592 5720 5598 5732
rect 5629 5729 5641 5732
rect 5675 5760 5687 5763
rect 7006 5760 7012 5772
rect 5675 5732 7012 5760
rect 5675 5729 5687 5732
rect 5629 5723 5687 5729
rect 7006 5720 7012 5732
rect 7064 5720 7070 5772
rect 7834 5760 7840 5772
rect 7795 5732 7840 5760
rect 7834 5720 7840 5732
rect 7892 5720 7898 5772
rect 9744 5763 9802 5769
rect 9744 5729 9756 5763
rect 9790 5760 9802 5763
rect 9950 5760 9956 5772
rect 9790 5732 9956 5760
rect 9790 5729 9802 5732
rect 9744 5723 9802 5729
rect 9950 5720 9956 5732
rect 10008 5720 10014 5772
rect 10042 5720 10048 5772
rect 10100 5760 10106 5772
rect 10137 5763 10195 5769
rect 10137 5760 10149 5763
rect 10100 5732 10149 5760
rect 10100 5720 10106 5732
rect 10137 5729 10149 5732
rect 10183 5729 10195 5763
rect 10137 5723 10195 5729
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 12492 5732 12537 5760
rect 12492 5720 12498 5732
rect 13906 5720 13912 5772
rect 13964 5760 13970 5772
rect 14220 5763 14278 5769
rect 14220 5760 14232 5763
rect 13964 5732 14232 5760
rect 13964 5720 13970 5732
rect 14220 5729 14232 5732
rect 14266 5729 14278 5763
rect 15746 5760 15752 5772
rect 15707 5732 15752 5760
rect 14220 5723 14278 5729
rect 15746 5720 15752 5732
rect 15804 5720 15810 5772
rect 7098 5652 7104 5704
rect 7156 5692 7162 5704
rect 7377 5695 7435 5701
rect 7377 5692 7389 5695
rect 7156 5664 7389 5692
rect 7156 5652 7162 5664
rect 7377 5661 7389 5664
rect 7423 5661 7435 5695
rect 7377 5655 7435 5661
rect 17589 5695 17647 5701
rect 17589 5661 17601 5695
rect 17635 5661 17647 5695
rect 17589 5655 17647 5661
rect 18233 5695 18291 5701
rect 18233 5661 18245 5695
rect 18279 5692 18291 5695
rect 18598 5692 18604 5704
rect 18279 5664 18604 5692
rect 18279 5661 18291 5664
rect 18233 5655 18291 5661
rect 1394 5584 1400 5636
rect 1452 5624 1458 5636
rect 1719 5627 1777 5633
rect 1719 5624 1731 5627
rect 1452 5596 1731 5624
rect 1452 5584 1458 5596
rect 1719 5593 1731 5596
rect 1765 5624 1777 5627
rect 2409 5627 2467 5633
rect 2409 5624 2421 5627
rect 1765 5596 2421 5624
rect 1765 5593 1777 5596
rect 1719 5587 1777 5593
rect 2409 5593 2421 5596
rect 2455 5593 2467 5627
rect 2409 5587 2467 5593
rect 14323 5627 14381 5633
rect 14323 5593 14335 5627
rect 14369 5624 14381 5627
rect 17604 5624 17632 5655
rect 18598 5652 18604 5664
rect 18656 5652 18662 5704
rect 19153 5695 19211 5701
rect 19153 5661 19165 5695
rect 19199 5692 19211 5695
rect 19334 5692 19340 5704
rect 19199 5664 19340 5692
rect 19199 5661 19211 5664
rect 19153 5655 19211 5661
rect 19334 5652 19340 5664
rect 19392 5652 19398 5704
rect 19426 5652 19432 5704
rect 19484 5692 19490 5704
rect 19484 5664 19529 5692
rect 19484 5652 19490 5664
rect 17678 5624 17684 5636
rect 14369 5596 17684 5624
rect 14369 5593 14381 5596
rect 14323 5587 14381 5593
rect 17678 5584 17684 5596
rect 17736 5584 17742 5636
rect 6546 5556 6552 5568
rect 6507 5528 6552 5556
rect 6546 5516 6552 5528
rect 6604 5516 6610 5568
rect 9030 5516 9036 5568
rect 9088 5556 9094 5568
rect 9401 5559 9459 5565
rect 9401 5556 9413 5559
rect 9088 5528 9413 5556
rect 9088 5516 9094 5528
rect 9401 5525 9413 5528
rect 9447 5556 9459 5559
rect 9858 5556 9864 5568
rect 9447 5528 9864 5556
rect 9447 5525 9459 5528
rect 9401 5519 9459 5525
rect 9858 5516 9864 5528
rect 9916 5516 9922 5568
rect 13357 5559 13415 5565
rect 13357 5525 13369 5559
rect 13403 5556 13415 5559
rect 13814 5556 13820 5568
rect 13403 5528 13820 5556
rect 13403 5525 13415 5528
rect 13357 5519 13415 5525
rect 13814 5516 13820 5528
rect 13872 5516 13878 5568
rect 18506 5556 18512 5568
rect 18467 5528 18512 5556
rect 18506 5516 18512 5528
rect 18564 5516 18570 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 4433 5355 4491 5361
rect 4433 5321 4445 5355
rect 4479 5352 4491 5355
rect 4706 5352 4712 5364
rect 4479 5324 4712 5352
rect 4479 5321 4491 5324
rect 4433 5315 4491 5321
rect 4706 5312 4712 5324
rect 4764 5312 4770 5364
rect 10321 5355 10379 5361
rect 10321 5321 10333 5355
rect 10367 5352 10379 5355
rect 11054 5352 11060 5364
rect 10367 5324 11060 5352
rect 10367 5321 10379 5324
rect 10321 5315 10379 5321
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 11885 5355 11943 5361
rect 11885 5321 11897 5355
rect 11931 5352 11943 5355
rect 12342 5352 12348 5364
rect 11931 5324 12348 5352
rect 11931 5321 11943 5324
rect 11885 5315 11943 5321
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 15473 5355 15531 5361
rect 15473 5321 15485 5355
rect 15519 5352 15531 5355
rect 15746 5352 15752 5364
rect 15519 5324 15752 5352
rect 15519 5321 15531 5324
rect 15473 5315 15531 5321
rect 15746 5312 15752 5324
rect 15804 5312 15810 5364
rect 15838 5312 15844 5364
rect 15896 5352 15902 5364
rect 17589 5355 17647 5361
rect 15896 5324 15941 5352
rect 15896 5312 15902 5324
rect 17589 5321 17601 5355
rect 17635 5352 17647 5355
rect 17770 5352 17776 5364
rect 17635 5324 17776 5352
rect 17635 5321 17647 5324
rect 17589 5315 17647 5321
rect 17770 5312 17776 5324
rect 17828 5312 17834 5364
rect 19153 5355 19211 5361
rect 19153 5321 19165 5355
rect 19199 5352 19211 5355
rect 19242 5352 19248 5364
rect 19199 5324 19248 5352
rect 19199 5321 19211 5324
rect 19153 5315 19211 5321
rect 19242 5312 19248 5324
rect 19300 5312 19306 5364
rect 19334 5312 19340 5364
rect 19392 5352 19398 5364
rect 19429 5355 19487 5361
rect 19429 5352 19441 5355
rect 19392 5324 19441 5352
rect 19392 5312 19398 5324
rect 19429 5321 19441 5324
rect 19475 5321 19487 5355
rect 19429 5315 19487 5321
rect 12253 5287 12311 5293
rect 12253 5253 12265 5287
rect 12299 5284 12311 5287
rect 12710 5284 12716 5296
rect 12299 5256 12716 5284
rect 12299 5253 12311 5256
rect 12253 5247 12311 5253
rect 12710 5244 12716 5256
rect 12768 5244 12774 5296
rect 16758 5244 16764 5296
rect 16816 5284 16822 5296
rect 17037 5287 17095 5293
rect 17037 5284 17049 5287
rect 16816 5256 17049 5284
rect 16816 5244 16822 5256
rect 17037 5253 17049 5256
rect 17083 5284 17095 5287
rect 17083 5256 18644 5284
rect 17083 5253 17095 5256
rect 17037 5247 17095 5253
rect 18616 5228 18644 5256
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5216 2743 5219
rect 3145 5219 3203 5225
rect 3145 5216 3157 5219
rect 2731 5188 3157 5216
rect 2731 5185 2743 5188
rect 2685 5179 2743 5185
rect 3145 5185 3157 5188
rect 3191 5216 3203 5219
rect 4430 5216 4436 5228
rect 3191 5188 4436 5216
rect 3191 5185 3203 5188
rect 3145 5179 3203 5185
rect 4430 5176 4436 5188
rect 4488 5176 4494 5228
rect 6270 5216 6276 5228
rect 5000 5188 6276 5216
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5148 1455 5151
rect 1443 5120 2084 5148
rect 1443 5117 1455 5120
rect 1397 5111 1455 5117
rect 2056 5024 2084 5120
rect 3053 5083 3111 5089
rect 3053 5049 3065 5083
rect 3099 5080 3111 5083
rect 3326 5080 3332 5092
rect 3099 5052 3332 5080
rect 3099 5049 3111 5052
rect 3053 5043 3111 5049
rect 3326 5040 3332 5052
rect 3384 5080 3390 5092
rect 3507 5083 3565 5089
rect 3507 5080 3519 5083
rect 3384 5052 3519 5080
rect 3384 5040 3390 5052
rect 3507 5049 3519 5052
rect 3553 5080 3565 5083
rect 5000 5080 5028 5188
rect 6270 5176 6276 5188
rect 6328 5216 6334 5228
rect 6825 5219 6883 5225
rect 6328 5188 6684 5216
rect 6328 5176 6334 5188
rect 5077 5151 5135 5157
rect 5077 5117 5089 5151
rect 5123 5148 5135 5151
rect 5813 5151 5871 5157
rect 5813 5148 5825 5151
rect 5123 5120 5825 5148
rect 5123 5117 5135 5120
rect 5077 5111 5135 5117
rect 5813 5117 5825 5120
rect 5859 5148 5871 5151
rect 6546 5148 6552 5160
rect 5859 5120 6552 5148
rect 5859 5117 5871 5120
rect 5813 5111 5871 5117
rect 6546 5108 6552 5120
rect 6604 5108 6610 5160
rect 6656 5157 6684 5188
rect 6825 5185 6837 5219
rect 6871 5216 6883 5219
rect 6914 5216 6920 5228
rect 6871 5188 6920 5216
rect 6871 5185 6883 5188
rect 6825 5179 6883 5185
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 9309 5219 9367 5225
rect 9309 5185 9321 5219
rect 9355 5216 9367 5219
rect 9674 5216 9680 5228
rect 9355 5188 9680 5216
rect 9355 5185 9367 5188
rect 9309 5179 9367 5185
rect 9674 5176 9680 5188
rect 9732 5176 9738 5228
rect 11514 5216 11520 5228
rect 11475 5188 11520 5216
rect 11514 5176 11520 5188
rect 11572 5176 11578 5228
rect 13078 5216 13084 5228
rect 13039 5188 13084 5216
rect 13078 5176 13084 5188
rect 13136 5216 13142 5228
rect 14185 5219 14243 5225
rect 14185 5216 14197 5219
rect 13136 5188 14197 5216
rect 13136 5176 13142 5188
rect 14185 5185 14197 5188
rect 14231 5185 14243 5219
rect 14185 5179 14243 5185
rect 14366 5176 14372 5228
rect 14424 5216 14430 5228
rect 14461 5219 14519 5225
rect 14461 5216 14473 5219
rect 14424 5188 14473 5216
rect 14424 5176 14430 5188
rect 14461 5185 14473 5188
rect 14507 5185 14519 5219
rect 14461 5179 14519 5185
rect 15286 5176 15292 5228
rect 15344 5216 15350 5228
rect 16482 5216 16488 5228
rect 15344 5188 16488 5216
rect 15344 5176 15350 5188
rect 16482 5176 16488 5188
rect 16540 5176 16546 5228
rect 18141 5219 18199 5225
rect 18141 5185 18153 5219
rect 18187 5216 18199 5219
rect 18506 5216 18512 5228
rect 18187 5188 18512 5216
rect 18187 5185 18199 5188
rect 18141 5179 18199 5185
rect 18506 5176 18512 5188
rect 18564 5176 18570 5228
rect 18598 5176 18604 5228
rect 18656 5216 18662 5228
rect 18656 5188 18701 5216
rect 18656 5176 18662 5188
rect 6641 5151 6699 5157
rect 6641 5117 6653 5151
rect 6687 5148 6699 5151
rect 8481 5151 8539 5157
rect 6687 5120 7189 5148
rect 6687 5117 6699 5120
rect 6641 5111 6699 5117
rect 3553 5052 5028 5080
rect 5905 5083 5963 5089
rect 3553 5049 3565 5052
rect 3507 5043 3565 5049
rect 5905 5049 5917 5083
rect 5951 5080 5963 5083
rect 6086 5080 6092 5092
rect 5951 5052 6092 5080
rect 5951 5049 5963 5052
rect 5905 5043 5963 5049
rect 6086 5040 6092 5052
rect 6144 5040 6150 5092
rect 7161 5089 7189 5120
rect 8481 5117 8493 5151
rect 8527 5148 8539 5151
rect 8662 5148 8668 5160
rect 8527 5120 8668 5148
rect 8527 5117 8539 5120
rect 8481 5111 8539 5117
rect 8662 5108 8668 5120
rect 8720 5108 8726 5160
rect 10689 5151 10747 5157
rect 10689 5117 10701 5151
rect 10735 5148 10747 5151
rect 10962 5148 10968 5160
rect 10735 5120 10968 5148
rect 10735 5117 10747 5120
rect 10689 5111 10747 5117
rect 10962 5108 10968 5120
rect 11020 5108 11026 5160
rect 11333 5151 11391 5157
rect 11333 5117 11345 5151
rect 11379 5148 11391 5151
rect 11422 5148 11428 5160
rect 11379 5120 11428 5148
rect 11379 5117 11391 5120
rect 11333 5111 11391 5117
rect 11422 5108 11428 5120
rect 11480 5108 11486 5160
rect 7161 5083 7245 5089
rect 7161 5052 7199 5083
rect 7187 5049 7199 5052
rect 7233 5080 7245 5083
rect 8110 5080 8116 5092
rect 7233 5052 8116 5080
rect 7233 5049 7245 5052
rect 7187 5043 7245 5049
rect 8110 5040 8116 5052
rect 8168 5040 8174 5092
rect 12621 5083 12679 5089
rect 12621 5049 12633 5083
rect 12667 5049 12679 5083
rect 12621 5043 12679 5049
rect 1578 5012 1584 5024
rect 1539 4984 1584 5012
rect 1578 4972 1584 4984
rect 1636 4972 1642 5024
rect 2038 5012 2044 5024
rect 1999 4984 2044 5012
rect 2038 4972 2044 4984
rect 2096 4972 2102 5024
rect 4065 5015 4123 5021
rect 4065 4981 4077 5015
rect 4111 5012 4123 5015
rect 4246 5012 4252 5024
rect 4111 4984 4252 5012
rect 4111 4981 4123 4984
rect 4065 4975 4123 4981
rect 4246 4972 4252 4984
rect 4304 4972 4310 5024
rect 7745 5015 7803 5021
rect 7745 4981 7757 5015
rect 7791 5012 7803 5015
rect 7834 5012 7840 5024
rect 7791 4984 7840 5012
rect 7791 4981 7803 4984
rect 7745 4975 7803 4981
rect 7834 4972 7840 4984
rect 7892 5012 7898 5024
rect 8021 5015 8079 5021
rect 8021 5012 8033 5015
rect 7892 4984 8033 5012
rect 7892 4972 7898 4984
rect 8021 4981 8033 4984
rect 8067 4981 8079 5015
rect 8021 4975 8079 4981
rect 9769 5015 9827 5021
rect 9769 4981 9781 5015
rect 9815 5012 9827 5015
rect 9858 5012 9864 5024
rect 9815 4984 9864 5012
rect 9815 4981 9827 4984
rect 9769 4975 9827 4981
rect 9858 4972 9864 4984
rect 9916 4972 9922 5024
rect 12636 5012 12664 5043
rect 12710 5040 12716 5092
rect 12768 5080 12774 5092
rect 12768 5052 12813 5080
rect 12768 5040 12774 5052
rect 13814 5040 13820 5092
rect 13872 5080 13878 5092
rect 14277 5083 14335 5089
rect 13872 5052 14136 5080
rect 13872 5040 13878 5052
rect 13630 5012 13636 5024
rect 12636 4984 13636 5012
rect 13630 4972 13636 4984
rect 13688 4972 13694 5024
rect 13906 5012 13912 5024
rect 13867 4984 13912 5012
rect 13906 4972 13912 4984
rect 13964 4972 13970 5024
rect 14108 5012 14136 5052
rect 14277 5049 14289 5083
rect 14323 5049 14335 5083
rect 14277 5043 14335 5049
rect 16301 5083 16359 5089
rect 16301 5049 16313 5083
rect 16347 5080 16359 5083
rect 16577 5083 16635 5089
rect 16577 5080 16589 5083
rect 16347 5052 16589 5080
rect 16347 5049 16359 5052
rect 16301 5043 16359 5049
rect 16577 5049 16589 5052
rect 16623 5049 16635 5083
rect 16577 5043 16635 5049
rect 14292 5012 14320 5043
rect 14108 4984 14320 5012
rect 16592 5012 16620 5043
rect 17954 5040 17960 5092
rect 18012 5080 18018 5092
rect 18233 5083 18291 5089
rect 18233 5080 18245 5083
rect 18012 5052 18245 5080
rect 18012 5040 18018 5052
rect 18233 5049 18245 5052
rect 18279 5049 18291 5083
rect 18233 5043 18291 5049
rect 19242 5012 19248 5024
rect 16592 4984 19248 5012
rect 19242 4972 19248 4984
rect 19300 4972 19306 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 2225 4811 2283 4817
rect 2225 4808 2237 4811
rect 1728 4780 2237 4808
rect 1728 4768 1734 4780
rect 2225 4777 2237 4780
rect 2271 4777 2283 4811
rect 2225 4771 2283 4777
rect 5534 4768 5540 4820
rect 5592 4808 5598 4820
rect 5629 4811 5687 4817
rect 5629 4808 5641 4811
rect 5592 4780 5641 4808
rect 5592 4768 5598 4780
rect 5629 4777 5641 4780
rect 5675 4777 5687 4811
rect 5629 4771 5687 4777
rect 10873 4811 10931 4817
rect 10873 4777 10885 4811
rect 10919 4808 10931 4811
rect 11422 4808 11428 4820
rect 10919 4780 11428 4808
rect 10919 4777 10931 4780
rect 10873 4771 10931 4777
rect 11422 4768 11428 4780
rect 11480 4768 11486 4820
rect 12621 4811 12679 4817
rect 12621 4777 12633 4811
rect 12667 4808 12679 4811
rect 12710 4808 12716 4820
rect 12667 4780 12716 4808
rect 12667 4777 12679 4780
rect 12621 4771 12679 4777
rect 12710 4768 12716 4780
rect 12768 4768 12774 4820
rect 13814 4768 13820 4820
rect 13872 4808 13878 4820
rect 14093 4811 14151 4817
rect 14093 4808 14105 4811
rect 13872 4780 14105 4808
rect 13872 4768 13878 4780
rect 14093 4777 14105 4780
rect 14139 4777 14151 4811
rect 16482 4808 16488 4820
rect 16443 4780 16488 4808
rect 14093 4771 14151 4777
rect 16482 4768 16488 4780
rect 16540 4768 16546 4820
rect 17678 4808 17684 4820
rect 17639 4780 17684 4808
rect 17678 4768 17684 4780
rect 17736 4768 17742 4820
rect 17954 4768 17960 4820
rect 18012 4808 18018 4820
rect 18049 4811 18107 4817
rect 18049 4808 18061 4811
rect 18012 4780 18061 4808
rect 18012 4768 18018 4780
rect 18049 4777 18061 4780
rect 18095 4777 18107 4811
rect 18049 4771 18107 4777
rect 18371 4811 18429 4817
rect 18371 4777 18383 4811
rect 18417 4808 18429 4811
rect 18506 4808 18512 4820
rect 18417 4780 18512 4808
rect 18417 4777 18429 4780
rect 18371 4771 18429 4777
rect 18506 4768 18512 4780
rect 18564 4768 18570 4820
rect 19334 4768 19340 4820
rect 19392 4817 19398 4820
rect 19392 4811 19441 4817
rect 19392 4777 19395 4811
rect 19429 4777 19441 4811
rect 19392 4771 19441 4777
rect 19392 4768 19398 4771
rect 20714 4768 20720 4820
rect 20772 4808 20778 4820
rect 21407 4811 21465 4817
rect 21407 4808 21419 4811
rect 20772 4780 21419 4808
rect 20772 4768 20778 4780
rect 21407 4777 21419 4780
rect 21453 4777 21465 4811
rect 21407 4771 21465 4777
rect 6086 4740 6092 4752
rect 6047 4712 6092 4740
rect 6086 4700 6092 4712
rect 6144 4700 6150 4752
rect 7653 4743 7711 4749
rect 7653 4709 7665 4743
rect 7699 4740 7711 4743
rect 7834 4740 7840 4752
rect 7699 4712 7840 4740
rect 7699 4709 7711 4712
rect 7653 4703 7711 4709
rect 7834 4700 7840 4712
rect 7892 4700 7898 4752
rect 11330 4740 11336 4752
rect 11291 4712 11336 4740
rect 11330 4700 11336 4712
rect 11388 4700 11394 4752
rect 12897 4743 12955 4749
rect 12897 4740 12909 4743
rect 12636 4712 12909 4740
rect 12636 4684 12664 4712
rect 12897 4709 12909 4712
rect 12943 4709 12955 4743
rect 12897 4703 12955 4709
rect 16574 4700 16580 4752
rect 16632 4740 16638 4752
rect 16853 4743 16911 4749
rect 16853 4740 16865 4743
rect 16632 4712 16865 4740
rect 16632 4700 16638 4712
rect 16853 4709 16865 4712
rect 16899 4709 16911 4743
rect 17402 4740 17408 4752
rect 17363 4712 17408 4740
rect 16853 4703 16911 4709
rect 17402 4700 17408 4712
rect 17460 4700 17466 4752
rect 1486 4681 1492 4684
rect 1464 4675 1492 4681
rect 1464 4672 1476 4675
rect 1399 4644 1476 4672
rect 1464 4641 1476 4644
rect 1544 4672 1550 4684
rect 2038 4672 2044 4684
rect 1544 4644 2044 4672
rect 1464 4635 1492 4641
rect 1486 4632 1492 4635
rect 1544 4632 1550 4644
rect 2038 4632 2044 4644
rect 2096 4632 2102 4684
rect 2498 4632 2504 4684
rect 2556 4672 2562 4684
rect 3053 4675 3111 4681
rect 3053 4672 3065 4675
rect 2556 4644 3065 4672
rect 2556 4632 2562 4644
rect 3053 4641 3065 4644
rect 3099 4672 3111 4675
rect 4246 4672 4252 4684
rect 3099 4644 4252 4672
rect 3099 4641 3111 4644
rect 3053 4635 3111 4641
rect 4246 4632 4252 4644
rect 4304 4632 4310 4684
rect 10045 4675 10103 4681
rect 10045 4641 10057 4675
rect 10091 4672 10103 4675
rect 10778 4672 10784 4684
rect 10091 4644 10784 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 12618 4632 12624 4684
rect 12676 4632 12682 4684
rect 14366 4632 14372 4684
rect 14424 4672 14430 4684
rect 15324 4675 15382 4681
rect 15324 4672 15336 4675
rect 14424 4644 15336 4672
rect 14424 4632 14430 4644
rect 15324 4641 15336 4644
rect 15370 4672 15382 4675
rect 15654 4672 15660 4684
rect 15370 4644 15660 4672
rect 15370 4641 15382 4644
rect 15324 4635 15382 4641
rect 15654 4632 15660 4644
rect 15712 4632 15718 4684
rect 18300 4675 18358 4681
rect 18300 4641 18312 4675
rect 18346 4672 18358 4675
rect 18414 4672 18420 4684
rect 18346 4644 18420 4672
rect 18346 4641 18358 4644
rect 18300 4635 18358 4641
rect 18414 4632 18420 4644
rect 18472 4632 18478 4684
rect 19334 4681 19340 4684
rect 19312 4675 19340 4681
rect 19312 4641 19324 4675
rect 19312 4635 19340 4641
rect 19334 4632 19340 4635
rect 19392 4632 19398 4684
rect 21358 4681 21364 4684
rect 21336 4675 21364 4681
rect 21336 4641 21348 4675
rect 21336 4635 21364 4641
rect 21358 4632 21364 4635
rect 21416 4632 21422 4684
rect 4893 4607 4951 4613
rect 4893 4573 4905 4607
rect 4939 4604 4951 4607
rect 5997 4607 6055 4613
rect 5997 4604 6009 4607
rect 4939 4576 6009 4604
rect 4939 4573 4951 4576
rect 4893 4567 4951 4573
rect 5997 4573 6009 4576
rect 6043 4604 6055 4607
rect 6270 4604 6276 4616
rect 6043 4576 6276 4604
rect 6043 4573 6055 4576
rect 5997 4567 6055 4573
rect 6270 4564 6276 4576
rect 6328 4564 6334 4616
rect 6641 4607 6699 4613
rect 6641 4573 6653 4607
rect 6687 4604 6699 4607
rect 6914 4604 6920 4616
rect 6687 4576 6920 4604
rect 6687 4573 6699 4576
rect 6641 4567 6699 4573
rect 6914 4564 6920 4576
rect 6972 4564 6978 4616
rect 7561 4607 7619 4613
rect 7561 4573 7573 4607
rect 7607 4604 7619 4607
rect 7650 4604 7656 4616
rect 7607 4576 7656 4604
rect 7607 4573 7619 4576
rect 7561 4567 7619 4573
rect 7650 4564 7656 4576
rect 7708 4564 7714 4616
rect 7837 4607 7895 4613
rect 7837 4573 7849 4607
rect 7883 4573 7895 4607
rect 7837 4567 7895 4573
rect 1535 4539 1593 4545
rect 1535 4505 1547 4539
rect 1581 4536 1593 4539
rect 4617 4539 4675 4545
rect 4617 4536 4629 4539
rect 1581 4508 4629 4536
rect 1581 4505 1593 4508
rect 1535 4499 1593 4505
rect 4617 4505 4629 4508
rect 4663 4536 4675 4539
rect 4706 4536 4712 4548
rect 4663 4508 4712 4536
rect 4663 4505 4675 4508
rect 4617 4499 4675 4505
rect 4706 4496 4712 4508
rect 4764 4496 4770 4548
rect 7374 4536 7380 4548
rect 7287 4508 7380 4536
rect 7374 4496 7380 4508
rect 7432 4536 7438 4548
rect 7852 4536 7880 4567
rect 10962 4564 10968 4616
rect 11020 4604 11026 4616
rect 11241 4607 11299 4613
rect 11241 4604 11253 4607
rect 11020 4576 11253 4604
rect 11020 4564 11026 4576
rect 11241 4573 11253 4576
rect 11287 4573 11299 4607
rect 11606 4604 11612 4616
rect 11567 4576 11612 4604
rect 11241 4567 11299 4573
rect 11606 4564 11612 4576
rect 11664 4604 11670 4616
rect 12434 4604 12440 4616
rect 11664 4576 12440 4604
rect 11664 4564 11670 4576
rect 12434 4564 12440 4576
rect 12492 4564 12498 4616
rect 12805 4607 12863 4613
rect 12805 4573 12817 4607
rect 12851 4573 12863 4607
rect 13078 4604 13084 4616
rect 13039 4576 13084 4604
rect 12805 4567 12863 4573
rect 7432 4508 7880 4536
rect 7432 4496 7438 4508
rect 12342 4496 12348 4548
rect 12400 4536 12406 4548
rect 12820 4536 12848 4567
rect 13078 4564 13084 4576
rect 13136 4604 13142 4616
rect 14461 4607 14519 4613
rect 14461 4604 14473 4607
rect 13136 4576 14473 4604
rect 13136 4564 13142 4576
rect 14461 4573 14473 4576
rect 14507 4573 14519 4607
rect 16758 4604 16764 4616
rect 16719 4576 16764 4604
rect 14461 4567 14519 4573
rect 16758 4564 16764 4576
rect 16816 4564 16822 4616
rect 13814 4536 13820 4548
rect 12400 4508 13820 4536
rect 12400 4496 12406 4508
rect 13814 4496 13820 4508
rect 13872 4496 13878 4548
rect 15427 4539 15485 4545
rect 15427 4505 15439 4539
rect 15473 4536 15485 4539
rect 16482 4536 16488 4548
rect 15473 4508 16488 4536
rect 15473 4505 15485 4508
rect 15427 4499 15485 4505
rect 16482 4496 16488 4508
rect 16540 4496 16546 4548
rect 1946 4468 1952 4480
rect 1907 4440 1952 4468
rect 1946 4428 1952 4440
rect 2004 4428 2010 4480
rect 2866 4468 2872 4480
rect 2827 4440 2872 4468
rect 2866 4428 2872 4440
rect 2924 4428 2930 4480
rect 6546 4428 6552 4480
rect 6604 4468 6610 4480
rect 7006 4468 7012 4480
rect 6604 4440 7012 4468
rect 6604 4428 6610 4440
rect 7006 4428 7012 4440
rect 7064 4428 7070 4480
rect 10229 4471 10287 4477
rect 10229 4437 10241 4471
rect 10275 4468 10287 4471
rect 10870 4468 10876 4480
rect 10275 4440 10876 4468
rect 10275 4437 10287 4440
rect 10229 4431 10287 4437
rect 10870 4428 10876 4440
rect 10928 4428 10934 4480
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 14458 4468 14464 4480
rect 11112 4440 14464 4468
rect 11112 4428 11118 4440
rect 14458 4428 14464 4440
rect 14516 4428 14522 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 2498 4264 2504 4276
rect 2459 4236 2504 4264
rect 2498 4224 2504 4236
rect 2556 4224 2562 4276
rect 2866 4264 2872 4276
rect 2827 4236 2872 4264
rect 2866 4224 2872 4236
rect 2924 4224 2930 4276
rect 5997 4267 6055 4273
rect 5997 4233 6009 4267
rect 6043 4264 6055 4267
rect 6086 4264 6092 4276
rect 6043 4236 6092 4264
rect 6043 4233 6055 4236
rect 5997 4227 6055 4233
rect 6086 4224 6092 4236
rect 6144 4224 6150 4276
rect 6270 4264 6276 4276
rect 6231 4236 6276 4264
rect 6270 4224 6276 4236
rect 6328 4224 6334 4276
rect 7834 4264 7840 4276
rect 7795 4236 7840 4264
rect 7834 4224 7840 4236
rect 7892 4224 7898 4276
rect 10137 4267 10195 4273
rect 10137 4233 10149 4267
rect 10183 4264 10195 4267
rect 11054 4264 11060 4276
rect 10183 4236 11060 4264
rect 10183 4233 10195 4236
rect 10137 4227 10195 4233
rect 2038 4196 2044 4208
rect 1951 4168 2044 4196
rect 2038 4156 2044 4168
rect 2096 4196 2102 4208
rect 8478 4196 8484 4208
rect 2096 4168 8484 4196
rect 2096 4156 2102 4168
rect 8478 4156 8484 4168
rect 8536 4156 8542 4208
rect 10152 4196 10180 4227
rect 11054 4224 11060 4236
rect 11112 4224 11118 4276
rect 11241 4267 11299 4273
rect 11241 4233 11253 4267
rect 11287 4264 11299 4267
rect 11330 4264 11336 4276
rect 11287 4236 11336 4264
rect 11287 4233 11299 4236
rect 11241 4227 11299 4233
rect 11330 4224 11336 4236
rect 11388 4264 11394 4276
rect 12069 4267 12127 4273
rect 12069 4264 12081 4267
rect 11388 4236 12081 4264
rect 11388 4224 11394 4236
rect 12069 4233 12081 4236
rect 12115 4264 12127 4267
rect 12161 4267 12219 4273
rect 12161 4264 12173 4267
rect 12115 4236 12173 4264
rect 12115 4233 12127 4236
rect 12069 4227 12127 4233
rect 12161 4233 12173 4236
rect 12207 4233 12219 4267
rect 13814 4264 13820 4276
rect 13775 4236 13820 4264
rect 12161 4227 12219 4233
rect 13814 4224 13820 4236
rect 13872 4224 13878 4276
rect 14553 4267 14611 4273
rect 14553 4233 14565 4267
rect 14599 4264 14611 4267
rect 14642 4264 14648 4276
rect 14599 4236 14648 4264
rect 14599 4233 14611 4236
rect 14553 4227 14611 4233
rect 14642 4224 14648 4236
rect 14700 4224 14706 4276
rect 15654 4264 15660 4276
rect 15615 4236 15660 4264
rect 15654 4224 15660 4236
rect 15712 4224 15718 4276
rect 16574 4224 16580 4276
rect 16632 4264 16638 4276
rect 16761 4267 16819 4273
rect 16761 4264 16773 4267
rect 16632 4236 16773 4264
rect 16632 4224 16638 4236
rect 16761 4233 16773 4236
rect 16807 4233 16819 4267
rect 16761 4227 16819 4233
rect 9651 4168 10180 4196
rect 11471 4199 11529 4205
rect 3878 4088 3884 4140
rect 3936 4128 3942 4140
rect 4430 4128 4436 4140
rect 3936 4100 4436 4128
rect 3936 4088 3942 4100
rect 4430 4088 4436 4100
rect 4488 4088 4494 4140
rect 4706 4128 4712 4140
rect 4667 4100 4712 4128
rect 4706 4088 4712 4100
rect 4764 4088 4770 4140
rect 4982 4128 4988 4140
rect 4943 4100 4988 4128
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 6917 4131 6975 4137
rect 6917 4097 6929 4131
rect 6963 4128 6975 4131
rect 7374 4128 7380 4140
rect 6963 4100 7380 4128
rect 6963 4097 6975 4100
rect 6917 4091 6975 4097
rect 7374 4088 7380 4100
rect 7432 4088 7438 4140
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4060 1455 4063
rect 1946 4060 1952 4072
rect 1443 4032 1952 4060
rect 1443 4029 1455 4032
rect 1397 4023 1455 4029
rect 1946 4020 1952 4032
rect 2004 4020 2010 4072
rect 9651 4069 9679 4168
rect 11471 4165 11483 4199
rect 11517 4196 11529 4199
rect 12342 4196 12348 4208
rect 11517 4168 12348 4196
rect 11517 4165 11529 4168
rect 11471 4159 11529 4165
rect 12342 4156 12348 4168
rect 12400 4156 12406 4208
rect 13078 4196 13084 4208
rect 13039 4168 13084 4196
rect 13078 4156 13084 4168
rect 13136 4156 13142 4208
rect 14660 4196 14688 4224
rect 17402 4196 17408 4208
rect 14660 4168 14780 4196
rect 9766 4137 9772 4140
rect 9723 4131 9772 4137
rect 9723 4097 9735 4131
rect 9769 4097 9772 4131
rect 9723 4091 9772 4097
rect 9766 4088 9772 4091
rect 9824 4088 9830 4140
rect 10873 4131 10931 4137
rect 10873 4097 10885 4131
rect 10919 4128 10931 4131
rect 10962 4128 10968 4140
rect 10919 4100 10968 4128
rect 10919 4097 10931 4100
rect 10873 4091 10931 4097
rect 10962 4088 10968 4100
rect 11020 4088 11026 4140
rect 12618 4088 12624 4140
rect 12676 4128 12682 4140
rect 13449 4131 13507 4137
rect 13449 4128 13461 4131
rect 12676 4100 13461 4128
rect 12676 4088 12682 4100
rect 13449 4097 13461 4100
rect 13495 4097 13507 4131
rect 13449 4091 13507 4097
rect 8640 4063 8698 4069
rect 8640 4029 8652 4063
rect 8686 4060 8698 4063
rect 9631 4063 9689 4069
rect 8686 4032 9168 4060
rect 8686 4029 8698 4032
rect 8640 4023 8698 4029
rect 3142 3992 3148 4004
rect 3103 3964 3148 3992
rect 3142 3952 3148 3964
rect 3200 3952 3206 4004
rect 3237 3995 3295 4001
rect 3237 3961 3249 3995
rect 3283 3961 3295 3995
rect 3237 3955 3295 3961
rect 3789 3995 3847 4001
rect 3789 3961 3801 3995
rect 3835 3992 3847 3995
rect 4522 3992 4528 4004
rect 3835 3964 4528 3992
rect 3835 3961 3847 3964
rect 3789 3955 3847 3961
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 2866 3884 2872 3936
rect 2924 3924 2930 3936
rect 3252 3924 3280 3955
rect 4522 3952 4528 3964
rect 4580 3952 4586 4004
rect 4801 3995 4859 4001
rect 4801 3961 4813 3995
rect 4847 3961 4859 3995
rect 7006 3992 7012 4004
rect 6967 3964 7012 3992
rect 4801 3955 4859 3961
rect 2924 3896 3280 3924
rect 2924 3884 2930 3896
rect 4430 3884 4436 3936
rect 4488 3924 4494 3936
rect 4816 3924 4844 3955
rect 7006 3952 7012 3964
rect 7064 3952 7070 4004
rect 7561 3995 7619 4001
rect 7561 3961 7573 3995
rect 7607 3961 7619 3995
rect 7561 3955 7619 3961
rect 4488 3896 4844 3924
rect 4488 3884 4494 3896
rect 6914 3884 6920 3936
rect 6972 3924 6978 3936
rect 7190 3924 7196 3936
rect 6972 3896 7196 3924
rect 6972 3884 6978 3896
rect 7190 3884 7196 3896
rect 7248 3924 7254 3936
rect 7576 3924 7604 3955
rect 7248 3896 7604 3924
rect 7248 3884 7254 3896
rect 7650 3884 7656 3936
rect 7708 3924 7714 3936
rect 8202 3924 8208 3936
rect 7708 3896 8208 3924
rect 7708 3884 7714 3896
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 8711 3927 8769 3933
rect 8711 3893 8723 3927
rect 8757 3924 8769 3927
rect 9030 3924 9036 3936
rect 8757 3896 9036 3924
rect 8757 3893 8769 3896
rect 8711 3887 8769 3893
rect 9030 3884 9036 3896
rect 9088 3884 9094 3936
rect 9140 3933 9168 4032
rect 9631 4029 9643 4063
rect 9677 4029 9689 4063
rect 9631 4023 9689 4029
rect 9651 3936 9679 4023
rect 11330 4020 11336 4072
rect 11388 4069 11394 4072
rect 11388 4063 11426 4069
rect 11414 4060 11426 4063
rect 11793 4063 11851 4069
rect 11793 4060 11805 4063
rect 11414 4032 11805 4060
rect 11414 4029 11426 4032
rect 11388 4023 11426 4029
rect 11793 4029 11805 4032
rect 11839 4060 11851 4063
rect 11974 4060 11980 4072
rect 11839 4032 11980 4060
rect 11839 4029 11851 4032
rect 11793 4023 11851 4029
rect 11388 4020 11394 4023
rect 11974 4020 11980 4032
rect 12032 4020 12038 4072
rect 14752 4069 14780 4168
rect 16592 4168 17408 4196
rect 16209 4131 16267 4137
rect 16209 4097 16221 4131
rect 16255 4128 16267 4131
rect 16592 4128 16620 4168
rect 17402 4156 17408 4168
rect 17460 4156 17466 4208
rect 16255 4100 16620 4128
rect 16255 4097 16267 4100
rect 16209 4091 16267 4097
rect 14737 4063 14795 4069
rect 14737 4029 14749 4063
rect 14783 4029 14795 4063
rect 15102 4060 15108 4072
rect 15063 4032 15108 4060
rect 14737 4023 14795 4029
rect 15102 4020 15108 4032
rect 15160 4020 15166 4072
rect 16408 4069 16436 4100
rect 16758 4088 16764 4140
rect 16816 4128 16822 4140
rect 17129 4131 17187 4137
rect 17129 4128 17141 4131
rect 16816 4100 17141 4128
rect 16816 4088 16822 4100
rect 17129 4097 17141 4100
rect 17175 4097 17187 4131
rect 17129 4091 17187 4097
rect 16368 4063 16436 4069
rect 16368 4029 16380 4063
rect 16414 4032 16436 4063
rect 16414 4029 16426 4032
rect 16368 4023 16426 4029
rect 12526 3992 12532 4004
rect 12487 3964 12532 3992
rect 12526 3952 12532 3964
rect 12584 3952 12590 4004
rect 12621 3995 12679 4001
rect 12621 3961 12633 3995
rect 12667 3961 12679 3995
rect 12621 3955 12679 3961
rect 9125 3927 9183 3933
rect 9125 3893 9137 3927
rect 9171 3924 9183 3927
rect 9398 3924 9404 3936
rect 9171 3896 9404 3924
rect 9171 3893 9183 3896
rect 9125 3887 9183 3893
rect 9398 3884 9404 3896
rect 9456 3884 9462 3936
rect 9651 3896 9680 3936
rect 9674 3884 9680 3896
rect 9732 3884 9738 3936
rect 10505 3927 10563 3933
rect 10505 3893 10517 3927
rect 10551 3924 10563 3927
rect 10778 3924 10784 3936
rect 10551 3896 10784 3924
rect 10551 3893 10563 3896
rect 10505 3887 10563 3893
rect 10778 3884 10784 3896
rect 10836 3884 10842 3936
rect 12069 3927 12127 3933
rect 12069 3893 12081 3927
rect 12115 3924 12127 3927
rect 12636 3924 12664 3955
rect 12115 3896 12664 3924
rect 12115 3893 12127 3896
rect 12069 3887 12127 3893
rect 14826 3884 14832 3936
rect 14884 3924 14890 3936
rect 14921 3927 14979 3933
rect 14921 3924 14933 3927
rect 14884 3896 14933 3924
rect 14884 3884 14890 3896
rect 14921 3893 14933 3896
rect 14967 3893 14979 3927
rect 14921 3887 14979 3893
rect 16206 3884 16212 3936
rect 16264 3924 16270 3936
rect 16439 3927 16497 3933
rect 16439 3924 16451 3927
rect 16264 3896 16451 3924
rect 16264 3884 16270 3896
rect 16439 3893 16451 3896
rect 16485 3893 16497 3927
rect 16439 3887 16497 3893
rect 18325 3927 18383 3933
rect 18325 3893 18337 3927
rect 18371 3924 18383 3927
rect 18414 3924 18420 3936
rect 18371 3896 18420 3924
rect 18371 3893 18383 3896
rect 18325 3887 18383 3893
rect 18414 3884 18420 3896
rect 18472 3924 18478 3936
rect 18874 3924 18880 3936
rect 18472 3896 18880 3924
rect 18472 3884 18478 3896
rect 18874 3884 18880 3896
rect 18932 3884 18938 3936
rect 19334 3924 19340 3936
rect 19295 3896 19340 3924
rect 19334 3884 19340 3896
rect 19392 3884 19398 3936
rect 21358 3924 21364 3936
rect 21319 3896 21364 3924
rect 21358 3884 21364 3896
rect 21416 3884 21422 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1394 3680 1400 3732
rect 1452 3720 1458 3732
rect 1673 3723 1731 3729
rect 1673 3720 1685 3723
rect 1452 3692 1685 3720
rect 1452 3680 1458 3692
rect 1673 3689 1685 3692
rect 1719 3720 1731 3723
rect 2222 3720 2228 3732
rect 1719 3692 2228 3720
rect 1719 3689 1731 3692
rect 1673 3683 1731 3689
rect 2222 3680 2228 3692
rect 2280 3680 2286 3732
rect 3878 3720 3884 3732
rect 2516 3692 3884 3720
rect 2516 3661 2544 3692
rect 3878 3680 3884 3692
rect 3936 3680 3942 3732
rect 5534 3680 5540 3732
rect 5592 3720 5598 3732
rect 5767 3723 5825 3729
rect 5767 3720 5779 3723
rect 5592 3692 5779 3720
rect 5592 3680 5598 3692
rect 5767 3689 5779 3692
rect 5813 3689 5825 3723
rect 5767 3683 5825 3689
rect 8711 3723 8769 3729
rect 8711 3689 8723 3723
rect 8757 3720 8769 3723
rect 9122 3720 9128 3732
rect 8757 3692 9128 3720
rect 8757 3689 8769 3692
rect 8711 3683 8769 3689
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 10091 3723 10149 3729
rect 10091 3689 10103 3723
rect 10137 3720 10149 3723
rect 10962 3720 10968 3732
rect 10137 3692 10968 3720
rect 10137 3689 10149 3692
rect 10091 3683 10149 3689
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 11563 3723 11621 3729
rect 11563 3689 11575 3723
rect 11609 3720 11621 3723
rect 12526 3720 12532 3732
rect 11609 3692 12532 3720
rect 11609 3689 11621 3692
rect 11563 3683 11621 3689
rect 12526 3680 12532 3692
rect 12584 3680 12590 3732
rect 14734 3720 14740 3732
rect 14647 3692 14740 3720
rect 14734 3680 14740 3692
rect 14792 3720 14798 3732
rect 15102 3720 15108 3732
rect 14792 3692 15108 3720
rect 14792 3680 14798 3692
rect 15102 3680 15108 3692
rect 15160 3680 15166 3732
rect 15286 3680 15292 3732
rect 15344 3720 15350 3732
rect 15427 3723 15485 3729
rect 15427 3720 15439 3723
rect 15344 3692 15439 3720
rect 15344 3680 15350 3692
rect 15427 3689 15439 3692
rect 15473 3689 15485 3723
rect 15427 3683 15485 3689
rect 2494 3655 2552 3661
rect 2494 3621 2506 3655
rect 2540 3621 2552 3655
rect 2494 3615 2552 3621
rect 3053 3655 3111 3661
rect 3053 3621 3065 3655
rect 3099 3652 3111 3655
rect 3142 3652 3148 3664
rect 3099 3624 3148 3652
rect 3099 3621 3111 3624
rect 3053 3615 3111 3621
rect 3142 3612 3148 3624
rect 3200 3652 3206 3664
rect 3329 3655 3387 3661
rect 3329 3652 3341 3655
rect 3200 3624 3341 3652
rect 3200 3612 3206 3624
rect 3329 3621 3341 3624
rect 3375 3621 3387 3655
rect 4246 3652 4252 3664
rect 4207 3624 4252 3652
rect 3329 3615 3387 3621
rect 4246 3612 4252 3624
rect 4304 3612 4310 3664
rect 4522 3612 4528 3664
rect 4580 3652 4586 3664
rect 4801 3655 4859 3661
rect 4801 3652 4813 3655
rect 4580 3624 4813 3652
rect 4580 3612 4586 3624
rect 4801 3621 4813 3624
rect 4847 3621 4859 3655
rect 7098 3652 7104 3664
rect 7059 3624 7104 3652
rect 4801 3615 4859 3621
rect 4816 3584 4844 3615
rect 7098 3612 7104 3624
rect 7156 3612 7162 3664
rect 12618 3612 12624 3664
rect 12676 3652 12682 3664
rect 12897 3655 12955 3661
rect 12897 3652 12909 3655
rect 12676 3624 12909 3652
rect 12676 3612 12682 3624
rect 12897 3621 12909 3624
rect 12943 3652 12955 3655
rect 13170 3652 13176 3664
rect 12943 3624 13176 3652
rect 12943 3621 12955 3624
rect 12897 3615 12955 3621
rect 13170 3612 13176 3624
rect 13228 3612 13234 3664
rect 5534 3584 5540 3596
rect 4816 3556 5540 3584
rect 5534 3544 5540 3556
rect 5592 3584 5598 3596
rect 5664 3587 5722 3593
rect 5664 3584 5676 3587
rect 5592 3556 5676 3584
rect 5592 3544 5598 3556
rect 5664 3553 5676 3556
rect 5710 3553 5722 3587
rect 5664 3547 5722 3553
rect 8640 3587 8698 3593
rect 8640 3553 8652 3587
rect 8686 3584 8698 3587
rect 8938 3584 8944 3596
rect 8686 3556 8944 3584
rect 8686 3553 8698 3556
rect 8640 3547 8698 3553
rect 8938 3544 8944 3556
rect 8996 3544 9002 3596
rect 9950 3544 9956 3596
rect 10008 3593 10014 3596
rect 10008 3587 10046 3593
rect 10034 3553 10046 3587
rect 10008 3547 10046 3553
rect 10008 3544 10014 3547
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 11460 3587 11518 3593
rect 11460 3584 11472 3587
rect 11296 3556 11472 3584
rect 11296 3544 11302 3556
rect 11460 3553 11472 3556
rect 11506 3553 11518 3587
rect 11460 3547 11518 3553
rect 15356 3587 15414 3593
rect 15356 3553 15368 3587
rect 15402 3584 15414 3587
rect 15654 3584 15660 3596
rect 15402 3556 15660 3584
rect 15402 3553 15414 3556
rect 15356 3547 15414 3553
rect 15654 3544 15660 3556
rect 15712 3544 15718 3596
rect 16574 3584 16580 3596
rect 16535 3556 16580 3584
rect 16574 3544 16580 3556
rect 16632 3544 16638 3596
rect 2225 3519 2283 3525
rect 2225 3485 2237 3519
rect 2271 3516 2283 3519
rect 2406 3516 2412 3528
rect 2271 3488 2412 3516
rect 2271 3485 2283 3488
rect 2225 3479 2283 3485
rect 2406 3476 2412 3488
rect 2464 3476 2470 3528
rect 4157 3519 4215 3525
rect 4157 3485 4169 3519
rect 4203 3516 4215 3519
rect 4982 3516 4988 3528
rect 4203 3488 4988 3516
rect 4203 3485 4215 3488
rect 4157 3479 4215 3485
rect 4982 3476 4988 3488
rect 5040 3476 5046 3528
rect 7006 3516 7012 3528
rect 6967 3488 7012 3516
rect 7006 3476 7012 3488
rect 7064 3476 7070 3528
rect 7374 3516 7380 3528
rect 7335 3488 7380 3516
rect 7374 3476 7380 3488
rect 7432 3476 7438 3528
rect 12802 3516 12808 3528
rect 12763 3488 12808 3516
rect 12802 3476 12808 3488
rect 12860 3476 12866 3528
rect 13081 3519 13139 3525
rect 13081 3485 13093 3519
rect 13127 3485 13139 3519
rect 13081 3479 13139 3485
rect 12434 3408 12440 3460
rect 12492 3448 12498 3460
rect 13096 3448 13124 3479
rect 12492 3420 13124 3448
rect 12492 3408 12498 3420
rect 16761 3383 16819 3389
rect 16761 3349 16773 3383
rect 16807 3380 16819 3383
rect 17862 3380 17868 3392
rect 16807 3352 17868 3380
rect 16807 3349 16819 3352
rect 16761 3343 16819 3349
rect 17862 3340 17868 3352
rect 17920 3340 17926 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 3789 3179 3847 3185
rect 3789 3145 3801 3179
rect 3835 3176 3847 3179
rect 3878 3176 3884 3188
rect 3835 3148 3884 3176
rect 3835 3145 3847 3148
rect 3789 3139 3847 3145
rect 3878 3136 3884 3148
rect 3936 3136 3942 3188
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 5629 3179 5687 3185
rect 5629 3176 5641 3179
rect 5592 3148 5641 3176
rect 5592 3136 5598 3148
rect 5629 3145 5641 3148
rect 5675 3145 5687 3179
rect 5629 3139 5687 3145
rect 6641 3179 6699 3185
rect 6641 3145 6653 3179
rect 6687 3176 6699 3179
rect 7006 3176 7012 3188
rect 6687 3148 7012 3176
rect 6687 3145 6699 3148
rect 6641 3139 6699 3145
rect 7006 3136 7012 3148
rect 7064 3176 7070 3188
rect 7975 3179 8033 3185
rect 7975 3176 7987 3179
rect 7064 3148 7987 3176
rect 7064 3136 7070 3148
rect 7975 3145 7987 3148
rect 8021 3145 8033 3179
rect 7975 3139 8033 3145
rect 8757 3179 8815 3185
rect 8757 3145 8769 3179
rect 8803 3176 8815 3179
rect 8938 3176 8944 3188
rect 8803 3148 8944 3176
rect 8803 3145 8815 3148
rect 8757 3139 8815 3145
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 11471 3179 11529 3185
rect 11471 3145 11483 3179
rect 11517 3176 11529 3179
rect 12802 3176 12808 3188
rect 11517 3148 12808 3176
rect 11517 3145 11529 3148
rect 11471 3139 11529 3145
rect 12802 3136 12808 3148
rect 12860 3176 12866 3188
rect 13725 3179 13783 3185
rect 13725 3176 13737 3179
rect 12860 3148 13737 3176
rect 12860 3136 12866 3148
rect 13725 3145 13737 3148
rect 13771 3145 13783 3179
rect 14550 3176 14556 3188
rect 14511 3148 14556 3176
rect 13725 3139 13783 3145
rect 14550 3136 14556 3148
rect 14608 3136 14614 3188
rect 15654 3176 15660 3188
rect 15615 3148 15660 3176
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 16574 3136 16580 3188
rect 16632 3176 16638 3188
rect 16669 3179 16727 3185
rect 16669 3176 16681 3179
rect 16632 3148 16681 3176
rect 16632 3136 16638 3148
rect 16669 3145 16681 3148
rect 16715 3145 16727 3179
rect 17034 3176 17040 3188
rect 16995 3148 17040 3176
rect 16669 3139 16727 3145
rect 17034 3136 17040 3148
rect 17092 3136 17098 3188
rect 18690 3185 18696 3188
rect 18647 3179 18696 3185
rect 18647 3145 18659 3179
rect 18693 3145 18696 3179
rect 18647 3139 18696 3145
rect 18690 3136 18696 3139
rect 18748 3136 18754 3188
rect 4893 3111 4951 3117
rect 4893 3077 4905 3111
rect 4939 3108 4951 3111
rect 4982 3108 4988 3120
rect 4939 3080 4988 3108
rect 4939 3077 4951 3080
rect 4893 3071 4951 3077
rect 4982 3068 4988 3080
rect 5040 3068 5046 3120
rect 7098 3068 7104 3120
rect 7156 3108 7162 3120
rect 7653 3111 7711 3117
rect 7653 3108 7665 3111
rect 7156 3080 7665 3108
rect 7156 3068 7162 3080
rect 7653 3077 7665 3080
rect 7699 3077 7711 3111
rect 9950 3108 9956 3120
rect 9911 3080 9956 3108
rect 7653 3071 7711 3077
rect 9950 3068 9956 3080
rect 10008 3068 10014 3120
rect 12158 3108 12164 3120
rect 12119 3080 12164 3108
rect 12158 3068 12164 3080
rect 12216 3068 12222 3120
rect 12621 3111 12679 3117
rect 12621 3077 12633 3111
rect 12667 3108 12679 3111
rect 13906 3108 13912 3120
rect 12667 3080 13912 3108
rect 12667 3077 12679 3080
rect 12621 3071 12679 3077
rect 13906 3068 13912 3080
rect 13964 3068 13970 3120
rect 14093 3111 14151 3117
rect 14093 3077 14105 3111
rect 14139 3108 14151 3111
rect 15930 3108 15936 3120
rect 14139 3080 15936 3108
rect 14139 3077 14151 3080
rect 14093 3071 14151 3077
rect 15930 3068 15936 3080
rect 15988 3068 15994 3120
rect 2225 3043 2283 3049
rect 2225 3009 2237 3043
rect 2271 3040 2283 3043
rect 2774 3040 2780 3052
rect 2271 3012 2780 3040
rect 2271 3009 2283 3012
rect 2225 3003 2283 3009
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 3142 3040 3148 3052
rect 3103 3012 3148 3040
rect 3142 3000 3148 3012
rect 3200 3000 3206 3052
rect 4338 3040 4344 3052
rect 4251 3012 4344 3040
rect 4338 3000 4344 3012
rect 4396 3040 4402 3052
rect 5261 3043 5319 3049
rect 5261 3040 5273 3043
rect 4396 3012 5273 3040
rect 4396 3000 4402 3012
rect 5261 3009 5273 3012
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 6963 3043 7021 3049
rect 6963 3009 6975 3043
rect 7009 3040 7021 3043
rect 8202 3040 8208 3052
rect 7009 3012 8208 3040
rect 7009 3009 7021 3012
rect 6963 3003 7021 3009
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 11882 3040 11888 3052
rect 11843 3012 11888 3040
rect 11882 3000 11888 3012
rect 11940 3000 11946 3052
rect 13170 3000 13176 3052
rect 13228 3040 13234 3052
rect 13357 3043 13415 3049
rect 13357 3040 13369 3043
rect 13228 3012 13369 3040
rect 13228 3000 13234 3012
rect 13357 3009 13369 3012
rect 13403 3009 13415 3043
rect 13357 3003 13415 3009
rect 1394 2972 1400 2984
rect 1355 2944 1400 2972
rect 1394 2932 1400 2944
rect 1452 2932 1458 2984
rect 6876 2975 6934 2981
rect 6876 2941 6888 2975
rect 6922 2972 6934 2975
rect 7374 2972 7380 2984
rect 6922 2944 7380 2972
rect 6922 2941 6934 2944
rect 6876 2935 6934 2941
rect 7374 2932 7380 2944
rect 7432 2932 7438 2984
rect 7904 2975 7962 2981
rect 7904 2941 7916 2975
rect 7950 2972 7962 2975
rect 11400 2975 11458 2981
rect 7950 2944 8432 2972
rect 7950 2941 7962 2944
rect 7904 2935 7962 2941
rect 8404 2913 8432 2944
rect 11400 2941 11412 2975
rect 11446 2972 11458 2975
rect 11900 2972 11928 3000
rect 11446 2944 11928 2972
rect 11446 2941 11458 2944
rect 11400 2935 11458 2941
rect 11974 2932 11980 2984
rect 12032 2972 12038 2984
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 12032 2944 12449 2972
rect 12032 2932 12038 2944
rect 12437 2941 12449 2944
rect 12483 2972 12495 2975
rect 12989 2975 13047 2981
rect 12989 2972 13001 2975
rect 12483 2944 13001 2972
rect 12483 2941 12495 2944
rect 12437 2935 12495 2941
rect 12989 2941 13001 2944
rect 13035 2941 13047 2975
rect 12989 2935 13047 2941
rect 13909 2975 13967 2981
rect 13909 2941 13921 2975
rect 13955 2972 13967 2975
rect 14550 2972 14556 2984
rect 13955 2944 14556 2972
rect 13955 2941 13967 2944
rect 13909 2935 13967 2941
rect 14550 2932 14556 2944
rect 14608 2932 14614 2984
rect 14921 2975 14979 2981
rect 14921 2941 14933 2975
rect 14967 2972 14979 2975
rect 15013 2975 15071 2981
rect 15013 2972 15025 2975
rect 14967 2944 15025 2972
rect 14967 2941 14979 2944
rect 14921 2935 14979 2941
rect 15013 2941 15025 2944
rect 15059 2941 15071 2975
rect 15013 2935 15071 2941
rect 16260 2975 16318 2981
rect 16260 2941 16272 2975
rect 16306 2972 16318 2975
rect 17034 2972 17040 2984
rect 16306 2944 17040 2972
rect 16306 2941 16318 2944
rect 16260 2935 16318 2941
rect 2869 2907 2927 2913
rect 2869 2873 2881 2907
rect 2915 2873 2927 2907
rect 2869 2867 2927 2873
rect 4157 2907 4215 2913
rect 4157 2873 4169 2907
rect 4203 2904 4215 2907
rect 4433 2907 4491 2913
rect 4433 2904 4445 2907
rect 4203 2876 4445 2904
rect 4203 2873 4215 2876
rect 4157 2867 4215 2873
rect 4433 2873 4445 2876
rect 4479 2873 4491 2907
rect 4433 2867 4491 2873
rect 8389 2907 8447 2913
rect 8389 2873 8401 2907
rect 8435 2904 8447 2907
rect 8754 2904 8760 2916
rect 8435 2876 8760 2904
rect 8435 2873 8447 2876
rect 8389 2867 8447 2873
rect 1578 2836 1584 2848
rect 1539 2808 1584 2836
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 2593 2839 2651 2845
rect 2593 2805 2605 2839
rect 2639 2836 2651 2839
rect 2884 2836 2912 2867
rect 3142 2836 3148 2848
rect 2639 2808 3148 2836
rect 2639 2805 2651 2808
rect 2593 2799 2651 2805
rect 3142 2796 3148 2808
rect 3200 2836 3206 2848
rect 4172 2836 4200 2867
rect 8754 2864 8760 2876
rect 8812 2864 8818 2916
rect 15028 2904 15056 2935
rect 17034 2932 17040 2944
rect 17092 2932 17098 2984
rect 18576 2975 18634 2981
rect 18576 2941 18588 2975
rect 18622 2972 18634 2975
rect 18622 2944 19104 2972
rect 18622 2941 18634 2944
rect 18576 2935 18634 2941
rect 19076 2916 19104 2944
rect 16347 2907 16405 2913
rect 16347 2904 16359 2907
rect 15028 2876 16359 2904
rect 16347 2873 16359 2876
rect 16393 2873 16405 2907
rect 19058 2904 19064 2916
rect 19019 2876 19064 2904
rect 16347 2867 16405 2873
rect 19058 2864 19064 2876
rect 19116 2864 19122 2916
rect 3200 2808 4200 2836
rect 3200 2796 3206 2808
rect 14918 2796 14924 2848
rect 14976 2836 14982 2848
rect 15197 2839 15255 2845
rect 15197 2836 15209 2839
rect 14976 2808 15209 2836
rect 14976 2796 14982 2808
rect 15197 2805 15209 2808
rect 15243 2805 15255 2839
rect 15197 2799 15255 2805
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 1535 2635 1593 2641
rect 1535 2601 1547 2635
rect 1581 2632 1593 2635
rect 2682 2632 2688 2644
rect 1581 2604 2688 2632
rect 1581 2601 1593 2604
rect 1535 2595 1593 2601
rect 2682 2592 2688 2604
rect 2740 2592 2746 2644
rect 2774 2592 2780 2644
rect 2832 2632 2838 2644
rect 4065 2635 4123 2641
rect 4065 2632 4077 2635
rect 2832 2604 4077 2632
rect 2832 2592 2838 2604
rect 4065 2601 4077 2604
rect 4111 2601 4123 2635
rect 4065 2595 4123 2601
rect 4246 2592 4252 2644
rect 4304 2632 4310 2644
rect 4525 2635 4583 2641
rect 4525 2632 4537 2635
rect 4304 2604 4537 2632
rect 4304 2592 4310 2604
rect 4525 2601 4537 2604
rect 4571 2601 4583 2635
rect 4982 2632 4988 2644
rect 4943 2604 4988 2632
rect 4525 2595 4583 2601
rect 4982 2592 4988 2604
rect 5040 2592 5046 2644
rect 5074 2592 5080 2644
rect 5132 2632 5138 2644
rect 5215 2635 5273 2641
rect 5215 2632 5227 2635
rect 5132 2604 5227 2632
rect 5132 2592 5138 2604
rect 5215 2601 5227 2604
rect 5261 2601 5273 2635
rect 5215 2595 5273 2601
rect 6914 2592 6920 2644
rect 6972 2632 6978 2644
rect 7055 2635 7113 2641
rect 7055 2632 7067 2635
rect 6972 2604 7067 2632
rect 6972 2592 6978 2604
rect 7055 2601 7067 2604
rect 7101 2601 7113 2635
rect 7055 2595 7113 2601
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 7377 2635 7435 2641
rect 7377 2632 7389 2635
rect 7248 2604 7389 2632
rect 7248 2592 7254 2604
rect 7377 2601 7389 2604
rect 7423 2601 7435 2635
rect 7377 2595 7435 2601
rect 13078 2592 13084 2644
rect 13136 2632 13142 2644
rect 13173 2635 13231 2641
rect 13173 2632 13185 2635
rect 13136 2604 13185 2632
rect 13136 2592 13142 2604
rect 13173 2601 13185 2604
rect 13219 2601 13231 2635
rect 14458 2632 14464 2644
rect 14419 2604 14464 2632
rect 13173 2595 13231 2601
rect 14458 2592 14464 2604
rect 14516 2592 14522 2644
rect 18322 2592 18328 2644
rect 18380 2632 18386 2644
rect 18923 2635 18981 2641
rect 18923 2632 18935 2635
rect 18380 2604 18935 2632
rect 18380 2592 18386 2604
rect 18923 2601 18935 2604
rect 18969 2601 18981 2635
rect 18923 2595 18981 2601
rect 24670 2592 24676 2644
rect 24728 2641 24734 2644
rect 24728 2635 24777 2641
rect 24728 2601 24731 2635
rect 24765 2601 24777 2635
rect 24728 2595 24777 2601
rect 24728 2592 24734 2595
rect 3142 2564 3148 2576
rect 3103 2536 3148 2564
rect 3142 2524 3148 2536
rect 3200 2524 3206 2576
rect 1464 2499 1522 2505
rect 1464 2465 1476 2499
rect 1510 2496 1522 2499
rect 1946 2496 1952 2508
rect 1510 2468 1952 2496
rect 1510 2465 1522 2468
rect 1464 2459 1522 2465
rect 1946 2456 1952 2468
rect 2004 2456 2010 2508
rect 2317 2499 2375 2505
rect 2317 2465 2329 2499
rect 2363 2496 2375 2499
rect 3053 2499 3111 2505
rect 3053 2496 3065 2499
rect 2363 2468 3065 2496
rect 2363 2465 2375 2468
rect 2317 2459 2375 2465
rect 3053 2465 3065 2468
rect 3099 2496 3111 2499
rect 3878 2496 3884 2508
rect 3099 2468 3884 2496
rect 3099 2465 3111 2468
rect 3053 2459 3111 2465
rect 3878 2456 3884 2468
rect 3936 2456 3942 2508
rect 4154 2456 4160 2508
rect 4212 2496 4218 2508
rect 5112 2499 5170 2505
rect 5112 2496 5124 2499
rect 4212 2468 5124 2496
rect 4212 2456 4218 2468
rect 5112 2465 5124 2468
rect 5158 2496 5170 2499
rect 5537 2499 5595 2505
rect 5537 2496 5549 2499
rect 5158 2468 5549 2496
rect 5158 2465 5170 2468
rect 5112 2459 5170 2465
rect 5537 2465 5549 2468
rect 5583 2465 5595 2499
rect 5537 2459 5595 2465
rect 6984 2499 7042 2505
rect 6984 2465 6996 2499
rect 7030 2496 7042 2499
rect 7208 2496 7236 2592
rect 7030 2468 7236 2496
rect 7030 2465 7042 2468
rect 6984 2459 7042 2465
rect 10042 2456 10048 2508
rect 10100 2496 10106 2508
rect 10597 2499 10655 2505
rect 10597 2496 10609 2499
rect 10100 2468 10609 2496
rect 10100 2456 10106 2468
rect 10597 2465 10609 2468
rect 10643 2496 10655 2499
rect 11149 2499 11207 2505
rect 11149 2496 11161 2499
rect 10643 2468 11161 2496
rect 10643 2465 10655 2468
rect 10597 2459 10655 2465
rect 11149 2465 11161 2468
rect 11195 2465 11207 2499
rect 11149 2459 11207 2465
rect 12621 2499 12679 2505
rect 12621 2465 12633 2499
rect 12667 2496 12679 2499
rect 13096 2496 13124 2592
rect 14274 2496 14280 2508
rect 12667 2468 13124 2496
rect 14235 2468 14280 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 14274 2456 14280 2468
rect 14332 2496 14338 2508
rect 14829 2499 14887 2505
rect 14829 2496 14841 2499
rect 14332 2468 14841 2496
rect 14332 2456 14338 2468
rect 14829 2465 14841 2468
rect 14875 2465 14887 2499
rect 16022 2496 16028 2508
rect 15935 2468 16028 2496
rect 14829 2459 14887 2465
rect 16022 2456 16028 2468
rect 16080 2496 16086 2508
rect 16577 2499 16635 2505
rect 16577 2496 16589 2499
rect 16080 2468 16589 2496
rect 16080 2456 16086 2468
rect 16577 2465 16589 2468
rect 16623 2465 16635 2499
rect 16577 2459 16635 2465
rect 18852 2499 18910 2505
rect 18852 2465 18864 2499
rect 18898 2496 18910 2499
rect 24648 2499 24706 2505
rect 18898 2468 19380 2496
rect 18898 2465 18910 2468
rect 18852 2459 18910 2465
rect 10781 2363 10839 2369
rect 10781 2329 10793 2363
rect 10827 2360 10839 2363
rect 11790 2360 11796 2372
rect 10827 2332 11796 2360
rect 10827 2329 10839 2332
rect 10781 2323 10839 2329
rect 11790 2320 11796 2332
rect 11848 2320 11854 2372
rect 16209 2363 16267 2369
rect 16209 2329 16221 2363
rect 16255 2360 16267 2363
rect 18046 2360 18052 2372
rect 16255 2332 18052 2360
rect 16255 2329 16267 2332
rect 16209 2323 16267 2329
rect 18046 2320 18052 2332
rect 18104 2320 18110 2372
rect 1946 2292 1952 2304
rect 1907 2264 1952 2292
rect 1946 2252 1952 2264
rect 2004 2252 2010 2304
rect 12805 2295 12863 2301
rect 12805 2261 12817 2295
rect 12851 2292 12863 2295
rect 12894 2292 12900 2304
rect 12851 2264 12900 2292
rect 12851 2261 12863 2264
rect 12805 2255 12863 2261
rect 12894 2252 12900 2264
rect 12952 2252 12958 2304
rect 19352 2301 19380 2468
rect 24648 2465 24660 2499
rect 24694 2496 24706 2499
rect 25130 2496 25136 2508
rect 24694 2468 25136 2496
rect 24694 2465 24706 2468
rect 24648 2459 24706 2465
rect 25130 2456 25136 2468
rect 25188 2456 25194 2508
rect 19337 2295 19395 2301
rect 19337 2261 19349 2295
rect 19383 2292 19395 2295
rect 21174 2292 21180 2304
rect 19383 2264 21180 2292
rect 19383 2261 19395 2264
rect 19337 2255 19395 2261
rect 21174 2252 21180 2264
rect 21232 2252 21238 2304
rect 25130 2292 25136 2304
rect 25091 2264 25136 2292
rect 25130 2252 25136 2264
rect 25188 2252 25194 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
<< via1 >>
rect 17500 26324 17552 26376
rect 24768 26324 24820 26376
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 13820 25347 13872 25356
rect 13820 25313 13864 25347
rect 13864 25313 13872 25347
rect 13820 25304 13872 25313
rect 14188 25100 14240 25152
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 2964 24828 3016 24880
rect 12532 24828 12584 24880
rect 16672 24803 16724 24812
rect 16672 24769 16681 24803
rect 16681 24769 16715 24803
rect 16715 24769 16724 24803
rect 16672 24760 16724 24769
rect 10692 24556 10744 24608
rect 14280 24692 14332 24744
rect 14740 24692 14792 24744
rect 13820 24667 13872 24676
rect 13820 24633 13829 24667
rect 13829 24633 13863 24667
rect 13863 24633 13872 24667
rect 13820 24624 13872 24633
rect 12072 24556 12124 24608
rect 14096 24599 14148 24608
rect 14096 24565 14105 24599
rect 14105 24565 14139 24599
rect 14139 24565 14148 24599
rect 14096 24556 14148 24565
rect 17040 24624 17092 24676
rect 16304 24556 16356 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 10140 24395 10192 24404
rect 10140 24361 10149 24395
rect 10149 24361 10183 24395
rect 10183 24361 10192 24395
rect 10140 24352 10192 24361
rect 12900 24352 12952 24404
rect 13728 24352 13780 24404
rect 14832 24352 14884 24404
rect 17868 24352 17920 24404
rect 13912 24284 13964 24336
rect 14280 24284 14332 24336
rect 15476 24327 15528 24336
rect 15476 24293 15485 24327
rect 15485 24293 15519 24327
rect 15519 24293 15528 24327
rect 15476 24284 15528 24293
rect 9956 24259 10008 24268
rect 9956 24225 9965 24259
rect 9965 24225 9999 24259
rect 9999 24225 10008 24259
rect 9956 24216 10008 24225
rect 11704 24259 11756 24268
rect 11704 24225 11713 24259
rect 11713 24225 11747 24259
rect 11747 24225 11756 24259
rect 11704 24216 11756 24225
rect 13544 24216 13596 24268
rect 14648 24216 14700 24268
rect 16580 24216 16632 24268
rect 18328 24259 18380 24268
rect 18328 24225 18346 24259
rect 18346 24225 18380 24259
rect 18328 24216 18380 24225
rect 16028 24191 16080 24200
rect 15292 24080 15344 24132
rect 12624 24055 12676 24064
rect 12624 24021 12633 24055
rect 12633 24021 12667 24055
rect 12667 24021 12676 24055
rect 12624 24012 12676 24021
rect 16028 24157 16037 24191
rect 16037 24157 16071 24191
rect 16071 24157 16080 24191
rect 16028 24148 16080 24157
rect 16396 24123 16448 24132
rect 16396 24089 16405 24123
rect 16405 24089 16439 24123
rect 16439 24089 16448 24123
rect 16396 24080 16448 24089
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 480 23604 532 23656
rect 2688 23604 2740 23656
rect 4620 23808 4672 23860
rect 8760 23808 8812 23860
rect 9588 23808 9640 23860
rect 10692 23851 10744 23860
rect 10692 23817 10701 23851
rect 10701 23817 10735 23851
rect 10735 23817 10744 23851
rect 10692 23808 10744 23817
rect 15476 23808 15528 23860
rect 19064 23808 19116 23860
rect 16028 23740 16080 23792
rect 18328 23740 18380 23792
rect 12256 23715 12308 23724
rect 12256 23681 12265 23715
rect 12265 23681 12299 23715
rect 12299 23681 12308 23715
rect 12256 23672 12308 23681
rect 14188 23715 14240 23724
rect 14188 23681 14197 23715
rect 14197 23681 14231 23715
rect 14231 23681 14240 23715
rect 14188 23672 14240 23681
rect 14280 23672 14332 23724
rect 16396 23672 16448 23724
rect 12716 23647 12768 23656
rect 12716 23613 12725 23647
rect 12725 23613 12759 23647
rect 12759 23613 12768 23647
rect 12716 23604 12768 23613
rect 12624 23536 12676 23588
rect 13268 23579 13320 23588
rect 13268 23545 13277 23579
rect 13277 23545 13311 23579
rect 13311 23545 13320 23579
rect 13268 23536 13320 23545
rect 15016 23536 15068 23588
rect 15844 23579 15896 23588
rect 15844 23545 15853 23579
rect 15853 23545 15887 23579
rect 15887 23545 15896 23579
rect 15844 23536 15896 23545
rect 22192 23808 22244 23860
rect 23480 23808 23532 23860
rect 26148 23808 26200 23860
rect 2872 23468 2924 23520
rect 7564 23468 7616 23520
rect 8852 23468 8904 23520
rect 9956 23511 10008 23520
rect 9956 23477 9965 23511
rect 9965 23477 9999 23511
rect 9999 23477 10008 23511
rect 9956 23468 10008 23477
rect 10784 23468 10836 23520
rect 11336 23468 11388 23520
rect 11704 23468 11756 23520
rect 12440 23468 12492 23520
rect 13544 23511 13596 23520
rect 13544 23477 13553 23511
rect 13553 23477 13587 23511
rect 13587 23477 13596 23511
rect 13544 23468 13596 23477
rect 14096 23468 14148 23520
rect 16580 23468 16632 23520
rect 19432 23468 19484 23520
rect 19984 23468 20036 23520
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 9864 23239 9916 23248
rect 9864 23205 9873 23239
rect 9873 23205 9907 23239
rect 9907 23205 9916 23239
rect 9864 23196 9916 23205
rect 11336 23239 11388 23248
rect 11336 23205 11345 23239
rect 11345 23205 11379 23239
rect 11379 23205 11388 23239
rect 11336 23196 11388 23205
rect 11428 23239 11480 23248
rect 11428 23205 11437 23239
rect 11437 23205 11471 23239
rect 11471 23205 11480 23239
rect 11428 23196 11480 23205
rect 9772 23103 9824 23112
rect 9772 23069 9781 23103
rect 9781 23069 9815 23103
rect 9815 23069 9824 23103
rect 9772 23060 9824 23069
rect 12992 23239 13044 23248
rect 12992 23205 13001 23239
rect 13001 23205 13035 23239
rect 13035 23205 13044 23239
rect 12992 23196 13044 23205
rect 13268 23264 13320 23316
rect 13636 23264 13688 23316
rect 14188 23307 14240 23316
rect 14188 23273 14197 23307
rect 14197 23273 14231 23307
rect 14231 23273 14240 23307
rect 14188 23264 14240 23273
rect 15108 23307 15160 23316
rect 15108 23273 15117 23307
rect 15117 23273 15151 23307
rect 15151 23273 15160 23307
rect 15108 23264 15160 23273
rect 14648 23239 14700 23248
rect 14648 23205 14657 23239
rect 14657 23205 14691 23239
rect 14691 23205 14700 23239
rect 15476 23239 15528 23248
rect 14648 23196 14700 23205
rect 15476 23205 15485 23239
rect 15485 23205 15519 23239
rect 15519 23205 15528 23239
rect 15476 23196 15528 23205
rect 18512 23196 18564 23248
rect 12900 23103 12952 23112
rect 12900 23069 12909 23103
rect 12909 23069 12943 23103
rect 12943 23069 12952 23103
rect 12900 23060 12952 23069
rect 16028 23060 16080 23112
rect 11244 22992 11296 23044
rect 14832 22992 14884 23044
rect 17132 23128 17184 23180
rect 21180 23128 21232 23180
rect 24676 23171 24728 23180
rect 24676 23137 24694 23171
rect 24694 23137 24728 23171
rect 24676 23128 24728 23137
rect 17868 23060 17920 23112
rect 19248 23035 19300 23044
rect 19248 23001 19257 23035
rect 19257 23001 19291 23035
rect 19291 23001 19300 23035
rect 19248 22992 19300 23001
rect 12716 22924 12768 22976
rect 13084 22924 13136 22976
rect 15844 22924 15896 22976
rect 23480 22924 23532 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 9772 22720 9824 22772
rect 12900 22720 12952 22772
rect 15476 22720 15528 22772
rect 12532 22652 12584 22704
rect 12716 22652 12768 22704
rect 15292 22695 15344 22704
rect 15292 22661 15301 22695
rect 15301 22661 15335 22695
rect 15335 22661 15344 22695
rect 15292 22652 15344 22661
rect 10876 22584 10928 22636
rect 10692 22516 10744 22568
rect 13636 22627 13688 22636
rect 12532 22559 12584 22568
rect 12532 22525 12550 22559
rect 12550 22525 12584 22559
rect 12532 22516 12584 22525
rect 11152 22448 11204 22500
rect 11428 22448 11480 22500
rect 13636 22593 13645 22627
rect 13645 22593 13679 22627
rect 13679 22593 13688 22627
rect 13636 22584 13688 22593
rect 16304 22720 16356 22772
rect 17132 22763 17184 22772
rect 17132 22729 17141 22763
rect 17141 22729 17175 22763
rect 17175 22729 17184 22763
rect 17132 22720 17184 22729
rect 17868 22763 17920 22772
rect 17868 22729 17877 22763
rect 17877 22729 17911 22763
rect 17911 22729 17920 22763
rect 17868 22720 17920 22729
rect 19800 22763 19852 22772
rect 19800 22729 19809 22763
rect 19809 22729 19843 22763
rect 19843 22729 19852 22763
rect 19800 22720 19852 22729
rect 20168 22763 20220 22772
rect 20168 22729 20177 22763
rect 20177 22729 20211 22763
rect 20211 22729 20220 22763
rect 20168 22720 20220 22729
rect 21180 22720 21232 22772
rect 24676 22763 24728 22772
rect 24676 22729 24685 22763
rect 24685 22729 24719 22763
rect 24719 22729 24728 22763
rect 24676 22720 24728 22729
rect 16028 22695 16080 22704
rect 16028 22661 16037 22695
rect 16037 22661 16071 22695
rect 16071 22661 16080 22695
rect 16028 22652 16080 22661
rect 19248 22627 19300 22636
rect 19248 22593 19257 22627
rect 19257 22593 19291 22627
rect 19291 22593 19300 22627
rect 19248 22584 19300 22593
rect 20168 22516 20220 22568
rect 13636 22448 13688 22500
rect 15292 22448 15344 22500
rect 18880 22491 18932 22500
rect 18880 22457 18889 22491
rect 18889 22457 18923 22491
rect 18923 22457 18932 22491
rect 18880 22448 18932 22457
rect 9864 22380 9916 22432
rect 11520 22423 11572 22432
rect 11520 22389 11529 22423
rect 11529 22389 11563 22423
rect 11563 22389 11572 22423
rect 11520 22380 11572 22389
rect 12716 22380 12768 22432
rect 18052 22380 18104 22432
rect 18512 22423 18564 22432
rect 18512 22389 18521 22423
rect 18521 22389 18555 22423
rect 18555 22389 18564 22423
rect 18512 22380 18564 22389
rect 19340 22380 19392 22432
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 12992 22176 13044 22228
rect 11244 22151 11296 22160
rect 11244 22117 11253 22151
rect 11253 22117 11287 22151
rect 11287 22117 11296 22151
rect 11244 22108 11296 22117
rect 11520 22108 11572 22160
rect 13728 22151 13780 22160
rect 13728 22117 13737 22151
rect 13737 22117 13771 22151
rect 13771 22117 13780 22151
rect 13728 22108 13780 22117
rect 16212 22151 16264 22160
rect 16212 22117 16221 22151
rect 16221 22117 16255 22151
rect 16255 22117 16264 22151
rect 16212 22108 16264 22117
rect 17500 22151 17552 22160
rect 17500 22117 17503 22151
rect 17503 22117 17537 22151
rect 17537 22117 17552 22151
rect 17500 22108 17552 22117
rect 18788 22151 18840 22160
rect 18788 22117 18797 22151
rect 18797 22117 18831 22151
rect 18831 22117 18840 22151
rect 18788 22108 18840 22117
rect 19064 22151 19116 22160
rect 19064 22117 19073 22151
rect 19073 22117 19107 22151
rect 19107 22117 19116 22151
rect 19064 22108 19116 22117
rect 14280 22083 14332 22092
rect 14280 22049 14289 22083
rect 14289 22049 14323 22083
rect 14323 22049 14332 22083
rect 14280 22040 14332 22049
rect 15384 22040 15436 22092
rect 16488 22040 16540 22092
rect 12072 21972 12124 22024
rect 12808 21972 12860 22024
rect 17132 22015 17184 22024
rect 17132 21981 17141 22015
rect 17141 21981 17175 22015
rect 17175 21981 17184 22015
rect 17132 21972 17184 21981
rect 18972 22015 19024 22024
rect 18972 21981 18981 22015
rect 18981 21981 19015 22015
rect 19015 21981 19024 22015
rect 18972 21972 19024 21981
rect 19248 21972 19300 22024
rect 19432 22015 19484 22024
rect 19432 21981 19441 22015
rect 19441 21981 19475 22015
rect 19475 21981 19484 22015
rect 19432 21972 19484 21981
rect 8944 21836 8996 21888
rect 9128 21836 9180 21888
rect 10692 21836 10744 21888
rect 14004 21836 14056 21888
rect 16488 21879 16540 21888
rect 16488 21845 16497 21879
rect 16497 21845 16531 21879
rect 16531 21845 16540 21879
rect 16488 21836 16540 21845
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 9864 21632 9916 21684
rect 11244 21632 11296 21684
rect 12808 21675 12860 21684
rect 12808 21641 12817 21675
rect 12817 21641 12851 21675
rect 12851 21641 12860 21675
rect 12808 21632 12860 21641
rect 13820 21675 13872 21684
rect 13820 21641 13829 21675
rect 13829 21641 13863 21675
rect 13863 21641 13872 21675
rect 13820 21632 13872 21641
rect 19064 21632 19116 21684
rect 9128 21539 9180 21548
rect 9128 21505 9137 21539
rect 9137 21505 9171 21539
rect 9171 21505 9180 21539
rect 9128 21496 9180 21505
rect 11520 21496 11572 21548
rect 14004 21539 14056 21548
rect 14004 21505 14013 21539
rect 14013 21505 14047 21539
rect 14047 21505 14056 21539
rect 14004 21496 14056 21505
rect 14372 21539 14424 21548
rect 14372 21505 14381 21539
rect 14381 21505 14415 21539
rect 14415 21505 14424 21539
rect 14372 21496 14424 21505
rect 17132 21496 17184 21548
rect 17960 21496 18012 21548
rect 18788 21496 18840 21548
rect 18972 21496 19024 21548
rect 8944 21471 8996 21480
rect 8944 21437 8953 21471
rect 8953 21437 8987 21471
rect 8987 21437 8996 21471
rect 8944 21428 8996 21437
rect 9680 21428 9732 21480
rect 12900 21428 12952 21480
rect 15752 21471 15804 21480
rect 10876 21360 10928 21412
rect 15752 21437 15761 21471
rect 15761 21437 15795 21471
rect 15795 21437 15804 21471
rect 15752 21428 15804 21437
rect 16488 21471 16540 21480
rect 16488 21437 16497 21471
rect 16497 21437 16531 21471
rect 16531 21437 16540 21471
rect 16488 21428 16540 21437
rect 14096 21403 14148 21412
rect 14096 21369 14105 21403
rect 14105 21369 14139 21403
rect 14139 21369 14148 21403
rect 14096 21360 14148 21369
rect 8300 21335 8352 21344
rect 8300 21301 8309 21335
rect 8309 21301 8343 21335
rect 8343 21301 8352 21335
rect 8300 21292 8352 21301
rect 13452 21335 13504 21344
rect 13452 21301 13461 21335
rect 13461 21301 13495 21335
rect 13495 21301 13504 21335
rect 13452 21292 13504 21301
rect 15384 21335 15436 21344
rect 15384 21301 15393 21335
rect 15393 21301 15427 21335
rect 15427 21301 15436 21335
rect 15384 21292 15436 21301
rect 16672 21292 16724 21344
rect 17500 21292 17552 21344
rect 18788 21403 18840 21412
rect 18788 21369 18797 21403
rect 18797 21369 18831 21403
rect 18831 21369 18840 21403
rect 18788 21360 18840 21369
rect 19340 21292 19392 21344
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 10968 21088 11020 21140
rect 12992 21088 13044 21140
rect 14096 21088 14148 21140
rect 10876 21020 10928 21072
rect 13084 21020 13136 21072
rect 13636 21020 13688 21072
rect 8300 20995 8352 21004
rect 8300 20961 8309 20995
rect 8309 20961 8343 20995
rect 8343 20961 8352 20995
rect 8300 20952 8352 20961
rect 8576 20995 8628 21004
rect 8576 20961 8585 20995
rect 8585 20961 8619 20995
rect 8619 20961 8628 20995
rect 8576 20952 8628 20961
rect 11888 20952 11940 21004
rect 13820 20952 13872 21004
rect 16120 20952 16172 21004
rect 17224 21088 17276 21140
rect 19340 21131 19392 21140
rect 19340 21097 19349 21131
rect 19349 21097 19383 21131
rect 19383 21097 19392 21131
rect 19340 21088 19392 21097
rect 16672 21020 16724 21072
rect 18052 21063 18104 21072
rect 18052 21029 18061 21063
rect 18061 21029 18095 21063
rect 18095 21029 18104 21063
rect 18052 21020 18104 21029
rect 18512 20995 18564 21004
rect 18512 20961 18521 20995
rect 18521 20961 18555 20995
rect 18555 20961 18564 20995
rect 18512 20952 18564 20961
rect 11060 20884 11112 20936
rect 13176 20927 13228 20936
rect 13176 20893 13185 20927
rect 13185 20893 13219 20927
rect 13219 20893 13228 20927
rect 13176 20884 13228 20893
rect 16580 20884 16632 20936
rect 17776 20884 17828 20936
rect 9680 20748 9732 20800
rect 12440 20748 12492 20800
rect 16028 20748 16080 20800
rect 16672 20748 16724 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 8576 20544 8628 20596
rect 10876 20544 10928 20596
rect 11060 20544 11112 20596
rect 11888 20544 11940 20596
rect 12348 20544 12400 20596
rect 14096 20544 14148 20596
rect 18512 20544 18564 20596
rect 9680 20408 9732 20460
rect 11060 20451 11112 20460
rect 11060 20417 11069 20451
rect 11069 20417 11103 20451
rect 11103 20417 11112 20451
rect 11060 20408 11112 20417
rect 16212 20451 16264 20460
rect 16212 20417 16221 20451
rect 16221 20417 16255 20451
rect 16255 20417 16264 20451
rect 16212 20408 16264 20417
rect 16580 20408 16632 20460
rect 17776 20451 17828 20460
rect 17776 20417 17785 20451
rect 17785 20417 17819 20451
rect 17819 20417 17828 20451
rect 17776 20408 17828 20417
rect 9128 20340 9180 20392
rect 12808 20340 12860 20392
rect 15200 20383 15252 20392
rect 15200 20349 15244 20383
rect 15244 20349 15252 20383
rect 15200 20340 15252 20349
rect 17868 20340 17920 20392
rect 19616 20383 19668 20392
rect 19616 20349 19660 20383
rect 19660 20349 19668 20383
rect 19616 20340 19668 20349
rect 20168 20340 20220 20392
rect 10140 20272 10192 20324
rect 8300 20204 8352 20256
rect 8760 20247 8812 20256
rect 8760 20213 8769 20247
rect 8769 20213 8803 20247
rect 8803 20213 8812 20247
rect 8760 20204 8812 20213
rect 10048 20247 10100 20256
rect 10048 20213 10057 20247
rect 10057 20213 10091 20247
rect 10091 20213 10100 20247
rect 10968 20272 11020 20324
rect 10048 20204 10100 20213
rect 13084 20204 13136 20256
rect 16672 20272 16724 20324
rect 18144 20315 18196 20324
rect 18144 20281 18153 20315
rect 18153 20281 18187 20315
rect 18187 20281 18196 20315
rect 18144 20272 18196 20281
rect 15568 20204 15620 20256
rect 16120 20247 16172 20256
rect 16120 20213 16129 20247
rect 16129 20213 16163 20247
rect 16163 20213 16172 20247
rect 16120 20204 16172 20213
rect 17040 20204 17092 20256
rect 18052 20204 18104 20256
rect 18972 20272 19024 20324
rect 19340 20204 19392 20256
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 13176 20043 13228 20052
rect 13176 20009 13185 20043
rect 13185 20009 13219 20043
rect 13219 20009 13228 20043
rect 13176 20000 13228 20009
rect 16212 20000 16264 20052
rect 17224 20043 17276 20052
rect 17224 20009 17233 20043
rect 17233 20009 17267 20043
rect 17267 20009 17276 20043
rect 17224 20000 17276 20009
rect 18052 20000 18104 20052
rect 19156 20000 19208 20052
rect 10968 19932 11020 19984
rect 12808 19975 12860 19984
rect 12808 19941 12817 19975
rect 12817 19941 12851 19975
rect 12851 19941 12860 19975
rect 12808 19932 12860 19941
rect 13820 19975 13872 19984
rect 13820 19941 13829 19975
rect 13829 19941 13863 19975
rect 13863 19941 13872 19975
rect 13820 19932 13872 19941
rect 16304 19975 16356 19984
rect 16304 19941 16313 19975
rect 16313 19941 16347 19975
rect 16347 19941 16356 19975
rect 16304 19932 16356 19941
rect 17776 19975 17828 19984
rect 17776 19941 17785 19975
rect 17785 19941 17819 19975
rect 17819 19941 17828 19975
rect 17776 19932 17828 19941
rect 17868 19975 17920 19984
rect 17868 19941 17877 19975
rect 17877 19941 17911 19975
rect 17911 19941 17920 19975
rect 19340 19975 19392 19984
rect 17868 19932 17920 19941
rect 19340 19941 19349 19975
rect 19349 19941 19383 19975
rect 19383 19941 19392 19975
rect 19340 19932 19392 19941
rect 8576 19907 8628 19916
rect 8576 19873 8620 19907
rect 8620 19873 8628 19907
rect 8576 19864 8628 19873
rect 11980 19864 12032 19916
rect 12624 19907 12676 19916
rect 12624 19873 12633 19907
rect 12633 19873 12667 19907
rect 12667 19873 12676 19907
rect 12624 19864 12676 19873
rect 8208 19796 8260 19848
rect 9128 19839 9180 19848
rect 9128 19805 9137 19839
rect 9137 19805 9171 19839
rect 9171 19805 9180 19839
rect 9128 19796 9180 19805
rect 11336 19796 11388 19848
rect 12440 19796 12492 19848
rect 13268 19796 13320 19848
rect 16028 19796 16080 19848
rect 16580 19796 16632 19848
rect 18972 19796 19024 19848
rect 9404 19703 9456 19712
rect 9404 19669 9413 19703
rect 9413 19669 9447 19703
rect 9447 19669 9456 19703
rect 9404 19660 9456 19669
rect 10232 19703 10284 19712
rect 10232 19669 10241 19703
rect 10241 19669 10275 19703
rect 10275 19669 10284 19703
rect 10232 19660 10284 19669
rect 18236 19728 18288 19780
rect 14372 19660 14424 19712
rect 16212 19660 16264 19712
rect 18144 19660 18196 19712
rect 19248 19660 19300 19712
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 8116 19456 8168 19508
rect 10048 19499 10100 19508
rect 10048 19465 10057 19499
rect 10057 19465 10091 19499
rect 10091 19465 10100 19499
rect 10048 19456 10100 19465
rect 13820 19456 13872 19508
rect 16304 19456 16356 19508
rect 17868 19456 17920 19508
rect 19156 19456 19208 19508
rect 19616 19499 19668 19508
rect 19616 19465 19625 19499
rect 19625 19465 19659 19499
rect 19659 19465 19668 19499
rect 19616 19456 19668 19465
rect 6644 19388 6696 19440
rect 9220 19388 9272 19440
rect 7748 19320 7800 19372
rect 7840 19320 7892 19372
rect 8576 19363 8628 19372
rect 8576 19329 8585 19363
rect 8585 19329 8619 19363
rect 8619 19329 8628 19363
rect 8576 19320 8628 19329
rect 9404 19320 9456 19372
rect 12256 19320 12308 19372
rect 12532 19320 12584 19372
rect 13176 19363 13228 19372
rect 13176 19329 13185 19363
rect 13185 19329 13219 19363
rect 13219 19329 13228 19363
rect 13176 19320 13228 19329
rect 14372 19363 14424 19372
rect 14372 19329 14381 19363
rect 14381 19329 14415 19363
rect 14415 19329 14424 19363
rect 14372 19320 14424 19329
rect 14832 19363 14884 19372
rect 14832 19329 14841 19363
rect 14841 19329 14875 19363
rect 14875 19329 14884 19363
rect 14832 19320 14884 19329
rect 16212 19363 16264 19372
rect 16212 19329 16221 19363
rect 16221 19329 16255 19363
rect 16255 19329 16264 19363
rect 16212 19320 16264 19329
rect 7932 19295 7984 19304
rect 7932 19261 7941 19295
rect 7941 19261 7975 19295
rect 7975 19261 7984 19295
rect 7932 19252 7984 19261
rect 8944 19252 8996 19304
rect 10416 19295 10468 19304
rect 10416 19261 10425 19295
rect 10425 19261 10459 19295
rect 10459 19261 10468 19295
rect 10416 19252 10468 19261
rect 12716 19295 12768 19304
rect 12716 19261 12725 19295
rect 12725 19261 12759 19295
rect 12759 19261 12768 19295
rect 12716 19252 12768 19261
rect 12900 19252 12952 19304
rect 20260 19295 20312 19304
rect 9864 19116 9916 19168
rect 11152 19184 11204 19236
rect 11336 19227 11388 19236
rect 11336 19193 11345 19227
rect 11345 19193 11379 19227
rect 11379 19193 11388 19227
rect 11336 19184 11388 19193
rect 12164 19184 12216 19236
rect 12532 19184 12584 19236
rect 20260 19261 20269 19295
rect 20269 19261 20303 19295
rect 20303 19261 20312 19295
rect 20260 19252 20312 19261
rect 20812 19295 20864 19304
rect 20812 19261 20821 19295
rect 20821 19261 20855 19295
rect 20855 19261 20864 19295
rect 20812 19252 20864 19261
rect 14464 19227 14516 19236
rect 14464 19193 14473 19227
rect 14473 19193 14507 19227
rect 14507 19193 14516 19227
rect 14464 19184 14516 19193
rect 15936 19227 15988 19236
rect 15936 19193 15945 19227
rect 15945 19193 15979 19227
rect 15979 19193 15988 19227
rect 15936 19184 15988 19193
rect 18328 19227 18380 19236
rect 11060 19116 11112 19168
rect 11980 19116 12032 19168
rect 15844 19116 15896 19168
rect 18328 19193 18337 19227
rect 18337 19193 18371 19227
rect 18371 19193 18380 19227
rect 18328 19184 18380 19193
rect 18420 19227 18472 19236
rect 18420 19193 18429 19227
rect 18429 19193 18463 19227
rect 18463 19193 18472 19227
rect 18420 19184 18472 19193
rect 18696 19184 18748 19236
rect 18972 19227 19024 19236
rect 18972 19193 18981 19227
rect 18981 19193 19015 19227
rect 19015 19193 19024 19227
rect 18972 19184 19024 19193
rect 19340 19184 19392 19236
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 9404 18912 9456 18964
rect 11152 18955 11204 18964
rect 11152 18921 11161 18955
rect 11161 18921 11195 18955
rect 11195 18921 11204 18955
rect 11152 18912 11204 18921
rect 13268 18955 13320 18964
rect 13268 18921 13277 18955
rect 13277 18921 13311 18955
rect 13311 18921 13320 18955
rect 13268 18912 13320 18921
rect 14464 18912 14516 18964
rect 15844 18912 15896 18964
rect 16028 18912 16080 18964
rect 16580 18912 16632 18964
rect 9864 18844 9916 18896
rect 11888 18887 11940 18896
rect 11888 18853 11897 18887
rect 11897 18853 11931 18887
rect 11931 18853 11940 18887
rect 11888 18844 11940 18853
rect 13084 18844 13136 18896
rect 16856 18844 16908 18896
rect 17040 18844 17092 18896
rect 18420 18844 18472 18896
rect 19064 18844 19116 18896
rect 7748 18776 7800 18828
rect 8484 18776 8536 18828
rect 9956 18776 10008 18828
rect 15384 18819 15436 18828
rect 15384 18785 15393 18819
rect 15393 18785 15427 18819
rect 15427 18785 15436 18819
rect 15384 18776 15436 18785
rect 16212 18776 16264 18828
rect 16488 18776 16540 18828
rect 10048 18708 10100 18760
rect 11336 18708 11388 18760
rect 11796 18751 11848 18760
rect 11796 18717 11805 18751
rect 11805 18717 11839 18751
rect 11839 18717 11848 18751
rect 11796 18708 11848 18717
rect 12072 18751 12124 18760
rect 12072 18717 12081 18751
rect 12081 18717 12115 18751
rect 12115 18717 12124 18751
rect 12072 18708 12124 18717
rect 13452 18751 13504 18760
rect 13452 18717 13461 18751
rect 13461 18717 13495 18751
rect 13495 18717 13504 18751
rect 13452 18708 13504 18717
rect 17316 18708 17368 18760
rect 18972 18708 19024 18760
rect 19432 18708 19484 18760
rect 19340 18683 19392 18692
rect 19340 18649 19349 18683
rect 19349 18649 19383 18683
rect 19383 18649 19392 18683
rect 19340 18640 19392 18649
rect 8668 18572 8720 18624
rect 8760 18572 8812 18624
rect 9588 18572 9640 18624
rect 9956 18615 10008 18624
rect 9956 18581 9965 18615
rect 9965 18581 9999 18615
rect 9999 18581 10008 18615
rect 9956 18572 10008 18581
rect 11704 18572 11756 18624
rect 12716 18615 12768 18624
rect 12716 18581 12725 18615
rect 12725 18581 12759 18615
rect 12759 18581 12768 18615
rect 12716 18572 12768 18581
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 7840 18411 7892 18420
rect 7840 18377 7849 18411
rect 7849 18377 7883 18411
rect 7883 18377 7892 18411
rect 7840 18368 7892 18377
rect 9864 18368 9916 18420
rect 11888 18411 11940 18420
rect 11888 18377 11897 18411
rect 11897 18377 11931 18411
rect 11931 18377 11940 18411
rect 11888 18368 11940 18377
rect 17316 18411 17368 18420
rect 17316 18377 17325 18411
rect 17325 18377 17359 18411
rect 17359 18377 17368 18411
rect 17316 18368 17368 18377
rect 19064 18411 19116 18420
rect 19064 18377 19073 18411
rect 19073 18377 19107 18411
rect 19107 18377 19116 18411
rect 19064 18368 19116 18377
rect 19432 18411 19484 18420
rect 19432 18377 19441 18411
rect 19441 18377 19475 18411
rect 19475 18377 19484 18411
rect 19432 18368 19484 18377
rect 14280 18300 14332 18352
rect 9956 18232 10008 18284
rect 12164 18275 12216 18284
rect 12164 18241 12173 18275
rect 12173 18241 12207 18275
rect 12207 18241 12216 18275
rect 12164 18232 12216 18241
rect 12624 18232 12676 18284
rect 13452 18275 13504 18284
rect 1860 18164 1912 18216
rect 7012 18207 7064 18216
rect 7012 18173 7056 18207
rect 7056 18173 7064 18207
rect 7012 18164 7064 18173
rect 9312 18207 9364 18216
rect 9312 18173 9321 18207
rect 9321 18173 9355 18207
rect 9355 18173 9364 18207
rect 9312 18164 9364 18173
rect 9588 18207 9640 18216
rect 9588 18173 9597 18207
rect 9597 18173 9631 18207
rect 9631 18173 9640 18207
rect 9588 18164 9640 18173
rect 12992 18207 13044 18216
rect 12992 18173 13001 18207
rect 13001 18173 13035 18207
rect 13035 18173 13044 18207
rect 12992 18164 13044 18173
rect 13452 18241 13461 18275
rect 13461 18241 13495 18275
rect 13495 18241 13504 18275
rect 13452 18232 13504 18241
rect 14648 18232 14700 18284
rect 14832 18275 14884 18284
rect 14832 18241 14841 18275
rect 14841 18241 14875 18275
rect 14875 18241 14884 18275
rect 14832 18232 14884 18241
rect 18236 18232 18288 18284
rect 19340 18232 19392 18284
rect 19616 18207 19668 18216
rect 19616 18173 19660 18207
rect 19660 18173 19668 18207
rect 19616 18164 19668 18173
rect 20260 18164 20312 18216
rect 8208 18096 8260 18148
rect 15936 18139 15988 18148
rect 2320 18028 2372 18080
rect 7196 18028 7248 18080
rect 8484 18028 8536 18080
rect 10692 18028 10744 18080
rect 13084 18028 13136 18080
rect 14280 18028 14332 18080
rect 15936 18105 15945 18139
rect 15945 18105 15979 18139
rect 15979 18105 15988 18139
rect 15936 18096 15988 18105
rect 16028 18139 16080 18148
rect 16028 18105 16037 18139
rect 16037 18105 16071 18139
rect 16071 18105 16080 18139
rect 16028 18096 16080 18105
rect 15384 18071 15436 18080
rect 15384 18037 15393 18071
rect 15393 18037 15427 18071
rect 15427 18037 15436 18071
rect 15384 18028 15436 18037
rect 16856 18028 16908 18080
rect 17776 18071 17828 18080
rect 17776 18037 17785 18071
rect 17785 18037 17819 18071
rect 17819 18037 17828 18071
rect 17776 18028 17828 18037
rect 19984 18028 20036 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 9312 17824 9364 17876
rect 10048 17824 10100 17876
rect 11060 17824 11112 17876
rect 1676 17756 1728 17808
rect 2688 17756 2740 17808
rect 7564 17799 7616 17808
rect 7564 17765 7573 17799
rect 7573 17765 7607 17799
rect 7607 17765 7616 17799
rect 7564 17756 7616 17765
rect 7840 17756 7892 17808
rect 12992 17824 13044 17876
rect 13452 17824 13504 17876
rect 14280 17824 14332 17876
rect 14648 17867 14700 17876
rect 14648 17833 14657 17867
rect 14657 17833 14691 17867
rect 14691 17833 14700 17867
rect 14648 17824 14700 17833
rect 15936 17824 15988 17876
rect 17776 17824 17828 17876
rect 18236 17824 18288 17876
rect 18328 17824 18380 17876
rect 11520 17756 11572 17808
rect 12072 17756 12124 17808
rect 13084 17756 13136 17808
rect 16856 17756 16908 17808
rect 2228 17688 2280 17740
rect 5448 17731 5500 17740
rect 5448 17697 5457 17731
rect 5457 17697 5491 17731
rect 5491 17697 5500 17731
rect 5448 17688 5500 17697
rect 6552 17731 6604 17740
rect 6552 17697 6570 17731
rect 6570 17697 6604 17731
rect 6552 17688 6604 17697
rect 6736 17688 6788 17740
rect 9956 17688 10008 17740
rect 15292 17731 15344 17740
rect 15292 17697 15336 17731
rect 15336 17697 15344 17731
rect 15292 17688 15344 17697
rect 8024 17663 8076 17672
rect 8024 17629 8033 17663
rect 8033 17629 8067 17663
rect 8067 17629 8076 17663
rect 8024 17620 8076 17629
rect 11796 17620 11848 17672
rect 13452 17663 13504 17672
rect 13452 17629 13461 17663
rect 13461 17629 13495 17663
rect 13495 17629 13504 17663
rect 13452 17620 13504 17629
rect 16764 17663 16816 17672
rect 16764 17629 16773 17663
rect 16773 17629 16807 17663
rect 16807 17629 16816 17663
rect 16764 17620 16816 17629
rect 16212 17552 16264 17604
rect 2136 17484 2188 17536
rect 2688 17527 2740 17536
rect 2688 17493 2697 17527
rect 2697 17493 2731 17527
rect 2731 17493 2740 17527
rect 2688 17484 2740 17493
rect 6184 17484 6236 17536
rect 6368 17484 6420 17536
rect 10140 17484 10192 17536
rect 10968 17484 11020 17536
rect 16304 17527 16356 17536
rect 16304 17493 16313 17527
rect 16313 17493 16347 17527
rect 16347 17493 16356 17527
rect 16304 17484 16356 17493
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 1676 17323 1728 17332
rect 1676 17289 1685 17323
rect 1685 17289 1719 17323
rect 1719 17289 1728 17323
rect 1676 17280 1728 17289
rect 2688 17323 2740 17332
rect 2688 17289 2697 17323
rect 2697 17289 2731 17323
rect 2731 17289 2740 17323
rect 2688 17280 2740 17289
rect 6276 17323 6328 17332
rect 6276 17289 6285 17323
rect 6285 17289 6319 17323
rect 6319 17289 6328 17323
rect 6276 17280 6328 17289
rect 11520 17323 11572 17332
rect 11520 17289 11529 17323
rect 11529 17289 11563 17323
rect 11563 17289 11572 17323
rect 11520 17280 11572 17289
rect 12624 17323 12676 17332
rect 12624 17289 12633 17323
rect 12633 17289 12667 17323
rect 12667 17289 12676 17323
rect 12624 17280 12676 17289
rect 14464 17323 14516 17332
rect 14464 17289 14473 17323
rect 14473 17289 14507 17323
rect 14507 17289 14516 17323
rect 14464 17280 14516 17289
rect 8024 17255 8076 17264
rect 8024 17221 8033 17255
rect 8033 17221 8067 17255
rect 8067 17221 8076 17255
rect 8024 17212 8076 17221
rect 2872 17187 2924 17196
rect 2872 17153 2881 17187
rect 2881 17153 2915 17187
rect 2915 17153 2924 17187
rect 2872 17144 2924 17153
rect 3056 17144 3108 17196
rect 5448 17144 5500 17196
rect 6644 17144 6696 17196
rect 7840 17144 7892 17196
rect 10968 17144 11020 17196
rect 13452 17144 13504 17196
rect 15292 17187 15344 17196
rect 15292 17153 15301 17187
rect 15301 17153 15335 17187
rect 15335 17153 15344 17187
rect 15292 17144 15344 17153
rect 18236 17144 18288 17196
rect 6276 17076 6328 17128
rect 2688 17008 2740 17060
rect 7472 17051 7524 17060
rect 1768 16983 1820 16992
rect 1768 16949 1777 16983
rect 1777 16949 1811 16983
rect 1811 16949 1820 16983
rect 1768 16940 1820 16949
rect 2228 16983 2280 16992
rect 2228 16949 2237 16983
rect 2237 16949 2271 16983
rect 2271 16949 2280 16983
rect 2228 16940 2280 16949
rect 7472 17017 7481 17051
rect 7481 17017 7515 17051
rect 7515 17017 7524 17051
rect 7472 17008 7524 17017
rect 4160 16940 4212 16992
rect 6736 16940 6788 16992
rect 7840 16940 7892 16992
rect 13360 17076 13412 17128
rect 13544 17119 13596 17128
rect 13544 17085 13553 17119
rect 13553 17085 13587 17119
rect 13587 17085 13596 17119
rect 13544 17076 13596 17085
rect 16304 17076 16356 17128
rect 10692 17008 10744 17060
rect 9956 16940 10008 16992
rect 13084 16983 13136 16992
rect 13084 16949 13093 16983
rect 13093 16949 13127 16983
rect 13127 16949 13136 16983
rect 13084 16940 13136 16949
rect 13360 16940 13412 16992
rect 18144 17051 18196 17060
rect 18144 17017 18153 17051
rect 18153 17017 18187 17051
rect 18187 17017 18196 17051
rect 18144 17008 18196 17017
rect 16856 16940 16908 16992
rect 18420 17008 18472 17060
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 2872 16736 2924 16788
rect 7840 16779 7892 16788
rect 7840 16745 7849 16779
rect 7849 16745 7883 16779
rect 7883 16745 7892 16779
rect 7840 16736 7892 16745
rect 11060 16736 11112 16788
rect 12624 16779 12676 16788
rect 12624 16745 12633 16779
rect 12633 16745 12667 16779
rect 12667 16745 12676 16779
rect 12624 16736 12676 16745
rect 18144 16779 18196 16788
rect 18144 16745 18153 16779
rect 18153 16745 18187 16779
rect 18187 16745 18196 16779
rect 18144 16736 18196 16745
rect 2136 16711 2188 16720
rect 2136 16677 2145 16711
rect 2145 16677 2179 16711
rect 2179 16677 2188 16711
rect 2136 16668 2188 16677
rect 2228 16711 2280 16720
rect 2228 16677 2237 16711
rect 2237 16677 2271 16711
rect 2271 16677 2280 16711
rect 2228 16668 2280 16677
rect 4160 16668 4212 16720
rect 7012 16668 7064 16720
rect 7472 16668 7524 16720
rect 10692 16668 10744 16720
rect 13084 16668 13136 16720
rect 6920 16643 6972 16652
rect 6920 16609 6929 16643
rect 6929 16609 6963 16643
rect 6963 16609 6972 16643
rect 6920 16600 6972 16609
rect 4252 16532 4304 16584
rect 4344 16532 4396 16584
rect 6460 16532 6512 16584
rect 10692 16532 10744 16584
rect 10876 16532 10928 16584
rect 11152 16600 11204 16652
rect 13544 16668 13596 16720
rect 16764 16711 16816 16720
rect 16764 16677 16773 16711
rect 16773 16677 16807 16711
rect 16807 16677 16816 16711
rect 16764 16668 16816 16677
rect 17960 16668 18012 16720
rect 14372 16643 14424 16652
rect 14372 16609 14381 16643
rect 14381 16609 14415 16643
rect 14415 16609 14424 16643
rect 14372 16600 14424 16609
rect 15660 16600 15712 16652
rect 16212 16643 16264 16652
rect 16212 16609 16221 16643
rect 16221 16609 16255 16643
rect 16255 16609 16264 16643
rect 16212 16600 16264 16609
rect 17316 16643 17368 16652
rect 17316 16609 17360 16643
rect 17360 16609 17368 16643
rect 17316 16600 17368 16609
rect 18328 16643 18380 16652
rect 18328 16609 18372 16643
rect 18372 16609 18380 16643
rect 18328 16600 18380 16609
rect 13636 16532 13688 16584
rect 2872 16464 2924 16516
rect 4436 16396 4488 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2228 16192 2280 16244
rect 4160 16235 4212 16244
rect 4160 16201 4169 16235
rect 4169 16201 4203 16235
rect 4203 16201 4212 16235
rect 4160 16192 4212 16201
rect 4252 16192 4304 16244
rect 8024 16235 8076 16244
rect 8024 16201 8033 16235
rect 8033 16201 8067 16235
rect 8067 16201 8076 16235
rect 8024 16192 8076 16201
rect 10600 16192 10652 16244
rect 18328 16192 18380 16244
rect 2780 16124 2832 16176
rect 3148 16099 3200 16108
rect 3148 16065 3157 16099
rect 3157 16065 3191 16099
rect 3191 16065 3200 16099
rect 3148 16056 3200 16065
rect 4436 16099 4488 16108
rect 4436 16065 4445 16099
rect 4445 16065 4479 16099
rect 4479 16065 4488 16099
rect 4436 16056 4488 16065
rect 4712 16099 4764 16108
rect 4712 16065 4721 16099
rect 4721 16065 4755 16099
rect 4755 16065 4764 16099
rect 4712 16056 4764 16065
rect 11060 16124 11112 16176
rect 11612 16124 11664 16176
rect 12716 16124 12768 16176
rect 15660 16124 15712 16176
rect 10140 16056 10192 16108
rect 13452 16056 13504 16108
rect 14372 16056 14424 16108
rect 14556 16099 14608 16108
rect 14556 16065 14565 16099
rect 14565 16065 14599 16099
rect 14599 16065 14608 16099
rect 14556 16056 14608 16065
rect 16304 16099 16356 16108
rect 16304 16065 16313 16099
rect 16313 16065 16347 16099
rect 16347 16065 16356 16099
rect 16304 16056 16356 16065
rect 17316 16099 17368 16108
rect 17316 16065 17325 16099
rect 17325 16065 17359 16099
rect 17359 16065 17368 16099
rect 17316 16056 17368 16065
rect 1584 15988 1636 16040
rect 1768 16031 1820 16040
rect 1768 15997 1812 16031
rect 1812 15997 1820 16031
rect 1768 15988 1820 15997
rect 8852 16031 8904 16040
rect 8852 15997 8861 16031
rect 8861 15997 8895 16031
rect 8895 15997 8904 16031
rect 8852 15988 8904 15997
rect 12716 16031 12768 16040
rect 12716 15997 12725 16031
rect 12725 15997 12759 16031
rect 12759 15997 12768 16031
rect 13084 16031 13136 16040
rect 12716 15988 12768 15997
rect 13084 15997 13093 16031
rect 13093 15997 13127 16031
rect 13127 15997 13136 16031
rect 13084 15988 13136 15997
rect 15752 16031 15804 16040
rect 15752 15997 15761 16031
rect 15761 15997 15795 16031
rect 15795 15997 15804 16031
rect 15752 15988 15804 15997
rect 16212 16031 16264 16040
rect 16212 15997 16221 16031
rect 16221 15997 16255 16031
rect 16255 15997 16264 16031
rect 16212 15988 16264 15997
rect 18052 16031 18104 16040
rect 18052 15997 18096 16031
rect 18096 15997 18104 16031
rect 18052 15988 18104 15997
rect 18604 15988 18656 16040
rect 2872 15963 2924 15972
rect 2872 15929 2881 15963
rect 2881 15929 2915 15963
rect 2915 15929 2924 15963
rect 2872 15920 2924 15929
rect 3240 15920 3292 15972
rect 4160 15920 4212 15972
rect 5080 15920 5132 15972
rect 6828 15920 6880 15972
rect 6092 15852 6144 15904
rect 7012 15920 7064 15972
rect 7104 15963 7156 15972
rect 7104 15929 7113 15963
rect 7113 15929 7147 15963
rect 7147 15929 7156 15963
rect 7104 15920 7156 15929
rect 7288 15920 7340 15972
rect 9496 15963 9548 15972
rect 9496 15929 9505 15963
rect 9505 15929 9539 15963
rect 9539 15929 9548 15963
rect 9496 15920 9548 15929
rect 10876 15920 10928 15972
rect 13636 15895 13688 15904
rect 13636 15861 13645 15895
rect 13645 15861 13679 15895
rect 13679 15861 13688 15895
rect 13636 15852 13688 15861
rect 14004 15895 14056 15904
rect 14004 15861 14013 15895
rect 14013 15861 14047 15895
rect 14047 15861 14056 15895
rect 15292 15895 15344 15904
rect 14004 15852 14056 15861
rect 15292 15861 15301 15895
rect 15301 15861 15335 15895
rect 15335 15861 15344 15895
rect 15292 15852 15344 15861
rect 15660 15895 15712 15904
rect 15660 15861 15669 15895
rect 15669 15861 15703 15895
rect 15703 15861 15712 15895
rect 15660 15852 15712 15861
rect 18144 15852 18196 15904
rect 18972 15852 19024 15904
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 2136 15691 2188 15700
rect 2136 15657 2145 15691
rect 2145 15657 2179 15691
rect 2179 15657 2188 15691
rect 2136 15648 2188 15657
rect 2872 15648 2924 15700
rect 4344 15648 4396 15700
rect 5080 15691 5132 15700
rect 5080 15657 5089 15691
rect 5089 15657 5123 15691
rect 5123 15657 5132 15691
rect 5080 15648 5132 15657
rect 10692 15691 10744 15700
rect 10692 15657 10701 15691
rect 10701 15657 10735 15691
rect 10735 15657 10744 15691
rect 10692 15648 10744 15657
rect 13084 15648 13136 15700
rect 15752 15691 15804 15700
rect 15752 15657 15761 15691
rect 15761 15657 15795 15691
rect 15795 15657 15804 15691
rect 15752 15648 15804 15657
rect 16028 15648 16080 15700
rect 2504 15623 2556 15632
rect 2504 15589 2513 15623
rect 2513 15589 2547 15623
rect 2547 15589 2556 15623
rect 2504 15580 2556 15589
rect 2596 15623 2648 15632
rect 2596 15589 2605 15623
rect 2605 15589 2639 15623
rect 2639 15589 2648 15623
rect 3148 15623 3200 15632
rect 2596 15580 2648 15589
rect 3148 15589 3157 15623
rect 3157 15589 3191 15623
rect 3191 15589 3200 15623
rect 3148 15580 3200 15589
rect 3240 15580 3292 15632
rect 6460 15623 6512 15632
rect 6460 15589 6469 15623
rect 6469 15589 6503 15623
rect 6503 15589 6512 15623
rect 6460 15580 6512 15589
rect 6552 15623 6604 15632
rect 6552 15589 6561 15623
rect 6561 15589 6595 15623
rect 6595 15589 6604 15623
rect 6552 15580 6604 15589
rect 9496 15580 9548 15632
rect 9772 15580 9824 15632
rect 13820 15623 13872 15632
rect 13820 15589 13829 15623
rect 13829 15589 13863 15623
rect 13863 15589 13872 15623
rect 13820 15580 13872 15589
rect 14556 15580 14608 15632
rect 16856 15580 16908 15632
rect 4160 15555 4212 15564
rect 4160 15521 4169 15555
rect 4169 15521 4203 15555
rect 4203 15521 4212 15555
rect 4160 15512 4212 15521
rect 7104 15512 7156 15564
rect 7840 15512 7892 15564
rect 11244 15555 11296 15564
rect 11244 15521 11253 15555
rect 11253 15521 11287 15555
rect 11287 15521 11296 15555
rect 11244 15512 11296 15521
rect 11796 15555 11848 15564
rect 11796 15521 11805 15555
rect 11805 15521 11839 15555
rect 11839 15521 11848 15555
rect 11796 15512 11848 15521
rect 17500 15580 17552 15632
rect 8944 15444 8996 15496
rect 9404 15444 9456 15496
rect 10048 15487 10100 15496
rect 10048 15453 10057 15487
rect 10057 15453 10091 15487
rect 10091 15453 10100 15487
rect 10048 15444 10100 15453
rect 13728 15487 13780 15496
rect 13728 15453 13737 15487
rect 13737 15453 13771 15487
rect 13771 15453 13780 15487
rect 13728 15444 13780 15453
rect 16488 15444 16540 15496
rect 18052 15487 18104 15496
rect 18052 15453 18061 15487
rect 18061 15453 18095 15487
rect 18095 15453 18104 15487
rect 18052 15444 18104 15453
rect 2044 15376 2096 15428
rect 3148 15376 3200 15428
rect 7288 15376 7340 15428
rect 17960 15376 18012 15428
rect 2412 15308 2464 15360
rect 8116 15308 8168 15360
rect 13176 15308 13228 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2596 15104 2648 15156
rect 4160 15147 4212 15156
rect 4160 15113 4169 15147
rect 4169 15113 4203 15147
rect 4203 15113 4212 15147
rect 4160 15104 4212 15113
rect 6552 15104 6604 15156
rect 7840 15104 7892 15156
rect 8852 15104 8904 15156
rect 9772 15147 9824 15156
rect 2780 15036 2832 15088
rect 4068 15036 4120 15088
rect 9772 15113 9781 15147
rect 9781 15113 9815 15147
rect 9815 15113 9824 15147
rect 9772 15104 9824 15113
rect 11796 15147 11848 15156
rect 11796 15113 11805 15147
rect 11805 15113 11839 15147
rect 11839 15113 11848 15147
rect 11796 15104 11848 15113
rect 13360 15104 13412 15156
rect 14648 15147 14700 15156
rect 14648 15113 14657 15147
rect 14657 15113 14691 15147
rect 14691 15113 14700 15147
rect 14648 15104 14700 15113
rect 15292 15147 15344 15156
rect 15292 15113 15301 15147
rect 15301 15113 15335 15147
rect 15335 15113 15344 15147
rect 15292 15104 15344 15113
rect 17500 15147 17552 15156
rect 17500 15113 17509 15147
rect 17509 15113 17543 15147
rect 17543 15113 17552 15147
rect 17500 15104 17552 15113
rect 18052 15104 18104 15156
rect 10508 15036 10560 15088
rect 13820 15036 13872 15088
rect 15476 15036 15528 15088
rect 2964 14968 3016 15020
rect 3976 14968 4028 15020
rect 5264 14968 5316 15020
rect 6092 14968 6144 15020
rect 3056 14900 3108 14952
rect 5356 14875 5408 14884
rect 5356 14841 5365 14875
rect 5365 14841 5399 14875
rect 5399 14841 5408 14875
rect 5356 14832 5408 14841
rect 6000 14832 6052 14884
rect 7104 14968 7156 15020
rect 10048 14968 10100 15020
rect 18144 15011 18196 15020
rect 18144 14977 18153 15011
rect 18153 14977 18187 15011
rect 18187 14977 18196 15011
rect 18144 14968 18196 14977
rect 9588 14900 9640 14952
rect 13176 14900 13228 14952
rect 8484 14832 8536 14884
rect 10416 14875 10468 14884
rect 10416 14841 10425 14875
rect 10425 14841 10459 14875
rect 10459 14841 10468 14875
rect 10416 14832 10468 14841
rect 10508 14875 10560 14884
rect 10508 14841 10517 14875
rect 10517 14841 10551 14875
rect 10551 14841 10560 14875
rect 10508 14832 10560 14841
rect 13452 14832 13504 14884
rect 1400 14764 1452 14816
rect 2688 14764 2740 14816
rect 2872 14764 2924 14816
rect 4620 14807 4672 14816
rect 4620 14773 4629 14807
rect 4629 14773 4663 14807
rect 4663 14773 4672 14807
rect 4620 14764 4672 14773
rect 10692 14764 10744 14816
rect 10784 14764 10836 14816
rect 11244 14764 11296 14816
rect 14832 14764 14884 14816
rect 16212 14943 16264 14952
rect 16212 14909 16221 14943
rect 16221 14909 16255 14943
rect 16255 14909 16264 14943
rect 16212 14900 16264 14909
rect 16856 14832 16908 14884
rect 17316 14764 17368 14816
rect 18788 14875 18840 14884
rect 18788 14841 18797 14875
rect 18797 14841 18831 14875
rect 18831 14841 18840 14875
rect 18788 14832 18840 14841
rect 19340 14764 19392 14816
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2044 14603 2096 14612
rect 2044 14569 2053 14603
rect 2053 14569 2087 14603
rect 2087 14569 2096 14603
rect 2044 14560 2096 14569
rect 2504 14603 2556 14612
rect 2504 14569 2513 14603
rect 2513 14569 2547 14603
rect 2547 14569 2556 14603
rect 2504 14560 2556 14569
rect 2688 14560 2740 14612
rect 6460 14560 6512 14612
rect 7840 14603 7892 14612
rect 7840 14569 7849 14603
rect 7849 14569 7883 14603
rect 7883 14569 7892 14603
rect 7840 14560 7892 14569
rect 9404 14603 9456 14612
rect 9404 14569 9413 14603
rect 9413 14569 9447 14603
rect 9447 14569 9456 14603
rect 9404 14560 9456 14569
rect 10692 14603 10744 14612
rect 10692 14569 10701 14603
rect 10701 14569 10735 14603
rect 10735 14569 10744 14603
rect 10692 14560 10744 14569
rect 16212 14560 16264 14612
rect 2964 14492 3016 14544
rect 6276 14492 6328 14544
rect 8116 14535 8168 14544
rect 8116 14501 8125 14535
rect 8125 14501 8159 14535
rect 8159 14501 8168 14535
rect 8116 14492 8168 14501
rect 8208 14535 8260 14544
rect 8208 14501 8217 14535
rect 8217 14501 8251 14535
rect 8251 14501 8260 14535
rect 8208 14492 8260 14501
rect 9956 14492 10008 14544
rect 13360 14535 13412 14544
rect 13360 14501 13363 14535
rect 13363 14501 13397 14535
rect 13397 14501 13412 14535
rect 13360 14492 13412 14501
rect 15476 14535 15528 14544
rect 15476 14501 15485 14535
rect 15485 14501 15519 14535
rect 15519 14501 15528 14535
rect 15476 14492 15528 14501
rect 17316 14535 17368 14544
rect 17316 14501 17325 14535
rect 17325 14501 17359 14535
rect 17359 14501 17368 14535
rect 17316 14492 17368 14501
rect 18144 14560 18196 14612
rect 2044 14424 2096 14476
rect 4528 14467 4580 14476
rect 4528 14433 4537 14467
rect 4537 14433 4571 14467
rect 4571 14433 4580 14467
rect 4528 14424 4580 14433
rect 11704 14467 11756 14476
rect 11704 14433 11713 14467
rect 11713 14433 11747 14467
rect 11747 14433 11756 14467
rect 11704 14424 11756 14433
rect 1952 14356 2004 14408
rect 2964 14399 3016 14408
rect 2964 14365 2973 14399
rect 2973 14365 3007 14399
rect 3007 14365 3016 14399
rect 2964 14356 3016 14365
rect 6000 14399 6052 14408
rect 6000 14365 6009 14399
rect 6009 14365 6043 14399
rect 6043 14365 6052 14399
rect 6000 14356 6052 14365
rect 8392 14399 8444 14408
rect 8392 14365 8401 14399
rect 8401 14365 8435 14399
rect 8435 14365 8444 14399
rect 8392 14356 8444 14365
rect 9772 14399 9824 14408
rect 9772 14365 9781 14399
rect 9781 14365 9815 14399
rect 9815 14365 9824 14399
rect 9772 14356 9824 14365
rect 11428 14356 11480 14408
rect 12900 14424 12952 14476
rect 18052 14424 18104 14476
rect 19248 14467 19300 14476
rect 12992 14399 13044 14408
rect 12992 14365 13001 14399
rect 13001 14365 13035 14399
rect 13035 14365 13044 14399
rect 12992 14356 13044 14365
rect 15752 14356 15804 14408
rect 16304 14356 16356 14408
rect 17224 14399 17276 14408
rect 17224 14365 17233 14399
rect 17233 14365 17267 14399
rect 17267 14365 17276 14399
rect 17224 14356 17276 14365
rect 17592 14356 17644 14408
rect 19248 14433 19257 14467
rect 19257 14433 19291 14467
rect 19291 14433 19300 14467
rect 19248 14424 19300 14433
rect 19064 14356 19116 14408
rect 4712 14263 4764 14272
rect 4712 14229 4721 14263
rect 4721 14229 4755 14263
rect 4755 14229 4764 14263
rect 4712 14220 4764 14229
rect 5080 14263 5132 14272
rect 5080 14229 5089 14263
rect 5089 14229 5123 14263
rect 5123 14229 5132 14263
rect 5080 14220 5132 14229
rect 5540 14220 5592 14272
rect 6920 14263 6972 14272
rect 6920 14229 6929 14263
rect 6929 14229 6963 14263
rect 6963 14229 6972 14263
rect 6920 14220 6972 14229
rect 7104 14220 7156 14272
rect 9036 14263 9088 14272
rect 9036 14229 9045 14263
rect 9045 14229 9079 14263
rect 9079 14229 9088 14263
rect 9036 14220 9088 14229
rect 12900 14220 12952 14272
rect 14004 14220 14056 14272
rect 14188 14263 14240 14272
rect 14188 14229 14197 14263
rect 14197 14229 14231 14263
rect 14231 14229 14240 14263
rect 14188 14220 14240 14229
rect 16580 14220 16632 14272
rect 18328 14220 18380 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 4160 14016 4212 14068
rect 5356 14016 5408 14068
rect 6920 14016 6972 14068
rect 8484 14059 8536 14068
rect 8484 14025 8493 14059
rect 8493 14025 8527 14059
rect 8527 14025 8536 14059
rect 8484 14016 8536 14025
rect 9772 14016 9824 14068
rect 13360 14016 13412 14068
rect 14004 14059 14056 14068
rect 14004 14025 14013 14059
rect 14013 14025 14047 14059
rect 14047 14025 14056 14059
rect 14004 14016 14056 14025
rect 17316 14016 17368 14068
rect 19064 14059 19116 14068
rect 1584 13991 1636 14000
rect 1584 13957 1593 13991
rect 1593 13957 1627 13991
rect 1627 13957 1636 13991
rect 1584 13948 1636 13957
rect 6276 13991 6328 14000
rect 6276 13957 6285 13991
rect 6285 13957 6319 13991
rect 6319 13957 6328 13991
rect 6276 13948 6328 13957
rect 10600 13991 10652 14000
rect 10600 13957 10609 13991
rect 10609 13957 10643 13991
rect 10643 13957 10652 13991
rect 10600 13948 10652 13957
rect 15476 13948 15528 14000
rect 16764 13948 16816 14000
rect 17224 13948 17276 14000
rect 8668 13923 8720 13932
rect 8668 13889 8677 13923
rect 8677 13889 8711 13923
rect 8711 13889 8720 13923
rect 8668 13880 8720 13889
rect 9036 13880 9088 13932
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 2044 13855 2096 13864
rect 2044 13821 2053 13855
rect 2053 13821 2087 13855
rect 2087 13821 2096 13855
rect 2044 13812 2096 13821
rect 4068 13812 4120 13864
rect 4528 13855 4580 13864
rect 4528 13821 4537 13855
rect 4537 13821 4571 13855
rect 4571 13821 4580 13855
rect 4528 13812 4580 13821
rect 5080 13812 5132 13864
rect 5264 13744 5316 13796
rect 6920 13855 6972 13864
rect 6920 13821 6929 13855
rect 6929 13821 6963 13855
rect 6963 13821 6972 13855
rect 6920 13812 6972 13821
rect 8208 13812 8260 13864
rect 10968 13880 11020 13932
rect 13176 13923 13228 13932
rect 10784 13855 10836 13864
rect 5724 13744 5776 13796
rect 8484 13744 8536 13796
rect 2872 13719 2924 13728
rect 2872 13685 2881 13719
rect 2881 13685 2915 13719
rect 2915 13685 2924 13719
rect 2872 13676 2924 13685
rect 6828 13676 6880 13728
rect 10784 13821 10793 13855
rect 10793 13821 10827 13855
rect 10827 13821 10836 13855
rect 10784 13812 10836 13821
rect 10876 13812 10928 13864
rect 11612 13812 11664 13864
rect 11980 13812 12032 13864
rect 12900 13855 12952 13864
rect 12900 13821 12909 13855
rect 12909 13821 12943 13855
rect 12943 13821 12952 13855
rect 12900 13812 12952 13821
rect 13176 13889 13185 13923
rect 13185 13889 13219 13923
rect 13219 13889 13228 13923
rect 13176 13880 13228 13889
rect 14188 13923 14240 13932
rect 14188 13889 14197 13923
rect 14197 13889 14231 13923
rect 14231 13889 14240 13923
rect 14188 13880 14240 13889
rect 15752 13923 15804 13932
rect 15752 13889 15761 13923
rect 15761 13889 15795 13923
rect 15795 13889 15804 13923
rect 15752 13880 15804 13889
rect 16580 13880 16632 13932
rect 17132 13923 17184 13932
rect 17132 13889 17141 13923
rect 17141 13889 17175 13923
rect 17175 13889 17184 13923
rect 17132 13880 17184 13889
rect 17684 13880 17736 13932
rect 13728 13812 13780 13864
rect 14004 13812 14056 13864
rect 15108 13812 15160 13864
rect 19064 14025 19073 14059
rect 19073 14025 19107 14059
rect 19107 14025 19116 14059
rect 19064 14016 19116 14025
rect 19248 14016 19300 14068
rect 18328 13880 18380 13932
rect 18420 13923 18472 13932
rect 18420 13889 18429 13923
rect 18429 13889 18463 13923
rect 18463 13889 18472 13923
rect 18420 13880 18472 13889
rect 19340 13880 19392 13932
rect 16304 13744 16356 13796
rect 16580 13787 16632 13796
rect 16580 13753 16589 13787
rect 16589 13753 16623 13787
rect 16623 13753 16632 13787
rect 19432 13812 19484 13864
rect 16580 13744 16632 13753
rect 18144 13744 18196 13796
rect 9772 13676 9824 13728
rect 9956 13719 10008 13728
rect 9956 13685 9965 13719
rect 9965 13685 9999 13719
rect 9999 13685 10008 13719
rect 9956 13676 10008 13685
rect 11704 13676 11756 13728
rect 12624 13676 12676 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 5724 13515 5776 13524
rect 5724 13481 5733 13515
rect 5733 13481 5767 13515
rect 5767 13481 5776 13515
rect 5724 13472 5776 13481
rect 8484 13515 8536 13524
rect 8484 13481 8493 13515
rect 8493 13481 8527 13515
rect 8527 13481 8536 13515
rect 8484 13472 8536 13481
rect 9956 13515 10008 13524
rect 9956 13481 9965 13515
rect 9965 13481 9999 13515
rect 9999 13481 10008 13515
rect 9956 13472 10008 13481
rect 10876 13515 10928 13524
rect 10876 13481 10885 13515
rect 10885 13481 10919 13515
rect 10919 13481 10928 13515
rect 10876 13472 10928 13481
rect 12992 13515 13044 13524
rect 12992 13481 13001 13515
rect 13001 13481 13035 13515
rect 13035 13481 13044 13515
rect 12992 13472 13044 13481
rect 15108 13515 15160 13524
rect 15108 13481 15117 13515
rect 15117 13481 15151 13515
rect 15151 13481 15160 13515
rect 15108 13472 15160 13481
rect 15200 13472 15252 13524
rect 16304 13472 16356 13524
rect 16580 13472 16632 13524
rect 18144 13515 18196 13524
rect 18144 13481 18153 13515
rect 18153 13481 18187 13515
rect 18187 13481 18196 13515
rect 18144 13472 18196 13481
rect 19340 13472 19392 13524
rect 2688 13404 2740 13456
rect 4252 13447 4304 13456
rect 4252 13413 4261 13447
rect 4261 13413 4295 13447
rect 4295 13413 4304 13447
rect 4252 13404 4304 13413
rect 6184 13379 6236 13388
rect 2044 13268 2096 13320
rect 4344 13268 4396 13320
rect 6184 13345 6193 13379
rect 6193 13345 6227 13379
rect 6227 13345 6236 13379
rect 6184 13336 6236 13345
rect 6368 13336 6420 13388
rect 9036 13404 9088 13456
rect 12900 13404 12952 13456
rect 7472 13336 7524 13388
rect 8760 13336 8812 13388
rect 9772 13336 9824 13388
rect 10876 13336 10928 13388
rect 11704 13379 11756 13388
rect 11704 13345 11713 13379
rect 11713 13345 11747 13379
rect 11747 13345 11756 13379
rect 11704 13336 11756 13345
rect 13636 13379 13688 13388
rect 13636 13345 13645 13379
rect 13645 13345 13679 13379
rect 13679 13345 13688 13379
rect 13636 13336 13688 13345
rect 15200 13336 15252 13388
rect 16856 13447 16908 13456
rect 16856 13413 16859 13447
rect 16859 13413 16893 13447
rect 16893 13413 16908 13447
rect 16856 13404 16908 13413
rect 18052 13404 18104 13456
rect 19064 13404 19116 13456
rect 1492 13132 1544 13184
rect 6092 13268 6144 13320
rect 11428 13311 11480 13320
rect 11428 13277 11437 13311
rect 11437 13277 11471 13311
rect 11471 13277 11480 13311
rect 11428 13268 11480 13277
rect 12440 13268 12492 13320
rect 16672 13336 16724 13388
rect 16580 13268 16632 13320
rect 19800 13379 19852 13388
rect 19800 13345 19844 13379
rect 19844 13345 19852 13379
rect 19800 13336 19852 13345
rect 18604 13268 18656 13320
rect 18788 13311 18840 13320
rect 18788 13277 18797 13311
rect 18797 13277 18831 13311
rect 18831 13277 18840 13311
rect 18788 13268 18840 13277
rect 16856 13200 16908 13252
rect 2228 13175 2280 13184
rect 2228 13141 2237 13175
rect 2237 13141 2271 13175
rect 2271 13141 2280 13175
rect 2228 13132 2280 13141
rect 3516 13175 3568 13184
rect 3516 13141 3525 13175
rect 3525 13141 3559 13175
rect 3559 13141 3568 13175
rect 3516 13132 3568 13141
rect 7380 13175 7432 13184
rect 7380 13141 7389 13175
rect 7389 13141 7423 13175
rect 7423 13141 7432 13175
rect 7380 13132 7432 13141
rect 7932 13132 7984 13184
rect 10140 13132 10192 13184
rect 15660 13132 15712 13184
rect 17776 13175 17828 13184
rect 17776 13141 17785 13175
rect 17785 13141 17819 13175
rect 17819 13141 17828 13175
rect 17776 13132 17828 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2044 12971 2096 12980
rect 2044 12937 2053 12971
rect 2053 12937 2087 12971
rect 2087 12937 2096 12971
rect 2044 12928 2096 12937
rect 3884 12971 3936 12980
rect 3884 12937 3893 12971
rect 3893 12937 3927 12971
rect 3927 12937 3936 12971
rect 4252 12971 4304 12980
rect 3884 12928 3936 12937
rect 4252 12937 4261 12971
rect 4261 12937 4295 12971
rect 4295 12937 4304 12971
rect 4252 12928 4304 12937
rect 4896 12971 4948 12980
rect 4896 12937 4905 12971
rect 4905 12937 4939 12971
rect 4939 12937 4948 12971
rect 4896 12928 4948 12937
rect 8760 12928 8812 12980
rect 9036 12971 9088 12980
rect 9036 12937 9045 12971
rect 9045 12937 9079 12971
rect 9079 12937 9088 12971
rect 9036 12928 9088 12937
rect 9772 12928 9824 12980
rect 11704 12971 11756 12980
rect 11704 12937 11713 12971
rect 11713 12937 11747 12971
rect 11747 12937 11756 12971
rect 11704 12928 11756 12937
rect 13636 12971 13688 12980
rect 13636 12937 13645 12971
rect 13645 12937 13679 12971
rect 13679 12937 13688 12971
rect 13636 12928 13688 12937
rect 14464 12928 14516 12980
rect 16120 12928 16172 12980
rect 17592 12928 17644 12980
rect 18604 12928 18656 12980
rect 19892 12928 19944 12980
rect 5908 12860 5960 12912
rect 6184 12860 6236 12912
rect 1584 12724 1636 12776
rect 2228 12724 2280 12776
rect 3516 12724 3568 12776
rect 4712 12767 4764 12776
rect 4712 12733 4721 12767
rect 4721 12733 4755 12767
rect 4755 12733 4764 12767
rect 4712 12724 4764 12733
rect 2596 12656 2648 12708
rect 2872 12656 2924 12708
rect 6460 12724 6512 12776
rect 6828 12767 6880 12776
rect 6828 12733 6837 12767
rect 6837 12733 6871 12767
rect 6871 12733 6880 12767
rect 6828 12724 6880 12733
rect 7380 12767 7432 12776
rect 7380 12733 7389 12767
rect 7389 12733 7423 12767
rect 7423 12733 7432 12767
rect 7380 12724 7432 12733
rect 7564 12724 7616 12776
rect 7932 12724 7984 12776
rect 6276 12699 6328 12708
rect 6276 12665 6285 12699
rect 6285 12665 6319 12699
rect 6319 12665 6328 12699
rect 6276 12656 6328 12665
rect 6552 12656 6604 12708
rect 8944 12724 8996 12776
rect 14832 12792 14884 12844
rect 16488 12860 16540 12912
rect 19064 12903 19116 12912
rect 19064 12869 19073 12903
rect 19073 12869 19107 12903
rect 19107 12869 19116 12903
rect 19064 12860 19116 12869
rect 19800 12903 19852 12912
rect 19800 12869 19809 12903
rect 19809 12869 19843 12903
rect 19843 12869 19852 12903
rect 19800 12860 19852 12869
rect 17776 12792 17828 12844
rect 18512 12792 18564 12844
rect 18788 12835 18840 12844
rect 18788 12801 18797 12835
rect 18797 12801 18831 12835
rect 18831 12801 18840 12835
rect 18788 12792 18840 12801
rect 9680 12724 9732 12776
rect 9864 12767 9916 12776
rect 9864 12733 9873 12767
rect 9873 12733 9907 12767
rect 9907 12733 9916 12767
rect 9864 12724 9916 12733
rect 10140 12767 10192 12776
rect 10140 12733 10149 12767
rect 10149 12733 10183 12767
rect 10183 12733 10192 12767
rect 10140 12724 10192 12733
rect 1400 12588 1452 12640
rect 2688 12588 2740 12640
rect 5172 12631 5224 12640
rect 5172 12597 5181 12631
rect 5181 12597 5215 12631
rect 5215 12597 5224 12631
rect 5172 12588 5224 12597
rect 6368 12588 6420 12640
rect 7104 12631 7156 12640
rect 7104 12597 7113 12631
rect 7113 12597 7147 12631
rect 7147 12597 7156 12631
rect 7104 12588 7156 12597
rect 9680 12588 9732 12640
rect 11980 12724 12032 12776
rect 13544 12724 13596 12776
rect 14188 12767 14240 12776
rect 14188 12733 14197 12767
rect 14197 12733 14231 12767
rect 14231 12733 14240 12767
rect 14188 12724 14240 12733
rect 15200 12724 15252 12776
rect 15384 12724 15436 12776
rect 15752 12724 15804 12776
rect 15844 12724 15896 12776
rect 16304 12724 16356 12776
rect 16488 12724 16540 12776
rect 19340 12724 19392 12776
rect 14004 12699 14056 12708
rect 12716 12631 12768 12640
rect 12716 12597 12725 12631
rect 12725 12597 12759 12631
rect 12759 12597 12768 12631
rect 12716 12588 12768 12597
rect 14004 12665 14013 12699
rect 14013 12665 14047 12699
rect 14047 12665 14056 12699
rect 14004 12656 14056 12665
rect 16764 12656 16816 12708
rect 14188 12588 14240 12640
rect 16580 12631 16632 12640
rect 16580 12597 16589 12631
rect 16589 12597 16623 12631
rect 16623 12597 16632 12631
rect 16580 12588 16632 12597
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1584 12384 1636 12436
rect 2780 12384 2832 12436
rect 3884 12427 3936 12436
rect 3884 12393 3893 12427
rect 3893 12393 3927 12427
rect 3927 12393 3936 12427
rect 3884 12384 3936 12393
rect 4344 12427 4396 12436
rect 4344 12393 4353 12427
rect 4353 12393 4387 12427
rect 4387 12393 4396 12427
rect 4344 12384 4396 12393
rect 4620 12384 4672 12436
rect 5540 12384 5592 12436
rect 5908 12427 5960 12436
rect 5908 12393 5917 12427
rect 5917 12393 5951 12427
rect 5951 12393 5960 12427
rect 5908 12384 5960 12393
rect 6184 12384 6236 12436
rect 7012 12384 7064 12436
rect 9864 12384 9916 12436
rect 10140 12384 10192 12436
rect 10876 12427 10928 12436
rect 10876 12393 10885 12427
rect 10885 12393 10919 12427
rect 10919 12393 10928 12427
rect 10876 12384 10928 12393
rect 12440 12384 12492 12436
rect 14372 12427 14424 12436
rect 1492 12291 1544 12300
rect 1492 12257 1510 12291
rect 1510 12257 1544 12291
rect 1492 12248 1544 12257
rect 5356 12248 5408 12300
rect 5540 12291 5592 12300
rect 5540 12257 5558 12291
rect 5558 12257 5592 12291
rect 5540 12248 5592 12257
rect 6460 12291 6512 12300
rect 4896 12223 4948 12232
rect 4896 12189 4905 12223
rect 4905 12189 4939 12223
rect 4939 12189 4948 12223
rect 4896 12180 4948 12189
rect 2872 12112 2924 12164
rect 5356 12112 5408 12164
rect 6460 12257 6469 12291
rect 6469 12257 6503 12291
rect 6503 12257 6512 12291
rect 6460 12248 6512 12257
rect 6644 12180 6696 12232
rect 7104 12248 7156 12300
rect 7932 12316 7984 12368
rect 9956 12316 10008 12368
rect 14372 12393 14381 12427
rect 14381 12393 14415 12427
rect 14415 12393 14424 12427
rect 14372 12384 14424 12393
rect 15568 12427 15620 12436
rect 15568 12393 15577 12427
rect 15577 12393 15611 12427
rect 15611 12393 15620 12427
rect 15568 12384 15620 12393
rect 16672 12384 16724 12436
rect 7656 12291 7708 12300
rect 7656 12257 7665 12291
rect 7665 12257 7699 12291
rect 7699 12257 7708 12291
rect 7656 12248 7708 12257
rect 9680 12248 9732 12300
rect 9864 12291 9916 12300
rect 9864 12257 9873 12291
rect 9873 12257 9907 12291
rect 9907 12257 9916 12291
rect 9864 12248 9916 12257
rect 10140 12291 10192 12300
rect 10140 12257 10149 12291
rect 10149 12257 10183 12291
rect 10183 12257 10192 12291
rect 10140 12248 10192 12257
rect 11796 12248 11848 12300
rect 7564 12180 7616 12232
rect 8576 12223 8628 12232
rect 8576 12189 8585 12223
rect 8585 12189 8619 12223
rect 8619 12189 8628 12223
rect 8576 12180 8628 12189
rect 10324 12223 10376 12232
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 12716 12248 12768 12300
rect 12164 12223 12216 12232
rect 12164 12189 12173 12223
rect 12173 12189 12207 12223
rect 12207 12189 12216 12223
rect 12164 12180 12216 12189
rect 13176 12248 13228 12300
rect 15200 12316 15252 12368
rect 19064 12316 19116 12368
rect 13544 12291 13596 12300
rect 13544 12257 13553 12291
rect 13553 12257 13587 12291
rect 13587 12257 13596 12291
rect 13544 12248 13596 12257
rect 15476 12291 15528 12300
rect 15476 12257 15485 12291
rect 15485 12257 15519 12291
rect 15519 12257 15528 12291
rect 15476 12248 15528 12257
rect 16672 12248 16724 12300
rect 16764 12223 16816 12232
rect 16764 12189 16773 12223
rect 16773 12189 16807 12223
rect 16807 12189 16816 12223
rect 16764 12180 16816 12189
rect 18788 12180 18840 12232
rect 19432 12180 19484 12232
rect 11704 12112 11756 12164
rect 12072 12112 12124 12164
rect 17132 12112 17184 12164
rect 2044 12044 2096 12096
rect 4068 12044 4120 12096
rect 7288 12044 7340 12096
rect 9128 12044 9180 12096
rect 13544 12044 13596 12096
rect 15292 12044 15344 12096
rect 15660 12044 15712 12096
rect 18236 12044 18288 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1584 11883 1636 11892
rect 1584 11849 1593 11883
rect 1593 11849 1627 11883
rect 1627 11849 1636 11883
rect 1584 11840 1636 11849
rect 5540 11883 5592 11892
rect 5540 11849 5549 11883
rect 5549 11849 5583 11883
rect 5583 11849 5592 11883
rect 5540 11840 5592 11849
rect 6276 11840 6328 11892
rect 7288 11883 7340 11892
rect 7288 11849 7297 11883
rect 7297 11849 7331 11883
rect 7331 11849 7340 11883
rect 7288 11840 7340 11849
rect 7656 11883 7708 11892
rect 7656 11849 7665 11883
rect 7665 11849 7699 11883
rect 7699 11849 7708 11883
rect 7656 11840 7708 11849
rect 9864 11883 9916 11892
rect 9864 11849 9873 11883
rect 9873 11849 9907 11883
rect 9907 11849 9916 11883
rect 9864 11840 9916 11849
rect 13544 11883 13596 11892
rect 13544 11849 13553 11883
rect 13553 11849 13587 11883
rect 13587 11849 13596 11883
rect 13544 11840 13596 11849
rect 19064 11883 19116 11892
rect 19064 11849 19073 11883
rect 19073 11849 19107 11883
rect 19107 11849 19116 11883
rect 19064 11840 19116 11849
rect 19340 11840 19392 11892
rect 19800 11883 19852 11892
rect 19800 11849 19809 11883
rect 19809 11849 19843 11883
rect 19843 11849 19852 11883
rect 19800 11840 19852 11849
rect 4160 11772 4212 11824
rect 5908 11815 5960 11824
rect 5908 11781 5917 11815
rect 5917 11781 5951 11815
rect 5951 11781 5960 11815
rect 5908 11772 5960 11781
rect 7932 11772 7984 11824
rect 12440 11772 12492 11824
rect 2228 11704 2280 11756
rect 5172 11704 5224 11756
rect 7472 11704 7524 11756
rect 7564 11704 7616 11756
rect 16764 11704 16816 11756
rect 18420 11704 18472 11756
rect 1952 11636 2004 11688
rect 2136 11636 2188 11688
rect 2412 11636 2464 11688
rect 3424 11679 3476 11688
rect 3424 11645 3433 11679
rect 3433 11645 3467 11679
rect 3467 11645 3476 11679
rect 3424 11636 3476 11645
rect 3884 11679 3936 11688
rect 3884 11645 3893 11679
rect 3893 11645 3927 11679
rect 3927 11645 3936 11679
rect 3884 11636 3936 11645
rect 4068 11679 4120 11688
rect 4068 11645 4077 11679
rect 4077 11645 4111 11679
rect 4111 11645 4120 11679
rect 4068 11636 4120 11645
rect 4528 11679 4580 11688
rect 4528 11645 4537 11679
rect 4537 11645 4571 11679
rect 4571 11645 4580 11679
rect 4528 11636 4580 11645
rect 5448 11636 5500 11688
rect 7656 11636 7708 11688
rect 8300 11679 8352 11688
rect 8300 11645 8309 11679
rect 8309 11645 8343 11679
rect 8343 11645 8352 11679
rect 8300 11636 8352 11645
rect 8576 11679 8628 11688
rect 8576 11645 8585 11679
rect 8585 11645 8619 11679
rect 8619 11645 8628 11679
rect 8576 11636 8628 11645
rect 9128 11679 9180 11688
rect 9128 11645 9137 11679
rect 9137 11645 9171 11679
rect 9171 11645 9180 11679
rect 9128 11636 9180 11645
rect 9496 11679 9548 11688
rect 9496 11645 9505 11679
rect 9505 11645 9539 11679
rect 9539 11645 9548 11679
rect 9496 11636 9548 11645
rect 10968 11679 11020 11688
rect 10968 11645 10977 11679
rect 10977 11645 11011 11679
rect 11011 11645 11020 11679
rect 10968 11636 11020 11645
rect 12716 11679 12768 11688
rect 8760 11568 8812 11620
rect 9956 11568 10008 11620
rect 11704 11568 11756 11620
rect 12716 11645 12725 11679
rect 12725 11645 12759 11679
rect 12759 11645 12768 11679
rect 12716 11636 12768 11645
rect 14924 11636 14976 11688
rect 15660 11679 15712 11688
rect 15660 11645 15669 11679
rect 15669 11645 15703 11679
rect 15703 11645 15712 11679
rect 15660 11636 15712 11645
rect 15844 11636 15896 11688
rect 18052 11679 18104 11688
rect 18052 11645 18061 11679
rect 18061 11645 18095 11679
rect 18095 11645 18104 11679
rect 18052 11636 18104 11645
rect 18236 11636 18288 11688
rect 19616 11679 19668 11688
rect 19616 11645 19625 11679
rect 19625 11645 19659 11679
rect 19659 11645 19668 11679
rect 19616 11636 19668 11645
rect 13176 11568 13228 11620
rect 14740 11611 14792 11620
rect 14740 11577 14749 11611
rect 14749 11577 14783 11611
rect 14783 11577 14792 11611
rect 14740 11568 14792 11577
rect 19248 11568 19300 11620
rect 6276 11543 6328 11552
rect 6276 11509 6285 11543
rect 6285 11509 6319 11543
rect 6319 11509 6328 11543
rect 6276 11500 6328 11509
rect 8668 11500 8720 11552
rect 10692 11543 10744 11552
rect 10692 11509 10701 11543
rect 10701 11509 10735 11543
rect 10735 11509 10744 11543
rect 10692 11500 10744 11509
rect 12072 11500 12124 11552
rect 12900 11543 12952 11552
rect 12900 11509 12909 11543
rect 12909 11509 12943 11543
rect 12943 11509 12952 11543
rect 12900 11500 12952 11509
rect 15476 11500 15528 11552
rect 16304 11500 16356 11552
rect 16672 11500 16724 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 2412 11296 2464 11348
rect 4528 11296 4580 11348
rect 5356 11339 5408 11348
rect 5356 11305 5365 11339
rect 5365 11305 5399 11339
rect 5399 11305 5408 11339
rect 5356 11296 5408 11305
rect 6000 11296 6052 11348
rect 8576 11296 8628 11348
rect 1768 11160 1820 11212
rect 3424 11228 3476 11280
rect 2228 11203 2280 11212
rect 2228 11169 2237 11203
rect 2237 11169 2271 11203
rect 2271 11169 2280 11203
rect 2228 11160 2280 11169
rect 2688 11203 2740 11212
rect 2688 11169 2697 11203
rect 2697 11169 2731 11203
rect 2731 11169 2740 11203
rect 2688 11160 2740 11169
rect 2872 11203 2924 11212
rect 2872 11169 2881 11203
rect 2881 11169 2915 11203
rect 2915 11169 2924 11203
rect 2872 11160 2924 11169
rect 4620 11160 4672 11212
rect 6000 11160 6052 11212
rect 6184 11203 6236 11212
rect 6184 11169 6193 11203
rect 6193 11169 6227 11203
rect 6227 11169 6236 11203
rect 6184 11160 6236 11169
rect 6368 11203 6420 11212
rect 6368 11169 6377 11203
rect 6377 11169 6411 11203
rect 6411 11169 6420 11203
rect 6368 11160 6420 11169
rect 6552 11160 6604 11212
rect 7564 11160 7616 11212
rect 7932 11160 7984 11212
rect 10140 11296 10192 11348
rect 11060 11296 11112 11348
rect 12716 11339 12768 11348
rect 12716 11305 12725 11339
rect 12725 11305 12759 11339
rect 12759 11305 12768 11339
rect 12716 11296 12768 11305
rect 13176 11296 13228 11348
rect 16856 11296 16908 11348
rect 19432 11339 19484 11348
rect 19432 11305 19441 11339
rect 19441 11305 19475 11339
rect 19475 11305 19484 11339
rect 19432 11296 19484 11305
rect 14372 11271 14424 11280
rect 14372 11237 14381 11271
rect 14381 11237 14415 11271
rect 14415 11237 14424 11271
rect 14372 11228 14424 11237
rect 10968 11160 11020 11212
rect 11704 11203 11756 11212
rect 3884 11024 3936 11076
rect 5356 11092 5408 11144
rect 9680 11092 9732 11144
rect 10692 11092 10744 11144
rect 10876 11135 10928 11144
rect 10876 11101 10885 11135
rect 10885 11101 10919 11135
rect 10919 11101 10928 11135
rect 10876 11092 10928 11101
rect 4252 11067 4304 11076
rect 4252 11033 4261 11067
rect 4261 11033 4295 11067
rect 4295 11033 4304 11067
rect 4252 11024 4304 11033
rect 6092 11024 6144 11076
rect 9956 11024 10008 11076
rect 4160 10956 4212 11008
rect 7012 10956 7064 11008
rect 8668 10956 8720 11008
rect 8944 10999 8996 11008
rect 8944 10965 8953 10999
rect 8953 10965 8987 10999
rect 8987 10965 8996 10999
rect 8944 10956 8996 10965
rect 11428 10956 11480 11008
rect 11704 11169 11713 11203
rect 11713 11169 11747 11203
rect 11747 11169 11756 11203
rect 11704 11160 11756 11169
rect 11980 11203 12032 11212
rect 11980 11169 11989 11203
rect 11989 11169 12023 11203
rect 12023 11169 12032 11203
rect 11980 11160 12032 11169
rect 13636 11203 13688 11212
rect 13636 11169 13645 11203
rect 13645 11169 13679 11203
rect 13679 11169 13688 11203
rect 13636 11160 13688 11169
rect 14004 11160 14056 11212
rect 14832 11228 14884 11280
rect 16488 11228 16540 11280
rect 14648 11160 14700 11212
rect 15384 11160 15436 11212
rect 16856 11203 16908 11212
rect 13820 11092 13872 11144
rect 14740 11092 14792 11144
rect 16856 11169 16865 11203
rect 16865 11169 16899 11203
rect 16899 11169 16908 11203
rect 16856 11160 16908 11169
rect 17132 11203 17184 11212
rect 17132 11169 17141 11203
rect 17141 11169 17175 11203
rect 17175 11169 17184 11203
rect 17132 11160 17184 11169
rect 18052 11203 18104 11212
rect 18052 11169 18061 11203
rect 18061 11169 18095 11203
rect 18095 11169 18104 11203
rect 18052 11160 18104 11169
rect 18972 11203 19024 11212
rect 18972 11169 18981 11203
rect 18981 11169 19015 11203
rect 19015 11169 19024 11203
rect 18972 11160 19024 11169
rect 18236 11092 18288 11144
rect 12072 11024 12124 11076
rect 14924 11024 14976 11076
rect 15936 11024 15988 11076
rect 16948 11067 17000 11076
rect 16948 11033 16957 11067
rect 16957 11033 16991 11067
rect 16991 11033 17000 11067
rect 16948 11024 17000 11033
rect 14556 10956 14608 11008
rect 16488 10999 16540 11008
rect 16488 10965 16497 10999
rect 16497 10965 16531 10999
rect 16531 10965 16540 10999
rect 16488 10956 16540 10965
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 3884 10752 3936 10804
rect 5356 10752 5408 10804
rect 6368 10752 6420 10804
rect 6644 10795 6696 10804
rect 6644 10761 6653 10795
rect 6653 10761 6687 10795
rect 6687 10761 6696 10795
rect 6644 10752 6696 10761
rect 7104 10795 7156 10804
rect 7104 10761 7113 10795
rect 7113 10761 7147 10795
rect 7147 10761 7156 10795
rect 7104 10752 7156 10761
rect 9588 10752 9640 10804
rect 9956 10752 10008 10804
rect 10968 10795 11020 10804
rect 10968 10761 10977 10795
rect 10977 10761 11011 10795
rect 11011 10761 11020 10795
rect 10968 10752 11020 10761
rect 11428 10795 11480 10804
rect 11428 10761 11437 10795
rect 11437 10761 11471 10795
rect 11471 10761 11480 10795
rect 11428 10752 11480 10761
rect 11980 10752 12032 10804
rect 12072 10795 12124 10804
rect 12072 10761 12081 10795
rect 12081 10761 12115 10795
rect 12115 10761 12124 10795
rect 12072 10752 12124 10761
rect 13636 10752 13688 10804
rect 14188 10752 14240 10804
rect 14648 10795 14700 10804
rect 14648 10761 14657 10795
rect 14657 10761 14691 10795
rect 14691 10761 14700 10795
rect 14648 10752 14700 10761
rect 15476 10752 15528 10804
rect 16856 10752 16908 10804
rect 19340 10795 19392 10804
rect 19340 10761 19349 10795
rect 19349 10761 19383 10795
rect 19383 10761 19392 10795
rect 19340 10752 19392 10761
rect 15384 10684 15436 10736
rect 15936 10727 15988 10736
rect 15936 10693 15945 10727
rect 15945 10693 15979 10727
rect 15979 10693 15988 10727
rect 15936 10684 15988 10693
rect 17408 10684 17460 10736
rect 2044 10591 2096 10600
rect 2044 10557 2053 10591
rect 2053 10557 2087 10591
rect 2087 10557 2096 10591
rect 2044 10548 2096 10557
rect 3424 10548 3476 10600
rect 6276 10616 6328 10668
rect 4068 10591 4120 10600
rect 4068 10557 4077 10591
rect 4077 10557 4111 10591
rect 4111 10557 4120 10591
rect 4068 10548 4120 10557
rect 4160 10548 4212 10600
rect 5264 10548 5316 10600
rect 6644 10548 6696 10600
rect 8300 10616 8352 10668
rect 8944 10616 8996 10668
rect 13176 10659 13228 10668
rect 13176 10625 13185 10659
rect 13185 10625 13219 10659
rect 13219 10625 13228 10659
rect 13176 10616 13228 10625
rect 14004 10616 14056 10668
rect 16304 10616 16356 10668
rect 8208 10591 8260 10600
rect 8208 10557 8217 10591
rect 8217 10557 8251 10591
rect 8251 10557 8260 10591
rect 8208 10548 8260 10557
rect 8668 10548 8720 10600
rect 9956 10591 10008 10600
rect 1492 10480 1544 10532
rect 6000 10480 6052 10532
rect 6552 10480 6604 10532
rect 6736 10480 6788 10532
rect 8300 10480 8352 10532
rect 9956 10557 9965 10591
rect 9965 10557 9999 10591
rect 9999 10557 10008 10591
rect 9956 10548 10008 10557
rect 12992 10591 13044 10600
rect 12992 10557 13001 10591
rect 13001 10557 13035 10591
rect 13035 10557 13044 10591
rect 12992 10548 13044 10557
rect 14556 10548 14608 10600
rect 15016 10591 15068 10600
rect 15016 10557 15025 10591
rect 15025 10557 15059 10591
rect 15059 10557 15068 10591
rect 15016 10548 15068 10557
rect 16396 10591 16448 10600
rect 9036 10523 9088 10532
rect 9036 10489 9045 10523
rect 9045 10489 9079 10523
rect 9079 10489 9088 10523
rect 9036 10480 9088 10489
rect 9864 10523 9916 10532
rect 9864 10489 9873 10523
rect 9873 10489 9907 10523
rect 9907 10489 9916 10523
rect 9864 10480 9916 10489
rect 13728 10480 13780 10532
rect 14740 10480 14792 10532
rect 16396 10557 16405 10591
rect 16405 10557 16439 10591
rect 16439 10557 16448 10591
rect 16396 10548 16448 10557
rect 16488 10548 16540 10600
rect 18052 10591 18104 10600
rect 18052 10557 18061 10591
rect 18061 10557 18095 10591
rect 18095 10557 18104 10591
rect 18052 10548 18104 10557
rect 19340 10616 19392 10668
rect 15568 10523 15620 10532
rect 15568 10489 15577 10523
rect 15577 10489 15611 10523
rect 15611 10489 15620 10523
rect 15568 10480 15620 10489
rect 17132 10480 17184 10532
rect 2688 10412 2740 10464
rect 2964 10412 3016 10464
rect 3056 10412 3108 10464
rect 5540 10412 5592 10464
rect 7012 10412 7064 10464
rect 16580 10412 16632 10464
rect 18144 10412 18196 10464
rect 18972 10455 19024 10464
rect 18972 10421 18981 10455
rect 18981 10421 19015 10455
rect 19015 10421 19024 10455
rect 18972 10412 19024 10421
rect 19340 10412 19392 10464
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 1768 10251 1820 10260
rect 1768 10217 1777 10251
rect 1777 10217 1811 10251
rect 1811 10217 1820 10251
rect 1768 10208 1820 10217
rect 2044 10208 2096 10260
rect 3424 10251 3476 10260
rect 3424 10217 3433 10251
rect 3433 10217 3467 10251
rect 3467 10217 3476 10251
rect 3424 10208 3476 10217
rect 4068 10208 4120 10260
rect 4620 10251 4672 10260
rect 4620 10217 4629 10251
rect 4629 10217 4663 10251
rect 4663 10217 4672 10251
rect 4620 10208 4672 10217
rect 2596 10140 2648 10192
rect 6092 10251 6144 10260
rect 6092 10217 6101 10251
rect 6101 10217 6135 10251
rect 6135 10217 6144 10251
rect 6092 10208 6144 10217
rect 7932 10251 7984 10260
rect 7932 10217 7941 10251
rect 7941 10217 7975 10251
rect 7975 10217 7984 10251
rect 7932 10208 7984 10217
rect 8576 10208 8628 10260
rect 11060 10251 11112 10260
rect 11060 10217 11069 10251
rect 11069 10217 11103 10251
rect 11103 10217 11112 10251
rect 11060 10208 11112 10217
rect 12440 10208 12492 10260
rect 13820 10251 13872 10260
rect 13820 10217 13829 10251
rect 13829 10217 13863 10251
rect 13863 10217 13872 10251
rect 13820 10208 13872 10217
rect 15108 10251 15160 10260
rect 15108 10217 15117 10251
rect 15117 10217 15151 10251
rect 15151 10217 15160 10251
rect 15108 10208 15160 10217
rect 18052 10251 18104 10260
rect 18052 10217 18061 10251
rect 18061 10217 18095 10251
rect 18095 10217 18104 10251
rect 18052 10208 18104 10217
rect 18604 10251 18656 10260
rect 18604 10217 18613 10251
rect 18613 10217 18647 10251
rect 18647 10217 18656 10251
rect 18604 10208 18656 10217
rect 9956 10140 10008 10192
rect 11428 10183 11480 10192
rect 11428 10149 11437 10183
rect 11437 10149 11471 10183
rect 11471 10149 11480 10183
rect 11428 10140 11480 10149
rect 14832 10140 14884 10192
rect 6276 10115 6328 10124
rect 6276 10081 6285 10115
rect 6285 10081 6319 10115
rect 6319 10081 6328 10115
rect 6276 10072 6328 10081
rect 6736 10115 6788 10124
rect 6736 10081 6745 10115
rect 6745 10081 6779 10115
rect 6779 10081 6788 10115
rect 6736 10072 6788 10081
rect 7012 10115 7064 10124
rect 7012 10081 7021 10115
rect 7021 10081 7055 10115
rect 7055 10081 7064 10115
rect 7012 10072 7064 10081
rect 7932 10072 7984 10124
rect 8668 10072 8720 10124
rect 9588 10072 9640 10124
rect 12624 10072 12676 10124
rect 2136 10047 2188 10056
rect 2136 10013 2145 10047
rect 2145 10013 2179 10047
rect 2179 10013 2188 10047
rect 2136 10004 2188 10013
rect 5356 9868 5408 9920
rect 6184 9868 6236 9920
rect 8300 9911 8352 9920
rect 8300 9877 8309 9911
rect 8309 9877 8343 9911
rect 8343 9877 8352 9911
rect 8300 9868 8352 9877
rect 8944 9868 8996 9920
rect 9128 9868 9180 9920
rect 10140 10047 10192 10056
rect 10140 10013 10149 10047
rect 10149 10013 10183 10047
rect 10183 10013 10192 10047
rect 10140 10004 10192 10013
rect 11060 10004 11112 10056
rect 12532 10004 12584 10056
rect 13636 10072 13688 10124
rect 15292 10115 15344 10124
rect 15292 10081 15301 10115
rect 15301 10081 15335 10115
rect 15335 10081 15344 10115
rect 15292 10072 15344 10081
rect 15660 10072 15712 10124
rect 16028 10115 16080 10124
rect 16028 10081 16037 10115
rect 16037 10081 16071 10115
rect 16071 10081 16080 10115
rect 16028 10072 16080 10081
rect 16856 10115 16908 10124
rect 16856 10081 16865 10115
rect 16865 10081 16899 10115
rect 16899 10081 16908 10115
rect 16856 10072 16908 10081
rect 17132 10115 17184 10124
rect 17132 10081 17141 10115
rect 17141 10081 17175 10115
rect 17175 10081 17184 10115
rect 17132 10072 17184 10081
rect 18420 10115 18472 10124
rect 18420 10081 18429 10115
rect 18429 10081 18463 10115
rect 18463 10081 18472 10115
rect 18420 10072 18472 10081
rect 19432 10115 19484 10124
rect 19432 10081 19441 10115
rect 19441 10081 19475 10115
rect 19475 10081 19484 10115
rect 19432 10072 19484 10081
rect 13544 10004 13596 10056
rect 15844 10004 15896 10056
rect 17408 10004 17460 10056
rect 16396 9936 16448 9988
rect 16764 9936 16816 9988
rect 18236 9936 18288 9988
rect 19616 9979 19668 9988
rect 19616 9945 19625 9979
rect 19625 9945 19659 9979
rect 19659 9945 19668 9979
rect 19616 9936 19668 9945
rect 12992 9868 13044 9920
rect 14740 9911 14792 9920
rect 14740 9877 14749 9911
rect 14749 9877 14783 9911
rect 14783 9877 14792 9911
rect 14740 9868 14792 9877
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 5540 9707 5592 9716
rect 5540 9673 5549 9707
rect 5549 9673 5583 9707
rect 5583 9673 5592 9707
rect 5540 9664 5592 9673
rect 2964 9596 3016 9648
rect 1676 9571 1728 9580
rect 1676 9537 1685 9571
rect 1685 9537 1719 9571
rect 1719 9537 1728 9571
rect 1676 9528 1728 9537
rect 2320 9571 2372 9580
rect 2320 9537 2329 9571
rect 2329 9537 2363 9571
rect 2363 9537 2372 9571
rect 2320 9528 2372 9537
rect 3424 9503 3476 9512
rect 3424 9469 3433 9503
rect 3433 9469 3467 9503
rect 3467 9469 3476 9503
rect 3424 9460 3476 9469
rect 3884 9503 3936 9512
rect 3884 9469 3893 9503
rect 3893 9469 3927 9503
rect 3927 9469 3936 9503
rect 3884 9460 3936 9469
rect 4528 9503 4580 9512
rect 4528 9469 4537 9503
rect 4537 9469 4571 9503
rect 4571 9469 4580 9503
rect 4528 9460 4580 9469
rect 6736 9664 6788 9716
rect 7748 9664 7800 9716
rect 9956 9664 10008 9716
rect 10968 9664 11020 9716
rect 7380 9528 7432 9580
rect 8760 9596 8812 9648
rect 9036 9528 9088 9580
rect 7104 9503 7156 9512
rect 7104 9469 7113 9503
rect 7113 9469 7147 9503
rect 7147 9469 7156 9503
rect 7104 9460 7156 9469
rect 7840 9503 7892 9512
rect 2044 9392 2096 9444
rect 2596 9367 2648 9376
rect 2596 9333 2605 9367
rect 2605 9333 2639 9367
rect 2639 9333 2648 9367
rect 2596 9324 2648 9333
rect 4436 9324 4488 9376
rect 6184 9324 6236 9376
rect 6828 9324 6880 9376
rect 7840 9469 7849 9503
rect 7849 9469 7883 9503
rect 7883 9469 7892 9503
rect 7840 9460 7892 9469
rect 7932 9460 7984 9512
rect 12532 9664 12584 9716
rect 13544 9707 13596 9716
rect 13544 9673 13553 9707
rect 13553 9673 13587 9707
rect 13587 9673 13596 9707
rect 13544 9664 13596 9673
rect 16396 9664 16448 9716
rect 16856 9664 16908 9716
rect 18420 9664 18472 9716
rect 19432 9707 19484 9716
rect 19432 9673 19441 9707
rect 19441 9673 19475 9707
rect 19475 9673 19484 9707
rect 19432 9664 19484 9673
rect 12900 9596 12952 9648
rect 11520 9571 11572 9580
rect 11520 9537 11529 9571
rect 11529 9537 11563 9571
rect 11563 9537 11572 9571
rect 11520 9528 11572 9537
rect 12532 9571 12584 9580
rect 12532 9537 12541 9571
rect 12541 9537 12575 9571
rect 12575 9537 12584 9571
rect 12532 9528 12584 9537
rect 15292 9528 15344 9580
rect 15200 9460 15252 9512
rect 16120 9503 16172 9512
rect 9496 9392 9548 9444
rect 10784 9392 10836 9444
rect 12624 9435 12676 9444
rect 12624 9401 12633 9435
rect 12633 9401 12667 9435
rect 12667 9401 12676 9435
rect 12624 9392 12676 9401
rect 12900 9392 12952 9444
rect 8024 9367 8076 9376
rect 8024 9333 8033 9367
rect 8033 9333 8067 9367
rect 8067 9333 8076 9367
rect 8024 9324 8076 9333
rect 16120 9469 16129 9503
rect 16129 9469 16163 9503
rect 16163 9469 16172 9503
rect 16120 9460 16172 9469
rect 16304 9460 16356 9512
rect 16488 9460 16540 9512
rect 15660 9392 15712 9444
rect 17132 9596 17184 9648
rect 17408 9639 17460 9648
rect 17408 9605 17417 9639
rect 17417 9605 17451 9639
rect 17451 9605 17460 9639
rect 17408 9596 17460 9605
rect 17960 9528 18012 9580
rect 20168 9639 20220 9648
rect 20168 9605 20177 9639
rect 20177 9605 20211 9639
rect 20211 9605 20220 9639
rect 20168 9596 20220 9605
rect 18236 9435 18288 9444
rect 18236 9401 18245 9435
rect 18245 9401 18279 9435
rect 18279 9401 18288 9435
rect 18236 9392 18288 9401
rect 18788 9435 18840 9444
rect 18788 9401 18797 9435
rect 18797 9401 18831 9435
rect 18831 9401 18840 9435
rect 18788 9392 18840 9401
rect 15752 9324 15804 9376
rect 16212 9367 16264 9376
rect 16212 9333 16221 9367
rect 16221 9333 16255 9367
rect 16255 9333 16264 9367
rect 16212 9324 16264 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2872 9120 2924 9172
rect 3884 9120 3936 9172
rect 4344 9163 4396 9172
rect 4344 9129 4353 9163
rect 4353 9129 4387 9163
rect 4387 9129 4396 9163
rect 4344 9120 4396 9129
rect 8668 9163 8720 9172
rect 8668 9129 8677 9163
rect 8677 9129 8711 9163
rect 8711 9129 8720 9163
rect 8668 9120 8720 9129
rect 8944 9163 8996 9172
rect 8944 9129 8953 9163
rect 8953 9129 8987 9163
rect 8987 9129 8996 9163
rect 8944 9120 8996 9129
rect 9036 9120 9088 9172
rect 11428 9120 11480 9172
rect 12624 9163 12676 9172
rect 12624 9129 12633 9163
rect 12633 9129 12667 9163
rect 12667 9129 12676 9163
rect 12624 9120 12676 9129
rect 15384 9120 15436 9172
rect 15844 9163 15896 9172
rect 15844 9129 15853 9163
rect 15853 9129 15887 9163
rect 15887 9129 15896 9163
rect 15844 9120 15896 9129
rect 16120 9163 16172 9172
rect 16120 9129 16129 9163
rect 16129 9129 16163 9163
rect 16163 9129 16172 9163
rect 16120 9120 16172 9129
rect 17960 9163 18012 9172
rect 17960 9129 17969 9163
rect 17969 9129 18003 9163
rect 18003 9129 18012 9163
rect 17960 9120 18012 9129
rect 1492 9052 1544 9104
rect 1768 9052 1820 9104
rect 2320 9052 2372 9104
rect 3700 9052 3752 9104
rect 4252 9052 4304 9104
rect 3516 8984 3568 9036
rect 4068 9027 4120 9036
rect 4068 8993 4077 9027
rect 4077 8993 4111 9027
rect 4111 8993 4120 9027
rect 4068 8984 4120 8993
rect 6460 9052 6512 9104
rect 9864 9095 9916 9104
rect 4988 9027 5040 9036
rect 4988 8993 4997 9027
rect 4997 8993 5031 9027
rect 5031 8993 5040 9027
rect 4988 8984 5040 8993
rect 5264 9027 5316 9036
rect 5264 8993 5273 9027
rect 5273 8993 5307 9027
rect 5307 8993 5316 9027
rect 5264 8984 5316 8993
rect 5356 8984 5408 9036
rect 6000 8984 6052 9036
rect 6828 9027 6880 9036
rect 6828 8993 6837 9027
rect 6837 8993 6871 9027
rect 6871 8993 6880 9027
rect 6828 8984 6880 8993
rect 9864 9061 9873 9095
rect 9873 9061 9907 9095
rect 9907 9061 9916 9095
rect 9864 9052 9916 9061
rect 11796 9052 11848 9104
rect 16672 9095 16724 9104
rect 16672 9061 16675 9095
rect 16675 9061 16709 9095
rect 16709 9061 16724 9095
rect 16672 9052 16724 9061
rect 17776 9052 17828 9104
rect 18788 9095 18840 9104
rect 18788 9061 18797 9095
rect 18797 9061 18831 9095
rect 18831 9061 18840 9095
rect 18788 9052 18840 9061
rect 1492 8959 1544 8968
rect 1492 8925 1501 8959
rect 1501 8925 1535 8959
rect 1535 8925 1544 8959
rect 1492 8916 1544 8925
rect 7932 8984 7984 9036
rect 11888 8984 11940 9036
rect 12348 8984 12400 9036
rect 13728 9027 13780 9036
rect 13728 8993 13737 9027
rect 13737 8993 13771 9027
rect 13771 8993 13780 9027
rect 13728 8984 13780 8993
rect 9772 8959 9824 8968
rect 9772 8925 9781 8959
rect 9781 8925 9815 8959
rect 9815 8925 9824 8959
rect 9772 8916 9824 8925
rect 10140 8959 10192 8968
rect 10140 8925 10149 8959
rect 10149 8925 10183 8959
rect 10183 8925 10192 8959
rect 10140 8916 10192 8925
rect 13636 8916 13688 8968
rect 14280 8984 14332 9036
rect 15292 9027 15344 9036
rect 15292 8993 15301 9027
rect 15301 8993 15335 9027
rect 15335 8993 15344 9027
rect 15292 8984 15344 8993
rect 16488 8984 16540 9036
rect 20076 8984 20128 9036
rect 14004 8959 14056 8968
rect 14004 8925 14013 8959
rect 14013 8925 14047 8959
rect 14047 8925 14056 8959
rect 14004 8916 14056 8925
rect 18144 8959 18196 8968
rect 18144 8925 18153 8959
rect 18153 8925 18187 8959
rect 18187 8925 18196 8959
rect 18144 8916 18196 8925
rect 4528 8848 4580 8900
rect 4896 8848 4948 8900
rect 6092 8848 6144 8900
rect 7012 8848 7064 8900
rect 2872 8823 2924 8832
rect 2872 8789 2881 8823
rect 2881 8789 2915 8823
rect 2915 8789 2924 8823
rect 2872 8780 2924 8789
rect 7104 8780 7156 8832
rect 8760 8780 8812 8832
rect 14740 8780 14792 8832
rect 16304 8780 16356 8832
rect 17776 8780 17828 8832
rect 19800 8823 19852 8832
rect 19800 8789 19809 8823
rect 19809 8789 19843 8823
rect 19843 8789 19852 8823
rect 19800 8780 19852 8789
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 1768 8576 1820 8628
rect 2872 8619 2924 8628
rect 2872 8585 2881 8619
rect 2881 8585 2915 8619
rect 2915 8585 2924 8619
rect 2872 8576 2924 8585
rect 3240 8619 3292 8628
rect 3240 8585 3249 8619
rect 3249 8585 3283 8619
rect 3283 8585 3292 8619
rect 3240 8576 3292 8585
rect 3516 8619 3568 8628
rect 3516 8585 3525 8619
rect 3525 8585 3559 8619
rect 3559 8585 3568 8619
rect 3516 8576 3568 8585
rect 5264 8576 5316 8628
rect 6092 8619 6144 8628
rect 6092 8585 6101 8619
rect 6101 8585 6135 8619
rect 6135 8585 6144 8619
rect 6092 8576 6144 8585
rect 6368 8619 6420 8628
rect 6368 8585 6377 8619
rect 6377 8585 6411 8619
rect 6411 8585 6420 8619
rect 6368 8576 6420 8585
rect 8760 8619 8812 8628
rect 8760 8585 8769 8619
rect 8769 8585 8803 8619
rect 8803 8585 8812 8619
rect 8760 8576 8812 8585
rect 9864 8619 9916 8628
rect 9864 8585 9873 8619
rect 9873 8585 9907 8619
rect 9907 8585 9916 8619
rect 9864 8576 9916 8585
rect 11428 8576 11480 8628
rect 13728 8576 13780 8628
rect 15292 8576 15344 8628
rect 17776 8619 17828 8628
rect 17776 8585 17785 8619
rect 17785 8585 17819 8619
rect 17819 8585 17828 8619
rect 17776 8576 17828 8585
rect 18144 8576 18196 8628
rect 19984 8576 20036 8628
rect 6276 8508 6328 8560
rect 18236 8508 18288 8560
rect 19248 8508 19300 8560
rect 1952 8372 2004 8424
rect 3240 8372 3292 8424
rect 4068 8372 4120 8424
rect 4252 8415 4304 8424
rect 4252 8381 4261 8415
rect 4261 8381 4295 8415
rect 4295 8381 4304 8415
rect 4252 8372 4304 8381
rect 4988 8440 5040 8492
rect 6828 8440 6880 8492
rect 4896 8415 4948 8424
rect 4896 8381 4905 8415
rect 4905 8381 4939 8415
rect 4939 8381 4948 8415
rect 4896 8372 4948 8381
rect 6000 8372 6052 8424
rect 7104 8372 7156 8424
rect 10600 8483 10652 8492
rect 10600 8449 10609 8483
rect 10609 8449 10643 8483
rect 10643 8449 10652 8483
rect 10600 8440 10652 8449
rect 7840 8415 7892 8424
rect 7840 8381 7849 8415
rect 7849 8381 7883 8415
rect 7883 8381 7892 8415
rect 7840 8372 7892 8381
rect 8300 8415 8352 8424
rect 8300 8381 8309 8415
rect 8309 8381 8343 8415
rect 8343 8381 8352 8415
rect 8300 8372 8352 8381
rect 9496 8372 9548 8424
rect 9404 8304 9456 8356
rect 13636 8372 13688 8424
rect 15568 8440 15620 8492
rect 18788 8440 18840 8492
rect 14096 8415 14148 8424
rect 14096 8381 14105 8415
rect 14105 8381 14139 8415
rect 14139 8381 14148 8415
rect 14096 8372 14148 8381
rect 14740 8372 14792 8424
rect 20076 8415 20128 8424
rect 20076 8381 20085 8415
rect 20085 8381 20119 8415
rect 20119 8381 20128 8415
rect 20076 8372 20128 8381
rect 11796 8347 11848 8356
rect 11796 8313 11805 8347
rect 11805 8313 11839 8347
rect 11839 8313 11848 8347
rect 11796 8304 11848 8313
rect 13176 8347 13228 8356
rect 13176 8313 13185 8347
rect 13185 8313 13219 8347
rect 13219 8313 13228 8347
rect 13176 8304 13228 8313
rect 14832 8347 14884 8356
rect 14832 8313 14841 8347
rect 14841 8313 14875 8347
rect 14875 8313 14884 8347
rect 14832 8304 14884 8313
rect 3792 8279 3844 8288
rect 3792 8245 3801 8279
rect 3801 8245 3835 8279
rect 3835 8245 3844 8279
rect 3792 8236 3844 8245
rect 7840 8236 7892 8288
rect 15292 8236 15344 8288
rect 16672 8304 16724 8356
rect 17500 8279 17552 8288
rect 17500 8245 17509 8279
rect 17509 8245 17543 8279
rect 17543 8245 17552 8279
rect 17500 8236 17552 8245
rect 18604 8304 18656 8356
rect 19156 8236 19208 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1492 8032 1544 8084
rect 2044 8032 2096 8084
rect 4160 8032 4212 8084
rect 4988 7964 5040 8016
rect 3056 7939 3108 7948
rect 3056 7905 3065 7939
rect 3065 7905 3099 7939
rect 3099 7905 3108 7939
rect 3056 7896 3108 7905
rect 4712 7939 4764 7948
rect 4712 7905 4730 7939
rect 4730 7905 4764 7939
rect 4712 7896 4764 7905
rect 7748 8032 7800 8084
rect 10692 8075 10744 8084
rect 10692 8041 10701 8075
rect 10701 8041 10735 8075
rect 10735 8041 10744 8075
rect 10692 8032 10744 8041
rect 11888 8075 11940 8084
rect 11888 8041 11897 8075
rect 11897 8041 11931 8075
rect 11931 8041 11940 8075
rect 11888 8032 11940 8041
rect 13636 8075 13688 8084
rect 13636 8041 13645 8075
rect 13645 8041 13679 8075
rect 13679 8041 13688 8075
rect 13636 8032 13688 8041
rect 15476 8075 15528 8084
rect 15476 8041 15485 8075
rect 15485 8041 15519 8075
rect 15519 8041 15528 8075
rect 15476 8032 15528 8041
rect 15568 8032 15620 8084
rect 16488 8032 16540 8084
rect 17500 8075 17552 8084
rect 17500 8041 17509 8075
rect 17509 8041 17543 8075
rect 17543 8041 17552 8075
rect 17500 8032 17552 8041
rect 6276 7964 6328 8016
rect 6000 7896 6052 7948
rect 6184 7939 6236 7948
rect 6184 7905 6193 7939
rect 6193 7905 6227 7939
rect 6227 7905 6236 7939
rect 6184 7896 6236 7905
rect 6368 7896 6420 7948
rect 11796 7964 11848 8016
rect 8208 7896 8260 7948
rect 8668 7939 8720 7948
rect 8668 7905 8677 7939
rect 8677 7905 8711 7939
rect 8711 7905 8720 7939
rect 8668 7896 8720 7905
rect 10048 7896 10100 7948
rect 11152 7939 11204 7948
rect 11152 7905 11161 7939
rect 11161 7905 11195 7939
rect 11195 7905 11204 7939
rect 11152 7896 11204 7905
rect 11428 7939 11480 7948
rect 11428 7905 11437 7939
rect 11437 7905 11471 7939
rect 11471 7905 11480 7939
rect 16672 7964 16724 8016
rect 17868 7964 17920 8016
rect 18788 7964 18840 8016
rect 14188 7939 14240 7948
rect 11428 7896 11480 7905
rect 14188 7905 14197 7939
rect 14197 7905 14231 7939
rect 14231 7905 14240 7939
rect 14188 7896 14240 7905
rect 15476 7896 15528 7948
rect 15752 7896 15804 7948
rect 16580 7939 16632 7948
rect 16580 7905 16589 7939
rect 16589 7905 16623 7939
rect 16623 7905 16632 7939
rect 16580 7896 16632 7905
rect 8116 7828 8168 7880
rect 9312 7828 9364 7880
rect 12348 7828 12400 7880
rect 13176 7828 13228 7880
rect 19156 7828 19208 7880
rect 5540 7760 5592 7812
rect 6920 7760 6972 7812
rect 14188 7760 14240 7812
rect 2688 7735 2740 7744
rect 2688 7701 2697 7735
rect 2697 7701 2731 7735
rect 2731 7701 2740 7735
rect 2688 7692 2740 7701
rect 9588 7692 9640 7744
rect 10140 7692 10192 7744
rect 14740 7692 14792 7744
rect 17960 7692 18012 7744
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 1584 7531 1636 7540
rect 1584 7497 1593 7531
rect 1593 7497 1627 7531
rect 1627 7497 1636 7531
rect 1584 7488 1636 7497
rect 2136 7531 2188 7540
rect 2136 7497 2145 7531
rect 2145 7497 2179 7531
rect 2179 7497 2188 7531
rect 2136 7488 2188 7497
rect 2780 7488 2832 7540
rect 3056 7488 3108 7540
rect 3884 7531 3936 7540
rect 3884 7497 3893 7531
rect 3893 7497 3927 7531
rect 3927 7497 3936 7531
rect 3884 7488 3936 7497
rect 6368 7488 6420 7540
rect 7104 7531 7156 7540
rect 7104 7497 7113 7531
rect 7113 7497 7147 7531
rect 7147 7497 7156 7531
rect 7104 7488 7156 7497
rect 8668 7531 8720 7540
rect 8668 7497 8677 7531
rect 8677 7497 8711 7531
rect 8711 7497 8720 7531
rect 8668 7488 8720 7497
rect 10048 7488 10100 7540
rect 11152 7488 11204 7540
rect 11796 7488 11848 7540
rect 13176 7488 13228 7540
rect 14096 7488 14148 7540
rect 17684 7488 17736 7540
rect 17868 7531 17920 7540
rect 17868 7497 17877 7531
rect 17877 7497 17911 7531
rect 17911 7497 17920 7531
rect 17868 7488 17920 7497
rect 18236 7488 18288 7540
rect 18512 7488 18564 7540
rect 19156 7531 19208 7540
rect 19156 7497 19165 7531
rect 19165 7497 19199 7531
rect 19199 7497 19208 7531
rect 19156 7488 19208 7497
rect 6276 7463 6328 7472
rect 6276 7429 6285 7463
rect 6285 7429 6319 7463
rect 6319 7429 6328 7463
rect 6276 7420 6328 7429
rect 2320 7352 2372 7404
rect 3792 7352 3844 7404
rect 4344 7352 4396 7404
rect 5080 7352 5132 7404
rect 8024 7352 8076 7404
rect 1400 7327 1452 7336
rect 1400 7293 1409 7327
rect 1409 7293 1443 7327
rect 1443 7293 1452 7327
rect 1400 7284 1452 7293
rect 9496 7420 9548 7472
rect 12900 7395 12952 7404
rect 12900 7361 12909 7395
rect 12909 7361 12943 7395
rect 12943 7361 12952 7395
rect 14096 7395 14148 7404
rect 12900 7352 12952 7361
rect 14096 7361 14105 7395
rect 14105 7361 14139 7395
rect 14139 7361 14148 7395
rect 14096 7352 14148 7361
rect 14372 7395 14424 7404
rect 14372 7361 14381 7395
rect 14381 7361 14415 7395
rect 14415 7361 14424 7395
rect 14372 7352 14424 7361
rect 16212 7395 16264 7404
rect 16212 7361 16221 7395
rect 16221 7361 16255 7395
rect 16255 7361 16264 7395
rect 16212 7352 16264 7361
rect 18604 7395 18656 7404
rect 18604 7361 18613 7395
rect 18613 7361 18647 7395
rect 18647 7361 18656 7395
rect 18604 7352 18656 7361
rect 8944 7284 8996 7336
rect 9220 7284 9272 7336
rect 15292 7284 15344 7336
rect 20260 7488 20312 7540
rect 2596 7216 2648 7268
rect 6276 7216 6328 7268
rect 8116 7259 8168 7268
rect 8116 7225 8119 7259
rect 8119 7225 8153 7259
rect 8153 7225 8168 7259
rect 8116 7216 8168 7225
rect 4712 7148 4764 7200
rect 5356 7148 5408 7200
rect 5448 7148 5500 7200
rect 9220 7148 9272 7200
rect 9496 7148 9548 7200
rect 9680 7259 9732 7268
rect 9680 7225 9689 7259
rect 9689 7225 9723 7259
rect 9723 7225 9732 7259
rect 9680 7216 9732 7225
rect 10692 7216 10744 7268
rect 12532 7259 12584 7268
rect 12532 7225 12541 7259
rect 12541 7225 12575 7259
rect 12575 7225 12584 7259
rect 12532 7216 12584 7225
rect 11796 7191 11848 7200
rect 11796 7157 11805 7191
rect 11805 7157 11839 7191
rect 11839 7157 11848 7191
rect 11796 7148 11848 7157
rect 12256 7148 12308 7200
rect 14188 7259 14240 7268
rect 14188 7225 14197 7259
rect 14197 7225 14231 7259
rect 14231 7225 14240 7259
rect 14188 7216 14240 7225
rect 18144 7259 18196 7268
rect 18144 7225 18153 7259
rect 18153 7225 18187 7259
rect 18187 7225 18196 7259
rect 18144 7216 18196 7225
rect 15476 7148 15528 7200
rect 17960 7148 18012 7200
rect 19340 7148 19392 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 1400 6944 1452 6996
rect 2504 6944 2556 6996
rect 5080 6987 5132 6996
rect 5080 6953 5089 6987
rect 5089 6953 5123 6987
rect 5123 6953 5132 6987
rect 5080 6944 5132 6953
rect 8024 6944 8076 6996
rect 9220 6944 9272 6996
rect 9680 6944 9732 6996
rect 11428 6944 11480 6996
rect 12532 6987 12584 6996
rect 12532 6953 12541 6987
rect 12541 6953 12575 6987
rect 12575 6953 12584 6987
rect 12532 6944 12584 6953
rect 14096 6944 14148 6996
rect 15384 6987 15436 6996
rect 15384 6953 15393 6987
rect 15393 6953 15427 6987
rect 15427 6953 15436 6987
rect 15384 6944 15436 6953
rect 16580 6987 16632 6996
rect 16580 6953 16589 6987
rect 16589 6953 16623 6987
rect 16623 6953 16632 6987
rect 16580 6944 16632 6953
rect 2688 6876 2740 6928
rect 3884 6876 3936 6928
rect 4252 6919 4304 6928
rect 4252 6885 4261 6919
rect 4261 6885 4295 6919
rect 4295 6885 4304 6919
rect 4252 6876 4304 6885
rect 6092 6876 6144 6928
rect 8116 6876 8168 6928
rect 9312 6876 9364 6928
rect 9864 6919 9916 6928
rect 9864 6885 9873 6919
rect 9873 6885 9907 6919
rect 9907 6885 9916 6919
rect 9864 6876 9916 6885
rect 11704 6876 11756 6928
rect 12348 6876 12400 6928
rect 13360 6919 13412 6928
rect 13360 6885 13369 6919
rect 13369 6885 13403 6919
rect 13403 6885 13412 6919
rect 13360 6876 13412 6885
rect 14372 6876 14424 6928
rect 17684 6919 17736 6928
rect 17684 6885 17693 6919
rect 17693 6885 17727 6919
rect 17727 6885 17736 6919
rect 17684 6876 17736 6885
rect 2320 6808 2372 6860
rect 3700 6851 3752 6860
rect 3700 6817 3709 6851
rect 3709 6817 3743 6851
rect 3743 6817 3752 6851
rect 3700 6808 3752 6817
rect 7840 6851 7892 6860
rect 7840 6817 7849 6851
rect 7849 6817 7883 6851
rect 7883 6817 7892 6851
rect 7840 6808 7892 6817
rect 14648 6808 14700 6860
rect 15568 6808 15620 6860
rect 16396 6808 16448 6860
rect 19064 6851 19116 6860
rect 19064 6817 19073 6851
rect 19073 6817 19107 6851
rect 19107 6817 19116 6851
rect 19064 6808 19116 6817
rect 19432 6808 19484 6860
rect 2136 6740 2188 6792
rect 4160 6783 4212 6792
rect 4160 6749 4169 6783
rect 4169 6749 4203 6783
rect 4203 6749 4212 6783
rect 4160 6740 4212 6749
rect 2688 6672 2740 6724
rect 3516 6672 3568 6724
rect 5540 6740 5592 6792
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 9404 6740 9456 6792
rect 10048 6740 10100 6792
rect 11520 6740 11572 6792
rect 11612 6740 11664 6792
rect 14004 6740 14056 6792
rect 17592 6783 17644 6792
rect 17592 6749 17601 6783
rect 17601 6749 17635 6783
rect 17635 6749 17644 6783
rect 17592 6740 17644 6749
rect 19616 6783 19668 6792
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 9312 6672 9364 6724
rect 18144 6715 18196 6724
rect 18144 6681 18153 6715
rect 18153 6681 18187 6715
rect 18187 6681 18196 6715
rect 18144 6672 18196 6681
rect 3700 6604 3752 6656
rect 6184 6604 6236 6656
rect 8668 6604 8720 6656
rect 9220 6604 9272 6656
rect 9496 6647 9548 6656
rect 9496 6613 9505 6647
rect 9505 6613 9539 6647
rect 9539 6613 9548 6647
rect 9496 6604 9548 6613
rect 11060 6604 11112 6656
rect 11796 6604 11848 6656
rect 12256 6604 12308 6656
rect 18052 6604 18104 6656
rect 18880 6647 18932 6656
rect 18880 6613 18889 6647
rect 18889 6613 18923 6647
rect 18923 6613 18932 6647
rect 18880 6604 18932 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 2136 6443 2188 6452
rect 2136 6409 2145 6443
rect 2145 6409 2179 6443
rect 2179 6409 2188 6443
rect 2136 6400 2188 6409
rect 2596 6400 2648 6452
rect 4252 6443 4304 6452
rect 4252 6409 4261 6443
rect 4261 6409 4295 6443
rect 4295 6409 4304 6443
rect 4252 6400 4304 6409
rect 5540 6400 5592 6452
rect 7840 6400 7892 6452
rect 9864 6400 9916 6452
rect 11704 6400 11756 6452
rect 13360 6443 13412 6452
rect 1584 6375 1636 6384
rect 1584 6341 1593 6375
rect 1593 6341 1627 6375
rect 1627 6341 1636 6375
rect 1584 6332 1636 6341
rect 4160 6332 4212 6384
rect 6000 6332 6052 6384
rect 8116 6332 8168 6384
rect 2964 6307 3016 6316
rect 2964 6273 2973 6307
rect 2973 6273 3007 6307
rect 3007 6273 3016 6307
rect 2964 6264 3016 6273
rect 5264 6307 5316 6316
rect 5264 6273 5273 6307
rect 5273 6273 5307 6307
rect 5307 6273 5316 6307
rect 5264 6264 5316 6273
rect 9036 6264 9088 6316
rect 10692 6307 10744 6316
rect 10692 6273 10701 6307
rect 10701 6273 10735 6307
rect 10735 6273 10744 6307
rect 10692 6264 10744 6273
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 3332 6171 3384 6180
rect 3332 6137 3335 6171
rect 3335 6137 3369 6171
rect 3369 6137 3384 6171
rect 3332 6128 3384 6137
rect 4712 6128 4764 6180
rect 5448 6128 5500 6180
rect 8760 6171 8812 6180
rect 8760 6137 8769 6171
rect 8769 6137 8803 6171
rect 8803 6137 8812 6171
rect 9312 6171 9364 6180
rect 8760 6128 8812 6137
rect 9312 6137 9321 6171
rect 9321 6137 9355 6171
rect 9355 6137 9364 6171
rect 9312 6128 9364 6137
rect 9864 6128 9916 6180
rect 13360 6409 13369 6443
rect 13369 6409 13403 6443
rect 13403 6409 13412 6443
rect 13360 6400 13412 6409
rect 14004 6443 14056 6452
rect 14004 6409 14013 6443
rect 14013 6409 14047 6443
rect 14047 6409 14056 6443
rect 14004 6400 14056 6409
rect 16396 6400 16448 6452
rect 17776 6443 17828 6452
rect 17776 6409 17785 6443
rect 17785 6409 17819 6443
rect 17819 6409 17828 6443
rect 17776 6400 17828 6409
rect 19064 6443 19116 6452
rect 19064 6409 19073 6443
rect 19073 6409 19107 6443
rect 19107 6409 19116 6443
rect 19064 6400 19116 6409
rect 19432 6443 19484 6452
rect 19432 6409 19441 6443
rect 19441 6409 19475 6443
rect 19475 6409 19484 6443
rect 19432 6400 19484 6409
rect 12348 6264 12400 6316
rect 14556 6332 14608 6384
rect 14832 6375 14884 6384
rect 14832 6341 14841 6375
rect 14841 6341 14875 6375
rect 14875 6341 14884 6375
rect 14832 6332 14884 6341
rect 17684 6332 17736 6384
rect 17960 6332 18012 6384
rect 14832 6196 14884 6248
rect 16580 6196 16632 6248
rect 18880 6196 18932 6248
rect 19432 6196 19484 6248
rect 3884 6103 3936 6112
rect 3884 6069 3893 6103
rect 3893 6069 3927 6103
rect 3927 6069 3936 6103
rect 3884 6060 3936 6069
rect 5816 6060 5868 6112
rect 6092 6060 6144 6112
rect 7380 6103 7432 6112
rect 7380 6069 7389 6103
rect 7389 6069 7423 6103
rect 7423 6069 7432 6103
rect 7380 6060 7432 6069
rect 9680 6060 9732 6112
rect 12716 6128 12768 6180
rect 15292 6128 15344 6180
rect 11520 6060 11572 6112
rect 15200 6103 15252 6112
rect 15200 6069 15209 6103
rect 15209 6069 15243 6103
rect 15243 6069 15252 6103
rect 15844 6128 15896 6180
rect 18144 6171 18196 6180
rect 18144 6137 18153 6171
rect 18153 6137 18187 6171
rect 18187 6137 18196 6171
rect 18144 6128 18196 6137
rect 15200 6060 15252 6069
rect 17776 6060 17828 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 2044 5899 2096 5908
rect 2044 5865 2053 5899
rect 2053 5865 2087 5899
rect 2087 5865 2096 5899
rect 2044 5856 2096 5865
rect 2136 5856 2188 5908
rect 2964 5856 3016 5908
rect 3516 5899 3568 5908
rect 3516 5865 3525 5899
rect 3525 5865 3559 5899
rect 3559 5865 3568 5899
rect 3516 5856 3568 5865
rect 5264 5899 5316 5908
rect 5264 5865 5273 5899
rect 5273 5865 5307 5899
rect 5307 5865 5316 5899
rect 5264 5856 5316 5865
rect 6920 5899 6972 5908
rect 6920 5865 6929 5899
rect 6929 5865 6963 5899
rect 6963 5865 6972 5899
rect 6920 5856 6972 5865
rect 8760 5856 8812 5908
rect 9036 5899 9088 5908
rect 9036 5865 9045 5899
rect 9045 5865 9079 5899
rect 9079 5865 9088 5899
rect 9036 5856 9088 5865
rect 9496 5856 9548 5908
rect 10140 5856 10192 5908
rect 15568 5899 15620 5908
rect 2504 5788 2556 5840
rect 5816 5788 5868 5840
rect 6276 5788 6328 5840
rect 15568 5865 15577 5899
rect 15577 5865 15611 5899
rect 15611 5865 15620 5899
rect 15568 5856 15620 5865
rect 17868 5856 17920 5908
rect 11060 5831 11112 5840
rect 11060 5797 11069 5831
rect 11069 5797 11103 5831
rect 11103 5797 11112 5831
rect 11612 5831 11664 5840
rect 11060 5788 11112 5797
rect 11612 5797 11621 5831
rect 11621 5797 11655 5831
rect 11655 5797 11664 5831
rect 11612 5788 11664 5797
rect 12716 5788 12768 5840
rect 15844 5788 15896 5840
rect 17592 5788 17644 5840
rect 17776 5788 17828 5840
rect 19248 5831 19300 5840
rect 19248 5797 19257 5831
rect 19257 5797 19291 5831
rect 19291 5797 19300 5831
rect 19248 5788 19300 5797
rect 1676 5763 1728 5772
rect 1676 5729 1694 5763
rect 1694 5729 1728 5763
rect 1676 5720 1728 5729
rect 4712 5763 4764 5772
rect 4712 5729 4721 5763
rect 4721 5729 4755 5763
rect 4755 5729 4764 5763
rect 4712 5720 4764 5729
rect 5540 5720 5592 5772
rect 7012 5720 7064 5772
rect 7840 5763 7892 5772
rect 7840 5729 7849 5763
rect 7849 5729 7883 5763
rect 7883 5729 7892 5763
rect 7840 5720 7892 5729
rect 9956 5720 10008 5772
rect 10048 5720 10100 5772
rect 12440 5763 12492 5772
rect 12440 5729 12449 5763
rect 12449 5729 12483 5763
rect 12483 5729 12492 5763
rect 12440 5720 12492 5729
rect 13912 5720 13964 5772
rect 15752 5763 15804 5772
rect 15752 5729 15761 5763
rect 15761 5729 15795 5763
rect 15795 5729 15804 5763
rect 15752 5720 15804 5729
rect 7104 5652 7156 5704
rect 1400 5584 1452 5636
rect 18604 5652 18656 5704
rect 19340 5652 19392 5704
rect 19432 5695 19484 5704
rect 19432 5661 19441 5695
rect 19441 5661 19475 5695
rect 19475 5661 19484 5695
rect 19432 5652 19484 5661
rect 17684 5584 17736 5636
rect 6552 5559 6604 5568
rect 6552 5525 6561 5559
rect 6561 5525 6595 5559
rect 6595 5525 6604 5559
rect 6552 5516 6604 5525
rect 9036 5516 9088 5568
rect 9864 5516 9916 5568
rect 13820 5516 13872 5568
rect 18512 5559 18564 5568
rect 18512 5525 18521 5559
rect 18521 5525 18555 5559
rect 18555 5525 18564 5559
rect 18512 5516 18564 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 4712 5312 4764 5364
rect 11060 5312 11112 5364
rect 12348 5312 12400 5364
rect 15752 5312 15804 5364
rect 15844 5355 15896 5364
rect 15844 5321 15853 5355
rect 15853 5321 15887 5355
rect 15887 5321 15896 5355
rect 15844 5312 15896 5321
rect 17776 5312 17828 5364
rect 19248 5312 19300 5364
rect 19340 5312 19392 5364
rect 12716 5244 12768 5296
rect 16764 5244 16816 5296
rect 4436 5176 4488 5228
rect 6276 5219 6328 5228
rect 3332 5040 3384 5092
rect 6276 5185 6285 5219
rect 6285 5185 6319 5219
rect 6319 5185 6328 5219
rect 6276 5176 6328 5185
rect 6552 5108 6604 5160
rect 6920 5176 6972 5228
rect 9680 5176 9732 5228
rect 11520 5219 11572 5228
rect 11520 5185 11529 5219
rect 11529 5185 11563 5219
rect 11563 5185 11572 5219
rect 11520 5176 11572 5185
rect 13084 5219 13136 5228
rect 13084 5185 13093 5219
rect 13093 5185 13127 5219
rect 13127 5185 13136 5219
rect 13084 5176 13136 5185
rect 14372 5176 14424 5228
rect 15292 5176 15344 5228
rect 16488 5219 16540 5228
rect 16488 5185 16497 5219
rect 16497 5185 16531 5219
rect 16531 5185 16540 5219
rect 16488 5176 16540 5185
rect 18512 5176 18564 5228
rect 18604 5219 18656 5228
rect 18604 5185 18613 5219
rect 18613 5185 18647 5219
rect 18647 5185 18656 5219
rect 18604 5176 18656 5185
rect 6092 5040 6144 5092
rect 8668 5151 8720 5160
rect 8668 5117 8677 5151
rect 8677 5117 8711 5151
rect 8711 5117 8720 5151
rect 8668 5108 8720 5117
rect 10968 5151 11020 5160
rect 10968 5117 10977 5151
rect 10977 5117 11011 5151
rect 11011 5117 11020 5151
rect 10968 5108 11020 5117
rect 11428 5108 11480 5160
rect 8116 5040 8168 5092
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 2044 5015 2096 5024
rect 2044 4981 2053 5015
rect 2053 4981 2087 5015
rect 2087 4981 2096 5015
rect 2044 4972 2096 4981
rect 4252 4972 4304 5024
rect 7840 4972 7892 5024
rect 9864 4972 9916 5024
rect 12716 5083 12768 5092
rect 12716 5049 12725 5083
rect 12725 5049 12759 5083
rect 12759 5049 12768 5083
rect 12716 5040 12768 5049
rect 13820 5040 13872 5092
rect 13636 5015 13688 5024
rect 13636 4981 13645 5015
rect 13645 4981 13679 5015
rect 13679 4981 13688 5015
rect 13636 4972 13688 4981
rect 13912 5015 13964 5024
rect 13912 4981 13921 5015
rect 13921 4981 13955 5015
rect 13955 4981 13964 5015
rect 13912 4972 13964 4981
rect 17960 5040 18012 5092
rect 19248 4972 19300 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1676 4768 1728 4820
rect 5540 4768 5592 4820
rect 11428 4768 11480 4820
rect 12716 4768 12768 4820
rect 13820 4768 13872 4820
rect 16488 4811 16540 4820
rect 16488 4777 16497 4811
rect 16497 4777 16531 4811
rect 16531 4777 16540 4811
rect 16488 4768 16540 4777
rect 17684 4811 17736 4820
rect 17684 4777 17693 4811
rect 17693 4777 17727 4811
rect 17727 4777 17736 4811
rect 17684 4768 17736 4777
rect 17960 4768 18012 4820
rect 18512 4768 18564 4820
rect 19340 4768 19392 4820
rect 20720 4768 20772 4820
rect 6092 4743 6144 4752
rect 6092 4709 6101 4743
rect 6101 4709 6135 4743
rect 6135 4709 6144 4743
rect 6092 4700 6144 4709
rect 7840 4700 7892 4752
rect 11336 4743 11388 4752
rect 11336 4709 11345 4743
rect 11345 4709 11379 4743
rect 11379 4709 11388 4743
rect 11336 4700 11388 4709
rect 16580 4700 16632 4752
rect 17408 4743 17460 4752
rect 17408 4709 17417 4743
rect 17417 4709 17451 4743
rect 17451 4709 17460 4743
rect 17408 4700 17460 4709
rect 1492 4675 1544 4684
rect 1492 4641 1510 4675
rect 1510 4641 1544 4675
rect 1492 4632 1544 4641
rect 2044 4632 2096 4684
rect 2504 4632 2556 4684
rect 4252 4632 4304 4684
rect 10784 4632 10836 4684
rect 12624 4632 12676 4684
rect 14372 4632 14424 4684
rect 15660 4632 15712 4684
rect 18420 4632 18472 4684
rect 19340 4675 19392 4684
rect 19340 4641 19358 4675
rect 19358 4641 19392 4675
rect 19340 4632 19392 4641
rect 21364 4675 21416 4684
rect 21364 4641 21382 4675
rect 21382 4641 21416 4675
rect 21364 4632 21416 4641
rect 6276 4564 6328 4616
rect 6920 4564 6972 4616
rect 7656 4564 7708 4616
rect 4712 4496 4764 4548
rect 7380 4539 7432 4548
rect 7380 4505 7389 4539
rect 7389 4505 7423 4539
rect 7423 4505 7432 4539
rect 10968 4564 11020 4616
rect 11612 4607 11664 4616
rect 11612 4573 11621 4607
rect 11621 4573 11655 4607
rect 11655 4573 11664 4607
rect 11612 4564 11664 4573
rect 12440 4564 12492 4616
rect 13084 4607 13136 4616
rect 7380 4496 7432 4505
rect 12348 4496 12400 4548
rect 13084 4573 13093 4607
rect 13093 4573 13127 4607
rect 13127 4573 13136 4607
rect 13084 4564 13136 4573
rect 16764 4607 16816 4616
rect 16764 4573 16773 4607
rect 16773 4573 16807 4607
rect 16807 4573 16816 4607
rect 16764 4564 16816 4573
rect 13820 4496 13872 4548
rect 16488 4496 16540 4548
rect 1952 4471 2004 4480
rect 1952 4437 1961 4471
rect 1961 4437 1995 4471
rect 1995 4437 2004 4471
rect 1952 4428 2004 4437
rect 2872 4471 2924 4480
rect 2872 4437 2881 4471
rect 2881 4437 2915 4471
rect 2915 4437 2924 4471
rect 2872 4428 2924 4437
rect 6552 4428 6604 4480
rect 7012 4471 7064 4480
rect 7012 4437 7021 4471
rect 7021 4437 7055 4471
rect 7055 4437 7064 4471
rect 7012 4428 7064 4437
rect 10876 4428 10928 4480
rect 11060 4428 11112 4480
rect 14464 4428 14516 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 2504 4267 2556 4276
rect 2504 4233 2513 4267
rect 2513 4233 2547 4267
rect 2547 4233 2556 4267
rect 2504 4224 2556 4233
rect 2872 4267 2924 4276
rect 2872 4233 2881 4267
rect 2881 4233 2915 4267
rect 2915 4233 2924 4267
rect 2872 4224 2924 4233
rect 6092 4224 6144 4276
rect 6276 4267 6328 4276
rect 6276 4233 6285 4267
rect 6285 4233 6319 4267
rect 6319 4233 6328 4267
rect 6276 4224 6328 4233
rect 7840 4267 7892 4276
rect 7840 4233 7849 4267
rect 7849 4233 7883 4267
rect 7883 4233 7892 4267
rect 7840 4224 7892 4233
rect 2044 4199 2096 4208
rect 2044 4165 2053 4199
rect 2053 4165 2087 4199
rect 2087 4165 2096 4199
rect 2044 4156 2096 4165
rect 8484 4156 8536 4208
rect 11060 4224 11112 4276
rect 11336 4224 11388 4276
rect 13820 4267 13872 4276
rect 13820 4233 13829 4267
rect 13829 4233 13863 4267
rect 13863 4233 13872 4267
rect 13820 4224 13872 4233
rect 14648 4224 14700 4276
rect 15660 4267 15712 4276
rect 15660 4233 15669 4267
rect 15669 4233 15703 4267
rect 15703 4233 15712 4267
rect 15660 4224 15712 4233
rect 16580 4224 16632 4276
rect 3884 4088 3936 4140
rect 4436 4131 4488 4140
rect 4436 4097 4445 4131
rect 4445 4097 4479 4131
rect 4479 4097 4488 4131
rect 4436 4088 4488 4097
rect 4712 4131 4764 4140
rect 4712 4097 4721 4131
rect 4721 4097 4755 4131
rect 4755 4097 4764 4131
rect 4712 4088 4764 4097
rect 4988 4131 5040 4140
rect 4988 4097 4997 4131
rect 4997 4097 5031 4131
rect 5031 4097 5040 4131
rect 4988 4088 5040 4097
rect 7380 4088 7432 4140
rect 1952 4020 2004 4072
rect 12348 4156 12400 4208
rect 13084 4199 13136 4208
rect 13084 4165 13093 4199
rect 13093 4165 13127 4199
rect 13127 4165 13136 4199
rect 13084 4156 13136 4165
rect 9772 4088 9824 4140
rect 10968 4088 11020 4140
rect 12624 4088 12676 4140
rect 3148 3995 3200 4004
rect 3148 3961 3157 3995
rect 3157 3961 3191 3995
rect 3191 3961 3200 3995
rect 3148 3952 3200 3961
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 2872 3884 2924 3936
rect 4528 3952 4580 4004
rect 7012 3995 7064 4004
rect 4436 3884 4488 3936
rect 7012 3961 7021 3995
rect 7021 3961 7055 3995
rect 7055 3961 7064 3995
rect 7012 3952 7064 3961
rect 6920 3884 6972 3936
rect 7196 3884 7248 3936
rect 7656 3884 7708 3936
rect 8208 3927 8260 3936
rect 8208 3893 8217 3927
rect 8217 3893 8251 3927
rect 8251 3893 8260 3927
rect 8208 3884 8260 3893
rect 9036 3884 9088 3936
rect 11336 4063 11388 4072
rect 11336 4029 11380 4063
rect 11380 4029 11388 4063
rect 11336 4020 11388 4029
rect 11980 4020 12032 4072
rect 17408 4156 17460 4208
rect 15108 4063 15160 4072
rect 15108 4029 15117 4063
rect 15117 4029 15151 4063
rect 15151 4029 15160 4063
rect 15108 4020 15160 4029
rect 16764 4088 16816 4140
rect 12532 3995 12584 4004
rect 12532 3961 12541 3995
rect 12541 3961 12575 3995
rect 12575 3961 12584 3995
rect 12532 3952 12584 3961
rect 9404 3884 9456 3936
rect 9680 3884 9732 3936
rect 10784 3884 10836 3936
rect 14832 3884 14884 3936
rect 16212 3884 16264 3936
rect 18420 3884 18472 3936
rect 18880 3884 18932 3936
rect 19340 3927 19392 3936
rect 19340 3893 19349 3927
rect 19349 3893 19383 3927
rect 19383 3893 19392 3927
rect 19340 3884 19392 3893
rect 21364 3927 21416 3936
rect 21364 3893 21373 3927
rect 21373 3893 21407 3927
rect 21407 3893 21416 3927
rect 21364 3884 21416 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1400 3680 1452 3732
rect 2228 3680 2280 3732
rect 3884 3680 3936 3732
rect 5540 3680 5592 3732
rect 9128 3680 9180 3732
rect 10968 3680 11020 3732
rect 12532 3723 12584 3732
rect 12532 3689 12541 3723
rect 12541 3689 12575 3723
rect 12575 3689 12584 3723
rect 12532 3680 12584 3689
rect 14740 3723 14792 3732
rect 14740 3689 14749 3723
rect 14749 3689 14783 3723
rect 14783 3689 14792 3723
rect 14740 3680 14792 3689
rect 15108 3680 15160 3732
rect 15292 3680 15344 3732
rect 3148 3612 3200 3664
rect 4252 3655 4304 3664
rect 4252 3621 4261 3655
rect 4261 3621 4295 3655
rect 4295 3621 4304 3655
rect 4252 3612 4304 3621
rect 4528 3612 4580 3664
rect 7104 3655 7156 3664
rect 7104 3621 7113 3655
rect 7113 3621 7147 3655
rect 7147 3621 7156 3655
rect 7104 3612 7156 3621
rect 12624 3612 12676 3664
rect 13176 3612 13228 3664
rect 5540 3544 5592 3596
rect 8944 3544 8996 3596
rect 9956 3587 10008 3596
rect 9956 3553 10000 3587
rect 10000 3553 10008 3587
rect 9956 3544 10008 3553
rect 11244 3544 11296 3596
rect 15660 3544 15712 3596
rect 16580 3587 16632 3596
rect 16580 3553 16589 3587
rect 16589 3553 16623 3587
rect 16623 3553 16632 3587
rect 16580 3544 16632 3553
rect 2412 3519 2464 3528
rect 2412 3485 2421 3519
rect 2421 3485 2455 3519
rect 2455 3485 2464 3519
rect 2412 3476 2464 3485
rect 4988 3476 5040 3528
rect 7012 3519 7064 3528
rect 7012 3485 7021 3519
rect 7021 3485 7055 3519
rect 7055 3485 7064 3519
rect 7012 3476 7064 3485
rect 7380 3519 7432 3528
rect 7380 3485 7389 3519
rect 7389 3485 7423 3519
rect 7423 3485 7432 3519
rect 7380 3476 7432 3485
rect 12808 3519 12860 3528
rect 12808 3485 12817 3519
rect 12817 3485 12851 3519
rect 12851 3485 12860 3519
rect 12808 3476 12860 3485
rect 12440 3408 12492 3460
rect 17868 3340 17920 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 3884 3136 3936 3188
rect 5540 3136 5592 3188
rect 7012 3136 7064 3188
rect 8944 3136 8996 3188
rect 12808 3136 12860 3188
rect 14556 3179 14608 3188
rect 14556 3145 14565 3179
rect 14565 3145 14599 3179
rect 14599 3145 14608 3179
rect 14556 3136 14608 3145
rect 15660 3179 15712 3188
rect 15660 3145 15669 3179
rect 15669 3145 15703 3179
rect 15703 3145 15712 3179
rect 15660 3136 15712 3145
rect 16580 3136 16632 3188
rect 17040 3179 17092 3188
rect 17040 3145 17049 3179
rect 17049 3145 17083 3179
rect 17083 3145 17092 3179
rect 17040 3136 17092 3145
rect 18696 3136 18748 3188
rect 4988 3068 5040 3120
rect 7104 3068 7156 3120
rect 9956 3111 10008 3120
rect 9956 3077 9965 3111
rect 9965 3077 9999 3111
rect 9999 3077 10008 3111
rect 9956 3068 10008 3077
rect 12164 3111 12216 3120
rect 12164 3077 12173 3111
rect 12173 3077 12207 3111
rect 12207 3077 12216 3111
rect 12164 3068 12216 3077
rect 13912 3068 13964 3120
rect 15936 3068 15988 3120
rect 2780 3043 2832 3052
rect 2780 3009 2789 3043
rect 2789 3009 2823 3043
rect 2823 3009 2832 3043
rect 2780 3000 2832 3009
rect 3148 3043 3200 3052
rect 3148 3009 3157 3043
rect 3157 3009 3191 3043
rect 3191 3009 3200 3043
rect 3148 3000 3200 3009
rect 4344 3043 4396 3052
rect 4344 3009 4353 3043
rect 4353 3009 4387 3043
rect 4387 3009 4396 3043
rect 4344 3000 4396 3009
rect 8208 3000 8260 3052
rect 11888 3043 11940 3052
rect 11888 3009 11897 3043
rect 11897 3009 11931 3043
rect 11931 3009 11940 3043
rect 11888 3000 11940 3009
rect 13176 3000 13228 3052
rect 1400 2975 1452 2984
rect 1400 2941 1409 2975
rect 1409 2941 1443 2975
rect 1443 2941 1452 2975
rect 1400 2932 1452 2941
rect 7380 2975 7432 2984
rect 7380 2941 7389 2975
rect 7389 2941 7423 2975
rect 7423 2941 7432 2975
rect 7380 2932 7432 2941
rect 11980 2932 12032 2984
rect 14556 2932 14608 2984
rect 1584 2839 1636 2848
rect 1584 2805 1593 2839
rect 1593 2805 1627 2839
rect 1627 2805 1636 2839
rect 1584 2796 1636 2805
rect 3148 2796 3200 2848
rect 8760 2864 8812 2916
rect 17040 2932 17092 2984
rect 19064 2907 19116 2916
rect 19064 2873 19073 2907
rect 19073 2873 19107 2907
rect 19107 2873 19116 2907
rect 19064 2864 19116 2873
rect 14924 2796 14976 2848
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 2688 2592 2740 2644
rect 2780 2592 2832 2644
rect 4252 2592 4304 2644
rect 4988 2635 5040 2644
rect 4988 2601 4997 2635
rect 4997 2601 5031 2635
rect 5031 2601 5040 2635
rect 4988 2592 5040 2601
rect 5080 2592 5132 2644
rect 6920 2592 6972 2644
rect 7196 2592 7248 2644
rect 13084 2592 13136 2644
rect 14464 2635 14516 2644
rect 14464 2601 14473 2635
rect 14473 2601 14507 2635
rect 14507 2601 14516 2635
rect 14464 2592 14516 2601
rect 18328 2592 18380 2644
rect 24676 2592 24728 2644
rect 3148 2567 3200 2576
rect 3148 2533 3157 2567
rect 3157 2533 3191 2567
rect 3191 2533 3200 2567
rect 3148 2524 3200 2533
rect 1952 2456 2004 2508
rect 3884 2456 3936 2508
rect 4160 2456 4212 2508
rect 10048 2456 10100 2508
rect 14280 2499 14332 2508
rect 14280 2465 14289 2499
rect 14289 2465 14323 2499
rect 14323 2465 14332 2499
rect 14280 2456 14332 2465
rect 16028 2499 16080 2508
rect 16028 2465 16037 2499
rect 16037 2465 16071 2499
rect 16071 2465 16080 2499
rect 16028 2456 16080 2465
rect 11796 2320 11848 2372
rect 18052 2320 18104 2372
rect 1952 2295 2004 2304
rect 1952 2261 1961 2295
rect 1961 2261 1995 2295
rect 1995 2261 2004 2295
rect 1952 2252 2004 2261
rect 12900 2252 12952 2304
rect 25136 2456 25188 2508
rect 21180 2252 21232 2304
rect 25136 2295 25188 2304
rect 25136 2261 25145 2295
rect 25145 2261 25179 2295
rect 25179 2261 25188 2295
rect 25136 2252 25188 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
<< metal2 >>
rect 478 27520 534 28000
rect 1490 27520 1546 28000
rect 2502 27520 2558 28000
rect 3514 27520 3570 28000
rect 4618 27520 4674 28000
rect 5630 27520 5686 28000
rect 6642 27520 6698 28000
rect 7654 27520 7710 28000
rect 8758 27520 8814 28000
rect 9770 27520 9826 28000
rect 10782 27520 10838 28000
rect 11794 27520 11850 28000
rect 12898 27520 12954 28000
rect 13910 27520 13966 28000
rect 14922 27520 14978 28000
rect 15934 27520 15990 28000
rect 17038 27520 17094 28000
rect 18050 27520 18106 28000
rect 19062 27520 19118 28000
rect 20074 27520 20130 28000
rect 21178 27520 21234 28000
rect 22190 27520 22246 28000
rect 23202 27520 23258 28000
rect 24214 27520 24270 28000
rect 25318 27520 25374 28000
rect 26330 27520 26386 28000
rect 27342 27520 27398 28000
rect 492 23662 520 27520
rect 1504 27418 1532 27520
rect 1504 27390 1624 27418
rect 480 23656 532 23662
rect 480 23598 532 23604
rect 1596 16046 1624 27390
rect 2516 23769 2544 27520
rect 2778 27296 2834 27305
rect 2778 27231 2834 27240
rect 2502 23760 2558 23769
rect 2502 23695 2558 23704
rect 2688 23656 2740 23662
rect 2686 23624 2688 23633
rect 2740 23624 2742 23633
rect 2686 23559 2742 23568
rect 1860 18216 1912 18222
rect 1860 18158 1912 18164
rect 1676 17808 1728 17814
rect 1676 17750 1728 17756
rect 1688 17338 1716 17750
rect 1676 17332 1728 17338
rect 1676 17274 1728 17280
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 1780 16697 1808 16934
rect 1766 16688 1822 16697
rect 1766 16623 1822 16632
rect 1584 16040 1636 16046
rect 1584 15982 1636 15988
rect 1768 16040 1820 16046
rect 1768 15982 1820 15988
rect 1400 14816 1452 14822
rect 1400 14758 1452 14764
rect 1412 13870 1440 14758
rect 1584 14000 1636 14006
rect 1584 13942 1636 13948
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1596 13297 1624 13942
rect 1582 13288 1638 13297
rect 1582 13223 1638 13232
rect 1492 13184 1544 13190
rect 1492 13126 1544 13132
rect 1400 12640 1452 12646
rect 1400 12582 1452 12588
rect 1412 10577 1440 12582
rect 1504 12306 1532 13126
rect 1584 12776 1636 12782
rect 1584 12718 1636 12724
rect 1596 12442 1624 12718
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1492 12300 1544 12306
rect 1492 12242 1544 12248
rect 1582 11928 1638 11937
rect 1582 11863 1584 11872
rect 1636 11863 1638 11872
rect 1584 11834 1636 11840
rect 1780 11370 1808 15982
rect 1872 11506 1900 18158
rect 2320 18080 2372 18086
rect 2320 18022 2372 18028
rect 2228 17740 2280 17746
rect 2228 17682 2280 17688
rect 2136 17536 2188 17542
rect 2136 17478 2188 17484
rect 2148 16726 2176 17478
rect 2240 16998 2268 17682
rect 2228 16992 2280 16998
rect 2228 16934 2280 16940
rect 2240 16726 2268 16934
rect 2136 16720 2188 16726
rect 2136 16662 2188 16668
rect 2228 16720 2280 16726
rect 2228 16662 2280 16668
rect 2148 15706 2176 16662
rect 2240 16250 2268 16662
rect 2228 16244 2280 16250
rect 2228 16186 2280 16192
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 2044 15428 2096 15434
rect 2044 15370 2096 15376
rect 2056 14618 2084 15370
rect 2044 14612 2096 14618
rect 2044 14554 2096 14560
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 1964 12209 1992 14350
rect 2056 13870 2084 14418
rect 2044 13864 2096 13870
rect 2042 13832 2044 13841
rect 2096 13832 2098 13841
rect 2042 13767 2098 13776
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 2056 12986 2084 13262
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2044 12980 2096 12986
rect 2044 12922 2096 12928
rect 2240 12782 2268 13126
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 1950 12200 2006 12209
rect 1950 12135 2006 12144
rect 1964 11694 1992 12135
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 1872 11478 1992 11506
rect 1596 11342 1808 11370
rect 1398 10568 1454 10577
rect 1398 10503 1454 10512
rect 1492 10532 1544 10538
rect 1492 10474 1544 10480
rect 1504 9110 1532 10474
rect 1596 9466 1624 11342
rect 1768 11212 1820 11218
rect 1768 11154 1820 11160
rect 1780 10266 1808 11154
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1674 9616 1730 9625
rect 1674 9551 1676 9560
rect 1728 9551 1730 9560
rect 1676 9522 1728 9528
rect 1596 9438 1716 9466
rect 1492 9104 1544 9110
rect 1492 9046 1544 9052
rect 1582 9072 1638 9081
rect 1582 9007 1638 9016
rect 1492 8968 1544 8974
rect 1492 8910 1544 8916
rect 1504 8090 1532 8910
rect 1596 8634 1624 9007
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1688 8514 1716 9438
rect 1768 9104 1820 9110
rect 1768 9046 1820 9052
rect 1780 8634 1808 9046
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1688 8486 1808 8514
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 1582 7712 1638 7721
rect 1582 7647 1638 7656
rect 1596 7546 1624 7647
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1412 7002 1440 7278
rect 1400 6996 1452 7002
rect 1400 6938 1452 6944
rect 1584 6384 1636 6390
rect 1582 6352 1584 6361
rect 1636 6352 1638 6361
rect 1582 6287 1638 6296
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1412 5642 1440 6190
rect 1674 6080 1730 6089
rect 1674 6015 1730 6024
rect 1688 5778 1716 6015
rect 1676 5772 1728 5778
rect 1676 5714 1728 5720
rect 1400 5636 1452 5642
rect 1400 5578 1452 5584
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 1596 4865 1624 4966
rect 1582 4856 1638 4865
rect 1688 4826 1716 5714
rect 1582 4791 1638 4800
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1492 4684 1544 4690
rect 1492 4626 1544 4632
rect 1400 3732 1452 3738
rect 1400 3674 1452 3680
rect 478 3088 534 3097
rect 478 3023 534 3032
rect 492 480 520 3023
rect 1412 2990 1440 3674
rect 1400 2984 1452 2990
rect 1400 2926 1452 2932
rect 1504 480 1532 4626
rect 1780 4185 1808 8486
rect 1964 8430 1992 11478
rect 2056 10606 2084 12038
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 2136 11688 2188 11694
rect 2136 11630 2188 11636
rect 2044 10600 2096 10606
rect 2044 10542 2096 10548
rect 2056 10266 2084 10542
rect 2148 10282 2176 11630
rect 2240 11218 2268 11698
rect 2228 11212 2280 11218
rect 2228 11154 2280 11160
rect 2044 10260 2096 10266
rect 2148 10254 2268 10282
rect 2044 10202 2096 10208
rect 2056 9450 2084 10202
rect 2134 10160 2190 10169
rect 2134 10095 2190 10104
rect 2148 10062 2176 10095
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2044 9444 2096 9450
rect 2044 9386 2096 9392
rect 1952 8424 2004 8430
rect 1952 8366 2004 8372
rect 1964 5896 1992 8366
rect 2056 8090 2084 9386
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 2148 7546 2176 9998
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 2148 6458 2176 6734
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 2148 5914 2176 6394
rect 2044 5908 2096 5914
rect 1964 5868 2044 5896
rect 2044 5850 2096 5856
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 2044 5024 2096 5030
rect 2042 4992 2044 5001
rect 2096 4992 2098 5001
rect 2042 4927 2098 4936
rect 2044 4684 2096 4690
rect 2044 4626 2096 4632
rect 1952 4480 2004 4486
rect 1952 4422 2004 4428
rect 1766 4176 1822 4185
rect 1766 4111 1822 4120
rect 1964 4078 1992 4422
rect 2056 4214 2084 4626
rect 2044 4208 2096 4214
rect 2044 4150 2096 4156
rect 1952 4072 2004 4078
rect 1950 4040 1952 4049
rect 2004 4040 2006 4049
rect 1950 3975 2006 3984
rect 1964 3949 1992 3975
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1596 3505 1624 3878
rect 2240 3738 2268 10254
rect 2332 9586 2360 18022
rect 2792 17898 2820 27231
rect 2962 25936 3018 25945
rect 2962 25871 3018 25880
rect 2976 24886 3004 25871
rect 2964 24880 3016 24886
rect 3528 24857 3556 27520
rect 2964 24822 3016 24828
rect 3514 24848 3570 24857
rect 3514 24783 3570 24792
rect 3330 24576 3386 24585
rect 3330 24511 3386 24520
rect 2872 23520 2924 23526
rect 2872 23462 2924 23468
rect 2700 17870 2820 17898
rect 2700 17814 2728 17870
rect 2688 17808 2740 17814
rect 2688 17750 2740 17756
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2700 17338 2728 17478
rect 2688 17332 2740 17338
rect 2688 17274 2740 17280
rect 2700 17066 2728 17274
rect 2884 17202 2912 23462
rect 3344 20505 3372 24511
rect 4632 23866 4660 27520
rect 5644 25242 5672 27520
rect 5552 25214 5672 25242
rect 4620 23860 4672 23866
rect 4620 23802 4672 23808
rect 3422 23080 3478 23089
rect 3422 23015 3478 23024
rect 3330 20496 3386 20505
rect 3330 20431 3386 20440
rect 3436 19281 3464 23015
rect 3882 20360 3938 20369
rect 3882 20295 3938 20304
rect 3422 19272 3478 19281
rect 3422 19207 3478 19216
rect 3896 18329 3924 20295
rect 3882 18320 3938 18329
rect 3882 18255 3938 18264
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5460 17202 5488 17682
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 3056 17196 3108 17202
rect 3056 17138 3108 17144
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 2688 17060 2740 17066
rect 2688 17002 2740 17008
rect 2884 16794 2912 17138
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2872 16516 2924 16522
rect 2872 16458 2924 16464
rect 2780 16176 2832 16182
rect 2780 16118 2832 16124
rect 2504 15632 2556 15638
rect 2502 15600 2504 15609
rect 2596 15632 2648 15638
rect 2556 15600 2558 15609
rect 2596 15574 2648 15580
rect 2502 15535 2558 15544
rect 2412 15360 2464 15366
rect 2412 15302 2464 15308
rect 2424 11694 2452 15302
rect 2516 14618 2544 15535
rect 2608 15162 2636 15574
rect 2596 15156 2648 15162
rect 2596 15098 2648 15104
rect 2792 15094 2820 16118
rect 2884 15978 2912 16458
rect 2872 15972 2924 15978
rect 2872 15914 2924 15920
rect 2884 15706 2912 15914
rect 2872 15700 2924 15706
rect 2872 15642 2924 15648
rect 3068 15609 3096 17138
rect 4160 16992 4212 16998
rect 4160 16934 4212 16940
rect 4172 16726 4200 16934
rect 4160 16720 4212 16726
rect 4160 16662 4212 16668
rect 4250 16688 4306 16697
rect 4172 16250 4200 16662
rect 4250 16623 4306 16632
rect 4264 16590 4292 16623
rect 4252 16584 4304 16590
rect 4252 16526 4304 16532
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 4264 16250 4292 16526
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 3148 16108 3200 16114
rect 3148 16050 3200 16056
rect 3160 15638 3188 16050
rect 3240 15972 3292 15978
rect 3240 15914 3292 15920
rect 4160 15972 4212 15978
rect 4160 15914 4212 15920
rect 3252 15638 3280 15914
rect 4172 15858 4200 15914
rect 4080 15830 4200 15858
rect 3148 15632 3200 15638
rect 3054 15600 3110 15609
rect 3148 15574 3200 15580
rect 3240 15632 3292 15638
rect 3240 15574 3292 15580
rect 3054 15535 3110 15544
rect 3160 15434 3188 15574
rect 3148 15428 3200 15434
rect 3148 15370 3200 15376
rect 4080 15094 4108 15830
rect 4356 15706 4384 16526
rect 4436 16448 4488 16454
rect 4436 16390 4488 16396
rect 4448 16114 4476 16390
rect 4436 16108 4488 16114
rect 4436 16050 4488 16056
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 4344 15700 4396 15706
rect 4344 15642 4396 15648
rect 4724 15609 4752 16050
rect 5080 15972 5132 15978
rect 5080 15914 5132 15920
rect 5092 15706 5120 15914
rect 5080 15700 5132 15706
rect 5080 15642 5132 15648
rect 4710 15600 4766 15609
rect 4160 15564 4212 15570
rect 4710 15535 4766 15544
rect 4160 15506 4212 15512
rect 4172 15162 4200 15506
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 2780 15088 2832 15094
rect 4068 15088 4120 15094
rect 2780 15030 2832 15036
rect 3974 15056 4030 15065
rect 2964 15020 3016 15026
rect 4068 15030 4120 15036
rect 3974 14991 3976 15000
rect 2964 14962 3016 14968
rect 4028 14991 4030 15000
rect 3976 14962 4028 14968
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 2700 14618 2728 14758
rect 2504 14612 2556 14618
rect 2504 14554 2556 14560
rect 2688 14612 2740 14618
rect 2688 14554 2740 14560
rect 2884 13734 2912 14758
rect 2976 14550 3004 14962
rect 3056 14952 3108 14958
rect 3056 14894 3108 14900
rect 2964 14544 3016 14550
rect 2964 14486 3016 14492
rect 2964 14408 3016 14414
rect 2962 14376 2964 14385
rect 3016 14376 3018 14385
rect 2962 14311 3018 14320
rect 2872 13728 2924 13734
rect 2872 13670 2924 13676
rect 2688 13456 2740 13462
rect 2688 13398 2740 13404
rect 2596 12708 2648 12714
rect 2596 12650 2648 12656
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2332 9110 2360 9522
rect 2320 9104 2372 9110
rect 2320 9046 2372 9052
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 2332 6866 2360 7346
rect 2424 6905 2452 11290
rect 2608 10198 2636 12650
rect 2700 12646 2728 13398
rect 2884 12714 2912 13670
rect 2872 12708 2924 12714
rect 2872 12650 2924 12656
rect 2688 12640 2740 12646
rect 2740 12600 2820 12628
rect 2688 12582 2740 12588
rect 2792 12442 2820 12600
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2872 12164 2924 12170
rect 2872 12106 2924 12112
rect 2884 11218 2912 12106
rect 2688 11212 2740 11218
rect 2688 11154 2740 11160
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2700 10470 2728 11154
rect 2688 10464 2740 10470
rect 2688 10406 2740 10412
rect 2596 10192 2648 10198
rect 2596 10134 2648 10140
rect 2608 9382 2636 10134
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2608 7274 2636 9318
rect 2884 9178 2912 11154
rect 3068 10470 3096 14894
rect 4172 14074 4200 15098
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4528 14476 4580 14482
rect 4528 14418 4580 14424
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4540 13870 4568 14418
rect 4068 13864 4120 13870
rect 4528 13864 4580 13870
rect 4120 13812 4200 13818
rect 4068 13806 4200 13812
rect 4528 13806 4580 13812
rect 4080 13790 4200 13806
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3528 12782 3556 13126
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3516 12776 3568 12782
rect 3514 12744 3516 12753
rect 3568 12744 3570 12753
rect 3514 12679 3570 12688
rect 3528 12653 3556 12679
rect 3896 12442 3924 12922
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 4080 11694 4108 12038
rect 4172 11830 4200 13790
rect 4540 13705 4568 13806
rect 4526 13696 4582 13705
rect 4526 13631 4582 13640
rect 4342 13560 4398 13569
rect 4342 13495 4398 13504
rect 4252 13456 4304 13462
rect 4252 13398 4304 13404
rect 4264 12986 4292 13398
rect 4356 13326 4384 13495
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4356 12442 4384 13262
rect 4632 12442 4660 14758
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 5080 14272 5132 14278
rect 5080 14214 5132 14220
rect 4724 13977 4752 14214
rect 4710 13968 4766 13977
rect 4710 13903 4766 13912
rect 5092 13870 5120 14214
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 5276 13802 5304 14962
rect 5356 14884 5408 14890
rect 5356 14826 5408 14832
rect 5368 14074 5396 14826
rect 5552 14362 5580 25214
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6550 24848 6606 24857
rect 6550 24783 6606 24792
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 6274 23760 6330 23769
rect 6274 23695 6330 23704
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 6184 17536 6236 17542
rect 6184 17478 6236 17484
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 6092 15904 6144 15910
rect 6092 15846 6144 15852
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 6104 15026 6132 15846
rect 6092 15020 6144 15026
rect 6092 14962 6144 14968
rect 6000 14884 6052 14890
rect 6000 14826 6052 14832
rect 6012 14414 6040 14826
rect 5460 14334 5580 14362
rect 6000 14408 6052 14414
rect 6000 14350 6052 14356
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5264 13796 5316 13802
rect 5264 13738 5316 13744
rect 4894 13288 4950 13297
rect 4894 13223 4950 13232
rect 4908 12986 4936 13223
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 4724 12345 4752 12718
rect 5172 12640 5224 12646
rect 5172 12582 5224 12588
rect 4710 12336 4766 12345
rect 4710 12271 4766 12280
rect 4896 12232 4948 12238
rect 4894 12200 4896 12209
rect 4948 12200 4950 12209
rect 4894 12135 4950 12144
rect 4160 11824 4212 11830
rect 4160 11766 4212 11772
rect 5184 11762 5212 12582
rect 5460 12322 5488 14334
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5552 12442 5580 14214
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 5724 13796 5776 13802
rect 5724 13738 5776 13744
rect 5736 13530 5764 13738
rect 6012 13569 6040 14350
rect 5998 13560 6054 13569
rect 5724 13524 5776 13530
rect 5998 13495 6054 13504
rect 5724 13466 5776 13472
rect 6196 13394 6224 17478
rect 6288 17377 6316 23695
rect 6564 17746 6592 24783
rect 6656 19446 6684 27520
rect 7564 23520 7616 23526
rect 7564 23462 7616 23468
rect 6644 19440 6696 19446
rect 6644 19382 6696 19388
rect 7010 18864 7066 18873
rect 7010 18799 7066 18808
rect 7024 18222 7052 18799
rect 7012 18216 7064 18222
rect 7012 18158 7064 18164
rect 7196 18080 7248 18086
rect 7196 18022 7248 18028
rect 6552 17740 6604 17746
rect 6552 17682 6604 17688
rect 6736 17740 6788 17746
rect 6736 17682 6788 17688
rect 6368 17536 6420 17542
rect 6368 17478 6420 17484
rect 6274 17368 6330 17377
rect 6274 17303 6276 17312
rect 6328 17303 6330 17312
rect 6276 17274 6328 17280
rect 6288 17134 6316 17274
rect 6276 17128 6328 17134
rect 6276 17070 6328 17076
rect 6380 14929 6408 17478
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6460 16584 6512 16590
rect 6460 16526 6512 16532
rect 6472 15638 6500 16526
rect 6460 15632 6512 15638
rect 6460 15574 6512 15580
rect 6552 15632 6604 15638
rect 6552 15574 6604 15580
rect 6366 14920 6422 14929
rect 6366 14855 6422 14864
rect 6472 14618 6500 15574
rect 6564 15162 6592 15574
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6276 14544 6328 14550
rect 6276 14486 6328 14492
rect 6288 14006 6316 14486
rect 6276 14000 6328 14006
rect 6276 13942 6328 13948
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6092 13320 6144 13326
rect 6092 13262 6144 13268
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5908 12912 5960 12918
rect 5908 12854 5960 12860
rect 5920 12442 5948 12854
rect 5998 12744 6054 12753
rect 5998 12679 6054 12688
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 5368 12306 5488 12322
rect 5356 12300 5488 12306
rect 5408 12294 5488 12300
rect 5356 12242 5408 12248
rect 5356 12164 5408 12170
rect 5356 12106 5408 12112
rect 5172 11756 5224 11762
rect 5172 11698 5224 11704
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 3436 11286 3464 11630
rect 3514 11384 3570 11393
rect 3514 11319 3570 11328
rect 3424 11280 3476 11286
rect 3424 11222 3476 11228
rect 3436 11121 3464 11222
rect 3422 11112 3478 11121
rect 3422 11047 3478 11056
rect 3436 10606 3464 11047
rect 3424 10600 3476 10606
rect 3424 10542 3476 10548
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 3056 10464 3108 10470
rect 3056 10406 3108 10412
rect 2976 9654 3004 10406
rect 3436 10266 3464 10542
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 3436 9518 3464 10202
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3238 9208 3294 9217
rect 2872 9172 2924 9178
rect 3238 9143 3294 9152
rect 2872 9114 2924 9120
rect 2872 8832 2924 8838
rect 2872 8774 2924 8780
rect 2884 8634 2912 8774
rect 3252 8634 3280 9143
rect 3528 9042 3556 11319
rect 3896 11082 3924 11630
rect 3884 11076 3936 11082
rect 3884 11018 3936 11024
rect 3896 10810 3924 11018
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 3896 9518 3924 10746
rect 4080 10713 4108 11630
rect 4540 11354 4568 11630
rect 5184 11393 5212 11698
rect 5170 11384 5226 11393
rect 4528 11348 4580 11354
rect 5368 11354 5396 12106
rect 5460 11694 5488 12294
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5552 11898 5580 12242
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5908 11824 5960 11830
rect 5908 11766 5960 11772
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5460 11393 5488 11630
rect 5446 11384 5502 11393
rect 5170 11319 5226 11328
rect 5356 11348 5408 11354
rect 4528 11290 4580 11296
rect 5446 11319 5502 11328
rect 5356 11290 5408 11296
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 4066 10704 4122 10713
rect 4066 10639 4122 10648
rect 4080 10606 4108 10639
rect 4172 10606 4200 10950
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 4080 10266 4108 10542
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 4264 9625 4292 11018
rect 4250 9616 4306 9625
rect 4250 9551 4306 9560
rect 4540 9518 4568 11290
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4632 10266 4660 11154
rect 5356 11144 5408 11150
rect 5920 11121 5948 11766
rect 6012 11354 6040 12679
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 6000 11212 6052 11218
rect 6104 11200 6132 13262
rect 6196 12918 6224 13330
rect 6184 12912 6236 12918
rect 6184 12854 6236 12860
rect 6274 12744 6330 12753
rect 6274 12679 6276 12688
rect 6328 12679 6330 12688
rect 6276 12650 6328 12656
rect 6380 12646 6408 13330
rect 6460 12776 6512 12782
rect 6460 12718 6512 12724
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6184 12436 6236 12442
rect 6184 12378 6236 12384
rect 6196 11218 6224 12378
rect 6274 12064 6330 12073
rect 6274 11999 6330 12008
rect 6288 11898 6316 11999
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 6288 11257 6316 11494
rect 6274 11248 6330 11257
rect 6052 11172 6132 11200
rect 6000 11154 6052 11160
rect 5356 11086 5408 11092
rect 5906 11112 5962 11121
rect 5368 10810 5396 11086
rect 6104 11082 6132 11172
rect 6184 11212 6236 11218
rect 6380 11218 6408 12582
rect 6472 12306 6500 12718
rect 6552 12708 6604 12714
rect 6552 12650 6604 12656
rect 6460 12300 6512 12306
rect 6460 12242 6512 12248
rect 6458 11384 6514 11393
rect 6458 11319 6514 11328
rect 6274 11183 6330 11192
rect 6368 11212 6420 11218
rect 6184 11154 6236 11160
rect 6368 11154 6420 11160
rect 5906 11047 5962 11056
rect 6092 11076 6144 11082
rect 6092 11018 6144 11024
rect 6104 10962 6132 11018
rect 6104 10934 6316 10962
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 4986 10704 5042 10713
rect 6288 10674 6316 10934
rect 6380 10810 6408 11154
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 4986 10639 5042 10648
rect 6276 10668 6328 10674
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 4528 9512 4580 9518
rect 4528 9454 4580 9460
rect 3896 9178 3924 9454
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 3700 9104 3752 9110
rect 3700 9046 3752 9052
rect 4252 9104 4304 9110
rect 4252 9046 4304 9052
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3528 8634 3556 8978
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3252 8430 3280 8570
rect 3240 8424 3292 8430
rect 3240 8366 3292 8372
rect 3056 7948 3108 7954
rect 3056 7890 3108 7896
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2596 7268 2648 7274
rect 2596 7210 2648 7216
rect 2504 6996 2556 7002
rect 2504 6938 2556 6944
rect 2410 6896 2466 6905
rect 2320 6860 2372 6866
rect 2410 6831 2466 6840
rect 2320 6802 2372 6808
rect 2516 5846 2544 6938
rect 2700 6934 2728 7686
rect 3068 7546 3096 7890
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 2688 6928 2740 6934
rect 2608 6876 2688 6882
rect 2608 6870 2740 6876
rect 2608 6854 2728 6870
rect 2608 6458 2636 6854
rect 2792 6746 2820 7482
rect 2962 6896 3018 6905
rect 3712 6866 3740 9046
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 4080 8430 4108 8978
rect 4264 8430 4292 9046
rect 4068 8424 4120 8430
rect 4252 8424 4304 8430
rect 4120 8372 4200 8378
rect 4068 8366 4200 8372
rect 4252 8366 4304 8372
rect 4080 8350 4200 8366
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3804 7410 3832 8230
rect 4172 8090 4200 8350
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 3884 7540 3936 7546
rect 3884 7482 3936 7488
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 3896 6934 3924 7482
rect 4356 7410 4384 9114
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 3884 6928 3936 6934
rect 3884 6870 3936 6876
rect 4252 6928 4304 6934
rect 4252 6870 4304 6876
rect 2962 6831 3018 6840
rect 3700 6860 3752 6866
rect 2700 6730 2820 6746
rect 2688 6724 2820 6730
rect 2740 6718 2820 6724
rect 2688 6666 2740 6672
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2976 6322 3004 6831
rect 3700 6802 3752 6808
rect 3516 6724 3568 6730
rect 3516 6666 3568 6672
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 2976 5914 3004 6258
rect 3332 6180 3384 6186
rect 3332 6122 3384 6128
rect 2964 5908 3016 5914
rect 2964 5850 3016 5856
rect 2504 5840 2556 5846
rect 2504 5782 2556 5788
rect 3344 5098 3372 6122
rect 3528 5914 3556 6666
rect 3712 6662 3740 6802
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 4172 6390 4200 6734
rect 4264 6458 4292 6870
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3332 5092 3384 5098
rect 3332 5034 3384 5040
rect 2504 4684 2556 4690
rect 2504 4626 2556 4632
rect 2516 4282 2544 4626
rect 2872 4480 2924 4486
rect 2872 4422 2924 4428
rect 2884 4282 2912 4422
rect 2504 4276 2556 4282
rect 2504 4218 2556 4224
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2884 3942 2912 4218
rect 3896 4146 3924 6054
rect 4448 5234 4476 9318
rect 4540 8906 4568 9454
rect 5000 9042 5028 10639
rect 6276 10610 6328 10616
rect 5264 10600 5316 10606
rect 5264 10542 5316 10548
rect 5276 9042 5304 10542
rect 6000 10532 6052 10538
rect 6000 10474 6052 10480
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5368 9042 5396 9862
rect 5552 9722 5580 10406
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 6012 9217 6040 10474
rect 6092 10260 6144 10266
rect 6092 10202 6144 10208
rect 6104 10169 6132 10202
rect 6090 10160 6146 10169
rect 6288 10130 6316 10610
rect 6090 10095 6146 10104
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6184 9920 6236 9926
rect 6184 9862 6236 9868
rect 6196 9382 6224 9862
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 5998 9208 6054 9217
rect 5998 9143 6054 9152
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 6000 9036 6052 9042
rect 6000 8978 6052 8984
rect 4528 8900 4580 8906
rect 4528 8842 4580 8848
rect 4896 8900 4948 8906
rect 4896 8842 4948 8848
rect 4908 8430 4936 8842
rect 5000 8498 5028 8978
rect 5276 8634 5304 8978
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 5000 8022 5028 8434
rect 6012 8430 6040 8978
rect 6092 8900 6144 8906
rect 6092 8842 6144 8848
rect 6104 8634 6132 8842
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 6000 8424 6052 8430
rect 6000 8366 6052 8372
rect 4988 8016 5040 8022
rect 4988 7958 5040 7964
rect 6012 7954 6040 8366
rect 6196 7954 6224 9318
rect 6380 9092 6408 10746
rect 6472 10418 6500 11319
rect 6564 11218 6592 12650
rect 6656 12238 6684 17138
rect 6748 16998 6776 17682
rect 6736 16992 6788 16998
rect 6736 16934 6788 16940
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6564 10538 6592 11154
rect 6642 10840 6698 10849
rect 6642 10775 6644 10784
rect 6696 10775 6698 10784
rect 6644 10746 6696 10752
rect 6656 10606 6684 10746
rect 6748 10690 6776 16934
rect 7012 16720 7064 16726
rect 7012 16662 7064 16668
rect 6920 16652 6972 16658
rect 6920 16594 6972 16600
rect 6828 15972 6880 15978
rect 6828 15914 6880 15920
rect 6840 15858 6868 15914
rect 6932 15858 6960 16594
rect 7024 15978 7052 16662
rect 7012 15972 7064 15978
rect 7012 15914 7064 15920
rect 7104 15972 7156 15978
rect 7104 15914 7156 15920
rect 6840 15830 7052 15858
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6932 14074 6960 14214
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 6932 13870 6960 14010
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6840 12782 6868 13670
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 7024 12442 7052 15830
rect 7116 15570 7144 15914
rect 7104 15564 7156 15570
rect 7104 15506 7156 15512
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 7116 14278 7144 14962
rect 7104 14272 7156 14278
rect 7104 14214 7156 14220
rect 7116 12646 7144 14214
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 6748 10662 6868 10690
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6552 10532 6604 10538
rect 6552 10474 6604 10480
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6472 10390 6592 10418
rect 6460 9104 6512 9110
rect 6380 9064 6460 9092
rect 6380 8634 6408 9064
rect 6460 9046 6512 9052
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6276 8560 6328 8566
rect 6276 8502 6328 8508
rect 6288 8022 6316 8502
rect 6276 8016 6328 8022
rect 6276 7958 6328 7964
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 4724 7206 4752 7890
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 5092 7002 5120 7346
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 4724 5778 4752 6122
rect 5276 5914 5304 6258
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 4724 5370 4752 5714
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 4264 4690 4292 4966
rect 4252 4684 4304 4690
rect 4252 4626 4304 4632
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 3160 3670 3188 3946
rect 3514 3768 3570 3777
rect 3896 3738 3924 4082
rect 3514 3703 3570 3712
rect 3884 3732 3936 3738
rect 3148 3664 3200 3670
rect 3148 3606 3200 3612
rect 2412 3528 2464 3534
rect 1582 3496 1638 3505
rect 1582 3431 1638 3440
rect 2410 3496 2412 3505
rect 2464 3496 2466 3505
rect 2410 3431 2466 3440
rect 3160 3058 3188 3606
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 2502 2816 2558 2825
rect 1596 2145 1624 2790
rect 2502 2751 2558 2760
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 1964 2310 1992 2450
rect 1952 2304 2004 2310
rect 1950 2272 1952 2281
rect 2004 2272 2006 2281
rect 1950 2207 2006 2216
rect 1582 2136 1638 2145
rect 1582 2071 1638 2080
rect 2516 480 2544 2751
rect 2686 2680 2742 2689
rect 2792 2650 2820 2994
rect 3148 2848 3200 2854
rect 3148 2790 3200 2796
rect 2686 2615 2688 2624
rect 2740 2615 2742 2624
rect 2780 2644 2832 2650
rect 2688 2586 2740 2592
rect 2780 2586 2832 2592
rect 3160 2582 3188 2790
rect 3148 2576 3200 2582
rect 3148 2518 3200 2524
rect 3528 480 3556 3703
rect 3884 3674 3936 3680
rect 3896 3194 3924 3674
rect 4264 3670 4292 4626
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 4724 4146 4752 4490
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4448 3942 4476 4082
rect 4528 4004 4580 4010
rect 4528 3946 4580 3952
rect 4436 3936 4488 3942
rect 4436 3878 4488 3884
rect 4540 3670 4568 3946
rect 4252 3664 4304 3670
rect 4252 3606 4304 3612
rect 4528 3664 4580 3670
rect 4528 3606 4580 3612
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3896 2514 3924 3130
rect 4264 2650 4292 3606
rect 5000 3534 5028 4082
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 5078 3496 5134 3505
rect 5000 3126 5028 3470
rect 5078 3431 5134 3440
rect 4988 3120 5040 3126
rect 4988 3062 5040 3068
rect 4344 3052 4396 3058
rect 4344 2994 4396 3000
rect 4356 2689 4384 2994
rect 4342 2680 4398 2689
rect 4252 2644 4304 2650
rect 5000 2650 5028 3062
rect 5092 2650 5120 3431
rect 4342 2615 4398 2624
rect 4988 2644 5040 2650
rect 4252 2586 4304 2592
rect 4988 2586 5040 2592
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 3884 2508 3936 2514
rect 3884 2450 3936 2456
rect 4160 2508 4212 2514
rect 4160 2450 4212 2456
rect 4172 2394 4200 2450
rect 4080 2366 4200 2394
rect 4080 785 4108 2366
rect 4618 2272 4674 2281
rect 4618 2207 4674 2216
rect 4066 776 4122 785
rect 4066 711 4122 720
rect 4632 480 4660 2207
rect 5368 1986 5396 7142
rect 5460 6186 5488 7142
rect 5552 6798 5580 7754
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 6092 6928 6144 6934
rect 6092 6870 6144 6876
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 5552 6458 5580 6734
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 6012 6390 6040 6734
rect 6000 6384 6052 6390
rect 6000 6326 6052 6332
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 6104 6118 6132 6870
rect 6196 6662 6224 7890
rect 6288 7478 6316 7958
rect 6380 7954 6408 8570
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6380 7546 6408 7890
rect 6368 7540 6420 7546
rect 6368 7482 6420 7488
rect 6276 7472 6328 7478
rect 6276 7414 6328 7420
rect 6276 7268 6328 7274
rect 6276 7210 6328 7216
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 5828 5846 5856 6054
rect 6288 5846 6316 7210
rect 6564 6361 6592 10390
rect 6748 10130 6776 10474
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 6748 9722 6776 10066
rect 6736 9716 6788 9722
rect 6736 9658 6788 9664
rect 6840 9466 6868 10662
rect 7024 10470 7052 10950
rect 7116 10810 7144 12242
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 7116 10713 7144 10746
rect 7102 10704 7158 10713
rect 7102 10639 7158 10648
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 7024 10130 7052 10406
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 6748 9438 6868 9466
rect 7104 9512 7156 9518
rect 7208 9489 7236 18022
rect 7576 17814 7604 23462
rect 7668 22114 7696 27520
rect 8772 23866 8800 27520
rect 9784 23882 9812 27520
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10138 24712 10194 24721
rect 10138 24647 10194 24656
rect 10152 24410 10180 24647
rect 10692 24608 10744 24614
rect 10692 24550 10744 24556
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 10140 24404 10192 24410
rect 10140 24346 10192 24352
rect 9956 24268 10008 24274
rect 9956 24210 10008 24216
rect 9600 23866 9812 23882
rect 8760 23860 8812 23866
rect 8760 23802 8812 23808
rect 9588 23860 9812 23866
rect 9640 23854 9812 23860
rect 9588 23802 9640 23808
rect 9770 23624 9826 23633
rect 9770 23559 9826 23568
rect 8852 23520 8904 23526
rect 8852 23462 8904 23468
rect 7668 22086 7880 22114
rect 7852 19378 7880 22086
rect 8300 21344 8352 21350
rect 8300 21286 8352 21292
rect 8312 21010 8340 21286
rect 8300 21004 8352 21010
rect 8300 20946 8352 20952
rect 8576 21004 8628 21010
rect 8576 20946 8628 20952
rect 8312 20262 8340 20946
rect 8588 20913 8616 20946
rect 8574 20904 8630 20913
rect 8574 20839 8630 20848
rect 8588 20602 8616 20839
rect 8576 20596 8628 20602
rect 8576 20538 8628 20544
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 8760 20256 8812 20262
rect 8760 20198 8812 20204
rect 8576 19916 8628 19922
rect 8576 19858 8628 19864
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 8114 19680 8170 19689
rect 8114 19615 8170 19624
rect 8128 19514 8156 19615
rect 8116 19508 8168 19514
rect 8116 19450 8168 19456
rect 8220 19417 8248 19790
rect 8206 19408 8262 19417
rect 7748 19372 7800 19378
rect 7668 19332 7748 19360
rect 7668 19009 7696 19332
rect 7748 19314 7800 19320
rect 7840 19372 7892 19378
rect 8588 19378 8616 19858
rect 8206 19343 8262 19352
rect 8576 19372 8628 19378
rect 7840 19314 7892 19320
rect 8576 19314 8628 19320
rect 7932 19304 7984 19310
rect 7746 19272 7802 19281
rect 8588 19281 8616 19314
rect 7932 19246 7984 19252
rect 8574 19272 8630 19281
rect 7746 19207 7802 19216
rect 7654 19000 7710 19009
rect 7654 18935 7710 18944
rect 7654 18864 7710 18873
rect 7760 18834 7788 19207
rect 7654 18799 7710 18808
rect 7748 18828 7800 18834
rect 7564 17808 7616 17814
rect 7564 17750 7616 17756
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 7484 16726 7512 17002
rect 7472 16720 7524 16726
rect 7472 16662 7524 16668
rect 7288 15972 7340 15978
rect 7288 15914 7340 15920
rect 7300 15434 7328 15914
rect 7288 15428 7340 15434
rect 7288 15370 7340 15376
rect 7300 15065 7328 15370
rect 7286 15056 7342 15065
rect 7286 14991 7342 15000
rect 7472 13388 7524 13394
rect 7472 13330 7524 13336
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7392 12782 7420 13126
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7378 12064 7434 12073
rect 7300 11898 7328 12038
rect 7378 11999 7434 12008
rect 7484 12050 7512 13330
rect 7564 12776 7616 12782
rect 7564 12718 7616 12724
rect 7576 12238 7604 12718
rect 7668 12458 7696 18799
rect 7748 18770 7800 18776
rect 7760 18714 7788 18770
rect 7760 18686 7880 18714
rect 7852 18426 7880 18686
rect 7840 18420 7892 18426
rect 7840 18362 7892 18368
rect 7840 17808 7892 17814
rect 7840 17750 7892 17756
rect 7852 17202 7880 17750
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 7840 16992 7892 16998
rect 7840 16934 7892 16940
rect 7852 16794 7880 16934
rect 7840 16788 7892 16794
rect 7840 16730 7892 16736
rect 7840 15564 7892 15570
rect 7840 15506 7892 15512
rect 7852 15162 7880 15506
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 7852 14618 7880 15098
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7944 14396 7972 19246
rect 8574 19207 8630 19216
rect 8484 18828 8536 18834
rect 8484 18770 8536 18776
rect 8206 18184 8262 18193
rect 8206 18119 8208 18128
rect 8260 18119 8262 18128
rect 8208 18090 8260 18096
rect 8496 18086 8524 18770
rect 8772 18630 8800 20198
rect 8668 18624 8720 18630
rect 8668 18566 8720 18572
rect 8760 18624 8812 18630
rect 8760 18566 8812 18572
rect 8484 18080 8536 18086
rect 8536 18028 8616 18034
rect 8484 18022 8616 18028
rect 8496 18006 8616 18022
rect 8024 17672 8076 17678
rect 8024 17614 8076 17620
rect 8036 17270 8064 17614
rect 8024 17264 8076 17270
rect 8024 17206 8076 17212
rect 8036 16250 8064 17206
rect 8024 16244 8076 16250
rect 8024 16186 8076 16192
rect 8114 15464 8170 15473
rect 8114 15399 8170 15408
rect 8128 15366 8156 15399
rect 8116 15360 8168 15366
rect 8116 15302 8168 15308
rect 8128 14550 8156 15302
rect 8484 14884 8536 14890
rect 8484 14826 8536 14832
rect 8116 14544 8168 14550
rect 8116 14486 8168 14492
rect 8208 14544 8260 14550
rect 8208 14486 8260 14492
rect 7944 14368 8156 14396
rect 7932 13184 7984 13190
rect 7932 13126 7984 13132
rect 7944 12889 7972 13126
rect 7930 12880 7986 12889
rect 7930 12815 7986 12824
rect 7944 12782 7972 12815
rect 7932 12776 7984 12782
rect 7932 12718 7984 12724
rect 7668 12430 7742 12458
rect 7714 12424 7742 12430
rect 7714 12396 7788 12424
rect 7656 12300 7708 12306
rect 7656 12242 7708 12248
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7668 12050 7696 12242
rect 7484 12022 7696 12050
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7392 11098 7420 11999
rect 7484 11762 7512 12022
rect 7654 11928 7710 11937
rect 7654 11863 7656 11872
rect 7708 11863 7710 11872
rect 7656 11834 7708 11840
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7576 11218 7604 11698
rect 7668 11694 7696 11834
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7392 11070 7604 11098
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7104 9454 7156 9460
rect 7194 9480 7250 9489
rect 6550 6352 6606 6361
rect 6550 6287 6606 6296
rect 5816 5840 5868 5846
rect 5816 5782 5868 5788
rect 6276 5840 6328 5846
rect 6276 5782 6328 5788
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5552 4826 5580 5714
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6288 5234 6316 5782
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 6564 5166 6592 5510
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 6092 5092 6144 5098
rect 6092 5034 6144 5040
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 6104 4758 6132 5034
rect 6092 4752 6144 4758
rect 6092 4694 6144 4700
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6104 4282 6132 4694
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6288 4282 6316 4558
rect 6564 4486 6592 5102
rect 6552 4480 6604 4486
rect 6552 4422 6604 4428
rect 6092 4276 6144 4282
rect 6092 4218 6144 4224
rect 6276 4276 6328 4282
rect 6276 4218 6328 4224
rect 6748 4049 6776 9438
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6840 9042 6868 9318
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6840 8498 6868 8978
rect 7012 8900 7064 8906
rect 7012 8842 7064 8848
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6932 5914 6960 7754
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6932 5234 6960 5850
rect 7024 5778 7052 8842
rect 7116 8838 7144 9454
rect 7194 9415 7250 9424
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7116 8430 7144 8774
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 7116 7546 7144 8366
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 7392 6118 7420 9522
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 7012 5772 7064 5778
rect 7012 5714 7064 5720
rect 7104 5704 7156 5710
rect 7392 5681 7420 6054
rect 7104 5646 7156 5652
rect 7378 5672 7434 5681
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6826 4992 6882 5001
rect 6826 4927 6882 4936
rect 5538 4040 5594 4049
rect 5538 3975 5594 3984
rect 6734 4040 6790 4049
rect 6734 3975 6790 3984
rect 5552 3738 5580 3975
rect 6642 3904 6698 3913
rect 6642 3839 6698 3848
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5552 3194 5580 3538
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 5368 1958 5672 1986
rect 5644 480 5672 1958
rect 6656 480 6684 3839
rect 6840 3754 6868 4927
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6932 3942 6960 4558
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 7024 4010 7052 4422
rect 7012 4004 7064 4010
rect 7012 3946 7064 3952
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6840 3726 6960 3754
rect 6932 2650 6960 3726
rect 7116 3670 7144 5646
rect 7378 5607 7434 5616
rect 7380 4548 7432 4554
rect 7380 4490 7432 4496
rect 7392 4146 7420 4490
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7104 3664 7156 3670
rect 7104 3606 7156 3612
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 7024 3194 7052 3470
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 7116 3126 7144 3606
rect 7104 3120 7156 3126
rect 7104 3062 7156 3068
rect 7208 2650 7236 3878
rect 7392 3534 7420 4082
rect 7576 3754 7604 11070
rect 7760 9722 7788 12396
rect 7944 12374 7972 12718
rect 7932 12368 7984 12374
rect 7932 12310 7984 12316
rect 7932 11824 7984 11830
rect 7932 11766 7984 11772
rect 7944 11218 7972 11766
rect 7932 11212 7984 11218
rect 7932 11154 7984 11160
rect 7944 10266 7972 11154
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 7748 9716 7800 9722
rect 7748 9658 7800 9664
rect 7944 9518 7972 10066
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7852 8430 7880 9454
rect 7944 9042 7972 9454
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 7840 8424 7892 8430
rect 7760 8372 7840 8378
rect 7760 8366 7892 8372
rect 7760 8350 7880 8366
rect 7760 8090 7788 8350
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7852 6866 7880 8230
rect 8036 7410 8064 9318
rect 8128 7886 8156 14368
rect 8220 13870 8248 14486
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8208 13864 8260 13870
rect 8404 13841 8432 14350
rect 8496 14074 8524 14826
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8208 13806 8260 13812
rect 8390 13832 8446 13841
rect 8496 13802 8524 14010
rect 8390 13767 8446 13776
rect 8484 13796 8536 13802
rect 8484 13738 8536 13744
rect 8482 13696 8538 13705
rect 8482 13631 8538 13640
rect 8496 13530 8524 13631
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8588 12594 8616 18006
rect 8680 14056 8708 18566
rect 8864 16130 8892 23462
rect 9784 23118 9812 23559
rect 9968 23526 9996 24210
rect 10704 23866 10732 24550
rect 10692 23860 10744 23866
rect 10692 23802 10744 23808
rect 10796 23526 10824 27520
rect 11808 24721 11836 27520
rect 12532 24880 12584 24886
rect 12532 24822 12584 24828
rect 11794 24712 11850 24721
rect 11794 24647 11850 24656
rect 12072 24608 12124 24614
rect 12072 24550 12124 24556
rect 11704 24268 11756 24274
rect 11704 24210 11756 24216
rect 11716 23526 11744 24210
rect 9956 23520 10008 23526
rect 9956 23462 10008 23468
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 11336 23520 11388 23526
rect 11336 23462 11388 23468
rect 11704 23520 11756 23526
rect 11704 23462 11756 23468
rect 9864 23248 9916 23254
rect 9864 23190 9916 23196
rect 9772 23112 9824 23118
rect 9772 23054 9824 23060
rect 9784 22778 9812 23054
rect 9772 22772 9824 22778
rect 9772 22714 9824 22720
rect 9876 22438 9904 23190
rect 9864 22432 9916 22438
rect 9864 22374 9916 22380
rect 8944 21888 8996 21894
rect 8944 21830 8996 21836
rect 9128 21888 9180 21894
rect 9128 21830 9180 21836
rect 8956 21486 8984 21830
rect 9140 21554 9168 21830
rect 9876 21690 9904 22374
rect 9864 21684 9916 21690
rect 9864 21626 9916 21632
rect 9128 21548 9180 21554
rect 9128 21490 9180 21496
rect 8944 21480 8996 21486
rect 8942 21448 8944 21457
rect 9680 21480 9732 21486
rect 8996 21448 8998 21457
rect 9680 21422 9732 21428
rect 8942 21383 8998 21392
rect 9692 20806 9720 21422
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9692 20466 9720 20742
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9128 20392 9180 20398
rect 9128 20334 9180 20340
rect 9140 19854 9168 20334
rect 9128 19848 9180 19854
rect 9126 19816 9128 19825
rect 9180 19816 9182 19825
rect 9126 19751 9182 19760
rect 9404 19712 9456 19718
rect 9404 19654 9456 19660
rect 9220 19440 9272 19446
rect 9220 19382 9272 19388
rect 8944 19304 8996 19310
rect 8942 19272 8944 19281
rect 8996 19272 8998 19281
rect 8942 19207 8998 19216
rect 8864 16102 8984 16130
rect 8852 16040 8904 16046
rect 8852 15982 8904 15988
rect 8864 15162 8892 15982
rect 8956 15502 8984 16102
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 8852 15156 8904 15162
rect 8852 15098 8904 15104
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 8680 14028 8892 14056
rect 8668 13932 8720 13938
rect 8668 13874 8720 13880
rect 8588 12566 8651 12594
rect 8623 12424 8651 12566
rect 8588 12396 8651 12424
rect 8588 12356 8616 12396
rect 8496 12328 8616 12356
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8206 10976 8262 10985
rect 8206 10911 8262 10920
rect 8220 10606 8248 10911
rect 8312 10674 8340 11630
rect 8300 10668 8352 10674
rect 8300 10610 8352 10616
rect 8208 10600 8260 10606
rect 8208 10542 8260 10548
rect 8300 10532 8352 10538
rect 8300 10474 8352 10480
rect 8312 9926 8340 10474
rect 8300 9920 8352 9926
rect 8300 9862 8352 9868
rect 8312 8430 8340 9862
rect 8300 8424 8352 8430
rect 8220 8372 8300 8378
rect 8220 8366 8352 8372
rect 8220 8350 8340 8366
rect 8220 7954 8248 8350
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 8036 7002 8064 7346
rect 8116 7268 8168 7274
rect 8116 7210 8168 7216
rect 8024 6996 8076 7002
rect 8024 6938 8076 6944
rect 8128 6934 8156 7210
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 7840 6860 7892 6866
rect 7840 6802 7892 6808
rect 7852 6458 7880 6802
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 8128 6390 8156 6870
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7852 5030 7880 5714
rect 8128 5098 8156 6326
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7852 4758 7880 4966
rect 7840 4752 7892 4758
rect 7840 4694 7892 4700
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7668 3942 7696 4558
rect 7852 4282 7880 4694
rect 7840 4276 7892 4282
rect 7840 4218 7892 4224
rect 8496 4214 8524 12328
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8588 11694 8616 12174
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8588 11354 8616 11630
rect 8680 11558 8708 13874
rect 8760 13388 8812 13394
rect 8760 13330 8812 13336
rect 8772 13025 8800 13330
rect 8758 13016 8814 13025
rect 8758 12951 8760 12960
rect 8812 12951 8814 12960
rect 8760 12922 8812 12928
rect 8760 11620 8812 11626
rect 8760 11562 8812 11568
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8588 10266 8616 11290
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 8680 10713 8708 10950
rect 8666 10704 8722 10713
rect 8666 10639 8722 10648
rect 8680 10606 8708 10639
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8668 10124 8720 10130
rect 8668 10066 8720 10072
rect 8680 9178 8708 10066
rect 8772 9654 8800 11562
rect 8864 10577 8892 14028
rect 9048 13938 9076 14214
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 9036 13456 9088 13462
rect 9232 13433 9260 19382
rect 9416 19378 9444 19654
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 9416 18970 9444 19314
rect 9876 19174 9904 21626
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 9404 18964 9456 18970
rect 9404 18906 9456 18912
rect 9876 18902 9904 19110
rect 9864 18896 9916 18902
rect 9864 18838 9916 18844
rect 9588 18624 9640 18630
rect 9588 18566 9640 18572
rect 9310 18456 9366 18465
rect 9310 18391 9366 18400
rect 9324 18222 9352 18391
rect 9600 18222 9628 18566
rect 9876 18426 9904 18838
rect 9968 18834 9996 23462
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 11348 23254 11376 23462
rect 11336 23248 11388 23254
rect 11336 23190 11388 23196
rect 11428 23248 11480 23254
rect 11428 23190 11480 23196
rect 11244 23044 11296 23050
rect 11244 22986 11296 22992
rect 10876 22636 10928 22642
rect 10876 22578 10928 22584
rect 10692 22568 10744 22574
rect 10692 22510 10744 22516
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10704 21894 10732 22510
rect 10692 21888 10744 21894
rect 10692 21830 10744 21836
rect 10888 21418 10916 22578
rect 11152 22500 11204 22506
rect 11152 22442 11204 22448
rect 10876 21412 10928 21418
rect 10876 21354 10928 21360
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10888 21078 10916 21354
rect 10968 21140 11020 21146
rect 10968 21082 11020 21088
rect 10876 21072 10928 21078
rect 10876 21014 10928 21020
rect 10888 20602 10916 21014
rect 10876 20596 10928 20602
rect 10876 20538 10928 20544
rect 10980 20330 11008 21082
rect 11060 20936 11112 20942
rect 11060 20878 11112 20884
rect 11072 20602 11100 20878
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 10140 20324 10192 20330
rect 10140 20266 10192 20272
rect 10968 20324 11020 20330
rect 10968 20266 11020 20272
rect 10048 20256 10100 20262
rect 10048 20198 10100 20204
rect 10060 19514 10088 20198
rect 10152 19938 10180 20266
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10980 19990 11008 20266
rect 10968 19984 11020 19990
rect 10152 19910 10272 19938
rect 10968 19926 11020 19932
rect 10244 19718 10272 19910
rect 10232 19712 10284 19718
rect 10230 19680 10232 19689
rect 10284 19680 10286 19689
rect 10230 19615 10286 19624
rect 10048 19508 10100 19514
rect 10048 19450 10100 19456
rect 10414 19408 10470 19417
rect 10414 19343 10470 19352
rect 10428 19310 10456 19343
rect 10416 19304 10468 19310
rect 10416 19246 10468 19252
rect 11072 19174 11100 20402
rect 11164 19242 11192 22442
rect 11256 22166 11284 22986
rect 11440 22506 11468 23190
rect 11428 22500 11480 22506
rect 11428 22442 11480 22448
rect 11520 22432 11572 22438
rect 11520 22374 11572 22380
rect 11532 22166 11560 22374
rect 11244 22160 11296 22166
rect 11244 22102 11296 22108
rect 11520 22160 11572 22166
rect 11520 22102 11572 22108
rect 11256 21690 11284 22102
rect 11244 21684 11296 21690
rect 11244 21626 11296 21632
rect 11532 21554 11560 22102
rect 12084 22030 12112 24550
rect 12254 23760 12310 23769
rect 12254 23695 12256 23704
rect 12308 23695 12310 23704
rect 12256 23666 12308 23672
rect 12440 23520 12492 23526
rect 12440 23462 12492 23468
rect 12452 22556 12480 23462
rect 12544 22710 12572 24822
rect 12912 24410 12940 27520
rect 13820 25356 13872 25362
rect 13820 25298 13872 25304
rect 13832 24682 13860 25298
rect 13820 24676 13872 24682
rect 13820 24618 13872 24624
rect 13924 24426 13952 27520
rect 14936 25242 14964 27520
rect 14844 25214 14964 25242
rect 14188 25152 14240 25158
rect 14188 25094 14240 25100
rect 14094 24848 14150 24857
rect 14094 24783 14150 24792
rect 14108 24614 14136 24783
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 13740 24410 13952 24426
rect 12900 24404 12952 24410
rect 12900 24346 12952 24352
rect 13728 24404 13952 24410
rect 13780 24398 13952 24404
rect 13728 24346 13780 24352
rect 13912 24336 13964 24342
rect 13912 24278 13964 24284
rect 13544 24268 13596 24274
rect 13544 24210 13596 24216
rect 12624 24064 12676 24070
rect 12624 24006 12676 24012
rect 12636 23594 12664 24006
rect 12716 23656 12768 23662
rect 12716 23598 12768 23604
rect 12624 23588 12676 23594
rect 12624 23530 12676 23536
rect 12532 22704 12584 22710
rect 12532 22646 12584 22652
rect 12532 22568 12584 22574
rect 12452 22528 12532 22556
rect 12532 22510 12584 22516
rect 12072 22024 12124 22030
rect 12072 21966 12124 21972
rect 11886 21584 11942 21593
rect 11520 21548 11572 21554
rect 11886 21519 11942 21528
rect 11520 21490 11572 21496
rect 11900 21010 11928 21519
rect 11888 21004 11940 21010
rect 11888 20946 11940 20952
rect 11900 20602 11928 20946
rect 11978 20904 12034 20913
rect 11978 20839 12034 20848
rect 11888 20596 11940 20602
rect 11888 20538 11940 20544
rect 11992 19922 12020 20839
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 11336 19848 11388 19854
rect 11336 19790 11388 19796
rect 11348 19242 11376 19790
rect 11152 19236 11204 19242
rect 11152 19178 11204 19184
rect 11336 19236 11388 19242
rect 11336 19178 11388 19184
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 9956 18828 10008 18834
rect 9956 18770 10008 18776
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 9956 18624 10008 18630
rect 9956 18566 10008 18572
rect 9864 18420 9916 18426
rect 9864 18362 9916 18368
rect 9968 18290 9996 18566
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 9312 18216 9364 18222
rect 9312 18158 9364 18164
rect 9588 18216 9640 18222
rect 10060 18193 10088 18702
rect 9588 18158 9640 18164
rect 10046 18184 10102 18193
rect 9324 17882 9352 18158
rect 9312 17876 9364 17882
rect 9312 17818 9364 17824
rect 9496 15972 9548 15978
rect 9496 15914 9548 15920
rect 9508 15638 9536 15914
rect 9496 15632 9548 15638
rect 9496 15574 9548 15580
rect 9404 15496 9456 15502
rect 9600 15450 9628 18158
rect 10046 18119 10102 18128
rect 10060 17882 10088 18119
rect 10692 18080 10744 18086
rect 10692 18022 10744 18028
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10048 17876 10100 17882
rect 10048 17818 10100 17824
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 9968 16998 9996 17682
rect 10140 17536 10192 17542
rect 10140 17478 10192 17484
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 9772 15632 9824 15638
rect 9772 15574 9824 15580
rect 9404 15438 9456 15444
rect 9416 14618 9444 15438
rect 9508 15422 9628 15450
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9508 13977 9536 15422
rect 9784 15162 9812 15574
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 9600 14804 9628 14894
rect 9600 14776 9720 14804
rect 9494 13968 9550 13977
rect 9494 13903 9550 13912
rect 9036 13398 9088 13404
rect 9218 13424 9274 13433
rect 9048 12986 9076 13398
rect 9218 13359 9274 13368
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8956 11014 8984 12718
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9140 11694 9168 12038
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 8944 11008 8996 11014
rect 8944 10950 8996 10956
rect 8956 10674 8984 10950
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8850 10568 8906 10577
rect 8850 10503 8906 10512
rect 8956 9926 8984 10610
rect 9036 10532 9088 10538
rect 9036 10474 9088 10480
rect 8944 9920 8996 9926
rect 8944 9862 8996 9868
rect 8760 9648 8812 9654
rect 8760 9590 8812 9596
rect 8956 9178 8984 9862
rect 9048 9586 9076 10474
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9036 9580 9088 9586
rect 9036 9522 9088 9528
rect 9048 9178 9076 9522
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8772 8634 8800 8774
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 8680 7546 8708 7890
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8680 6848 8708 7482
rect 8944 7336 8996 7342
rect 8944 7278 8996 7284
rect 8680 6820 8800 6848
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8680 5166 8708 6598
rect 8772 6186 8800 6820
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8772 5914 8800 6122
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8484 4208 8536 4214
rect 8484 4150 8536 4156
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 7576 3726 7696 3754
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7378 3224 7434 3233
rect 7378 3159 7434 3168
rect 7392 2990 7420 3159
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 7392 2825 7420 2926
rect 7378 2816 7434 2825
rect 7378 2751 7434 2760
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7668 480 7696 3726
rect 8220 3058 8248 3878
rect 8956 3602 8984 7278
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 9048 5914 9076 6258
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 9048 3942 9076 5510
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 9140 3738 9168 9862
rect 9232 7342 9260 13359
rect 9692 12782 9720 14776
rect 9968 14770 9996 16934
rect 10152 16114 10180 17478
rect 10704 17066 10732 18022
rect 11072 17882 11100 19110
rect 11164 18970 11192 19178
rect 11152 18964 11204 18970
rect 11152 18906 11204 18912
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10980 17202 11008 17478
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 10692 17060 10744 17066
rect 10692 17002 10744 17008
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10704 16726 10732 17002
rect 10692 16720 10744 16726
rect 10612 16680 10692 16708
rect 10612 16250 10640 16680
rect 10692 16662 10744 16668
rect 10692 16584 10744 16590
rect 10692 16526 10744 16532
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 10600 16244 10652 16250
rect 10600 16186 10652 16192
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10704 15706 10732 16526
rect 10888 15978 10916 16526
rect 10876 15972 10928 15978
rect 10876 15914 10928 15920
rect 10692 15700 10744 15706
rect 10692 15642 10744 15648
rect 10048 15496 10100 15502
rect 10046 15464 10048 15473
rect 10100 15464 10102 15473
rect 10046 15399 10102 15408
rect 10060 15026 10088 15399
rect 10508 15088 10560 15094
rect 10508 15030 10560 15036
rect 10048 15020 10100 15026
rect 10048 14962 10100 14968
rect 10414 14920 10470 14929
rect 10520 14890 10548 15030
rect 10414 14855 10416 14864
rect 10468 14855 10470 14864
rect 10508 14884 10560 14890
rect 10416 14826 10468 14832
rect 10508 14826 10560 14832
rect 10692 14816 10744 14822
rect 10046 14784 10102 14793
rect 9968 14742 10046 14770
rect 10692 14758 10744 14764
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10046 14719 10102 14728
rect 9956 14544 10008 14550
rect 9956 14486 10008 14492
rect 9772 14408 9824 14414
rect 9770 14376 9772 14385
rect 9824 14376 9826 14385
rect 9770 14311 9826 14320
rect 9784 14074 9812 14311
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9968 13734 9996 14486
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 9784 13394 9812 13670
rect 9968 13530 9996 13670
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9692 12306 9720 12582
rect 9784 12322 9812 12922
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 9876 12442 9904 12718
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9956 12368 10008 12374
rect 9784 12306 9904 12322
rect 9956 12310 10008 12316
rect 9680 12300 9732 12306
rect 9784 12300 9916 12306
rect 9784 12294 9864 12300
rect 9680 12242 9732 12248
rect 9864 12242 9916 12248
rect 9876 11898 9904 12242
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9496 11688 9548 11694
rect 9494 11656 9496 11665
rect 9548 11656 9550 11665
rect 9968 11626 9996 12310
rect 9494 11591 9550 11600
rect 9956 11620 10008 11626
rect 9956 11562 10008 11568
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9692 10826 9720 11086
rect 9968 11082 9996 11562
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 9600 10810 9720 10826
rect 9968 10810 9996 11018
rect 9588 10804 9720 10810
rect 9640 10798 9720 10804
rect 9956 10804 10008 10810
rect 9588 10746 9640 10752
rect 9956 10746 10008 10752
rect 9600 10130 9628 10746
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9864 10532 9916 10538
rect 9864 10474 9916 10480
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9508 8430 9536 9386
rect 9876 9110 9904 10474
rect 9968 10198 9996 10542
rect 9956 10192 10008 10198
rect 9956 10134 10008 10140
rect 9968 9722 9996 10134
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9220 7200 9272 7206
rect 9220 7142 9272 7148
rect 9232 7002 9260 7142
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 9232 6662 9260 6938
rect 9324 6934 9352 7822
rect 9312 6928 9364 6934
rect 9312 6870 9364 6876
rect 9416 6798 9444 8298
rect 9508 7478 9536 8366
rect 9588 7744 9640 7750
rect 9784 7732 9812 8910
rect 9876 8634 9904 9046
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 10060 7954 10088 14719
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10704 14618 10732 14758
rect 10692 14612 10744 14618
rect 10692 14554 10744 14560
rect 10600 14000 10652 14006
rect 10598 13968 10600 13977
rect 10652 13968 10654 13977
rect 10598 13903 10654 13912
rect 10796 13870 10824 14758
rect 10980 13938 11008 17138
rect 11072 16794 11100 17818
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 11072 16182 11100 16730
rect 11164 16658 11192 18906
rect 11348 18766 11376 19178
rect 11992 19174 12020 19858
rect 11980 19168 12032 19174
rect 11980 19110 12032 19116
rect 11888 18896 11940 18902
rect 11888 18838 11940 18844
rect 11336 18760 11388 18766
rect 11336 18702 11388 18708
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11520 17808 11572 17814
rect 11520 17750 11572 17756
rect 11532 17338 11560 17750
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 11612 16176 11664 16182
rect 11612 16118 11664 16124
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11256 14822 11284 15506
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11428 14408 11480 14414
rect 11428 14350 11480 14356
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10876 13864 10928 13870
rect 10876 13806 10928 13812
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10888 13530 10916 13806
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 10152 12782 10180 13126
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 10152 12442 10180 12718
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10888 12442 10916 13330
rect 11440 13326 11468 14350
rect 11624 13870 11652 16118
rect 11716 14482 11744 18566
rect 11808 17678 11836 18702
rect 11900 18426 11928 18838
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11796 17672 11848 17678
rect 11796 17614 11848 17620
rect 11794 15736 11850 15745
rect 11794 15671 11850 15680
rect 11808 15570 11836 15671
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 11808 15162 11836 15506
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11612 13864 11664 13870
rect 11612 13806 11664 13812
rect 11716 13734 11744 14418
rect 11992 13870 12020 19110
rect 12084 18766 12112 21966
rect 12440 20800 12492 20806
rect 12440 20742 12492 20748
rect 12348 20596 12400 20602
rect 12348 20538 12400 20544
rect 12256 19372 12308 19378
rect 12256 19314 12308 19320
rect 12164 19236 12216 19242
rect 12164 19178 12216 19184
rect 12072 18760 12124 18766
rect 12072 18702 12124 18708
rect 12084 17814 12112 18702
rect 12176 18290 12204 19178
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 12072 17808 12124 17814
rect 12072 17750 12124 17756
rect 11980 13864 12032 13870
rect 11980 13806 12032 13812
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11428 13320 11480 13326
rect 11426 13288 11428 13297
rect 11480 13288 11482 13297
rect 11426 13223 11482 13232
rect 11518 13016 11574 13025
rect 11716 12986 11744 13330
rect 11518 12951 11574 12960
rect 11704 12980 11756 12986
rect 11058 12744 11114 12753
rect 11058 12679 11114 12688
rect 10140 12436 10192 12442
rect 10140 12378 10192 12384
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10322 12336 10378 12345
rect 10140 12300 10192 12306
rect 10322 12271 10378 12280
rect 10140 12242 10192 12248
rect 10152 11354 10180 12242
rect 10336 12238 10364 12271
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10966 11792 11022 11801
rect 10966 11727 11022 11736
rect 10980 11694 11008 11727
rect 10968 11688 11020 11694
rect 10888 11648 10968 11676
rect 10692 11552 10744 11558
rect 10692 11494 10744 11500
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10704 11150 10732 11494
rect 10888 11234 10916 11648
rect 10968 11630 11020 11636
rect 11072 11354 11100 12679
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 10796 11206 10916 11234
rect 10966 11248 11022 11257
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 10796 10985 10824 11206
rect 10966 11183 10968 11192
rect 11020 11183 11022 11192
rect 10968 11154 11020 11160
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10782 10976 10838 10985
rect 10782 10911 10838 10920
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 10152 9625 10180 9998
rect 10138 9616 10194 9625
rect 10138 9551 10194 9560
rect 10152 8974 10180 9551
rect 10796 9450 10824 10911
rect 10784 9444 10836 9450
rect 10784 9386 10836 9392
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10598 8528 10654 8537
rect 10598 8463 10600 8472
rect 10652 8463 10654 8472
rect 10600 8434 10652 8440
rect 10612 8378 10640 8434
rect 10888 8401 10916 11086
rect 10980 10810 11008 11154
rect 11428 11008 11480 11014
rect 11428 10950 11480 10956
rect 11440 10810 11468 10950
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 10980 9722 11008 10746
rect 11058 10568 11114 10577
rect 11058 10503 11114 10512
rect 11072 10266 11100 10503
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 11072 10062 11100 10202
rect 11428 10192 11480 10198
rect 11428 10134 11480 10140
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 10966 9208 11022 9217
rect 11440 9178 11468 10134
rect 11532 9586 11560 12951
rect 11704 12922 11756 12928
rect 11716 12753 11744 12922
rect 11980 12776 12032 12782
rect 11702 12744 11758 12753
rect 11980 12718 12032 12724
rect 11702 12679 11758 12688
rect 11716 12170 11744 12679
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11704 12164 11756 12170
rect 11704 12106 11756 12112
rect 11808 12050 11836 12242
rect 11716 12022 11836 12050
rect 11716 11626 11744 12022
rect 11704 11620 11756 11626
rect 11704 11562 11756 11568
rect 11716 11218 11744 11562
rect 11992 11218 12020 12718
rect 12164 12232 12216 12238
rect 12164 12174 12216 12180
rect 12072 12164 12124 12170
rect 12072 12106 12124 12112
rect 12084 11558 12112 12106
rect 12176 11937 12204 12174
rect 12162 11928 12218 11937
rect 12162 11863 12218 11872
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 11704 11212 11756 11218
rect 11704 11154 11756 11160
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 11992 10810 12020 11154
rect 12084 11082 12112 11494
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 12084 10810 12112 11018
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 10966 9143 11022 9152
rect 11428 9172 11480 9178
rect 10874 8392 10930 8401
rect 10612 8350 10732 8378
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10704 8090 10732 8350
rect 10874 8327 10930 8336
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10048 7948 10100 7954
rect 10048 7890 10100 7896
rect 9640 7704 9812 7732
rect 9588 7686 9640 7692
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9680 7268 9732 7274
rect 9680 7210 9732 7216
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9312 6724 9364 6730
rect 9312 6666 9364 6672
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9324 6186 9352 6666
rect 9508 6662 9536 7142
rect 9692 7002 9720 7210
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9312 6180 9364 6186
rect 9312 6122 9364 6128
rect 9324 6089 9352 6122
rect 9310 6080 9366 6089
rect 9310 6015 9366 6024
rect 9508 5914 9536 6598
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9692 5234 9720 6054
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9784 4146 9812 7704
rect 10060 7546 10088 7890
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 9864 6928 9916 6934
rect 9864 6870 9916 6876
rect 9876 6458 9904 6870
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9954 6216 10010 6225
rect 9864 6180 9916 6186
rect 9954 6151 10010 6160
rect 9864 6122 9916 6128
rect 9876 5574 9904 6122
rect 9968 5778 9996 6151
rect 10060 5778 10088 6734
rect 10152 5914 10180 7686
rect 10692 7268 10744 7274
rect 10692 7210 10744 7216
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10704 6322 10732 7210
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 9968 5386 9996 5714
rect 9876 5358 9996 5386
rect 9876 5030 9904 5358
rect 10980 5166 11008 9143
rect 11428 9114 11480 9120
rect 11440 8634 11468 9114
rect 11796 9104 11848 9110
rect 11796 9046 11848 9052
rect 11428 8628 11480 8634
rect 11428 8570 11480 8576
rect 11150 8256 11206 8265
rect 11150 8191 11206 8200
rect 11164 7954 11192 8191
rect 11440 8106 11468 8570
rect 11808 8362 11836 9046
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11796 8356 11848 8362
rect 11796 8298 11848 8304
rect 11348 8078 11468 8106
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 11164 7546 11192 7890
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11072 5846 11100 6598
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 11072 5370 11100 5782
rect 11242 5672 11298 5681
rect 11242 5607 11298 5616
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 10968 5160 11020 5166
rect 11072 5137 11100 5306
rect 10968 5102 11020 5108
rect 11058 5128 11114 5137
rect 11058 5063 11114 5072
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9404 3936 9456 3942
rect 9680 3936 9732 3942
rect 9404 3878 9456 3884
rect 9678 3904 9680 3913
rect 9732 3904 9734 3913
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 8956 3194 8984 3538
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8956 2961 8984 3130
rect 8942 2952 8998 2961
rect 8760 2916 8812 2922
rect 8942 2887 8998 2896
rect 8760 2858 8812 2864
rect 8772 480 8800 2858
rect 9416 2530 9444 3878
rect 9678 3839 9734 3848
rect 9876 3777 9904 4966
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 10046 4176 10102 4185
rect 10046 4111 10102 4120
rect 9862 3768 9918 3777
rect 9862 3703 9918 3712
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9968 3126 9996 3538
rect 9956 3120 10008 3126
rect 9954 3088 9956 3097
rect 10008 3088 10010 3097
rect 9954 3023 10010 3032
rect 9416 2502 9812 2530
rect 10060 2514 10088 4111
rect 10796 3942 10824 4626
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 10876 4480 10928 4486
rect 10876 4422 10928 4428
rect 10784 3936 10836 3942
rect 10782 3904 10784 3913
rect 10836 3904 10838 3913
rect 10289 3836 10585 3856
rect 10782 3839 10838 3848
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 9784 480 9812 2502
rect 10048 2508 10100 2514
rect 10048 2450 10100 2456
rect 10888 2258 10916 4422
rect 10980 4146 11008 4558
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11072 4282 11100 4422
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 10980 3738 11008 4082
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 11256 3641 11284 5607
rect 11348 4758 11376 8078
rect 11808 8022 11836 8298
rect 11900 8090 11928 8978
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11796 8016 11848 8022
rect 11796 7958 11848 7964
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 11440 7002 11468 7890
rect 11808 7546 11836 7958
rect 11796 7540 11848 7546
rect 11716 7500 11796 7528
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11440 5166 11468 6938
rect 11716 6934 11744 7500
rect 11796 7482 11848 7488
rect 12268 7290 12296 19314
rect 12360 16833 12388 20538
rect 12452 19854 12480 20742
rect 12440 19848 12492 19854
rect 12440 19790 12492 19796
rect 12544 19378 12572 22510
rect 12636 19922 12664 23530
rect 12728 22982 12756 23598
rect 13268 23588 13320 23594
rect 13268 23530 13320 23536
rect 13280 23322 13308 23530
rect 13556 23526 13584 24210
rect 13544 23520 13596 23526
rect 13544 23462 13596 23468
rect 13268 23316 13320 23322
rect 13268 23258 13320 23264
rect 12992 23248 13044 23254
rect 12898 23216 12954 23225
rect 12992 23190 13044 23196
rect 12898 23151 12954 23160
rect 12912 23118 12940 23151
rect 12900 23112 12952 23118
rect 12900 23054 12952 23060
rect 12716 22976 12768 22982
rect 12716 22918 12768 22924
rect 12912 22778 12940 23054
rect 12900 22772 12952 22778
rect 12900 22714 12952 22720
rect 12716 22704 12768 22710
rect 12768 22652 12940 22658
rect 12716 22646 12940 22652
rect 12728 22630 12940 22646
rect 12716 22432 12768 22438
rect 12716 22374 12768 22380
rect 12728 22012 12756 22374
rect 12808 22024 12860 22030
rect 12728 21984 12808 22012
rect 12808 21966 12860 21972
rect 12820 21690 12848 21966
rect 12808 21684 12860 21690
rect 12808 21626 12860 21632
rect 12912 21486 12940 22630
rect 13004 22234 13032 23190
rect 13084 22976 13136 22982
rect 13084 22918 13136 22924
rect 12992 22228 13044 22234
rect 12992 22170 13044 22176
rect 12900 21480 12952 21486
rect 12900 21422 12952 21428
rect 13004 21146 13032 22170
rect 13096 21457 13124 22918
rect 13082 21448 13138 21457
rect 13082 21383 13138 21392
rect 13452 21344 13504 21350
rect 13450 21312 13452 21321
rect 13504 21312 13506 21321
rect 13450 21247 13506 21256
rect 12992 21140 13044 21146
rect 12992 21082 13044 21088
rect 13084 21072 13136 21078
rect 13084 21014 13136 21020
rect 12808 20392 12860 20398
rect 12808 20334 12860 20340
rect 12820 19990 12848 20334
rect 13096 20262 13124 21014
rect 13176 20936 13228 20942
rect 13176 20878 13228 20884
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 12808 19984 12860 19990
rect 12808 19926 12860 19932
rect 12624 19916 12676 19922
rect 12624 19858 12676 19864
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 12532 19236 12584 19242
rect 12636 19224 12664 19858
rect 12898 19816 12954 19825
rect 12898 19751 12954 19760
rect 12806 19408 12862 19417
rect 12806 19343 12862 19352
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 12584 19196 12664 19224
rect 12532 19178 12584 19184
rect 12728 18630 12756 19246
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 12636 17338 12664 18226
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 12346 16824 12402 16833
rect 12636 16794 12664 17274
rect 12346 16759 12402 16768
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12716 16176 12768 16182
rect 12716 16118 12768 16124
rect 12728 16046 12756 16118
rect 12716 16040 12768 16046
rect 12716 15982 12768 15988
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12452 12442 12480 13262
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12452 11830 12480 12378
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12348 9036 12400 9042
rect 12452 9024 12480 10202
rect 12636 10130 12664 13670
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12728 12306 12756 12582
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12728 11694 12756 12242
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12728 11354 12756 11630
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12544 9722 12572 9998
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12544 9489 12572 9522
rect 12530 9480 12586 9489
rect 12530 9415 12586 9424
rect 12624 9444 12676 9450
rect 12624 9386 12676 9392
rect 12636 9178 12664 9386
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12400 8996 12480 9024
rect 12348 8978 12400 8984
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12084 7262 12296 7290
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11704 6928 11756 6934
rect 11704 6870 11756 6876
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11532 6118 11560 6734
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11532 5234 11560 6054
rect 11624 5846 11652 6734
rect 11716 6458 11744 6870
rect 11808 6662 11836 7142
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11612 5840 11664 5846
rect 11612 5782 11664 5788
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11428 5160 11480 5166
rect 11428 5102 11480 5108
rect 11440 4826 11468 5102
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11336 4752 11388 4758
rect 11336 4694 11388 4700
rect 11348 4282 11376 4694
rect 11624 4622 11652 5782
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 11336 4072 11388 4078
rect 11334 4040 11336 4049
rect 11980 4072 12032 4078
rect 11388 4040 11390 4049
rect 11980 4014 12032 4020
rect 11334 3975 11390 3984
rect 11242 3632 11298 3641
rect 11242 3567 11244 3576
rect 11296 3567 11298 3576
rect 11244 3538 11296 3544
rect 11256 3507 11284 3538
rect 11886 3088 11942 3097
rect 11886 3023 11888 3032
rect 11940 3023 11942 3032
rect 11888 2994 11940 3000
rect 11992 2990 12020 4014
rect 12084 3233 12112 7262
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12268 6662 12296 7142
rect 12360 6934 12388 7822
rect 12532 7268 12584 7274
rect 12532 7210 12584 7216
rect 12544 7002 12572 7210
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12348 6928 12400 6934
rect 12348 6870 12400 6876
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12360 6322 12388 6870
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12438 5808 12494 5817
rect 12438 5743 12440 5752
rect 12492 5743 12494 5752
rect 12440 5714 12492 5720
rect 12452 5556 12480 5714
rect 12360 5528 12480 5556
rect 12360 5370 12388 5528
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12636 4690 12664 9114
rect 12820 6225 12848 19343
rect 12912 19310 12940 19751
rect 12900 19304 12952 19310
rect 12900 19246 12952 19252
rect 13096 18902 13124 20198
rect 13188 20058 13216 20878
rect 13556 20369 13584 23462
rect 13818 23352 13874 23361
rect 13636 23316 13688 23322
rect 13818 23287 13874 23296
rect 13636 23258 13688 23264
rect 13648 22642 13676 23258
rect 13636 22636 13688 22642
rect 13636 22578 13688 22584
rect 13636 22500 13688 22506
rect 13636 22442 13688 22448
rect 13648 21078 13676 22442
rect 13728 22160 13780 22166
rect 13832 22114 13860 23287
rect 13780 22108 13860 22114
rect 13728 22102 13860 22108
rect 13740 22086 13860 22102
rect 13832 21690 13860 22086
rect 13820 21684 13872 21690
rect 13820 21626 13872 21632
rect 13726 21448 13782 21457
rect 13726 21383 13782 21392
rect 13636 21072 13688 21078
rect 13636 21014 13688 21020
rect 13542 20360 13598 20369
rect 13542 20295 13598 20304
rect 13176 20052 13228 20058
rect 13176 19994 13228 20000
rect 13188 19378 13216 19994
rect 13268 19848 13320 19854
rect 13268 19790 13320 19796
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 13280 18970 13308 19790
rect 13556 19417 13584 20295
rect 13542 19408 13598 19417
rect 13542 19343 13598 19352
rect 13268 18964 13320 18970
rect 13268 18906 13320 18912
rect 13084 18896 13136 18902
rect 13084 18838 13136 18844
rect 12990 18456 13046 18465
rect 12990 18391 13046 18400
rect 13004 18222 13032 18391
rect 12992 18216 13044 18222
rect 12990 18184 12992 18193
rect 13044 18184 13046 18193
rect 12990 18119 13046 18128
rect 13004 17882 13032 18119
rect 13096 18086 13124 18838
rect 13452 18760 13504 18766
rect 13452 18702 13504 18708
rect 13464 18290 13492 18702
rect 13452 18284 13504 18290
rect 13452 18226 13504 18232
rect 13084 18080 13136 18086
rect 13084 18022 13136 18028
rect 12992 17876 13044 17882
rect 12992 17818 13044 17824
rect 13096 17814 13124 18022
rect 13464 17882 13492 18226
rect 13452 17876 13504 17882
rect 13452 17818 13504 17824
rect 13084 17808 13136 17814
rect 13084 17750 13136 17756
rect 13096 16998 13124 17750
rect 13452 17672 13504 17678
rect 13452 17614 13504 17620
rect 13266 17368 13322 17377
rect 13266 17303 13322 17312
rect 13084 16992 13136 16998
rect 13084 16934 13136 16940
rect 13084 16720 13136 16726
rect 13084 16662 13136 16668
rect 13096 16046 13124 16662
rect 13084 16040 13136 16046
rect 13084 15982 13136 15988
rect 13096 15706 13124 15982
rect 13084 15700 13136 15706
rect 13084 15642 13136 15648
rect 13176 15360 13228 15366
rect 13176 15302 13228 15308
rect 13188 14958 13216 15302
rect 13176 14952 13228 14958
rect 13176 14894 13228 14900
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 12912 14278 12940 14418
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 12900 14272 12952 14278
rect 12900 14214 12952 14220
rect 12912 13870 12940 14214
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 12912 13462 12940 13806
rect 13004 13530 13032 14350
rect 13188 13938 13216 14894
rect 13280 14793 13308 17303
rect 13464 17202 13492 17614
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13360 17128 13412 17134
rect 13358 17096 13360 17105
rect 13412 17096 13414 17105
rect 13358 17031 13414 17040
rect 13360 16992 13412 16998
rect 13360 16934 13412 16940
rect 13372 15162 13400 16934
rect 13464 16114 13492 17138
rect 13544 17128 13596 17134
rect 13544 17070 13596 17076
rect 13556 16726 13584 17070
rect 13544 16720 13596 16726
rect 13544 16662 13596 16668
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 13648 15910 13676 16526
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 13648 15745 13676 15846
rect 13634 15736 13690 15745
rect 13634 15671 13690 15680
rect 13740 15586 13768 21383
rect 13832 21010 13860 21626
rect 13820 21004 13872 21010
rect 13820 20946 13872 20952
rect 13832 19990 13860 20946
rect 13820 19984 13872 19990
rect 13820 19926 13872 19932
rect 13832 19514 13860 19926
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13924 19281 13952 24278
rect 14200 23730 14228 25094
rect 14280 24744 14332 24750
rect 14280 24686 14332 24692
rect 14740 24744 14792 24750
rect 14740 24686 14792 24692
rect 14292 24342 14320 24686
rect 14280 24336 14332 24342
rect 14280 24278 14332 24284
rect 14648 24268 14700 24274
rect 14648 24210 14700 24216
rect 14188 23724 14240 23730
rect 14188 23666 14240 23672
rect 14280 23724 14332 23730
rect 14280 23666 14332 23672
rect 14096 23520 14148 23526
rect 14096 23462 14148 23468
rect 14004 21888 14056 21894
rect 14004 21830 14056 21836
rect 14016 21554 14044 21830
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 14108 21418 14136 23462
rect 14200 23322 14228 23666
rect 14188 23316 14240 23322
rect 14188 23258 14240 23264
rect 14292 22098 14320 23666
rect 14660 23254 14688 24210
rect 14648 23248 14700 23254
rect 14648 23190 14700 23196
rect 14280 22092 14332 22098
rect 14280 22034 14332 22040
rect 14096 21412 14148 21418
rect 14096 21354 14148 21360
rect 14108 21146 14136 21354
rect 14096 21140 14148 21146
rect 14096 21082 14148 21088
rect 14108 20602 14136 21082
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 13910 19272 13966 19281
rect 13910 19207 13966 19216
rect 14292 18358 14320 22034
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 14384 19718 14412 21490
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14384 19378 14412 19654
rect 14372 19372 14424 19378
rect 14372 19314 14424 19320
rect 14464 19236 14516 19242
rect 14464 19178 14516 19184
rect 14476 18970 14504 19178
rect 14464 18964 14516 18970
rect 14464 18906 14516 18912
rect 14280 18352 14332 18358
rect 14280 18294 14332 18300
rect 14648 18284 14700 18290
rect 14648 18226 14700 18232
rect 14280 18080 14332 18086
rect 14280 18022 14332 18028
rect 14462 18048 14518 18057
rect 14292 17882 14320 18022
rect 14462 17983 14518 17992
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 14476 17338 14504 17983
rect 14660 17882 14688 18226
rect 14648 17876 14700 17882
rect 14648 17818 14700 17824
rect 14464 17332 14516 17338
rect 14464 17274 14516 17280
rect 14370 16688 14426 16697
rect 14370 16623 14372 16632
rect 14424 16623 14426 16632
rect 14372 16594 14424 16600
rect 14384 16114 14412 16594
rect 14372 16108 14424 16114
rect 14372 16050 14424 16056
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 14004 15904 14056 15910
rect 14004 15846 14056 15852
rect 13648 15558 13768 15586
rect 13820 15632 13872 15638
rect 13820 15574 13872 15580
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 13372 14872 13400 15098
rect 13452 14884 13504 14890
rect 13372 14844 13452 14872
rect 13266 14784 13322 14793
rect 13266 14719 13322 14728
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 12900 13456 12952 13462
rect 12900 13398 12952 13404
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 13188 11626 13216 12242
rect 13176 11620 13228 11626
rect 13176 11562 13228 11568
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12912 10849 12940 11494
rect 13188 11354 13216 11562
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 12898 10840 12954 10849
rect 12898 10775 12954 10784
rect 13188 10674 13216 11290
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 13004 9926 13032 10542
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 12900 9648 12952 9654
rect 12900 9590 12952 9596
rect 12912 9450 12940 9590
rect 12900 9444 12952 9450
rect 12900 9386 12952 9392
rect 12912 7410 12940 9386
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 12806 6216 12862 6225
rect 12716 6180 12768 6186
rect 12806 6151 12862 6160
rect 12716 6122 12768 6128
rect 12728 5846 12756 6122
rect 12716 5840 12768 5846
rect 12716 5782 12768 5788
rect 12728 5302 12756 5782
rect 12716 5296 12768 5302
rect 12716 5238 12768 5244
rect 12714 5128 12770 5137
rect 12714 5063 12716 5072
rect 12768 5063 12770 5072
rect 12716 5034 12768 5040
rect 12728 4826 12756 5034
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12624 4684 12676 4690
rect 12624 4626 12676 4632
rect 12440 4616 12492 4622
rect 12440 4558 12492 4564
rect 12348 4548 12400 4554
rect 12348 4490 12400 4496
rect 12360 4214 12388 4490
rect 12348 4208 12400 4214
rect 12348 4150 12400 4156
rect 12162 3632 12218 3641
rect 12162 3567 12218 3576
rect 12070 3224 12126 3233
rect 12070 3159 12126 3168
rect 12176 3126 12204 3567
rect 12452 3466 12480 4558
rect 12636 4146 12664 4626
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12532 4004 12584 4010
rect 12532 3946 12584 3952
rect 12544 3738 12572 3946
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12636 3670 12664 4082
rect 12624 3664 12676 3670
rect 12624 3606 12676 3612
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 12820 3194 12848 3470
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 12164 3120 12216 3126
rect 12164 3062 12216 3068
rect 11980 2984 12032 2990
rect 11980 2926 12032 2932
rect 11796 2372 11848 2378
rect 11796 2314 11848 2320
rect 10796 2230 10916 2258
rect 10796 480 10824 2230
rect 11808 480 11836 2314
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 12912 480 12940 2246
rect 13004 1601 13032 9862
rect 13280 9636 13308 14719
rect 13372 14550 13400 14844
rect 13452 14826 13504 14832
rect 13360 14544 13412 14550
rect 13360 14486 13412 14492
rect 13372 14074 13400 14486
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13648 13394 13676 15558
rect 13728 15496 13780 15502
rect 13726 15464 13728 15473
rect 13780 15464 13782 15473
rect 13726 15399 13782 15408
rect 13832 15094 13860 15574
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 14016 14385 14044 15846
rect 14568 15638 14596 16050
rect 14556 15632 14608 15638
rect 14554 15600 14556 15609
rect 14608 15600 14610 15609
rect 14554 15535 14610 15544
rect 14646 15464 14702 15473
rect 14646 15399 14702 15408
rect 14660 15162 14688 15399
rect 14648 15156 14700 15162
rect 14648 15098 14700 15104
rect 14002 14376 14058 14385
rect 14002 14311 14058 14320
rect 14016 14278 14044 14311
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 14188 14272 14240 14278
rect 14188 14214 14240 14220
rect 14016 14074 14044 14214
rect 14004 14068 14056 14074
rect 14004 14010 14056 14016
rect 14016 13870 14044 14010
rect 14200 13977 14228 14214
rect 14186 13968 14242 13977
rect 14186 13903 14188 13912
rect 14240 13903 14242 13912
rect 14188 13874 14240 13880
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 13636 13388 13688 13394
rect 13636 13330 13688 13336
rect 13648 12986 13676 13330
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13556 12306 13584 12718
rect 13544 12300 13596 12306
rect 13544 12242 13596 12248
rect 13556 12102 13584 12242
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 13556 11898 13584 12038
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13634 11656 13690 11665
rect 13634 11591 13690 11600
rect 13648 11218 13676 11591
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13648 10810 13676 11154
rect 13636 10804 13688 10810
rect 13636 10746 13688 10752
rect 13740 10538 13768 13806
rect 14752 13784 14780 24686
rect 14844 24410 14872 25214
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15948 24857 15976 27520
rect 15934 24848 15990 24857
rect 15934 24783 15990 24792
rect 16670 24848 16726 24857
rect 16670 24783 16672 24792
rect 16724 24783 16726 24792
rect 16672 24754 16724 24760
rect 17052 24682 17080 27520
rect 17500 26376 17552 26382
rect 17500 26318 17552 26324
rect 17040 24676 17092 24682
rect 17040 24618 17092 24624
rect 16304 24608 16356 24614
rect 16304 24550 16356 24556
rect 14832 24404 14884 24410
rect 14832 24346 14884 24352
rect 15476 24336 15528 24342
rect 15476 24278 15528 24284
rect 15292 24132 15344 24138
rect 15292 24074 15344 24080
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15304 23746 15332 24074
rect 15488 23866 15516 24278
rect 16028 24200 16080 24206
rect 16028 24142 16080 24148
rect 15476 23860 15528 23866
rect 15476 23802 15528 23808
rect 15120 23718 15332 23746
rect 15016 23588 15068 23594
rect 15016 23530 15068 23536
rect 15028 23066 15056 23530
rect 15120 23322 15148 23718
rect 15488 23361 15516 23802
rect 16040 23798 16068 24142
rect 16028 23792 16080 23798
rect 16028 23734 16080 23740
rect 15844 23588 15896 23594
rect 15844 23530 15896 23536
rect 15474 23352 15530 23361
rect 15108 23316 15160 23322
rect 15474 23287 15530 23296
rect 15108 23258 15160 23264
rect 15476 23248 15528 23254
rect 15476 23190 15528 23196
rect 14832 23044 14884 23050
rect 15028 23038 15332 23066
rect 14832 22986 14884 22992
rect 14844 19378 14872 22986
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15304 22710 15332 23038
rect 15488 22778 15516 23190
rect 15856 22982 15884 23530
rect 16040 23118 16068 23734
rect 16028 23112 16080 23118
rect 16028 23054 16080 23060
rect 15844 22976 15896 22982
rect 15844 22918 15896 22924
rect 15476 22772 15528 22778
rect 15476 22714 15528 22720
rect 15292 22704 15344 22710
rect 15292 22646 15344 22652
rect 15304 22506 15332 22646
rect 15292 22500 15344 22506
rect 15292 22442 15344 22448
rect 15384 22092 15436 22098
rect 15384 22034 15436 22040
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15396 21350 15424 22034
rect 15752 21480 15804 21486
rect 15750 21448 15752 21457
rect 15804 21448 15806 21457
rect 15750 21383 15806 21392
rect 15384 21344 15436 21350
rect 15384 21286 15436 21292
rect 15396 20913 15424 21286
rect 15382 20904 15438 20913
rect 15382 20839 15438 20848
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 15200 20392 15252 20398
rect 15198 20360 15200 20369
rect 15252 20360 15254 20369
rect 15198 20295 15254 20304
rect 15568 20256 15620 20262
rect 15568 20198 15620 20204
rect 15580 19961 15608 20198
rect 15566 19952 15622 19961
rect 15566 19887 15622 19896
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14844 18290 14872 19314
rect 15856 19174 15884 22918
rect 16040 22710 16068 23054
rect 16316 22778 16344 24550
rect 16580 24268 16632 24274
rect 16580 24210 16632 24216
rect 16394 24168 16450 24177
rect 16394 24103 16396 24112
rect 16448 24103 16450 24112
rect 16396 24074 16448 24080
rect 16408 23730 16436 24074
rect 16396 23724 16448 23730
rect 16396 23666 16448 23672
rect 16592 23526 16620 24210
rect 16580 23520 16632 23526
rect 16580 23462 16632 23468
rect 16304 22772 16356 22778
rect 16304 22714 16356 22720
rect 16028 22704 16080 22710
rect 16028 22646 16080 22652
rect 16212 22160 16264 22166
rect 16212 22102 16264 22108
rect 16120 21004 16172 21010
rect 16120 20946 16172 20952
rect 16028 20800 16080 20806
rect 16028 20742 16080 20748
rect 16040 19854 16068 20742
rect 16132 20262 16160 20946
rect 16224 20466 16252 22102
rect 16488 22092 16540 22098
rect 16488 22034 16540 22040
rect 16500 21894 16528 22034
rect 16488 21888 16540 21894
rect 16488 21830 16540 21836
rect 16500 21486 16528 21830
rect 16488 21480 16540 21486
rect 16488 21422 16540 21428
rect 16212 20460 16264 20466
rect 16212 20402 16264 20408
rect 16120 20256 16172 20262
rect 16120 20198 16172 20204
rect 16028 19848 16080 19854
rect 16028 19790 16080 19796
rect 15934 19272 15990 19281
rect 15934 19207 15936 19216
rect 15988 19207 15990 19216
rect 15936 19178 15988 19184
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15856 18970 15884 19110
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 16028 18964 16080 18970
rect 16028 18906 16080 18912
rect 15384 18828 15436 18834
rect 15384 18770 15436 18776
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 15396 18193 15424 18770
rect 15382 18184 15438 18193
rect 16040 18154 16068 18906
rect 15382 18119 15438 18128
rect 15936 18148 15988 18154
rect 15396 18086 15424 18119
rect 15936 18090 15988 18096
rect 16028 18148 16080 18154
rect 16028 18090 16080 18096
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 15292 17740 15344 17746
rect 15292 17682 15344 17688
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15304 17241 15332 17682
rect 15290 17232 15346 17241
rect 15290 17167 15292 17176
rect 15344 17167 15346 17176
rect 15292 17138 15344 17144
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 15304 15162 15332 15846
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 14568 13756 14780 13784
rect 14186 13016 14242 13025
rect 14186 12951 14242 12960
rect 14464 12980 14516 12986
rect 14200 12782 14228 12951
rect 14464 12922 14516 12928
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14004 12708 14056 12714
rect 14004 12650 14056 12656
rect 14016 12617 14044 12650
rect 14188 12640 14240 12646
rect 14002 12608 14058 12617
rect 14188 12582 14240 12588
rect 14370 12608 14426 12617
rect 14002 12543 14058 12552
rect 14094 11384 14150 11393
rect 14094 11319 14150 11328
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13728 10532 13780 10538
rect 13728 10474 13780 10480
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13556 9722 13584 9998
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 13096 9608 13308 9636
rect 13096 5352 13124 9608
rect 13648 8974 13676 10066
rect 13740 9042 13768 10474
rect 13832 10266 13860 11086
rect 14016 10674 14044 11154
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13648 8430 13676 8910
rect 13740 8634 13768 8978
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 14016 8537 14044 8910
rect 14002 8528 14058 8537
rect 14002 8463 14058 8472
rect 14108 8430 14136 11319
rect 14200 10810 14228 12582
rect 14370 12543 14426 12552
rect 14384 12442 14412 12543
rect 14372 12436 14424 12442
rect 14372 12378 14424 12384
rect 14278 12336 14334 12345
rect 14278 12271 14334 12280
rect 14292 12073 14320 12271
rect 14278 12064 14334 12073
rect 14278 11999 14334 12008
rect 14476 11778 14504 12922
rect 14292 11750 14504 11778
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14292 10305 14320 11750
rect 14568 11676 14596 13756
rect 14844 12850 14872 14758
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 15120 13530 15148 13806
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15212 13394 15240 13466
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 15396 12782 15424 18022
rect 15948 17882 15976 18090
rect 16040 18057 16068 18090
rect 16026 18048 16082 18057
rect 16026 17983 16082 17992
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 15566 17096 15622 17105
rect 15566 17031 15622 17040
rect 15476 15088 15528 15094
rect 15476 15030 15528 15036
rect 15488 14550 15516 15030
rect 15476 14544 15528 14550
rect 15476 14486 15528 14492
rect 15488 14006 15516 14486
rect 15476 14000 15528 14006
rect 15476 13942 15528 13948
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15212 12374 15240 12718
rect 15580 12442 15608 17031
rect 15660 16652 15712 16658
rect 15660 16594 15712 16600
rect 15672 16182 15700 16594
rect 15660 16176 15712 16182
rect 15660 16118 15712 16124
rect 15672 15910 15700 16118
rect 15752 16040 15804 16046
rect 15752 15982 15804 15988
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15672 13190 15700 15846
rect 15764 15745 15792 15982
rect 15750 15736 15806 15745
rect 15750 15671 15752 15680
rect 15804 15671 15806 15680
rect 16028 15700 16080 15706
rect 15752 15642 15804 15648
rect 16028 15642 16080 15648
rect 15764 15611 15792 15642
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 16040 14362 16068 15642
rect 16132 14498 16160 20198
rect 16224 20058 16252 20402
rect 16500 20346 16528 21422
rect 16592 20942 16620 23462
rect 17132 23180 17184 23186
rect 17132 23122 17184 23128
rect 17144 22778 17172 23122
rect 17132 22772 17184 22778
rect 17132 22714 17184 22720
rect 17512 22166 17540 26318
rect 18064 24426 18092 27520
rect 17880 24410 18092 24426
rect 17868 24404 18092 24410
rect 17920 24398 18092 24404
rect 17868 24346 17920 24352
rect 18326 24304 18382 24313
rect 18326 24239 18328 24248
rect 18380 24239 18382 24248
rect 18328 24210 18380 24216
rect 18340 23798 18368 24210
rect 19076 23866 19104 27520
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 20088 24313 20116 27520
rect 20074 24304 20130 24313
rect 20074 24239 20130 24248
rect 19064 23860 19116 23866
rect 19064 23802 19116 23808
rect 18328 23792 18380 23798
rect 18328 23734 18380 23740
rect 19432 23520 19484 23526
rect 19432 23462 19484 23468
rect 19984 23520 20036 23526
rect 19984 23462 20036 23468
rect 18512 23248 18564 23254
rect 18512 23190 18564 23196
rect 17868 23112 17920 23118
rect 17868 23054 17920 23060
rect 17880 22778 17908 23054
rect 17868 22772 17920 22778
rect 17868 22714 17920 22720
rect 18524 22438 18552 23190
rect 19248 23044 19300 23050
rect 19248 22986 19300 22992
rect 19260 22642 19288 22986
rect 19248 22636 19300 22642
rect 19248 22578 19300 22584
rect 18880 22500 18932 22506
rect 18880 22442 18932 22448
rect 18052 22432 18104 22438
rect 18052 22374 18104 22380
rect 18512 22432 18564 22438
rect 18512 22374 18564 22380
rect 17500 22160 17552 22166
rect 17500 22102 17552 22108
rect 17132 22024 17184 22030
rect 17132 21966 17184 21972
rect 17144 21554 17172 21966
rect 17132 21548 17184 21554
rect 17132 21490 17184 21496
rect 17512 21350 17540 22102
rect 17960 21548 18012 21554
rect 17960 21490 18012 21496
rect 16672 21344 16724 21350
rect 16672 21286 16724 21292
rect 17500 21344 17552 21350
rect 17500 21286 17552 21292
rect 16684 21078 16712 21286
rect 17224 21140 17276 21146
rect 17224 21082 17276 21088
rect 16672 21072 16724 21078
rect 16672 21014 16724 21020
rect 16580 20936 16632 20942
rect 16580 20878 16632 20884
rect 16684 20806 16712 21014
rect 16672 20800 16724 20806
rect 16672 20742 16724 20748
rect 16580 20460 16632 20466
rect 16580 20402 16632 20408
rect 16592 20346 16620 20402
rect 16500 20318 16620 20346
rect 16684 20330 16712 20742
rect 16672 20324 16724 20330
rect 16212 20052 16264 20058
rect 16212 19994 16264 20000
rect 16304 19984 16356 19990
rect 16304 19926 16356 19932
rect 16212 19712 16264 19718
rect 16212 19654 16264 19660
rect 16224 19378 16252 19654
rect 16316 19514 16344 19926
rect 16304 19508 16356 19514
rect 16304 19450 16356 19456
rect 16212 19372 16264 19378
rect 16212 19314 16264 19320
rect 16500 18834 16528 20318
rect 16672 20266 16724 20272
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 16580 19848 16632 19854
rect 16580 19790 16632 19796
rect 16592 18970 16620 19790
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 17052 18902 17080 20198
rect 17236 20058 17264 21082
rect 17776 20936 17828 20942
rect 17776 20878 17828 20884
rect 17788 20466 17816 20878
rect 17776 20460 17828 20466
rect 17776 20402 17828 20408
rect 17868 20392 17920 20398
rect 17868 20334 17920 20340
rect 17880 20210 17908 20334
rect 17972 20210 18000 21490
rect 18064 21078 18092 22374
rect 18892 22250 18920 22442
rect 18800 22222 18920 22250
rect 18800 22166 18828 22222
rect 18788 22160 18840 22166
rect 18788 22102 18840 22108
rect 19064 22160 19116 22166
rect 19064 22102 19116 22108
rect 18800 21706 18828 22102
rect 18972 22024 19024 22030
rect 18972 21966 19024 21972
rect 18708 21678 18828 21706
rect 18602 21312 18658 21321
rect 18602 21247 18658 21256
rect 18052 21072 18104 21078
rect 18052 21014 18104 21020
rect 18064 20262 18092 21014
rect 18512 21004 18564 21010
rect 18512 20946 18564 20952
rect 18524 20602 18552 20946
rect 18512 20596 18564 20602
rect 18512 20538 18564 20544
rect 18144 20324 18196 20330
rect 18144 20266 18196 20272
rect 17880 20182 18000 20210
rect 18052 20256 18104 20262
rect 18052 20198 18104 20204
rect 17774 20088 17830 20097
rect 17224 20052 17276 20058
rect 17774 20023 17830 20032
rect 17224 19994 17276 20000
rect 17788 19990 17816 20023
rect 17880 19990 17908 20182
rect 18064 20058 18092 20198
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 17776 19984 17828 19990
rect 17776 19926 17828 19932
rect 17868 19984 17920 19990
rect 17868 19926 17920 19932
rect 17880 19514 17908 19926
rect 18156 19718 18184 20266
rect 18524 19825 18552 20538
rect 18510 19816 18566 19825
rect 18236 19780 18288 19786
rect 18510 19751 18566 19760
rect 18236 19722 18288 19728
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 17868 19508 17920 19514
rect 17868 19450 17920 19456
rect 16856 18896 16908 18902
rect 16856 18838 16908 18844
rect 17040 18896 17092 18902
rect 17040 18838 17092 18844
rect 16212 18828 16264 18834
rect 16212 18770 16264 18776
rect 16488 18828 16540 18834
rect 16488 18770 16540 18776
rect 16224 17610 16252 18770
rect 16868 18086 16896 18838
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 17328 18426 17356 18702
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 18248 18290 18276 19722
rect 18328 19236 18380 19242
rect 18328 19178 18380 19184
rect 18420 19236 18472 19242
rect 18420 19178 18472 19184
rect 18236 18284 18288 18290
rect 18236 18226 18288 18232
rect 16856 18080 16908 18086
rect 16856 18022 16908 18028
rect 17776 18080 17828 18086
rect 17776 18022 17828 18028
rect 16868 17814 16896 18022
rect 17788 17882 17816 18022
rect 18248 17882 18276 18226
rect 18340 17882 18368 19178
rect 18432 18902 18460 19178
rect 18420 18896 18472 18902
rect 18420 18838 18472 18844
rect 17776 17876 17828 17882
rect 17776 17818 17828 17824
rect 18236 17876 18288 17882
rect 18236 17818 18288 17824
rect 18328 17876 18380 17882
rect 18328 17818 18380 17824
rect 16856 17808 16908 17814
rect 16856 17750 16908 17756
rect 16764 17672 16816 17678
rect 16764 17614 16816 17620
rect 16212 17604 16264 17610
rect 16212 17546 16264 17552
rect 16224 16658 16252 17546
rect 16304 17536 16356 17542
rect 16304 17478 16356 17484
rect 16316 17134 16344 17478
rect 16304 17128 16356 17134
rect 16304 17070 16356 17076
rect 16212 16652 16264 16658
rect 16212 16594 16264 16600
rect 16224 16046 16252 16594
rect 16316 16114 16344 17070
rect 16776 16726 16804 17614
rect 16868 16998 16896 17750
rect 18050 17232 18106 17241
rect 18248 17202 18276 17818
rect 18050 17167 18106 17176
rect 18236 17196 18288 17202
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16764 16720 16816 16726
rect 16764 16662 16816 16668
rect 16304 16108 16356 16114
rect 16304 16050 16356 16056
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 16868 15638 16896 16934
rect 17960 16720 18012 16726
rect 17958 16688 17960 16697
rect 18012 16688 18014 16697
rect 17316 16652 17368 16658
rect 17958 16623 18014 16632
rect 17316 16594 17368 16600
rect 17328 16153 17356 16594
rect 17314 16144 17370 16153
rect 17314 16079 17316 16088
rect 17368 16079 17370 16088
rect 17316 16050 17368 16056
rect 16856 15632 16908 15638
rect 16856 15574 16908 15580
rect 16488 15496 16540 15502
rect 16488 15438 16540 15444
rect 16212 14952 16264 14958
rect 16212 14894 16264 14900
rect 16224 14618 16252 14894
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 16132 14470 16252 14498
rect 15764 13938 15792 14350
rect 16040 14334 16160 14362
rect 15752 13932 15804 13938
rect 15752 13874 15804 13880
rect 15764 13705 15792 13874
rect 15750 13696 15806 13705
rect 15750 13631 15806 13640
rect 15660 13184 15712 13190
rect 15660 13126 15712 13132
rect 15568 12436 15620 12442
rect 15568 12378 15620 12384
rect 15200 12368 15252 12374
rect 15200 12310 15252 12316
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15290 12200 15346 12209
rect 15290 12135 15346 12144
rect 15304 12102 15332 12135
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14370 11656 14426 11665
rect 14370 11591 14426 11600
rect 14476 11648 14596 11676
rect 14924 11688 14976 11694
rect 14384 11286 14412 11591
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 14278 10296 14334 10305
rect 14278 10231 14334 10240
rect 14476 9908 14504 11648
rect 14924 11630 14976 11636
rect 14740 11620 14792 11626
rect 14740 11562 14792 11568
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 14556 11008 14608 11014
rect 14556 10950 14608 10956
rect 14568 10606 14596 10950
rect 14660 10810 14688 11154
rect 14752 11150 14780 11562
rect 14832 11280 14884 11286
rect 14832 11222 14884 11228
rect 14740 11144 14792 11150
rect 14738 11112 14740 11121
rect 14792 11112 14794 11121
rect 14738 11047 14794 11056
rect 14752 11021 14780 11047
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14740 10532 14792 10538
rect 14740 10474 14792 10480
rect 14646 10296 14702 10305
rect 14646 10231 14702 10240
rect 14292 9880 14504 9908
rect 14292 9704 14320 9880
rect 14292 9676 14504 9704
rect 14186 9072 14242 9081
rect 14186 9007 14242 9016
rect 14280 9036 14332 9042
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 13176 8356 13228 8362
rect 13176 8298 13228 8304
rect 13188 7886 13216 8298
rect 13648 8090 13676 8366
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 14200 7970 14228 9007
rect 14280 8978 14332 8984
rect 14292 8537 14320 8978
rect 14278 8528 14334 8537
rect 14278 8463 14334 8472
rect 14108 7954 14228 7970
rect 14108 7948 14240 7954
rect 14108 7942 14188 7948
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13188 7546 13216 7822
rect 14108 7546 14136 7942
rect 14188 7890 14240 7896
rect 14188 7812 14240 7818
rect 14188 7754 14240 7760
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 14108 7002 14136 7346
rect 14200 7274 14228 7754
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14188 7268 14240 7274
rect 14188 7210 14240 7216
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 14384 6934 14412 7346
rect 13360 6928 13412 6934
rect 13360 6870 13412 6876
rect 14372 6928 14424 6934
rect 14372 6870 14424 6876
rect 13372 6458 13400 6870
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 14016 6458 14044 6734
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 14004 6452 14056 6458
rect 14004 6394 14056 6400
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13096 5324 13216 5352
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 13096 4622 13124 5170
rect 13084 4616 13136 4622
rect 13084 4558 13136 4564
rect 13096 4214 13124 4558
rect 13084 4208 13136 4214
rect 13084 4150 13136 4156
rect 13188 3754 13216 5324
rect 13832 5098 13860 5510
rect 13820 5092 13872 5098
rect 13820 5034 13872 5040
rect 13636 5024 13688 5030
rect 13634 4992 13636 5001
rect 13688 4992 13690 5001
rect 13634 4927 13690 4936
rect 13832 4826 13860 5034
rect 13924 5030 13952 5714
rect 14384 5234 14412 6870
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 13912 5024 13964 5030
rect 13912 4966 13964 4972
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13820 4548 13872 4554
rect 13820 4490 13872 4496
rect 13832 4282 13860 4490
rect 13820 4276 13872 4282
rect 13820 4218 13872 4224
rect 13924 4185 13952 4966
rect 14384 4690 14412 5170
rect 14372 4684 14424 4690
rect 14372 4626 14424 4632
rect 14476 4486 14504 9676
rect 14660 6866 14688 10231
rect 14752 9926 14780 10474
rect 14844 10198 14872 11222
rect 14936 11082 14964 11630
rect 15488 11558 15516 12242
rect 15672 12102 15700 13126
rect 16132 12986 16160 14334
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 15752 12776 15804 12782
rect 15752 12718 15804 12724
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15672 11694 15700 12038
rect 15764 11937 15792 12718
rect 15750 11928 15806 11937
rect 15750 11863 15806 11872
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15474 11248 15530 11257
rect 15384 11212 15436 11218
rect 15304 11172 15384 11200
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15304 10690 15332 11172
rect 15474 11183 15530 11192
rect 15384 11154 15436 11160
rect 15488 11098 15516 11183
rect 15396 11070 15516 11098
rect 15396 10742 15424 11070
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15120 10662 15332 10690
rect 15384 10736 15436 10742
rect 15384 10678 15436 10684
rect 15016 10600 15068 10606
rect 15016 10542 15068 10548
rect 15028 10441 15056 10542
rect 15014 10432 15070 10441
rect 15014 10367 15070 10376
rect 15120 10266 15148 10662
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 14832 10192 14884 10198
rect 14832 10134 14884 10140
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14752 8838 14780 9862
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15304 9704 15332 10066
rect 15212 9676 15332 9704
rect 15212 9518 15240 9676
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 15200 9512 15252 9518
rect 15200 9454 15252 9460
rect 15304 9042 15332 9522
rect 15396 9178 15424 10678
rect 15384 9172 15436 9178
rect 15384 9114 15436 9120
rect 15292 9036 15344 9042
rect 15292 8978 15344 8984
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14752 8430 14780 8774
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15304 8634 15332 8978
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 14740 8424 14792 8430
rect 14740 8366 14792 8372
rect 14752 7750 14780 8366
rect 14832 8356 14884 8362
rect 14832 8298 14884 8304
rect 14844 7993 14872 8298
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 14830 7984 14886 7993
rect 14830 7919 14886 7928
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14752 7177 14780 7686
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 15304 7342 15332 8230
rect 15488 8090 15516 10746
rect 15672 10588 15700 11630
rect 15764 11393 15792 11863
rect 15856 11694 15884 12718
rect 15844 11688 15896 11694
rect 15844 11630 15896 11636
rect 15750 11384 15806 11393
rect 15750 11319 15806 11328
rect 15936 11076 15988 11082
rect 15936 11018 15988 11024
rect 15948 10742 15976 11018
rect 15936 10736 15988 10742
rect 15936 10678 15988 10684
rect 15672 10560 15976 10588
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15580 8498 15608 10474
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15672 9450 15700 10066
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15660 9444 15712 9450
rect 15660 9386 15712 9392
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15568 8492 15620 8498
rect 15568 8434 15620 8440
rect 15580 8090 15608 8434
rect 15476 8084 15528 8090
rect 15476 8026 15528 8032
rect 15568 8084 15620 8090
rect 15568 8026 15620 8032
rect 15764 7954 15792 9318
rect 15856 9178 15884 9998
rect 15844 9172 15896 9178
rect 15844 9114 15896 9120
rect 15948 8265 15976 10560
rect 16026 10160 16082 10169
rect 16026 10095 16028 10104
rect 16080 10095 16082 10104
rect 16028 10066 16080 10072
rect 16132 9518 16160 12922
rect 16224 12345 16252 14470
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16316 13841 16344 14350
rect 16500 14226 16528 15438
rect 16868 14890 16896 15574
rect 17328 15337 17356 16050
rect 18064 16046 18092 17167
rect 18236 17138 18288 17144
rect 18432 17066 18460 18838
rect 18144 17060 18196 17066
rect 18144 17002 18196 17008
rect 18420 17060 18472 17066
rect 18420 17002 18472 17008
rect 18156 16794 18184 17002
rect 18326 16824 18382 16833
rect 18144 16788 18196 16794
rect 18326 16759 18382 16768
rect 18144 16730 18196 16736
rect 18340 16658 18368 16759
rect 18328 16652 18380 16658
rect 18328 16594 18380 16600
rect 18340 16250 18368 16594
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 18616 16046 18644 21247
rect 18708 19242 18736 21678
rect 18984 21554 19012 21966
rect 19076 21690 19104 22102
rect 19260 22030 19288 22578
rect 19340 22432 19392 22438
rect 19340 22374 19392 22380
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 19064 21684 19116 21690
rect 19064 21626 19116 21632
rect 18788 21548 18840 21554
rect 18788 21490 18840 21496
rect 18972 21548 19024 21554
rect 18972 21490 19024 21496
rect 18800 21418 18828 21490
rect 18788 21412 18840 21418
rect 18788 21354 18840 21360
rect 19352 21350 19380 22374
rect 19444 22030 19472 23462
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19996 23225 20024 23462
rect 19982 23216 20038 23225
rect 21192 23186 21220 27520
rect 22204 23866 22232 27520
rect 23216 24857 23244 27520
rect 23202 24848 23258 24857
rect 23202 24783 23258 24792
rect 23478 24168 23534 24177
rect 23478 24103 23534 24112
rect 23492 23866 23520 24103
rect 22192 23860 22244 23866
rect 22192 23802 22244 23808
rect 23480 23860 23532 23866
rect 23480 23802 23532 23808
rect 19982 23151 20038 23160
rect 21180 23180 21232 23186
rect 21180 23122 21232 23128
rect 20166 23080 20222 23089
rect 20166 23015 20222 23024
rect 19798 22808 19854 22817
rect 20180 22778 20208 23015
rect 21192 22778 21220 23122
rect 24228 23089 24256 27520
rect 24766 26480 24822 26489
rect 24766 26415 24822 26424
rect 24780 26382 24808 26415
rect 24768 26376 24820 26382
rect 24768 26318 24820 26324
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24674 24440 24730 24449
rect 24674 24375 24730 24384
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24688 23186 24716 24375
rect 25332 23769 25360 27520
rect 26344 23882 26372 27520
rect 27356 24449 27384 27520
rect 27342 24440 27398 24449
rect 27342 24375 27398 24384
rect 26160 23866 26372 23882
rect 26148 23860 26372 23866
rect 26200 23854 26372 23860
rect 26148 23802 26200 23808
rect 25318 23760 25374 23769
rect 25318 23695 25374 23704
rect 24676 23180 24728 23186
rect 24676 23122 24728 23128
rect 24214 23080 24270 23089
rect 24214 23015 24270 23024
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23492 22817 23520 22918
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 23478 22808 23534 22817
rect 19798 22743 19800 22752
rect 19852 22743 19854 22752
rect 20168 22772 20220 22778
rect 19800 22714 19852 22720
rect 20168 22714 20220 22720
rect 21180 22772 21232 22778
rect 24289 22800 24585 22820
rect 24688 22778 24716 23122
rect 23478 22743 23534 22752
rect 24676 22772 24728 22778
rect 21180 22714 21232 22720
rect 24676 22714 24728 22720
rect 20180 22574 20208 22714
rect 20168 22568 20220 22574
rect 20168 22510 20220 22516
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19352 21146 19380 21286
rect 19340 21140 19392 21146
rect 19340 21082 19392 21088
rect 18972 20324 19024 20330
rect 18972 20266 19024 20272
rect 18984 19854 19012 20266
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 19352 20097 19380 20198
rect 19338 20088 19394 20097
rect 19156 20052 19208 20058
rect 19338 20023 19394 20032
rect 19156 19994 19208 20000
rect 18972 19848 19024 19854
rect 18972 19790 19024 19796
rect 18984 19242 19012 19790
rect 19168 19514 19196 19994
rect 19340 19984 19392 19990
rect 19338 19952 19340 19961
rect 19392 19952 19394 19961
rect 19338 19887 19394 19896
rect 19248 19712 19300 19718
rect 19300 19660 19380 19666
rect 19248 19654 19380 19660
rect 19260 19638 19380 19654
rect 19156 19508 19208 19514
rect 19156 19450 19208 19456
rect 19352 19242 19380 19638
rect 18696 19236 18748 19242
rect 18696 19178 18748 19184
rect 18972 19236 19024 19242
rect 18972 19178 19024 19184
rect 19340 19236 19392 19242
rect 19340 19178 19392 19184
rect 18984 18766 19012 19178
rect 19444 19122 19472 21966
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 19614 20496 19670 20505
rect 19614 20431 19670 20440
rect 19628 20398 19656 20431
rect 19616 20392 19668 20398
rect 19616 20334 19668 20340
rect 20168 20392 20220 20398
rect 20168 20334 20220 20340
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19614 19952 19670 19961
rect 19614 19887 19670 19896
rect 19628 19514 19656 19887
rect 19616 19508 19668 19514
rect 19616 19450 19668 19456
rect 19352 19094 19472 19122
rect 19064 18896 19116 18902
rect 19064 18838 19116 18844
rect 18972 18760 19024 18766
rect 18972 18702 19024 18708
rect 19076 18426 19104 18838
rect 19352 18698 19380 19094
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 19340 18692 19392 18698
rect 19340 18634 19392 18640
rect 19064 18420 19116 18426
rect 19064 18362 19116 18368
rect 19352 18290 19380 18634
rect 19444 18426 19472 18702
rect 19432 18420 19484 18426
rect 19432 18362 19484 18368
rect 19614 18320 19670 18329
rect 19340 18284 19392 18290
rect 19614 18255 19670 18264
rect 19340 18226 19392 18232
rect 19628 18222 19656 18255
rect 19616 18216 19668 18222
rect 19616 18158 19668 18164
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 18052 16040 18104 16046
rect 18052 15982 18104 15988
rect 18604 16040 18656 16046
rect 18604 15982 18656 15988
rect 18144 15904 18196 15910
rect 18144 15846 18196 15852
rect 18972 15904 19024 15910
rect 18972 15846 19024 15852
rect 17500 15632 17552 15638
rect 17500 15574 17552 15580
rect 18050 15600 18106 15609
rect 17314 15328 17370 15337
rect 17314 15263 17370 15272
rect 17512 15162 17540 15574
rect 18050 15535 18106 15544
rect 18064 15502 18092 15535
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 17500 15156 17552 15162
rect 17500 15098 17552 15104
rect 16856 14884 16908 14890
rect 16856 14826 16908 14832
rect 16580 14272 16632 14278
rect 16500 14220 16580 14226
rect 16500 14214 16632 14220
rect 16500 14198 16620 14214
rect 16302 13832 16358 13841
rect 16302 13767 16304 13776
rect 16356 13767 16358 13776
rect 16304 13738 16356 13744
rect 16302 13560 16358 13569
rect 16302 13495 16304 13504
rect 16356 13495 16358 13504
rect 16304 13466 16356 13472
rect 16316 12782 16344 13466
rect 16500 12918 16528 14198
rect 16764 14000 16816 14006
rect 16764 13942 16816 13948
rect 16580 13932 16632 13938
rect 16580 13874 16632 13880
rect 16592 13802 16620 13874
rect 16580 13796 16632 13802
rect 16580 13738 16632 13744
rect 16592 13530 16620 13738
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16488 12912 16540 12918
rect 16488 12854 16540 12860
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16210 12336 16266 12345
rect 16210 12271 16266 12280
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16316 10674 16344 11494
rect 16500 11286 16528 12718
rect 16592 12646 16620 13262
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16592 12288 16620 12582
rect 16684 12442 16712 13330
rect 16776 12714 16804 13942
rect 16868 13462 16896 14826
rect 17316 14816 17368 14822
rect 17316 14758 17368 14764
rect 17328 14550 17356 14758
rect 17316 14544 17368 14550
rect 17222 14512 17278 14521
rect 17316 14486 17368 14492
rect 17222 14447 17278 14456
rect 17236 14414 17264 14447
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 17236 14006 17264 14350
rect 17328 14074 17356 14486
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 17224 14000 17276 14006
rect 17224 13942 17276 13948
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 16856 13456 16908 13462
rect 16856 13398 16908 13404
rect 16856 13252 16908 13258
rect 16856 13194 16908 13200
rect 16764 12708 16816 12714
rect 16764 12650 16816 12656
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 16672 12300 16724 12306
rect 16592 12260 16672 12288
rect 16672 12242 16724 12248
rect 16684 11558 16712 12242
rect 16764 12232 16816 12238
rect 16762 12200 16764 12209
rect 16816 12200 16818 12209
rect 16762 12135 16818 12144
rect 16776 11762 16804 12135
rect 16764 11756 16816 11762
rect 16764 11698 16816 11704
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16488 11280 16540 11286
rect 16488 11222 16540 11228
rect 16488 11008 16540 11014
rect 16488 10950 16540 10956
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 16500 10606 16528 10950
rect 16396 10600 16448 10606
rect 16396 10542 16448 10548
rect 16488 10600 16540 10606
rect 16488 10542 16540 10548
rect 16408 9994 16436 10542
rect 16396 9988 16448 9994
rect 16396 9930 16448 9936
rect 16408 9722 16436 9930
rect 16396 9716 16448 9722
rect 16396 9658 16448 9664
rect 16500 9518 16528 10542
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16120 9512 16172 9518
rect 16120 9454 16172 9460
rect 16304 9512 16356 9518
rect 16304 9454 16356 9460
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 16132 9217 16160 9454
rect 16212 9376 16264 9382
rect 16212 9318 16264 9324
rect 16118 9208 16174 9217
rect 16118 9143 16120 9152
rect 16172 9143 16174 9152
rect 16120 9114 16172 9120
rect 15934 8256 15990 8265
rect 15934 8191 15990 8200
rect 15476 7948 15528 7954
rect 15476 7890 15528 7896
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 14738 7168 14794 7177
rect 14738 7103 14794 7112
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14556 6384 14608 6390
rect 14556 6326 14608 6332
rect 14464 4480 14516 4486
rect 14464 4422 14516 4428
rect 13910 4176 13966 4185
rect 13910 4111 13966 4120
rect 13096 3726 13216 3754
rect 13096 2650 13124 3726
rect 13176 3664 13228 3670
rect 13176 3606 13228 3612
rect 13188 3058 13216 3606
rect 14568 3194 14596 6326
rect 14660 4282 14688 6802
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 14752 3738 14780 7103
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15304 6440 15332 7278
rect 15488 7206 15516 7890
rect 16224 7410 16252 9318
rect 16316 8838 16344 9454
rect 16488 9036 16540 9042
rect 16592 9024 16620 10406
rect 16684 9110 16712 11494
rect 16868 11354 16896 13194
rect 17144 12170 17172 13874
rect 17604 12986 17632 14350
rect 17972 13954 18000 15370
rect 18064 15162 18092 15438
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 18064 14482 18092 15098
rect 18156 15026 18184 15846
rect 18984 15473 19012 15846
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 18970 15464 19026 15473
rect 18970 15399 19026 15408
rect 18144 15020 18196 15026
rect 18144 14962 18196 14968
rect 18156 14618 18184 14962
rect 18788 14884 18840 14890
rect 18788 14826 18840 14832
rect 18144 14612 18196 14618
rect 18144 14554 18196 14560
rect 18052 14476 18104 14482
rect 18052 14418 18104 14424
rect 18050 14376 18106 14385
rect 18050 14311 18106 14320
rect 17696 13938 18000 13954
rect 17684 13932 18000 13938
rect 17736 13926 18000 13932
rect 17684 13874 17736 13880
rect 18064 13462 18092 14311
rect 18328 14272 18380 14278
rect 18328 14214 18380 14220
rect 18340 13938 18368 14214
rect 18328 13932 18380 13938
rect 18328 13874 18380 13880
rect 18420 13932 18472 13938
rect 18420 13874 18472 13880
rect 18144 13796 18196 13802
rect 18144 13738 18196 13744
rect 18156 13530 18184 13738
rect 18144 13524 18196 13530
rect 18144 13466 18196 13472
rect 18052 13456 18104 13462
rect 18052 13398 18104 13404
rect 17776 13184 17828 13190
rect 17776 13126 17828 13132
rect 17592 12980 17644 12986
rect 17592 12922 17644 12928
rect 17788 12850 17816 13126
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17132 12164 17184 12170
rect 17132 12106 17184 12112
rect 17144 11370 17172 12106
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 18248 11694 18276 12038
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 18236 11688 18288 11694
rect 18236 11630 18288 11636
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 17052 11342 17172 11370
rect 16856 11212 16908 11218
rect 16856 11154 16908 11160
rect 16868 10810 16896 11154
rect 16946 11112 17002 11121
rect 16946 11047 16948 11056
rect 17000 11047 17002 11056
rect 16948 11018 17000 11024
rect 16856 10804 16908 10810
rect 16856 10746 16908 10752
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16762 10024 16818 10033
rect 16762 9959 16764 9968
rect 16816 9959 16818 9968
rect 16764 9930 16816 9936
rect 16868 9722 16896 10066
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16672 9104 16724 9110
rect 16672 9046 16724 9052
rect 16540 8996 16620 9024
rect 16488 8978 16540 8984
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 16394 8528 16450 8537
rect 16394 8463 16450 8472
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 15384 6996 15436 7002
rect 15384 6938 15436 6944
rect 15212 6412 15332 6440
rect 14832 6384 14884 6390
rect 14830 6352 14832 6361
rect 14884 6352 14886 6361
rect 14830 6287 14886 6296
rect 14832 6248 14884 6254
rect 14832 6190 14884 6196
rect 14844 3942 14872 6190
rect 15212 6118 15240 6412
rect 15292 6180 15344 6186
rect 15292 6122 15344 6128
rect 15200 6112 15252 6118
rect 15200 6054 15252 6060
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15304 5234 15332 6122
rect 15396 5817 15424 6938
rect 15382 5808 15438 5817
rect 15382 5743 15438 5752
rect 15292 5228 15344 5234
rect 15292 5170 15344 5176
rect 15290 4992 15346 5001
rect 15290 4927 15346 4936
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 15120 3738 15148 4014
rect 15304 3738 15332 4927
rect 15488 4185 15516 7142
rect 16408 6866 16436 8463
rect 16500 8090 16528 8978
rect 16684 8362 16712 9046
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16684 8022 16712 8298
rect 16672 8016 16724 8022
rect 16578 7984 16634 7993
rect 16672 7958 16724 7964
rect 16578 7919 16580 7928
rect 16632 7919 16634 7928
rect 16580 7890 16632 7896
rect 16592 7002 16620 7890
rect 16580 6996 16632 7002
rect 16580 6938 16632 6944
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 15580 5914 15608 6802
rect 16408 6458 16436 6802
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 16580 6248 16632 6254
rect 15750 6216 15806 6225
rect 16580 6190 16632 6196
rect 15750 6151 15806 6160
rect 15844 6180 15896 6186
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15764 5778 15792 6151
rect 15844 6122 15896 6128
rect 15856 5846 15884 6122
rect 15844 5840 15896 5846
rect 15844 5782 15896 5788
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15764 5370 15792 5714
rect 15856 5370 15884 5782
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15844 5364 15896 5370
rect 15844 5306 15896 5312
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 16500 4826 16528 5170
rect 16488 4820 16540 4826
rect 16488 4762 16540 4768
rect 16592 4758 16620 6190
rect 16764 5296 16816 5302
rect 16764 5238 16816 5244
rect 16580 4752 16632 4758
rect 16580 4694 16632 4700
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15672 4282 15700 4626
rect 16488 4548 16540 4554
rect 16488 4490 16540 4496
rect 15660 4276 15712 4282
rect 15660 4218 15712 4224
rect 15474 4176 15530 4185
rect 16500 4162 16528 4490
rect 16592 4282 16620 4694
rect 16776 4622 16804 5238
rect 16764 4616 16816 4622
rect 16764 4558 16816 4564
rect 16580 4276 16632 4282
rect 16580 4218 16632 4224
rect 16500 4134 16620 4162
rect 16776 4146 16804 4558
rect 15474 4111 15530 4120
rect 16212 3936 16264 3942
rect 16210 3904 16212 3913
rect 16264 3904 16266 3913
rect 16210 3839 16266 3848
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 15108 3732 15160 3738
rect 15108 3674 15160 3680
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 16026 3632 16082 3641
rect 15660 3596 15712 3602
rect 16592 3602 16620 4134
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16026 3567 16082 3576
rect 16580 3596 16632 3602
rect 15660 3538 15712 3544
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15672 3233 15700 3538
rect 15658 3224 15714 3233
rect 14556 3188 14608 3194
rect 15658 3159 15660 3168
rect 14556 3130 14608 3136
rect 15712 3159 15714 3168
rect 15660 3130 15712 3136
rect 13912 3120 13964 3126
rect 13912 3062 13964 3068
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 13084 2644 13136 2650
rect 13084 2586 13136 2592
rect 12990 1592 13046 1601
rect 12990 1527 13046 1536
rect 13924 480 13952 3062
rect 14568 2990 14596 3130
rect 15936 3120 15988 3126
rect 15936 3062 15988 3068
rect 14556 2984 14608 2990
rect 14278 2952 14334 2961
rect 14556 2926 14608 2932
rect 14278 2887 14334 2896
rect 14292 2514 14320 2887
rect 14924 2848 14976 2854
rect 14462 2816 14518 2825
rect 14924 2790 14976 2796
rect 14462 2751 14518 2760
rect 14476 2650 14504 2751
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 14936 2394 14964 2790
rect 14844 2366 14964 2394
rect 14844 1442 14872 2366
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 14844 1414 14964 1442
rect 14936 480 14964 1414
rect 15948 480 15976 3062
rect 16040 2514 16068 3567
rect 16580 3538 16632 3544
rect 16592 3194 16620 3538
rect 17052 3194 17080 11342
rect 18064 11257 18092 11630
rect 18050 11248 18106 11257
rect 17132 11212 17184 11218
rect 18050 11183 18052 11192
rect 17132 11154 17184 11160
rect 18104 11183 18106 11192
rect 18052 11154 18104 11160
rect 17144 10538 17172 11154
rect 18248 11150 18276 11630
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 17408 10736 17460 10742
rect 17408 10678 17460 10684
rect 18050 10704 18106 10713
rect 17420 10577 17448 10678
rect 18050 10639 18106 10648
rect 18064 10606 18092 10639
rect 18052 10600 18104 10606
rect 17406 10568 17462 10577
rect 17132 10532 17184 10538
rect 18052 10542 18104 10548
rect 17406 10503 17462 10512
rect 17132 10474 17184 10480
rect 17144 10130 17172 10474
rect 17132 10124 17184 10130
rect 17132 10066 17184 10072
rect 17144 9654 17172 10066
rect 17420 10062 17448 10503
rect 18064 10266 18092 10542
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 17408 10056 17460 10062
rect 17408 9998 17460 10004
rect 17420 9654 17448 9998
rect 17132 9648 17184 9654
rect 17132 9590 17184 9596
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 17972 9178 18000 9522
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 17776 9104 17828 9110
rect 18156 9081 18184 10406
rect 18236 9988 18288 9994
rect 18236 9930 18288 9936
rect 18248 9450 18276 9930
rect 18236 9444 18288 9450
rect 18236 9386 18288 9392
rect 17776 9046 17828 9052
rect 18142 9072 18198 9081
rect 17788 8838 17816 9046
rect 18142 9007 18198 9016
rect 18144 8968 18196 8974
rect 18144 8910 18196 8916
rect 17776 8832 17828 8838
rect 17776 8774 17828 8780
rect 17788 8634 17816 8774
rect 18156 8634 18184 8910
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 17500 8288 17552 8294
rect 17500 8230 17552 8236
rect 17512 8090 17540 8230
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17590 7032 17646 7041
rect 17590 6967 17646 6976
rect 17604 6798 17632 6967
rect 17696 6934 17724 7482
rect 17684 6928 17736 6934
rect 17684 6870 17736 6876
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17604 5846 17632 6734
rect 17696 6390 17724 6870
rect 17788 6458 17816 8570
rect 18248 8566 18276 9386
rect 18236 8560 18288 8566
rect 18236 8502 18288 8508
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17880 7546 17908 7958
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17868 7540 17920 7546
rect 17868 7482 17920 7488
rect 17972 7206 18000 7686
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18144 7268 18196 7274
rect 18144 7210 18196 7216
rect 17960 7200 18012 7206
rect 17880 7160 17960 7188
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17684 6384 17736 6390
rect 17684 6326 17736 6332
rect 17788 6118 17816 6394
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 17788 5846 17816 6054
rect 17880 5914 17908 7160
rect 17960 7142 18012 7148
rect 18156 6730 18184 7210
rect 18144 6724 18196 6730
rect 18144 6666 18196 6672
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 17960 6384 18012 6390
rect 17960 6326 18012 6332
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17592 5840 17644 5846
rect 17592 5782 17644 5788
rect 17776 5840 17828 5846
rect 17776 5782 17828 5788
rect 17684 5636 17736 5642
rect 17684 5578 17736 5584
rect 17406 4856 17462 4865
rect 17696 4826 17724 5578
rect 17788 5370 17816 5782
rect 17776 5364 17828 5370
rect 17776 5306 17828 5312
rect 17972 5098 18000 6326
rect 18064 6168 18092 6598
rect 18144 6180 18196 6186
rect 18064 6140 18144 6168
rect 18144 6122 18196 6128
rect 18156 5817 18184 6122
rect 18142 5808 18198 5817
rect 18142 5743 18198 5752
rect 17960 5092 18012 5098
rect 17960 5034 18012 5040
rect 17972 4826 18000 5034
rect 17406 4791 17462 4800
rect 17684 4820 17736 4826
rect 17420 4758 17448 4791
rect 17684 4762 17736 4768
rect 17960 4820 18012 4826
rect 17960 4762 18012 4768
rect 17408 4752 17460 4758
rect 17408 4694 17460 4700
rect 17420 4214 17448 4694
rect 17408 4208 17460 4214
rect 17408 4150 17460 4156
rect 17868 3392 17920 3398
rect 17868 3334 17920 3340
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 17052 2990 17080 3130
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 17880 2825 17908 3334
rect 17038 2816 17094 2825
rect 17038 2751 17094 2760
rect 17866 2816 17922 2825
rect 17866 2751 17922 2760
rect 16028 2508 16080 2514
rect 16028 2450 16080 2456
rect 17052 480 17080 2751
rect 18248 2553 18276 7482
rect 18340 2650 18368 13874
rect 18432 13841 18460 13874
rect 18418 13832 18474 13841
rect 18418 13767 18474 13776
rect 18800 13326 18828 14826
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19430 14784 19486 14793
rect 19352 14521 19380 14758
rect 19430 14719 19486 14728
rect 19338 14512 19394 14521
rect 19248 14476 19300 14482
rect 19338 14447 19394 14456
rect 19248 14418 19300 14424
rect 19064 14408 19116 14414
rect 19064 14350 19116 14356
rect 19076 14074 19104 14350
rect 19260 14074 19288 14418
rect 19064 14068 19116 14074
rect 19064 14010 19116 14016
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19260 13569 19288 14010
rect 19338 13968 19394 13977
rect 19338 13903 19340 13912
rect 19392 13903 19394 13912
rect 19340 13874 19392 13880
rect 19444 13870 19472 14719
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19338 13696 19394 13705
rect 19338 13631 19394 13640
rect 19246 13560 19302 13569
rect 19352 13530 19380 13631
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19246 13495 19302 13504
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19064 13456 19116 13462
rect 19064 13398 19116 13404
rect 19798 13424 19854 13433
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 18788 13320 18840 13326
rect 18788 13262 18840 13268
rect 18616 12986 18644 13262
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 18432 10713 18460 11698
rect 18418 10704 18474 10713
rect 18418 10639 18474 10648
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 18432 9722 18460 10066
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 18524 7546 18552 12786
rect 18616 12764 18644 12922
rect 18800 12850 18828 13262
rect 19076 12918 19104 13398
rect 19798 13359 19800 13368
rect 19852 13359 19854 13368
rect 19800 13330 19852 13336
rect 19812 13002 19840 13330
rect 19812 12986 19932 13002
rect 19812 12980 19944 12986
rect 19812 12974 19892 12980
rect 19892 12922 19944 12928
rect 19064 12912 19116 12918
rect 19800 12912 19852 12918
rect 19064 12854 19116 12860
rect 19798 12880 19800 12889
rect 19852 12880 19854 12889
rect 18788 12844 18840 12850
rect 19798 12815 19854 12824
rect 18788 12786 18840 12792
rect 18616 12736 18736 12764
rect 18602 10432 18658 10441
rect 18602 10367 18658 10376
rect 18616 10266 18644 10367
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18604 8356 18656 8362
rect 18604 8298 18656 8304
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 18616 7410 18644 8298
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18616 5794 18644 7346
rect 18432 5766 18644 5794
rect 18432 4865 18460 5766
rect 18604 5704 18656 5710
rect 18604 5646 18656 5652
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 18524 5234 18552 5510
rect 18616 5234 18644 5646
rect 18512 5228 18564 5234
rect 18512 5170 18564 5176
rect 18604 5228 18656 5234
rect 18604 5170 18656 5176
rect 18418 4856 18474 4865
rect 18524 4826 18552 5170
rect 18418 4791 18474 4800
rect 18512 4820 18564 4826
rect 18512 4762 18564 4768
rect 18420 4684 18472 4690
rect 18420 4626 18472 4632
rect 18432 3942 18460 4626
rect 18420 3936 18472 3942
rect 18420 3878 18472 3884
rect 18708 3194 18736 12736
rect 18800 12238 18828 12786
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 19352 12617 19380 12718
rect 19338 12608 19394 12617
rect 19338 12543 19394 12552
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19064 12368 19116 12374
rect 19064 12310 19116 12316
rect 18788 12232 18840 12238
rect 18788 12174 18840 12180
rect 19076 11898 19104 12310
rect 19432 12232 19484 12238
rect 19338 12200 19394 12209
rect 19432 12174 19484 12180
rect 19338 12135 19394 12144
rect 19352 11898 19380 12135
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19248 11620 19300 11626
rect 19248 11562 19300 11568
rect 18972 11212 19024 11218
rect 18972 11154 19024 11160
rect 18984 10470 19012 11154
rect 19260 10656 19288 11562
rect 19444 11354 19472 12174
rect 19798 11928 19854 11937
rect 19798 11863 19800 11872
rect 19852 11863 19854 11872
rect 19800 11834 19852 11840
rect 19616 11688 19668 11694
rect 19614 11656 19616 11665
rect 19668 11656 19670 11665
rect 19614 11591 19670 11600
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19338 11112 19394 11121
rect 19338 11047 19394 11056
rect 19352 10810 19380 11047
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19340 10668 19392 10674
rect 19260 10628 19340 10656
rect 19340 10610 19392 10616
rect 18972 10464 19024 10470
rect 18972 10406 19024 10412
rect 19340 10464 19392 10470
rect 19340 10406 19392 10412
rect 18788 9444 18840 9450
rect 18788 9386 18840 9392
rect 18800 9110 18828 9386
rect 18788 9104 18840 9110
rect 18788 9046 18840 9052
rect 18800 8498 18828 9046
rect 18788 8492 18840 8498
rect 18788 8434 18840 8440
rect 18800 8022 18828 8434
rect 18788 8016 18840 8022
rect 18984 7993 19012 10406
rect 19352 10305 19380 10406
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19338 10296 19394 10305
rect 19622 10288 19918 10308
rect 19338 10231 19394 10240
rect 19430 10160 19486 10169
rect 19430 10095 19432 10104
rect 19484 10095 19486 10104
rect 19432 10066 19484 10072
rect 19444 9722 19472 10066
rect 19614 10024 19670 10033
rect 19614 9959 19616 9968
rect 19668 9959 19670 9968
rect 19616 9930 19668 9936
rect 19432 9716 19484 9722
rect 19432 9658 19484 9664
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19800 8832 19852 8838
rect 19800 8774 19852 8780
rect 19248 8560 19300 8566
rect 19812 8537 19840 8774
rect 19996 8634 20024 18022
rect 20180 9654 20208 20334
rect 24122 20224 24178 20233
rect 24122 20159 24178 20168
rect 20260 19304 20312 19310
rect 20812 19304 20864 19310
rect 20260 19246 20312 19252
rect 20810 19272 20812 19281
rect 20864 19272 20866 19281
rect 20272 18222 20300 19246
rect 20810 19207 20866 19216
rect 20260 18216 20312 18222
rect 20260 18158 20312 18164
rect 23570 17096 23626 17105
rect 23570 17031 23626 17040
rect 20258 15328 20314 15337
rect 20258 15263 20314 15272
rect 20168 9648 20220 9654
rect 20168 9590 20220 9596
rect 20076 9036 20128 9042
rect 20076 8978 20128 8984
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 19248 8502 19300 8508
rect 19798 8528 19854 8537
rect 19156 8288 19208 8294
rect 19062 8256 19118 8265
rect 19156 8230 19208 8236
rect 19062 8191 19118 8200
rect 18788 7958 18840 7964
rect 18970 7984 19026 7993
rect 18970 7919 19026 7928
rect 19076 6866 19104 8191
rect 19168 7886 19196 8230
rect 19156 7880 19208 7886
rect 19156 7822 19208 7828
rect 19168 7546 19196 7822
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 19064 6860 19116 6866
rect 19064 6802 19116 6808
rect 18880 6656 18932 6662
rect 18880 6598 18932 6604
rect 18892 6254 18920 6598
rect 19076 6458 19104 6802
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 18880 6248 18932 6254
rect 18880 6190 18932 6196
rect 19260 5846 19288 8502
rect 19798 8463 19854 8472
rect 20088 8430 20116 8978
rect 20076 8424 20128 8430
rect 20074 8392 20076 8401
rect 20128 8392 20130 8401
rect 20074 8327 20130 8336
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 20272 7546 20300 15263
rect 23478 13968 23534 13977
rect 23478 13903 23534 13912
rect 23492 12345 23520 13903
rect 23584 12753 23612 17031
rect 23570 12744 23626 12753
rect 23570 12679 23626 12688
rect 23478 12336 23534 12345
rect 23478 12271 23534 12280
rect 24136 11801 24164 20159
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24122 11792 24178 11801
rect 24122 11727 24178 11736
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 20260 7540 20312 7546
rect 20260 7482 20312 7488
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 19430 7168 19486 7177
rect 19352 7041 19380 7142
rect 19430 7103 19486 7112
rect 19338 7032 19394 7041
rect 19338 6967 19394 6976
rect 19444 6866 19472 7103
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19444 6458 19472 6802
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 19432 6248 19484 6254
rect 19628 6225 19656 6734
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 19432 6190 19484 6196
rect 19614 6216 19670 6225
rect 19248 5840 19300 5846
rect 19248 5782 19300 5788
rect 19260 5370 19288 5782
rect 19444 5710 19472 6190
rect 19614 6151 19670 6160
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 20718 5808 20774 5817
rect 20718 5743 20774 5752
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 19352 5370 19380 5646
rect 19248 5364 19300 5370
rect 19248 5306 19300 5312
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19260 5030 19288 5306
rect 19248 5024 19300 5030
rect 19248 4966 19300 4972
rect 19352 4826 19380 5306
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 20732 4826 20760 5743
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 19340 4684 19392 4690
rect 19340 4626 19392 4632
rect 21364 4684 21416 4690
rect 21364 4626 21416 4632
rect 19352 3942 19380 4626
rect 21376 3942 21404 4626
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 19340 3936 19392 3942
rect 21364 3936 21416 3942
rect 19340 3878 19392 3884
rect 21362 3904 21364 3913
rect 21416 3904 21418 3913
rect 18892 3369 18920 3878
rect 19352 3641 19380 3878
rect 19622 3836 19918 3856
rect 21362 3839 21418 3848
rect 23202 3904 23258 3913
rect 23202 3839 23258 3848
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19622 3760 19918 3780
rect 19338 3632 19394 3641
rect 19338 3567 19394 3576
rect 18878 3360 18934 3369
rect 18878 3295 18934 3304
rect 20074 3360 20130 3369
rect 20074 3295 20130 3304
rect 18696 3188 18748 3194
rect 18696 3130 18748 3136
rect 19062 2952 19118 2961
rect 19062 2887 19064 2896
rect 19116 2887 19118 2896
rect 19064 2858 19116 2864
rect 19062 2816 19118 2825
rect 19062 2751 19118 2760
rect 18328 2644 18380 2650
rect 18328 2586 18380 2592
rect 18234 2544 18290 2553
rect 18234 2479 18290 2488
rect 18052 2372 18104 2378
rect 18052 2314 18104 2320
rect 18064 480 18092 2314
rect 19076 480 19104 2751
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 20088 480 20116 3295
rect 22190 3224 22246 3233
rect 22190 3159 22246 3168
rect 21180 2304 21232 2310
rect 21180 2246 21232 2252
rect 21192 480 21220 2246
rect 22204 480 22232 3159
rect 23216 480 23244 3839
rect 26330 3632 26386 3641
rect 26330 3567 26386 3576
rect 25318 3496 25374 3505
rect 25318 3431 25374 3440
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24214 2952 24270 2961
rect 24214 2887 24270 2896
rect 24228 480 24256 2887
rect 24676 2644 24728 2650
rect 24676 2586 24728 2592
rect 24688 2553 24716 2586
rect 24674 2544 24730 2553
rect 24674 2479 24730 2488
rect 25136 2508 25188 2514
rect 25136 2450 25188 2456
rect 25148 2310 25176 2450
rect 25136 2304 25188 2310
rect 25134 2272 25136 2281
rect 25188 2272 25190 2281
rect 24289 2204 24585 2224
rect 25134 2207 25190 2216
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 25332 480 25360 3431
rect 26344 480 26372 3567
rect 27342 2272 27398 2281
rect 27342 2207 27398 2216
rect 27356 480 27384 2207
rect 478 0 534 480
rect 1490 0 1546 480
rect 2502 0 2558 480
rect 3514 0 3570 480
rect 4618 0 4674 480
rect 5630 0 5686 480
rect 6642 0 6698 480
rect 7654 0 7710 480
rect 8758 0 8814 480
rect 9770 0 9826 480
rect 10782 0 10838 480
rect 11794 0 11850 480
rect 12898 0 12954 480
rect 13910 0 13966 480
rect 14922 0 14978 480
rect 15934 0 15990 480
rect 17038 0 17094 480
rect 18050 0 18106 480
rect 19062 0 19118 480
rect 20074 0 20130 480
rect 21178 0 21234 480
rect 22190 0 22246 480
rect 23202 0 23258 480
rect 24214 0 24270 480
rect 25318 0 25374 480
rect 26330 0 26386 480
rect 27342 0 27398 480
<< via2 >>
rect 2778 27240 2834 27296
rect 2502 23704 2558 23760
rect 2686 23604 2688 23624
rect 2688 23604 2740 23624
rect 2740 23604 2742 23624
rect 2686 23568 2742 23604
rect 1766 16632 1822 16688
rect 1582 13232 1638 13288
rect 1582 11892 1638 11928
rect 1582 11872 1584 11892
rect 1584 11872 1636 11892
rect 1636 11872 1638 11892
rect 2042 13812 2044 13832
rect 2044 13812 2096 13832
rect 2096 13812 2098 13832
rect 2042 13776 2098 13812
rect 1950 12144 2006 12200
rect 1398 10512 1454 10568
rect 1674 9580 1730 9616
rect 1674 9560 1676 9580
rect 1676 9560 1728 9580
rect 1728 9560 1730 9580
rect 1582 9016 1638 9072
rect 1582 7656 1638 7712
rect 1582 6332 1584 6352
rect 1584 6332 1636 6352
rect 1636 6332 1638 6352
rect 1582 6296 1638 6332
rect 1674 6024 1730 6080
rect 1582 4800 1638 4856
rect 478 3032 534 3088
rect 2134 10104 2190 10160
rect 2042 4972 2044 4992
rect 2044 4972 2096 4992
rect 2096 4972 2098 4992
rect 2042 4936 2098 4972
rect 1766 4120 1822 4176
rect 1950 4020 1952 4040
rect 1952 4020 2004 4040
rect 2004 4020 2006 4040
rect 1950 3984 2006 4020
rect 2962 25880 3018 25936
rect 3514 24792 3570 24848
rect 3330 24520 3386 24576
rect 3422 23024 3478 23080
rect 3330 20440 3386 20496
rect 3882 20304 3938 20360
rect 3422 19216 3478 19272
rect 3882 18264 3938 18320
rect 2502 15580 2504 15600
rect 2504 15580 2556 15600
rect 2556 15580 2558 15600
rect 2502 15544 2558 15580
rect 4250 16632 4306 16688
rect 3054 15544 3110 15600
rect 4710 15544 4766 15600
rect 3974 15020 4030 15056
rect 3974 15000 3976 15020
rect 3976 15000 4028 15020
rect 4028 15000 4030 15020
rect 2962 14356 2964 14376
rect 2964 14356 3016 14376
rect 3016 14356 3018 14376
rect 2962 14320 3018 14356
rect 3514 12724 3516 12744
rect 3516 12724 3568 12744
rect 3568 12724 3570 12744
rect 3514 12688 3570 12724
rect 4526 13640 4582 13696
rect 4342 13504 4398 13560
rect 4710 13912 4766 13968
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 6550 24792 6606 24848
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 6274 23704 6330 23760
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 4894 13232 4950 13288
rect 4710 12280 4766 12336
rect 4894 12180 4896 12200
rect 4896 12180 4948 12200
rect 4948 12180 4950 12200
rect 4894 12144 4950 12180
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5998 13504 6054 13560
rect 7010 18808 7066 18864
rect 6274 17332 6330 17368
rect 6274 17312 6276 17332
rect 6276 17312 6328 17332
rect 6328 17312 6330 17332
rect 6366 14864 6422 14920
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5998 12688 6054 12744
rect 3514 11328 3570 11384
rect 3422 11056 3478 11112
rect 3238 9152 3294 9208
rect 5170 11328 5226 11384
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5446 11328 5502 11384
rect 4066 10648 4122 10704
rect 4250 9560 4306 9616
rect 6274 12708 6330 12744
rect 6274 12688 6276 12708
rect 6276 12688 6328 12708
rect 6328 12688 6330 12708
rect 6274 12008 6330 12064
rect 5906 11056 5962 11112
rect 6274 11192 6330 11248
rect 6458 11328 6514 11384
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 4986 10648 5042 10704
rect 2410 6840 2466 6896
rect 2962 6840 3018 6896
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 6090 10104 6146 10160
rect 5998 9152 6054 9208
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 6642 10804 6698 10840
rect 6642 10784 6644 10804
rect 6644 10784 6696 10804
rect 6696 10784 6698 10804
rect 3514 3712 3570 3768
rect 1582 3440 1638 3496
rect 2410 3476 2412 3496
rect 2412 3476 2464 3496
rect 2464 3476 2466 3496
rect 2410 3440 2466 3476
rect 2502 2760 2558 2816
rect 1950 2252 1952 2272
rect 1952 2252 2004 2272
rect 2004 2252 2006 2272
rect 1950 2216 2006 2252
rect 1582 2080 1638 2136
rect 2686 2644 2742 2680
rect 2686 2624 2688 2644
rect 2688 2624 2740 2644
rect 2740 2624 2742 2644
rect 5078 3440 5134 3496
rect 4342 2624 4398 2680
rect 4618 2216 4674 2272
rect 4066 720 4122 776
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 7102 10648 7158 10704
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10138 24656 10194 24712
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 9770 23568 9826 23624
rect 8574 20848 8630 20904
rect 8114 19624 8170 19680
rect 8206 19352 8262 19408
rect 7746 19216 7802 19272
rect 7654 18944 7710 19000
rect 7654 18808 7710 18864
rect 7286 15000 7342 15056
rect 7378 12008 7434 12064
rect 8574 19216 8630 19272
rect 8206 18148 8262 18184
rect 8206 18128 8208 18148
rect 8208 18128 8260 18148
rect 8260 18128 8262 18148
rect 8114 15408 8170 15464
rect 7930 12824 7986 12880
rect 7654 11892 7710 11928
rect 7654 11872 7656 11892
rect 7656 11872 7708 11892
rect 7708 11872 7710 11892
rect 6550 6296 6606 6352
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 7194 9424 7250 9480
rect 6826 4936 6882 4992
rect 5538 3984 5594 4040
rect 6734 3984 6790 4040
rect 6642 3848 6698 3904
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 7378 5616 7434 5672
rect 8390 13776 8446 13832
rect 8482 13640 8538 13696
rect 11794 24656 11850 24712
rect 8942 21428 8944 21448
rect 8944 21428 8996 21448
rect 8996 21428 8998 21448
rect 8942 21392 8998 21428
rect 9126 19796 9128 19816
rect 9128 19796 9180 19816
rect 9180 19796 9182 19816
rect 9126 19760 9182 19796
rect 8942 19252 8944 19272
rect 8944 19252 8996 19272
rect 8996 19252 8998 19272
rect 8942 19216 8998 19252
rect 8206 10920 8262 10976
rect 8758 12980 8814 13016
rect 8758 12960 8760 12980
rect 8760 12960 8812 12980
rect 8812 12960 8814 12980
rect 8666 10648 8722 10704
rect 9310 18400 9366 18456
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10230 19660 10232 19680
rect 10232 19660 10284 19680
rect 10284 19660 10286 19680
rect 10230 19624 10286 19660
rect 10414 19352 10470 19408
rect 12254 23724 12310 23760
rect 12254 23704 12256 23724
rect 12256 23704 12308 23724
rect 12308 23704 12310 23724
rect 14094 24792 14150 24848
rect 11886 21528 11942 21584
rect 11978 20848 12034 20904
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10046 18128 10102 18184
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 9494 13912 9550 13968
rect 9218 13368 9274 13424
rect 8850 10512 8906 10568
rect 7378 3168 7434 3224
rect 7378 2760 7434 2816
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10046 15444 10048 15464
rect 10048 15444 10100 15464
rect 10100 15444 10102 15464
rect 10046 15408 10102 15444
rect 10414 14884 10470 14920
rect 10414 14864 10416 14884
rect 10416 14864 10468 14884
rect 10468 14864 10470 14884
rect 10046 14728 10102 14784
rect 9770 14356 9772 14376
rect 9772 14356 9824 14376
rect 9824 14356 9826 14376
rect 9770 14320 9826 14356
rect 9494 11636 9496 11656
rect 9496 11636 9548 11656
rect 9548 11636 9550 11656
rect 9494 11600 9550 11636
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10598 13948 10600 13968
rect 10600 13948 10652 13968
rect 10652 13948 10654 13968
rect 10598 13912 10654 13948
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 11794 15680 11850 15736
rect 11426 13268 11428 13288
rect 11428 13268 11480 13288
rect 11480 13268 11482 13288
rect 11426 13232 11482 13268
rect 11518 12960 11574 13016
rect 11058 12688 11114 12744
rect 10322 12280 10378 12336
rect 10966 11736 11022 11792
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10966 11212 11022 11248
rect 10966 11192 10968 11212
rect 10968 11192 11020 11212
rect 11020 11192 11022 11212
rect 10782 10920 10838 10976
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10138 9560 10194 9616
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10598 8492 10654 8528
rect 10598 8472 10600 8492
rect 10600 8472 10652 8492
rect 10652 8472 10654 8492
rect 11058 10512 11114 10568
rect 10966 9152 11022 9208
rect 11702 12688 11758 12744
rect 12162 11872 12218 11928
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10874 8336 10930 8392
rect 9310 6024 9366 6080
rect 9954 6160 10010 6216
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 11150 8200 11206 8256
rect 11242 5616 11298 5672
rect 11058 5072 11114 5128
rect 9678 3884 9680 3904
rect 9680 3884 9732 3904
rect 9732 3884 9734 3904
rect 8942 2896 8998 2952
rect 9678 3848 9734 3884
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10046 4120 10102 4176
rect 9862 3712 9918 3768
rect 9954 3068 9956 3088
rect 9956 3068 10008 3088
rect 10008 3068 10010 3088
rect 9954 3032 10010 3068
rect 10782 3884 10784 3904
rect 10784 3884 10836 3904
rect 10836 3884 10838 3904
rect 10782 3848 10838 3884
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 12898 23160 12954 23216
rect 13082 21392 13138 21448
rect 13450 21292 13452 21312
rect 13452 21292 13504 21312
rect 13504 21292 13506 21312
rect 13450 21256 13506 21292
rect 12898 19760 12954 19816
rect 12806 19352 12862 19408
rect 12346 16768 12402 16824
rect 12530 9424 12586 9480
rect 11334 4020 11336 4040
rect 11336 4020 11388 4040
rect 11388 4020 11390 4040
rect 11334 3984 11390 4020
rect 11242 3596 11298 3632
rect 11242 3576 11244 3596
rect 11244 3576 11296 3596
rect 11296 3576 11298 3596
rect 11886 3052 11942 3088
rect 11886 3032 11888 3052
rect 11888 3032 11940 3052
rect 11940 3032 11942 3052
rect 12438 5772 12494 5808
rect 12438 5752 12440 5772
rect 12440 5752 12492 5772
rect 12492 5752 12494 5772
rect 13818 23296 13874 23352
rect 13726 21392 13782 21448
rect 13542 20304 13598 20360
rect 13542 19352 13598 19408
rect 12990 18400 13046 18456
rect 12990 18164 12992 18184
rect 12992 18164 13044 18184
rect 13044 18164 13046 18184
rect 12990 18128 13046 18164
rect 13266 17312 13322 17368
rect 13358 17076 13360 17096
rect 13360 17076 13412 17096
rect 13412 17076 13414 17096
rect 13358 17040 13414 17076
rect 13634 15680 13690 15736
rect 13910 19216 13966 19272
rect 14462 17992 14518 18048
rect 14370 16652 14426 16688
rect 14370 16632 14372 16652
rect 14372 16632 14424 16652
rect 14424 16632 14426 16652
rect 13266 14728 13322 14784
rect 12898 10784 12954 10840
rect 12806 6160 12862 6216
rect 12714 5092 12770 5128
rect 12714 5072 12716 5092
rect 12716 5072 12768 5092
rect 12768 5072 12770 5092
rect 12162 3576 12218 3632
rect 12070 3168 12126 3224
rect 13726 15444 13728 15464
rect 13728 15444 13780 15464
rect 13780 15444 13782 15464
rect 13726 15408 13782 15444
rect 14554 15580 14556 15600
rect 14556 15580 14608 15600
rect 14608 15580 14610 15600
rect 14554 15544 14610 15580
rect 14646 15408 14702 15464
rect 14002 14320 14058 14376
rect 14186 13932 14242 13968
rect 14186 13912 14188 13932
rect 14188 13912 14240 13932
rect 14240 13912 14242 13932
rect 13634 11600 13690 11656
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 15934 24792 15990 24848
rect 16670 24812 16726 24848
rect 16670 24792 16672 24812
rect 16672 24792 16724 24812
rect 16724 24792 16726 24812
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 15474 23296 15530 23352
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 15750 21428 15752 21448
rect 15752 21428 15804 21448
rect 15804 21428 15806 21448
rect 15750 21392 15806 21428
rect 15382 20848 15438 20904
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 15198 20340 15200 20360
rect 15200 20340 15252 20360
rect 15252 20340 15254 20360
rect 15198 20304 15254 20340
rect 15566 19896 15622 19952
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 16394 24132 16450 24168
rect 16394 24112 16396 24132
rect 16396 24112 16448 24132
rect 16448 24112 16450 24132
rect 15934 19236 15990 19272
rect 15934 19216 15936 19236
rect 15936 19216 15988 19236
rect 15988 19216 15990 19236
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 15382 18128 15438 18184
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 15290 17196 15346 17232
rect 15290 17176 15292 17196
rect 15292 17176 15344 17196
rect 15344 17176 15346 17196
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14186 12960 14242 13016
rect 14002 12552 14058 12608
rect 14094 11328 14150 11384
rect 14002 8472 14058 8528
rect 14370 12552 14426 12608
rect 14278 12280 14334 12336
rect 14278 12008 14334 12064
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 16026 17992 16082 18048
rect 15566 17040 15622 17096
rect 15750 15700 15806 15736
rect 15750 15680 15752 15700
rect 15752 15680 15804 15700
rect 15804 15680 15806 15700
rect 18326 24268 18382 24304
rect 18326 24248 18328 24268
rect 18328 24248 18380 24268
rect 18380 24248 18382 24268
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 20074 24248 20130 24304
rect 18602 21256 18658 21312
rect 17774 20032 17830 20088
rect 18510 19760 18566 19816
rect 18050 17176 18106 17232
rect 17958 16668 17960 16688
rect 17960 16668 18012 16688
rect 18012 16668 18014 16688
rect 17958 16632 18014 16668
rect 17314 16108 17370 16144
rect 17314 16088 17316 16108
rect 17316 16088 17368 16108
rect 17368 16088 17370 16108
rect 15750 13640 15806 13696
rect 15290 12144 15346 12200
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14370 11600 14426 11656
rect 14278 10240 14334 10296
rect 14738 11092 14740 11112
rect 14740 11092 14792 11112
rect 14792 11092 14794 11112
rect 14738 11056 14794 11092
rect 14646 10240 14702 10296
rect 14186 9016 14242 9072
rect 14278 8472 14334 8528
rect 13634 4972 13636 4992
rect 13636 4972 13688 4992
rect 13688 4972 13690 4992
rect 13634 4936 13690 4972
rect 15750 11872 15806 11928
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 15474 11192 15530 11248
rect 15014 10376 15070 10432
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14830 7928 14886 7984
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 15750 11328 15806 11384
rect 16026 10124 16082 10160
rect 16026 10104 16028 10124
rect 16028 10104 16080 10124
rect 16080 10104 16082 10124
rect 18326 16768 18382 16824
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 19982 23160 20038 23216
rect 23202 24792 23258 24848
rect 23478 24112 23534 24168
rect 20166 23024 20222 23080
rect 19798 22772 19854 22808
rect 24766 26424 24822 26480
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24674 24384 24730 24440
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 27342 24384 27398 24440
rect 25318 23704 25374 23760
rect 24214 23024 24270 23080
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 19798 22752 19800 22772
rect 19800 22752 19852 22772
rect 19852 22752 19854 22772
rect 23478 22752 23534 22808
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19338 20032 19394 20088
rect 19338 19932 19340 19952
rect 19340 19932 19392 19952
rect 19392 19932 19394 19952
rect 19338 19896 19394 19932
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 19614 20440 19670 20496
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19614 19896 19670 19952
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19614 18264 19670 18320
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 17314 15272 17370 15328
rect 18050 15544 18106 15600
rect 16302 13796 16358 13832
rect 16302 13776 16304 13796
rect 16304 13776 16356 13796
rect 16356 13776 16358 13796
rect 16302 13524 16358 13560
rect 16302 13504 16304 13524
rect 16304 13504 16356 13524
rect 16356 13504 16358 13524
rect 16210 12280 16266 12336
rect 17222 14456 17278 14512
rect 16762 12180 16764 12200
rect 16764 12180 16816 12200
rect 16816 12180 16818 12200
rect 16762 12144 16818 12180
rect 16118 9172 16174 9208
rect 16118 9152 16120 9172
rect 16120 9152 16172 9172
rect 16172 9152 16174 9172
rect 15934 8200 15990 8256
rect 14738 7112 14794 7168
rect 13910 4120 13966 4176
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 18970 15408 19026 15464
rect 18050 14320 18106 14376
rect 16946 11076 17002 11112
rect 16946 11056 16948 11076
rect 16948 11056 17000 11076
rect 17000 11056 17002 11076
rect 16762 9988 16818 10024
rect 16762 9968 16764 9988
rect 16764 9968 16816 9988
rect 16816 9968 16818 9988
rect 16394 8472 16450 8528
rect 14830 6332 14832 6352
rect 14832 6332 14884 6352
rect 14884 6332 14886 6352
rect 14830 6296 14886 6332
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 15382 5752 15438 5808
rect 15290 4936 15346 4992
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 16578 7948 16634 7984
rect 16578 7928 16580 7948
rect 16580 7928 16632 7948
rect 16632 7928 16634 7948
rect 15750 6160 15806 6216
rect 15474 4120 15530 4176
rect 16210 3884 16212 3904
rect 16212 3884 16264 3904
rect 16264 3884 16266 3904
rect 16210 3848 16266 3884
rect 16026 3576 16082 3632
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 15658 3188 15714 3224
rect 15658 3168 15660 3188
rect 15660 3168 15712 3188
rect 15712 3168 15714 3188
rect 12990 1536 13046 1592
rect 14278 2896 14334 2952
rect 14462 2760 14518 2816
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 18050 11212 18106 11248
rect 18050 11192 18052 11212
rect 18052 11192 18104 11212
rect 18104 11192 18106 11212
rect 18050 10648 18106 10704
rect 17406 10512 17462 10568
rect 18142 9016 18198 9072
rect 17590 6976 17646 7032
rect 17406 4800 17462 4856
rect 18142 5752 18198 5808
rect 17038 2760 17094 2816
rect 17866 2760 17922 2816
rect 18418 13776 18474 13832
rect 19430 14728 19486 14784
rect 19338 14456 19394 14512
rect 19338 13932 19394 13968
rect 19338 13912 19340 13932
rect 19340 13912 19392 13932
rect 19392 13912 19394 13932
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19338 13640 19394 13696
rect 19246 13504 19302 13560
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 18418 10648 18474 10704
rect 19798 13388 19854 13424
rect 19798 13368 19800 13388
rect 19800 13368 19852 13388
rect 19852 13368 19854 13388
rect 19798 12860 19800 12880
rect 19800 12860 19852 12880
rect 19852 12860 19854 12880
rect 19798 12824 19854 12860
rect 18602 10376 18658 10432
rect 18418 4800 18474 4856
rect 19338 12552 19394 12608
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19338 12144 19394 12200
rect 19798 11892 19854 11928
rect 19798 11872 19800 11892
rect 19800 11872 19852 11892
rect 19852 11872 19854 11892
rect 19614 11636 19616 11656
rect 19616 11636 19668 11656
rect 19668 11636 19670 11656
rect 19614 11600 19670 11636
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19338 11056 19394 11112
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19338 10240 19394 10296
rect 19430 10124 19486 10160
rect 19430 10104 19432 10124
rect 19432 10104 19484 10124
rect 19484 10104 19486 10124
rect 19614 9988 19670 10024
rect 19614 9968 19616 9988
rect 19616 9968 19668 9988
rect 19668 9968 19670 9988
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 24122 20168 24178 20224
rect 20810 19252 20812 19272
rect 20812 19252 20864 19272
rect 20864 19252 20866 19272
rect 20810 19216 20866 19252
rect 23570 17040 23626 17096
rect 20258 15272 20314 15328
rect 19062 8200 19118 8256
rect 18970 7928 19026 7984
rect 19798 8472 19854 8528
rect 20074 8372 20076 8392
rect 20076 8372 20128 8392
rect 20128 8372 20130 8392
rect 20074 8336 20130 8372
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 23478 13912 23534 13968
rect 23570 12688 23626 12744
rect 23478 12280 23534 12336
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24122 11736 24178 11792
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 19430 7112 19486 7168
rect 19338 6976 19394 7032
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 19614 6160 19670 6216
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 20718 5752 20774 5808
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 21362 3884 21364 3904
rect 21364 3884 21416 3904
rect 21416 3884 21418 3904
rect 21362 3848 21418 3884
rect 23202 3848 23258 3904
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19338 3576 19394 3632
rect 18878 3304 18934 3360
rect 20074 3304 20130 3360
rect 19062 2916 19118 2952
rect 19062 2896 19064 2916
rect 19064 2896 19116 2916
rect 19116 2896 19118 2916
rect 19062 2760 19118 2816
rect 18234 2488 18290 2544
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 22190 3168 22246 3224
rect 26330 3576 26386 3632
rect 25318 3440 25374 3496
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24214 2896 24270 2952
rect 24674 2488 24730 2544
rect 25134 2252 25136 2272
rect 25136 2252 25188 2272
rect 25188 2252 25190 2272
rect 25134 2216 25190 2252
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 27342 2216 27398 2272
<< metal3 >>
rect 0 27298 480 27328
rect 2773 27298 2839 27301
rect 0 27296 2839 27298
rect 0 27240 2778 27296
rect 2834 27240 2839 27296
rect 0 27238 2839 27240
rect 0 27208 480 27238
rect 2773 27235 2839 27238
rect 24761 26482 24827 26485
rect 27520 26482 28000 26512
rect 24761 26480 28000 26482
rect 24761 26424 24766 26480
rect 24822 26424 28000 26480
rect 24761 26422 28000 26424
rect 24761 26419 24827 26422
rect 27520 26392 28000 26422
rect 0 25938 480 25968
rect 2957 25938 3023 25941
rect 0 25936 3023 25938
rect 0 25880 2962 25936
rect 3018 25880 3023 25936
rect 0 25878 3023 25880
rect 0 25848 480 25878
rect 2957 25875 3023 25878
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 3509 24850 3575 24853
rect 6545 24850 6611 24853
rect 3509 24848 6611 24850
rect 3509 24792 3514 24848
rect 3570 24792 6550 24848
rect 6606 24792 6611 24848
rect 3509 24790 6611 24792
rect 3509 24787 3575 24790
rect 6545 24787 6611 24790
rect 14089 24850 14155 24853
rect 15929 24850 15995 24853
rect 14089 24848 15995 24850
rect 14089 24792 14094 24848
rect 14150 24792 15934 24848
rect 15990 24792 15995 24848
rect 14089 24790 15995 24792
rect 14089 24787 14155 24790
rect 15929 24787 15995 24790
rect 16665 24850 16731 24853
rect 23197 24850 23263 24853
rect 16665 24848 23263 24850
rect 16665 24792 16670 24848
rect 16726 24792 23202 24848
rect 23258 24792 23263 24848
rect 16665 24790 23263 24792
rect 16665 24787 16731 24790
rect 23197 24787 23263 24790
rect 10133 24714 10199 24717
rect 11789 24714 11855 24717
rect 10133 24712 11855 24714
rect 10133 24656 10138 24712
rect 10194 24656 11794 24712
rect 11850 24656 11855 24712
rect 10133 24654 11855 24656
rect 10133 24651 10199 24654
rect 11789 24651 11855 24654
rect 0 24578 480 24608
rect 3325 24578 3391 24581
rect 0 24576 3391 24578
rect 0 24520 3330 24576
rect 3386 24520 3391 24576
rect 0 24518 3391 24520
rect 0 24488 480 24518
rect 3325 24515 3391 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 24669 24442 24735 24445
rect 27337 24442 27403 24445
rect 24669 24440 27403 24442
rect 24669 24384 24674 24440
rect 24730 24384 27342 24440
rect 27398 24384 27403 24440
rect 24669 24382 27403 24384
rect 24669 24379 24735 24382
rect 27337 24379 27403 24382
rect 18321 24306 18387 24309
rect 20069 24306 20135 24309
rect 18321 24304 20135 24306
rect 18321 24248 18326 24304
rect 18382 24248 20074 24304
rect 20130 24248 20135 24304
rect 18321 24246 20135 24248
rect 18321 24243 18387 24246
rect 20069 24243 20135 24246
rect 16389 24170 16455 24173
rect 23473 24170 23539 24173
rect 16389 24168 23539 24170
rect 16389 24112 16394 24168
rect 16450 24112 23478 24168
rect 23534 24112 23539 24168
rect 16389 24110 23539 24112
rect 16389 24107 16455 24110
rect 23473 24107 23539 24110
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 2497 23762 2563 23765
rect 6269 23762 6335 23765
rect 2497 23760 6335 23762
rect 2497 23704 2502 23760
rect 2558 23704 6274 23760
rect 6330 23704 6335 23760
rect 2497 23702 6335 23704
rect 2497 23699 2563 23702
rect 6269 23699 6335 23702
rect 12249 23762 12315 23765
rect 25313 23762 25379 23765
rect 12249 23760 25379 23762
rect 12249 23704 12254 23760
rect 12310 23704 25318 23760
rect 25374 23704 25379 23760
rect 12249 23702 25379 23704
rect 12249 23699 12315 23702
rect 25313 23699 25379 23702
rect 2681 23626 2747 23629
rect 9765 23626 9831 23629
rect 2681 23624 9831 23626
rect 2681 23568 2686 23624
rect 2742 23568 9770 23624
rect 9826 23568 9831 23624
rect 2681 23566 9831 23568
rect 2681 23563 2747 23566
rect 9765 23563 9831 23566
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 13813 23354 13879 23357
rect 15469 23354 15535 23357
rect 13813 23352 15535 23354
rect 13813 23296 13818 23352
rect 13874 23296 15474 23352
rect 15530 23296 15535 23352
rect 13813 23294 15535 23296
rect 13813 23291 13879 23294
rect 15469 23291 15535 23294
rect 23974 23292 23980 23356
rect 24044 23354 24050 23356
rect 27520 23354 28000 23384
rect 24044 23294 28000 23354
rect 24044 23292 24050 23294
rect 27520 23264 28000 23294
rect 12893 23218 12959 23221
rect 19977 23218 20043 23221
rect 12893 23216 20043 23218
rect 12893 23160 12898 23216
rect 12954 23160 19982 23216
rect 20038 23160 20043 23216
rect 12893 23158 20043 23160
rect 12893 23155 12959 23158
rect 19977 23155 20043 23158
rect 0 23082 480 23112
rect 3417 23082 3483 23085
rect 0 23080 3483 23082
rect 0 23024 3422 23080
rect 3478 23024 3483 23080
rect 0 23022 3483 23024
rect 0 22992 480 23022
rect 3417 23019 3483 23022
rect 20161 23082 20227 23085
rect 24209 23082 24275 23085
rect 20161 23080 24275 23082
rect 20161 23024 20166 23080
rect 20222 23024 24214 23080
rect 24270 23024 24275 23080
rect 20161 23022 24275 23024
rect 20161 23019 20227 23022
rect 24209 23019 24275 23022
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 19793 22810 19859 22813
rect 23473 22810 23539 22813
rect 19793 22808 23539 22810
rect 19793 22752 19798 22808
rect 19854 22752 23478 22808
rect 23534 22752 23539 22808
rect 19793 22750 23539 22752
rect 19793 22747 19859 22750
rect 23473 22747 23539 22750
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 5610 21792 5930 21793
rect 0 21722 480 21752
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 0 21662 2698 21722
rect 0 21632 480 21662
rect 2638 21586 2698 21662
rect 11881 21586 11947 21589
rect 2638 21552 2744 21586
rect 2822 21584 11947 21586
rect 2822 21552 11886 21584
rect 2638 21528 11886 21552
rect 11942 21528 11947 21584
rect 2638 21526 11947 21528
rect 2684 21492 2882 21526
rect 11881 21523 11947 21526
rect 8937 21450 9003 21453
rect 13077 21450 13143 21453
rect 13721 21450 13787 21453
rect 15745 21450 15811 21453
rect 8937 21448 15811 21450
rect 8937 21392 8942 21448
rect 8998 21392 13082 21448
rect 13138 21392 13726 21448
rect 13782 21392 15750 21448
rect 15806 21392 15811 21448
rect 8937 21390 15811 21392
rect 8937 21387 9003 21390
rect 13077 21387 13143 21390
rect 13721 21387 13787 21390
rect 15745 21387 15811 21390
rect 13445 21314 13511 21317
rect 18597 21314 18663 21317
rect 13445 21312 18663 21314
rect 13445 21256 13450 21312
rect 13506 21256 18602 21312
rect 18658 21256 18663 21312
rect 13445 21254 18663 21256
rect 13445 21251 13511 21254
rect 18597 21251 18663 21254
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 8569 20906 8635 20909
rect 11973 20906 12039 20909
rect 15377 20906 15443 20909
rect 8569 20904 15443 20906
rect 8569 20848 8574 20904
rect 8630 20848 11978 20904
rect 12034 20848 15382 20904
rect 15438 20848 15443 20904
rect 8569 20846 15443 20848
rect 8569 20843 8635 20846
rect 11973 20843 12039 20846
rect 15377 20843 15443 20846
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 3325 20498 3391 20501
rect 19609 20498 19675 20501
rect 3325 20496 19675 20498
rect 3325 20440 3330 20496
rect 3386 20440 19614 20496
rect 19670 20440 19675 20496
rect 3325 20438 19675 20440
rect 3325 20435 3391 20438
rect 19609 20435 19675 20438
rect 0 20362 480 20392
rect 3877 20362 3943 20365
rect 0 20360 3943 20362
rect 0 20304 3882 20360
rect 3938 20304 3943 20360
rect 0 20302 3943 20304
rect 0 20272 480 20302
rect 3877 20299 3943 20302
rect 13537 20362 13603 20365
rect 15193 20362 15259 20365
rect 13537 20360 15259 20362
rect 13537 20304 13542 20360
rect 13598 20304 15198 20360
rect 15254 20304 15259 20360
rect 13537 20302 15259 20304
rect 13537 20299 13603 20302
rect 15193 20299 15259 20302
rect 24117 20226 24183 20229
rect 27520 20226 28000 20256
rect 24117 20224 28000 20226
rect 24117 20168 24122 20224
rect 24178 20168 28000 20224
rect 24117 20166 28000 20168
rect 24117 20163 24183 20166
rect 10277 20160 10597 20161
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 27520 20136 28000 20166
rect 19610 20095 19930 20096
rect 17769 20090 17835 20093
rect 19333 20090 19399 20093
rect 17769 20088 19399 20090
rect 17769 20032 17774 20088
rect 17830 20032 19338 20088
rect 19394 20032 19399 20088
rect 17769 20030 19399 20032
rect 17769 20027 17835 20030
rect 19333 20027 19399 20030
rect 15561 19954 15627 19957
rect 19333 19954 19399 19957
rect 19609 19954 19675 19957
rect 15561 19952 19675 19954
rect 15561 19896 15566 19952
rect 15622 19896 19338 19952
rect 19394 19896 19614 19952
rect 19670 19896 19675 19952
rect 15561 19894 19675 19896
rect 15561 19891 15627 19894
rect 19333 19891 19399 19894
rect 19609 19891 19675 19894
rect 9121 19818 9187 19821
rect 12893 19818 12959 19821
rect 18505 19818 18571 19821
rect 9121 19816 18571 19818
rect 9121 19760 9126 19816
rect 9182 19760 12898 19816
rect 12954 19760 18510 19816
rect 18566 19760 18571 19816
rect 9121 19758 18571 19760
rect 9121 19755 9187 19758
rect 12893 19755 12959 19758
rect 18505 19755 18571 19758
rect 8109 19682 8175 19685
rect 10225 19682 10291 19685
rect 8109 19680 10291 19682
rect 8109 19624 8114 19680
rect 8170 19624 10230 19680
rect 10286 19624 10291 19680
rect 8109 19622 10291 19624
rect 8109 19619 8175 19622
rect 10225 19619 10291 19622
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 8201 19410 8267 19413
rect 10409 19410 10475 19413
rect 8201 19408 10475 19410
rect 8201 19352 8206 19408
rect 8262 19352 10414 19408
rect 10470 19352 10475 19408
rect 8201 19350 10475 19352
rect 8201 19347 8267 19350
rect 10409 19347 10475 19350
rect 12801 19410 12867 19413
rect 13537 19410 13603 19413
rect 12801 19408 13603 19410
rect 12801 19352 12806 19408
rect 12862 19352 13542 19408
rect 13598 19352 13603 19408
rect 12801 19350 13603 19352
rect 12801 19347 12867 19350
rect 13537 19347 13603 19350
rect 3417 19274 3483 19277
rect 7741 19274 7807 19277
rect 8569 19274 8635 19277
rect 3417 19272 8635 19274
rect 3417 19216 3422 19272
rect 3478 19216 7746 19272
rect 7802 19216 8574 19272
rect 8630 19216 8635 19272
rect 3417 19214 8635 19216
rect 3417 19211 3483 19214
rect 7741 19211 7807 19214
rect 8569 19211 8635 19214
rect 8937 19274 9003 19277
rect 13905 19274 13971 19277
rect 8937 19272 13971 19274
rect 8937 19216 8942 19272
rect 8998 19216 13910 19272
rect 13966 19216 13971 19272
rect 8937 19214 13971 19216
rect 8937 19211 9003 19214
rect 13905 19211 13971 19214
rect 15929 19274 15995 19277
rect 20805 19274 20871 19277
rect 15929 19272 20871 19274
rect 15929 19216 15934 19272
rect 15990 19216 20810 19272
rect 20866 19216 20871 19272
rect 15929 19214 20871 19216
rect 15929 19211 15995 19214
rect 20805 19211 20871 19214
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 7649 19000 7715 19005
rect 7649 18944 7654 19000
rect 7710 18944 7715 19000
rect 7649 18939 7715 18944
rect 0 18866 480 18896
rect 7652 18869 7712 18939
rect 7005 18866 7071 18869
rect 0 18864 7071 18866
rect 0 18808 7010 18864
rect 7066 18808 7071 18864
rect 0 18806 7071 18808
rect 0 18776 480 18806
rect 7005 18803 7071 18806
rect 7649 18864 7715 18869
rect 7649 18808 7654 18864
rect 7710 18808 7715 18864
rect 7649 18803 7715 18808
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 9305 18458 9371 18461
rect 12985 18458 13051 18461
rect 9305 18456 13051 18458
rect 9305 18400 9310 18456
rect 9366 18400 12990 18456
rect 13046 18400 13051 18456
rect 9305 18398 13051 18400
rect 9305 18395 9371 18398
rect 12985 18395 13051 18398
rect 3877 18322 3943 18325
rect 19609 18322 19675 18325
rect 3877 18320 19675 18322
rect 3877 18264 3882 18320
rect 3938 18264 19614 18320
rect 19670 18264 19675 18320
rect 3877 18262 19675 18264
rect 3877 18259 3943 18262
rect 19609 18259 19675 18262
rect 8201 18186 8267 18189
rect 10041 18186 10107 18189
rect 8201 18184 10107 18186
rect 8201 18128 8206 18184
rect 8262 18128 10046 18184
rect 10102 18128 10107 18184
rect 8201 18126 10107 18128
rect 8201 18123 8267 18126
rect 10041 18123 10107 18126
rect 12985 18186 13051 18189
rect 15377 18186 15443 18189
rect 12985 18184 15443 18186
rect 12985 18128 12990 18184
rect 13046 18128 15382 18184
rect 15438 18128 15443 18184
rect 12985 18126 15443 18128
rect 12985 18123 13051 18126
rect 15377 18123 15443 18126
rect 14457 18050 14523 18053
rect 16021 18050 16087 18053
rect 14457 18048 16087 18050
rect 14457 17992 14462 18048
rect 14518 17992 16026 18048
rect 16082 17992 16087 18048
rect 14457 17990 16087 17992
rect 14457 17987 14523 17990
rect 16021 17987 16087 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 0 17506 480 17536
rect 0 17446 2698 17506
rect 0 17416 480 17446
rect 2638 17370 2698 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 6269 17370 6335 17373
rect 13261 17370 13327 17373
rect 2638 17310 2882 17370
rect 2822 17234 2882 17310
rect 6269 17368 13327 17370
rect 6269 17312 6274 17368
rect 6330 17312 13266 17368
rect 13322 17312 13327 17368
rect 6269 17310 13327 17312
rect 6269 17307 6335 17310
rect 13261 17307 13327 17310
rect 15285 17234 15351 17237
rect 18045 17234 18111 17237
rect 2822 17232 18111 17234
rect 2822 17176 15290 17232
rect 15346 17176 18050 17232
rect 18106 17176 18111 17232
rect 2822 17174 18111 17176
rect 15285 17171 15351 17174
rect 18045 17171 18111 17174
rect 13353 17098 13419 17101
rect 15561 17098 15627 17101
rect 13353 17096 15627 17098
rect 13353 17040 13358 17096
rect 13414 17040 15566 17096
rect 15622 17040 15627 17096
rect 13353 17038 15627 17040
rect 13353 17035 13419 17038
rect 15561 17035 15627 17038
rect 23565 17098 23631 17101
rect 27520 17098 28000 17128
rect 23565 17096 28000 17098
rect 23565 17040 23570 17096
rect 23626 17040 28000 17096
rect 23565 17038 28000 17040
rect 23565 17035 23631 17038
rect 27520 17008 28000 17038
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 12341 16826 12407 16829
rect 18321 16826 18387 16829
rect 12341 16824 18387 16826
rect 12341 16768 12346 16824
rect 12402 16768 18326 16824
rect 18382 16768 18387 16824
rect 12341 16766 18387 16768
rect 12341 16763 12407 16766
rect 18321 16763 18387 16766
rect 1761 16690 1827 16693
rect 4245 16690 4311 16693
rect 1761 16688 4311 16690
rect 1761 16632 1766 16688
rect 1822 16632 4250 16688
rect 4306 16632 4311 16688
rect 1761 16630 4311 16632
rect 1761 16627 1827 16630
rect 4245 16627 4311 16630
rect 14365 16690 14431 16693
rect 17953 16690 18019 16693
rect 14365 16688 18019 16690
rect 14365 16632 14370 16688
rect 14426 16632 17958 16688
rect 18014 16632 18019 16688
rect 14365 16630 18019 16632
rect 14365 16627 14431 16630
rect 17953 16627 18019 16630
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 0 16146 480 16176
rect 9262 16146 9506 16180
rect 17309 16146 17375 16149
rect 0 16144 17375 16146
rect 0 16120 17314 16144
rect 0 16086 9322 16120
rect 9446 16088 17314 16120
rect 17370 16088 17375 16144
rect 9446 16086 17375 16088
rect 0 16056 480 16086
rect 17309 16083 17375 16086
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 11789 15738 11855 15741
rect 13629 15738 13695 15741
rect 15745 15738 15811 15741
rect 11789 15736 15811 15738
rect 11789 15680 11794 15736
rect 11850 15680 13634 15736
rect 13690 15680 15750 15736
rect 15806 15680 15811 15736
rect 11789 15678 15811 15680
rect 11789 15675 11855 15678
rect 13629 15675 13695 15678
rect 15745 15675 15811 15678
rect 2497 15602 2563 15605
rect 3049 15602 3115 15605
rect 4705 15602 4771 15605
rect 2497 15600 4771 15602
rect 2497 15544 2502 15600
rect 2558 15544 3054 15600
rect 3110 15544 4710 15600
rect 4766 15544 4771 15600
rect 2497 15542 4771 15544
rect 2497 15539 2563 15542
rect 3049 15539 3115 15542
rect 4705 15539 4771 15542
rect 14549 15602 14615 15605
rect 18045 15602 18111 15605
rect 14549 15600 18111 15602
rect 14549 15544 14554 15600
rect 14610 15544 18050 15600
rect 18106 15544 18111 15600
rect 14549 15542 18111 15544
rect 14549 15539 14615 15542
rect 18045 15539 18111 15542
rect 8109 15466 8175 15469
rect 10041 15466 10107 15469
rect 8109 15464 10107 15466
rect 8109 15408 8114 15464
rect 8170 15408 10046 15464
rect 10102 15408 10107 15464
rect 8109 15406 10107 15408
rect 8109 15403 8175 15406
rect 10041 15403 10107 15406
rect 13721 15466 13787 15469
rect 14641 15466 14707 15469
rect 18965 15466 19031 15469
rect 13721 15464 19031 15466
rect 13721 15408 13726 15464
rect 13782 15408 14646 15464
rect 14702 15408 18970 15464
rect 19026 15408 19031 15464
rect 13721 15406 19031 15408
rect 13721 15403 13787 15406
rect 14641 15403 14707 15406
rect 18965 15403 19031 15406
rect 17309 15330 17375 15333
rect 20253 15330 20319 15333
rect 17309 15328 20319 15330
rect 17309 15272 17314 15328
rect 17370 15272 20258 15328
rect 20314 15272 20319 15328
rect 17309 15270 20319 15272
rect 17309 15267 17375 15270
rect 20253 15267 20319 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 3969 15058 4035 15061
rect 7281 15058 7347 15061
rect 3969 15056 7347 15058
rect 3969 15000 3974 15056
rect 4030 15000 7286 15056
rect 7342 15000 7347 15056
rect 3969 14998 7347 15000
rect 3969 14995 4035 14998
rect 7281 14995 7347 14998
rect 6361 14922 6427 14925
rect 10409 14922 10475 14925
rect 6361 14920 10475 14922
rect 6361 14864 6366 14920
rect 6422 14864 10414 14920
rect 10470 14864 10475 14920
rect 6361 14862 10475 14864
rect 6361 14859 6427 14862
rect 10409 14859 10475 14862
rect 0 14786 480 14816
rect 10041 14786 10107 14789
rect 0 14784 10107 14786
rect 0 14728 10046 14784
rect 10102 14728 10107 14784
rect 0 14726 10107 14728
rect 0 14696 480 14726
rect 10041 14723 10107 14726
rect 13261 14786 13327 14789
rect 19425 14786 19491 14789
rect 13261 14784 19491 14786
rect 13261 14728 13266 14784
rect 13322 14728 19430 14784
rect 19486 14728 19491 14784
rect 13261 14726 19491 14728
rect 13261 14723 13327 14726
rect 19425 14723 19491 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 17217 14514 17283 14517
rect 19333 14514 19399 14517
rect 17217 14512 19399 14514
rect 17217 14456 17222 14512
rect 17278 14456 19338 14512
rect 19394 14456 19399 14512
rect 17217 14454 19399 14456
rect 17217 14451 17283 14454
rect 19333 14451 19399 14454
rect 2957 14378 3023 14381
rect 9765 14378 9831 14381
rect 2957 14376 9831 14378
rect 2957 14320 2962 14376
rect 3018 14320 9770 14376
rect 9826 14320 9831 14376
rect 2957 14318 9831 14320
rect 2957 14315 3023 14318
rect 9765 14315 9831 14318
rect 13997 14378 14063 14381
rect 18045 14378 18111 14381
rect 13997 14376 18111 14378
rect 13997 14320 14002 14376
rect 14058 14320 18050 14376
rect 18106 14320 18111 14376
rect 13997 14318 18111 14320
rect 13997 14315 14063 14318
rect 18045 14315 18111 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 4705 13970 4771 13973
rect 9489 13970 9555 13973
rect 10593 13970 10659 13973
rect 4705 13968 10659 13970
rect 4705 13912 4710 13968
rect 4766 13912 9494 13968
rect 9550 13912 10598 13968
rect 10654 13912 10659 13968
rect 4705 13910 10659 13912
rect 4705 13907 4771 13910
rect 9489 13907 9555 13910
rect 10593 13907 10659 13910
rect 14181 13970 14247 13973
rect 19333 13970 19399 13973
rect 14181 13968 19399 13970
rect 14181 13912 14186 13968
rect 14242 13912 19338 13968
rect 19394 13912 19399 13968
rect 14181 13910 19399 13912
rect 14181 13907 14247 13910
rect 19333 13907 19399 13910
rect 23473 13970 23539 13973
rect 27520 13970 28000 14000
rect 23473 13968 28000 13970
rect 23473 13912 23478 13968
rect 23534 13912 28000 13968
rect 23473 13910 28000 13912
rect 23473 13907 23539 13910
rect 27520 13880 28000 13910
rect 2037 13834 2103 13837
rect 8385 13834 8451 13837
rect 2037 13832 8451 13834
rect 2037 13776 2042 13832
rect 2098 13776 8390 13832
rect 8446 13776 8451 13832
rect 2037 13774 8451 13776
rect 2037 13771 2103 13774
rect 8385 13771 8451 13774
rect 16297 13834 16363 13837
rect 18413 13834 18479 13837
rect 16297 13832 18479 13834
rect 16297 13776 16302 13832
rect 16358 13776 18418 13832
rect 18474 13776 18479 13832
rect 16297 13774 18479 13776
rect 16297 13771 16363 13774
rect 18413 13771 18479 13774
rect 4521 13698 4587 13701
rect 8477 13698 8543 13701
rect 4521 13696 8543 13698
rect 4521 13640 4526 13696
rect 4582 13640 8482 13696
rect 8538 13640 8543 13696
rect 4521 13638 8543 13640
rect 4521 13635 4587 13638
rect 8477 13635 8543 13638
rect 15745 13698 15811 13701
rect 19333 13698 19399 13701
rect 15745 13696 19399 13698
rect 15745 13640 15750 13696
rect 15806 13640 19338 13696
rect 19394 13640 19399 13696
rect 15745 13638 19399 13640
rect 15745 13635 15811 13638
rect 19333 13635 19399 13638
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 4337 13562 4403 13565
rect 5993 13562 6059 13565
rect 4337 13560 6059 13562
rect 4337 13504 4342 13560
rect 4398 13504 5998 13560
rect 6054 13504 6059 13560
rect 4337 13502 6059 13504
rect 4337 13499 4403 13502
rect 5993 13499 6059 13502
rect 16297 13562 16363 13565
rect 19241 13562 19307 13565
rect 16297 13560 19307 13562
rect 16297 13504 16302 13560
rect 16358 13504 19246 13560
rect 19302 13504 19307 13560
rect 16297 13502 19307 13504
rect 16297 13499 16363 13502
rect 19241 13499 19307 13502
rect 9213 13426 9279 13429
rect 19793 13426 19859 13429
rect 9213 13424 19859 13426
rect 9213 13368 9218 13424
rect 9274 13368 19798 13424
rect 19854 13368 19859 13424
rect 9213 13366 19859 13368
rect 9213 13363 9279 13366
rect 19793 13363 19859 13366
rect 0 13290 480 13320
rect 1577 13290 1643 13293
rect 0 13288 1643 13290
rect 0 13232 1582 13288
rect 1638 13232 1643 13288
rect 0 13230 1643 13232
rect 0 13200 480 13230
rect 1577 13227 1643 13230
rect 4889 13290 4955 13293
rect 11421 13290 11487 13293
rect 4889 13288 11487 13290
rect 4889 13232 4894 13288
rect 4950 13232 11426 13288
rect 11482 13232 11487 13288
rect 4889 13230 11487 13232
rect 4889 13227 4955 13230
rect 11421 13227 11487 13230
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 8753 13018 8819 13021
rect 11513 13018 11579 13021
rect 14181 13018 14247 13021
rect 8753 13016 14247 13018
rect 8753 12960 8758 13016
rect 8814 12960 11518 13016
rect 11574 12960 14186 13016
rect 14242 12960 14247 13016
rect 8753 12958 14247 12960
rect 8753 12955 8819 12958
rect 11513 12955 11579 12958
rect 14181 12955 14247 12958
rect 7925 12882 7991 12885
rect 19793 12882 19859 12885
rect 7925 12880 19859 12882
rect 7925 12824 7930 12880
rect 7986 12824 19798 12880
rect 19854 12824 19859 12880
rect 7925 12822 19859 12824
rect 7925 12819 7991 12822
rect 19793 12819 19859 12822
rect 3509 12746 3575 12749
rect 5993 12746 6059 12749
rect 3509 12744 6059 12746
rect 3509 12688 3514 12744
rect 3570 12688 5998 12744
rect 6054 12688 6059 12744
rect 3509 12686 6059 12688
rect 3509 12683 3575 12686
rect 5993 12683 6059 12686
rect 6269 12746 6335 12749
rect 11053 12746 11119 12749
rect 6269 12744 11119 12746
rect 6269 12688 6274 12744
rect 6330 12688 11058 12744
rect 11114 12688 11119 12744
rect 6269 12686 11119 12688
rect 6269 12683 6335 12686
rect 11053 12683 11119 12686
rect 11697 12746 11763 12749
rect 23565 12746 23631 12749
rect 11697 12744 23631 12746
rect 11697 12688 11702 12744
rect 11758 12688 23570 12744
rect 23626 12688 23631 12744
rect 11697 12686 23631 12688
rect 11697 12683 11763 12686
rect 23565 12683 23631 12686
rect 13997 12610 14063 12613
rect 14365 12610 14431 12613
rect 19333 12610 19399 12613
rect 13997 12608 19399 12610
rect 13997 12552 14002 12608
rect 14058 12552 14370 12608
rect 14426 12552 19338 12608
rect 19394 12552 19399 12608
rect 13997 12550 19399 12552
rect 13997 12547 14063 12550
rect 14365 12547 14431 12550
rect 19333 12547 19399 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 4705 12338 4771 12341
rect 10317 12338 10383 12341
rect 4705 12336 10383 12338
rect 4705 12280 4710 12336
rect 4766 12280 10322 12336
rect 10378 12280 10383 12336
rect 4705 12278 10383 12280
rect 4705 12275 4771 12278
rect 10317 12275 10383 12278
rect 14273 12338 14339 12341
rect 16205 12338 16271 12341
rect 23473 12338 23539 12341
rect 14273 12336 16271 12338
rect 14273 12280 14278 12336
rect 14334 12280 16210 12336
rect 16266 12280 16271 12336
rect 14273 12278 16271 12280
rect 14273 12275 14339 12278
rect 16205 12275 16271 12278
rect 16438 12336 23539 12338
rect 16438 12280 23478 12336
rect 23534 12280 23539 12336
rect 16438 12278 23539 12280
rect 1945 12202 2011 12205
rect 4889 12202 4955 12205
rect 1945 12200 4955 12202
rect 1945 12144 1950 12200
rect 2006 12144 4894 12200
rect 4950 12144 4955 12200
rect 1945 12142 4955 12144
rect 1945 12139 2011 12142
rect 4889 12139 4955 12142
rect 15285 12202 15351 12205
rect 16438 12202 16498 12278
rect 23473 12275 23539 12278
rect 15285 12200 16498 12202
rect 15285 12144 15290 12200
rect 15346 12144 16498 12200
rect 15285 12142 16498 12144
rect 16757 12202 16823 12205
rect 19333 12202 19399 12205
rect 16757 12200 19399 12202
rect 16757 12144 16762 12200
rect 16818 12144 19338 12200
rect 19394 12144 19399 12200
rect 16757 12142 19399 12144
rect 15285 12139 15351 12142
rect 16757 12139 16823 12142
rect 19333 12139 19399 12142
rect 6269 12066 6335 12069
rect 7373 12066 7439 12069
rect 14273 12066 14339 12069
rect 6269 12064 14339 12066
rect 6269 12008 6274 12064
rect 6330 12008 7378 12064
rect 7434 12008 14278 12064
rect 14334 12008 14339 12064
rect 6269 12006 14339 12008
rect 6269 12003 6335 12006
rect 7373 12003 7439 12006
rect 14273 12003 14339 12006
rect 5610 12000 5930 12001
rect 0 11930 480 11960
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 1577 11930 1643 11933
rect 0 11928 1643 11930
rect 0 11872 1582 11928
rect 1638 11872 1643 11928
rect 0 11870 1643 11872
rect 0 11840 480 11870
rect 1577 11867 1643 11870
rect 7649 11930 7715 11933
rect 12157 11930 12223 11933
rect 7649 11928 12223 11930
rect 7649 11872 7654 11928
rect 7710 11872 12162 11928
rect 12218 11872 12223 11928
rect 7649 11870 12223 11872
rect 7649 11867 7715 11870
rect 12157 11867 12223 11870
rect 15745 11930 15811 11933
rect 19793 11930 19859 11933
rect 15745 11928 19859 11930
rect 15745 11872 15750 11928
rect 15806 11872 19798 11928
rect 19854 11872 19859 11928
rect 15745 11870 19859 11872
rect 15745 11867 15811 11870
rect 19793 11867 19859 11870
rect 10961 11794 11027 11797
rect 24117 11794 24183 11797
rect 10961 11792 24183 11794
rect 10961 11736 10966 11792
rect 11022 11736 24122 11792
rect 24178 11736 24183 11792
rect 10961 11734 24183 11736
rect 10961 11731 11027 11734
rect 24117 11731 24183 11734
rect 9489 11658 9555 11661
rect 13629 11658 13695 11661
rect 9489 11656 13695 11658
rect 9489 11600 9494 11656
rect 9550 11600 13634 11656
rect 13690 11600 13695 11656
rect 9489 11598 13695 11600
rect 9489 11595 9555 11598
rect 13629 11595 13695 11598
rect 14365 11658 14431 11661
rect 19609 11658 19675 11661
rect 14365 11656 19675 11658
rect 14365 11600 14370 11656
rect 14426 11600 19614 11656
rect 19670 11600 19675 11656
rect 14365 11598 19675 11600
rect 14365 11595 14431 11598
rect 19609 11595 19675 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 3509 11386 3575 11389
rect 5165 11386 5231 11389
rect 3509 11384 5231 11386
rect 3509 11328 3514 11384
rect 3570 11328 5170 11384
rect 5226 11328 5231 11384
rect 3509 11326 5231 11328
rect 3509 11323 3575 11326
rect 5165 11323 5231 11326
rect 5441 11386 5507 11389
rect 6453 11386 6519 11389
rect 5441 11384 6519 11386
rect 5441 11328 5446 11384
rect 5502 11328 6458 11384
rect 6514 11328 6519 11384
rect 5441 11326 6519 11328
rect 5441 11323 5507 11326
rect 6453 11323 6519 11326
rect 14089 11386 14155 11389
rect 15745 11386 15811 11389
rect 14089 11384 15811 11386
rect 14089 11328 14094 11384
rect 14150 11328 15750 11384
rect 15806 11328 15811 11384
rect 14089 11326 15811 11328
rect 14089 11323 14155 11326
rect 15745 11323 15811 11326
rect 6269 11250 6335 11253
rect 10961 11252 11027 11253
rect 10910 11250 10916 11252
rect 6269 11248 10916 11250
rect 10980 11250 11027 11252
rect 15469 11250 15535 11253
rect 18045 11250 18111 11253
rect 10980 11248 11072 11250
rect 6269 11192 6274 11248
rect 6330 11192 10916 11248
rect 11022 11192 11072 11248
rect 6269 11190 10916 11192
rect 6269 11187 6335 11190
rect 10910 11188 10916 11190
rect 10980 11190 11072 11192
rect 15469 11248 18111 11250
rect 15469 11192 15474 11248
rect 15530 11192 18050 11248
rect 18106 11192 18111 11248
rect 15469 11190 18111 11192
rect 10980 11188 11027 11190
rect 10961 11187 11027 11188
rect 15469 11187 15535 11190
rect 18045 11187 18111 11190
rect 3417 11114 3483 11117
rect 5901 11114 5967 11117
rect 3417 11112 5967 11114
rect 3417 11056 3422 11112
rect 3478 11056 5906 11112
rect 5962 11056 5967 11112
rect 3417 11054 5967 11056
rect 3417 11051 3483 11054
rect 5901 11051 5967 11054
rect 14733 11114 14799 11117
rect 16941 11114 17007 11117
rect 19333 11114 19399 11117
rect 14733 11112 19399 11114
rect 14733 11056 14738 11112
rect 14794 11056 16946 11112
rect 17002 11056 19338 11112
rect 19394 11056 19399 11112
rect 14733 11054 19399 11056
rect 14733 11051 14799 11054
rect 16941 11051 17007 11054
rect 19333 11051 19399 11054
rect 8201 10978 8267 10981
rect 10777 10978 10843 10981
rect 8201 10976 10843 10978
rect 8201 10920 8206 10976
rect 8262 10920 10782 10976
rect 10838 10920 10843 10976
rect 8201 10918 10843 10920
rect 8201 10915 8267 10918
rect 10777 10915 10843 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 6637 10842 6703 10845
rect 12893 10842 12959 10845
rect 27520 10842 28000 10872
rect 6637 10840 12959 10842
rect 6637 10784 6642 10840
rect 6698 10784 12898 10840
rect 12954 10784 12959 10840
rect 6637 10782 12959 10784
rect 6637 10779 6703 10782
rect 12893 10779 12959 10782
rect 24718 10782 28000 10842
rect 4061 10706 4127 10709
rect 4981 10706 5047 10709
rect 7097 10706 7163 10709
rect 4061 10704 7163 10706
rect 4061 10648 4066 10704
rect 4122 10648 4986 10704
rect 5042 10648 7102 10704
rect 7158 10648 7163 10704
rect 4061 10646 7163 10648
rect 4061 10643 4127 10646
rect 4981 10643 5047 10646
rect 7097 10643 7163 10646
rect 8661 10706 8727 10709
rect 18045 10706 18111 10709
rect 18413 10706 18479 10709
rect 24718 10706 24778 10782
rect 27520 10752 28000 10782
rect 8661 10704 18111 10706
rect 8661 10648 8666 10704
rect 8722 10648 18050 10704
rect 18106 10648 18111 10704
rect 8661 10646 18111 10648
rect 8661 10643 8727 10646
rect 18045 10643 18111 10646
rect 18232 10704 24778 10706
rect 18232 10648 18418 10704
rect 18474 10648 24778 10704
rect 18232 10646 24778 10648
rect 0 10570 480 10600
rect 1393 10570 1459 10573
rect 0 10568 1459 10570
rect 0 10512 1398 10568
rect 1454 10512 1459 10568
rect 0 10510 1459 10512
rect 0 10480 480 10510
rect 1393 10507 1459 10510
rect 8845 10570 8911 10573
rect 11053 10570 11119 10573
rect 8845 10568 11119 10570
rect 8845 10512 8850 10568
rect 8906 10512 11058 10568
rect 11114 10512 11119 10568
rect 8845 10510 11119 10512
rect 8845 10507 8911 10510
rect 11053 10507 11119 10510
rect 17401 10570 17467 10573
rect 18232 10570 18292 10646
rect 18413 10643 18479 10646
rect 17401 10568 18292 10570
rect 17401 10512 17406 10568
rect 17462 10512 18292 10568
rect 17401 10510 18292 10512
rect 17401 10507 17467 10510
rect 15009 10434 15075 10437
rect 18597 10434 18663 10437
rect 15009 10432 18663 10434
rect 15009 10376 15014 10432
rect 15070 10376 18602 10432
rect 18658 10376 18663 10432
rect 15009 10374 18663 10376
rect 15009 10371 15075 10374
rect 18597 10371 18663 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 14273 10298 14339 10301
rect 14641 10298 14707 10301
rect 19333 10298 19399 10301
rect 14273 10296 19399 10298
rect 14273 10240 14278 10296
rect 14334 10240 14646 10296
rect 14702 10240 19338 10296
rect 19394 10240 19399 10296
rect 14273 10238 19399 10240
rect 14273 10235 14339 10238
rect 14641 10235 14707 10238
rect 19333 10235 19399 10238
rect 2129 10162 2195 10165
rect 6085 10162 6151 10165
rect 2129 10160 6151 10162
rect 2129 10104 2134 10160
rect 2190 10104 6090 10160
rect 6146 10104 6151 10160
rect 2129 10102 6151 10104
rect 2129 10099 2195 10102
rect 6085 10099 6151 10102
rect 16021 10162 16087 10165
rect 19425 10162 19491 10165
rect 16021 10160 19491 10162
rect 16021 10104 16026 10160
rect 16082 10104 19430 10160
rect 19486 10104 19491 10160
rect 16021 10102 19491 10104
rect 16021 10099 16087 10102
rect 19425 10099 19491 10102
rect 16757 10026 16823 10029
rect 19609 10026 19675 10029
rect 16757 10024 19675 10026
rect 16757 9968 16762 10024
rect 16818 9968 19614 10024
rect 19670 9968 19675 10024
rect 16757 9966 19675 9968
rect 16757 9963 16823 9966
rect 19609 9963 19675 9966
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 1669 9618 1735 9621
rect 4245 9618 4311 9621
rect 10133 9618 10199 9621
rect 1669 9616 10199 9618
rect 1669 9560 1674 9616
rect 1730 9560 4250 9616
rect 4306 9560 10138 9616
rect 10194 9560 10199 9616
rect 1669 9558 10199 9560
rect 1669 9555 1735 9558
rect 4245 9555 4311 9558
rect 10133 9555 10199 9558
rect 7189 9482 7255 9485
rect 12525 9482 12591 9485
rect 7189 9480 12591 9482
rect 7189 9424 7194 9480
rect 7250 9424 12530 9480
rect 12586 9424 12591 9480
rect 7189 9422 12591 9424
rect 7189 9419 7255 9422
rect 12525 9419 12591 9422
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 3233 9210 3299 9213
rect 5993 9210 6059 9213
rect 3233 9208 6059 9210
rect 3233 9152 3238 9208
rect 3294 9152 5998 9208
rect 6054 9152 6059 9208
rect 3233 9150 6059 9152
rect 3233 9147 3299 9150
rect 5993 9147 6059 9150
rect 10961 9210 11027 9213
rect 16113 9210 16179 9213
rect 10961 9208 16179 9210
rect 10961 9152 10966 9208
rect 11022 9152 16118 9208
rect 16174 9152 16179 9208
rect 10961 9150 16179 9152
rect 10961 9147 11027 9150
rect 16113 9147 16179 9150
rect 0 9074 480 9104
rect 1577 9074 1643 9077
rect 0 9072 1643 9074
rect 0 9016 1582 9072
rect 1638 9016 1643 9072
rect 0 9014 1643 9016
rect 0 8984 480 9014
rect 1577 9011 1643 9014
rect 14181 9074 14247 9077
rect 18137 9074 18203 9077
rect 14181 9072 18203 9074
rect 14181 9016 14186 9072
rect 14242 9016 18142 9072
rect 18198 9016 18203 9072
rect 14181 9014 18203 9016
rect 14181 9011 14247 9014
rect 18137 9011 18203 9014
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 10593 8530 10659 8533
rect 13997 8530 14063 8533
rect 10593 8528 14063 8530
rect 10593 8472 10598 8528
rect 10654 8472 14002 8528
rect 14058 8472 14063 8528
rect 10593 8470 14063 8472
rect 10593 8467 10659 8470
rect 13997 8467 14063 8470
rect 14273 8530 14339 8533
rect 16389 8530 16455 8533
rect 19793 8530 19859 8533
rect 14273 8528 19859 8530
rect 14273 8472 14278 8528
rect 14334 8472 16394 8528
rect 16450 8472 19798 8528
rect 19854 8472 19859 8528
rect 14273 8470 19859 8472
rect 14273 8467 14339 8470
rect 16389 8467 16455 8470
rect 19793 8467 19859 8470
rect 10869 8394 10935 8397
rect 20069 8394 20135 8397
rect 10869 8392 20135 8394
rect 10869 8336 10874 8392
rect 10930 8336 20074 8392
rect 20130 8336 20135 8392
rect 10869 8334 20135 8336
rect 10869 8331 10935 8334
rect 20069 8331 20135 8334
rect 11145 8258 11211 8261
rect 15929 8258 15995 8261
rect 19057 8258 19123 8261
rect 11145 8256 19123 8258
rect 11145 8200 11150 8256
rect 11206 8200 15934 8256
rect 15990 8200 19062 8256
rect 19118 8200 19123 8256
rect 11145 8198 19123 8200
rect 11145 8195 11211 8198
rect 15929 8195 15995 8198
rect 19057 8195 19123 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 14825 7986 14891 7989
rect 16573 7986 16639 7989
rect 14825 7984 16639 7986
rect 14825 7928 14830 7984
rect 14886 7928 16578 7984
rect 16634 7928 16639 7984
rect 14825 7926 16639 7928
rect 14825 7923 14891 7926
rect 16573 7923 16639 7926
rect 18965 7986 19031 7989
rect 18965 7984 24778 7986
rect 18965 7928 18970 7984
rect 19026 7928 24778 7984
rect 18965 7926 24778 7928
rect 18965 7923 19031 7926
rect 0 7714 480 7744
rect 1577 7714 1643 7717
rect 0 7712 1643 7714
rect 0 7656 1582 7712
rect 1638 7656 1643 7712
rect 0 7654 1643 7656
rect 24718 7714 24778 7926
rect 27520 7714 28000 7744
rect 24718 7654 28000 7714
rect 0 7624 480 7654
rect 1577 7651 1643 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 27520 7624 28000 7654
rect 24277 7583 24597 7584
rect 14733 7170 14799 7173
rect 19425 7170 19491 7173
rect 14733 7168 19491 7170
rect 14733 7112 14738 7168
rect 14794 7112 19430 7168
rect 19486 7112 19491 7168
rect 14733 7110 19491 7112
rect 14733 7107 14799 7110
rect 19425 7107 19491 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 17585 7034 17651 7037
rect 19333 7034 19399 7037
rect 17585 7032 19399 7034
rect 17585 6976 17590 7032
rect 17646 6976 19338 7032
rect 19394 6976 19399 7032
rect 17585 6974 19399 6976
rect 17585 6971 17651 6974
rect 19333 6971 19399 6974
rect 2405 6898 2471 6901
rect 2957 6898 3023 6901
rect 2405 6896 3023 6898
rect 2405 6840 2410 6896
rect 2466 6840 2962 6896
rect 3018 6840 3023 6896
rect 2405 6838 3023 6840
rect 2405 6835 2471 6838
rect 2957 6835 3023 6838
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 0 6354 480 6384
rect 1577 6354 1643 6357
rect 0 6352 1643 6354
rect 0 6296 1582 6352
rect 1638 6296 1643 6352
rect 0 6294 1643 6296
rect 0 6264 480 6294
rect 1577 6291 1643 6294
rect 6545 6354 6611 6357
rect 14825 6354 14891 6357
rect 6545 6352 14891 6354
rect 6545 6296 6550 6352
rect 6606 6296 14830 6352
rect 14886 6296 14891 6352
rect 6545 6294 14891 6296
rect 6545 6291 6611 6294
rect 14825 6291 14891 6294
rect 9949 6218 10015 6221
rect 12801 6218 12867 6221
rect 9949 6216 12867 6218
rect 9949 6160 9954 6216
rect 10010 6160 12806 6216
rect 12862 6160 12867 6216
rect 9949 6158 12867 6160
rect 9949 6155 10015 6158
rect 12801 6155 12867 6158
rect 15745 6218 15811 6221
rect 19609 6218 19675 6221
rect 15745 6216 19675 6218
rect 15745 6160 15750 6216
rect 15806 6160 19614 6216
rect 19670 6160 19675 6216
rect 15745 6158 19675 6160
rect 15745 6155 15811 6158
rect 19609 6155 19675 6158
rect 1669 6082 1735 6085
rect 9305 6082 9371 6085
rect 1669 6080 9371 6082
rect 1669 6024 1674 6080
rect 1730 6024 9310 6080
rect 9366 6024 9371 6080
rect 1669 6022 9371 6024
rect 1669 6019 1735 6022
rect 9305 6019 9371 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 12433 5810 12499 5813
rect 15377 5810 15443 5813
rect 12433 5808 15443 5810
rect 12433 5752 12438 5808
rect 12494 5752 15382 5808
rect 15438 5752 15443 5808
rect 12433 5750 15443 5752
rect 12433 5747 12499 5750
rect 15377 5747 15443 5750
rect 18137 5810 18203 5813
rect 20713 5810 20779 5813
rect 18137 5808 20779 5810
rect 18137 5752 18142 5808
rect 18198 5752 20718 5808
rect 20774 5752 20779 5808
rect 18137 5750 20779 5752
rect 18137 5747 18203 5750
rect 20713 5747 20779 5750
rect 7373 5674 7439 5677
rect 11237 5674 11303 5677
rect 7373 5672 11303 5674
rect 7373 5616 7378 5672
rect 7434 5616 11242 5672
rect 11298 5616 11303 5672
rect 7373 5614 11303 5616
rect 7373 5611 7439 5614
rect 11237 5611 11303 5614
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 11053 5130 11119 5133
rect 12709 5130 12775 5133
rect 11053 5128 12775 5130
rect 11053 5072 11058 5128
rect 11114 5072 12714 5128
rect 12770 5072 12775 5128
rect 11053 5070 12775 5072
rect 11053 5067 11119 5070
rect 12709 5067 12775 5070
rect 2037 4994 2103 4997
rect 6821 4994 6887 4997
rect 2037 4992 6887 4994
rect 2037 4936 2042 4992
rect 2098 4936 6826 4992
rect 6882 4936 6887 4992
rect 2037 4934 6887 4936
rect 2037 4931 2103 4934
rect 6821 4931 6887 4934
rect 13629 4994 13695 4997
rect 15285 4994 15351 4997
rect 13629 4992 15351 4994
rect 13629 4936 13634 4992
rect 13690 4936 15290 4992
rect 15346 4936 15351 4992
rect 13629 4934 15351 4936
rect 13629 4931 13695 4934
rect 15285 4931 15351 4934
rect 10277 4928 10597 4929
rect 0 4858 480 4888
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 1577 4858 1643 4861
rect 0 4856 1643 4858
rect 0 4800 1582 4856
rect 1638 4800 1643 4856
rect 0 4798 1643 4800
rect 0 4768 480 4798
rect 1577 4795 1643 4798
rect 17401 4858 17467 4861
rect 18413 4858 18479 4861
rect 17401 4856 18479 4858
rect 17401 4800 17406 4856
rect 17462 4800 18418 4856
rect 18474 4800 18479 4856
rect 17401 4798 18479 4800
rect 17401 4795 17467 4798
rect 18413 4795 18479 4798
rect 27520 4586 28000 4616
rect 27478 4496 28000 4586
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 1761 4178 1827 4181
rect 10041 4178 10107 4181
rect 13905 4178 13971 4181
rect 1761 4176 13971 4178
rect 1761 4120 1766 4176
rect 1822 4120 10046 4176
rect 10102 4120 13910 4176
rect 13966 4120 13971 4176
rect 1761 4118 13971 4120
rect 1761 4115 1827 4118
rect 10041 4115 10107 4118
rect 13905 4115 13971 4118
rect 15469 4178 15535 4181
rect 27478 4178 27538 4496
rect 15469 4176 27538 4178
rect 15469 4120 15474 4176
rect 15530 4120 27538 4176
rect 15469 4118 27538 4120
rect 15469 4115 15535 4118
rect 1945 4042 2011 4045
rect 5533 4042 5599 4045
rect 1945 4040 5599 4042
rect 1945 3984 1950 4040
rect 2006 3984 5538 4040
rect 5594 3984 5599 4040
rect 1945 3982 5599 3984
rect 1945 3979 2011 3982
rect 5533 3979 5599 3982
rect 6729 4042 6795 4045
rect 11329 4042 11395 4045
rect 6729 4040 11395 4042
rect 6729 3984 6734 4040
rect 6790 3984 11334 4040
rect 11390 3984 11395 4040
rect 6729 3982 11395 3984
rect 6729 3979 6795 3982
rect 11329 3979 11395 3982
rect 6637 3906 6703 3909
rect 9673 3906 9739 3909
rect 6637 3904 9739 3906
rect 6637 3848 6642 3904
rect 6698 3848 9678 3904
rect 9734 3848 9739 3904
rect 6637 3846 9739 3848
rect 6637 3843 6703 3846
rect 9673 3843 9739 3846
rect 10777 3906 10843 3909
rect 16205 3906 16271 3909
rect 10777 3904 16271 3906
rect 10777 3848 10782 3904
rect 10838 3848 16210 3904
rect 16266 3848 16271 3904
rect 10777 3846 16271 3848
rect 10777 3843 10843 3846
rect 16205 3843 16271 3846
rect 21357 3906 21423 3909
rect 23197 3906 23263 3909
rect 21357 3904 23263 3906
rect 21357 3848 21362 3904
rect 21418 3848 23202 3904
rect 23258 3848 23263 3904
rect 21357 3846 23263 3848
rect 21357 3843 21423 3846
rect 23197 3843 23263 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 3509 3770 3575 3773
rect 9857 3770 9923 3773
rect 3509 3768 9923 3770
rect 3509 3712 3514 3768
rect 3570 3712 9862 3768
rect 9918 3712 9923 3768
rect 3509 3710 9923 3712
rect 3509 3707 3575 3710
rect 9857 3707 9923 3710
rect 11237 3634 11303 3637
rect 12157 3634 12223 3637
rect 16021 3634 16087 3637
rect 11237 3632 16087 3634
rect 11237 3576 11242 3632
rect 11298 3576 12162 3632
rect 12218 3576 16026 3632
rect 16082 3576 16087 3632
rect 11237 3574 16087 3576
rect 11237 3571 11303 3574
rect 12157 3571 12223 3574
rect 16021 3571 16087 3574
rect 19333 3634 19399 3637
rect 26325 3634 26391 3637
rect 19333 3632 26391 3634
rect 19333 3576 19338 3632
rect 19394 3576 26330 3632
rect 26386 3576 26391 3632
rect 19333 3574 26391 3576
rect 19333 3571 19399 3574
rect 26325 3571 26391 3574
rect 0 3498 480 3528
rect 1577 3498 1643 3501
rect 0 3496 1643 3498
rect 0 3440 1582 3496
rect 1638 3440 1643 3496
rect 0 3438 1643 3440
rect 0 3408 480 3438
rect 1577 3435 1643 3438
rect 2405 3498 2471 3501
rect 5073 3498 5139 3501
rect 25313 3498 25379 3501
rect 2405 3496 5139 3498
rect 2405 3440 2410 3496
rect 2466 3440 5078 3496
rect 5134 3440 5139 3496
rect 2405 3438 5139 3440
rect 2405 3435 2471 3438
rect 5073 3435 5139 3438
rect 15334 3496 25379 3498
rect 15334 3440 25318 3496
rect 25374 3440 25379 3496
rect 15334 3438 25379 3440
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 7373 3226 7439 3229
rect 12065 3226 12131 3229
rect 7373 3224 12131 3226
rect 7373 3168 7378 3224
rect 7434 3168 12070 3224
rect 12126 3168 12131 3224
rect 7373 3166 12131 3168
rect 7373 3163 7439 3166
rect 12065 3163 12131 3166
rect 473 3090 539 3093
rect 9949 3090 10015 3093
rect 473 3088 10015 3090
rect 473 3032 478 3088
rect 534 3032 9954 3088
rect 10010 3032 10015 3088
rect 473 3030 10015 3032
rect 473 3027 539 3030
rect 9949 3027 10015 3030
rect 11881 3090 11947 3093
rect 15334 3090 15394 3438
rect 25313 3435 25379 3438
rect 18873 3362 18939 3365
rect 20069 3362 20135 3365
rect 18873 3360 20135 3362
rect 18873 3304 18878 3360
rect 18934 3304 20074 3360
rect 20130 3304 20135 3360
rect 18873 3302 20135 3304
rect 18873 3299 18939 3302
rect 20069 3299 20135 3302
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 15653 3226 15719 3229
rect 22185 3226 22251 3229
rect 15653 3224 22251 3226
rect 15653 3168 15658 3224
rect 15714 3168 22190 3224
rect 22246 3168 22251 3224
rect 15653 3166 22251 3168
rect 15653 3163 15719 3166
rect 22185 3163 22251 3166
rect 11881 3088 15394 3090
rect 11881 3032 11886 3088
rect 11942 3032 15394 3088
rect 11881 3030 15394 3032
rect 11881 3027 11947 3030
rect 8937 2954 9003 2957
rect 14273 2954 14339 2957
rect 8937 2952 14339 2954
rect 8937 2896 8942 2952
rect 8998 2896 14278 2952
rect 14334 2896 14339 2952
rect 8937 2894 14339 2896
rect 8937 2891 9003 2894
rect 14273 2891 14339 2894
rect 19057 2954 19123 2957
rect 24209 2954 24275 2957
rect 19057 2952 24275 2954
rect 19057 2896 19062 2952
rect 19118 2896 24214 2952
rect 24270 2896 24275 2952
rect 19057 2894 24275 2896
rect 19057 2891 19123 2894
rect 24209 2891 24275 2894
rect 2497 2818 2563 2821
rect 7373 2818 7439 2821
rect 2497 2816 7439 2818
rect 2497 2760 2502 2816
rect 2558 2760 7378 2816
rect 7434 2760 7439 2816
rect 2497 2758 7439 2760
rect 2497 2755 2563 2758
rect 7373 2755 7439 2758
rect 14457 2818 14523 2821
rect 17033 2818 17099 2821
rect 14457 2816 17099 2818
rect 14457 2760 14462 2816
rect 14518 2760 17038 2816
rect 17094 2760 17099 2816
rect 14457 2758 17099 2760
rect 14457 2755 14523 2758
rect 17033 2755 17099 2758
rect 17861 2818 17927 2821
rect 19057 2818 19123 2821
rect 17861 2816 19123 2818
rect 17861 2760 17866 2816
rect 17922 2760 19062 2816
rect 19118 2760 19123 2816
rect 17861 2758 19123 2760
rect 17861 2755 17927 2758
rect 19057 2755 19123 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 2681 2682 2747 2685
rect 4337 2682 4403 2685
rect 2681 2680 4403 2682
rect 2681 2624 2686 2680
rect 2742 2624 4342 2680
rect 4398 2624 4403 2680
rect 2681 2622 4403 2624
rect 2681 2619 2747 2622
rect 4337 2619 4403 2622
rect 18229 2546 18295 2549
rect 24669 2546 24735 2549
rect 18229 2544 24735 2546
rect 18229 2488 18234 2544
rect 18290 2488 24674 2544
rect 24730 2488 24735 2544
rect 18229 2486 24735 2488
rect 18229 2483 18295 2486
rect 24669 2483 24735 2486
rect 1945 2274 2011 2277
rect 4613 2274 4679 2277
rect 1945 2272 4679 2274
rect 1945 2216 1950 2272
rect 2006 2216 4618 2272
rect 4674 2216 4679 2272
rect 1945 2214 4679 2216
rect 1945 2211 2011 2214
rect 4613 2211 4679 2214
rect 25129 2274 25195 2277
rect 27337 2274 27403 2277
rect 25129 2272 27403 2274
rect 25129 2216 25134 2272
rect 25190 2216 27342 2272
rect 27398 2216 27403 2272
rect 25129 2214 27403 2216
rect 25129 2211 25195 2214
rect 27337 2211 27403 2214
rect 5610 2208 5930 2209
rect 0 2138 480 2168
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 1577 2138 1643 2141
rect 0 2136 1643 2138
rect 0 2080 1582 2136
rect 1638 2080 1643 2136
rect 0 2078 1643 2080
rect 0 2048 480 2078
rect 1577 2075 1643 2078
rect 12985 1594 13051 1597
rect 27520 1594 28000 1624
rect 12985 1592 28000 1594
rect 12985 1536 12990 1592
rect 13046 1536 28000 1592
rect 12985 1534 28000 1536
rect 12985 1531 13051 1534
rect 27520 1504 28000 1534
rect 0 778 480 808
rect 4061 778 4127 781
rect 0 776 4127 778
rect 0 720 4066 776
rect 4122 720 4127 776
rect 0 718 4127 720
rect 0 688 480 718
rect 4061 715 4127 718
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 23980 23292 24044 23356
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 10916 11248 10980 11252
rect 10916 11192 10966 11248
rect 10966 11192 10980 11248
rect 10916 11188 10980 11192
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 23979 23356 24045 23357
rect 23979 23292 23980 23356
rect 24044 23292 24045 23356
rect 23979 23291 24045 23292
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 23982 11338 24042 23291
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 10830 11252 11066 11338
rect 10830 11188 10916 11252
rect 10916 11188 10980 11252
rect 10980 11188 11066 11252
rect 10830 11102 11066 11188
rect 23894 11102 24130 11338
<< metal5 >>
rect 10788 11338 24172 11380
rect 10788 11102 10830 11338
rect 11066 11102 23894 11338
rect 24130 11102 24172 11338
rect 10788 11060 24172 11102
use scs8hd_decap_4  FILLER_1_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_6 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_2  _230_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_13
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__192__A
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2668 0 1 2720
box -38 -48 866 592
use scs8hd_inv_8  _192_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_conb_1  _215_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_23 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_35
timestamp 1586364061
transform 1 0 4324 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_26
timestamp 1586364061
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_30
timestamp 1586364061
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_43
timestamp 1586364061
transform 1 0 5060 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_39
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_1_51
timestamp 1586364061
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_47
timestamp 1586364061
transform 1 0 5428 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_46
timestamp 1586364061
transform 1 0 5336 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5612 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5244 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5520 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_50 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5704 0 -1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_69
timestamp 1586364061
transform 1 0 7452 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_65
timestamp 1586364061
transform 1 0 7084 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_66
timestamp 1586364061
transform 1 0 7176 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7360 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_5.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_0_70
timestamp 1586364061
transform 1 0 7544 0 -1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_5.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_82
timestamp 1586364061
transform 1 0 8648 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_76
timestamp 1586364061
transform 1 0 8096 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_80
timestamp 1586364061
transform 1 0 8464 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_84
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _238_
timestamp 1586364061
transform 1 0 10580 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9936 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_90
timestamp 1586364061
transform 1 0 9384 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_0_94
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_1  FILLER_0_102 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_107
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_1_98
timestamp 1586364061
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_114
timestamp 1586364061
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_110
timestamp 1586364061
transform 1 0 11224 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__238__A
timestamp 1586364061
transform 1 0 11132 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_118
timestamp 1586364061
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_123
timestamp 1586364061
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _236_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_0_111
timestamp 1586364061
transform 1 0 11316 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_1_131
timestamp 1586364061
transform 1 0 13156 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_127
timestamp 1586364061
transform 1 0 12788 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_133
timestamp 1586364061
transform 1 0 13340 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_129
timestamp 1586364061
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13340 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__236__A
timestamp 1586364061
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__237__A
timestamp 1586364061
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _237_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_135
timestamp 1586364061
transform 1 0 13524 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_141
timestamp 1586364061
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13708 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _234_
timestamp 1586364061
transform 1 0 13892 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_143
timestamp 1586364061
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_147
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__235__A
timestamp 1586364061
transform 1 0 14812 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__233__A
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__234__A
timestamp 1586364061
transform 1 0 14444 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _233_
timestamp 1586364061
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_155
timestamp 1586364061
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_156 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_4  FILLER_0_151
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _235_
timestamp 1586364061
transform 1 0 14996 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_159
timestamp 1586364061
transform 1 0 15732 0 1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15548 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_167
timestamp 1586364061
transform 1 0 16468 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_163
timestamp 1586364061
transform 1 0 16100 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_166
timestamp 1586364061
transform 1 0 16376 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__231__A
timestamp 1586364061
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__232__A
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16192 0 1 2720
box -38 -48 314 592
use scs8hd_buf_2  _232_
timestamp 1586364061
transform 1 0 16008 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_170
timestamp 1586364061
transform 1 0 16744 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_187
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_0_182
timestamp 1586364061
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_192
timestamp 1586364061
transform 1 0 18768 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_188
timestamp 1586364061
transform 1 0 18400 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_195
timestamp 1586364061
transform 1 0 19044 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_191
timestamp 1586364061
transform 1 0 18676 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18952 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18492 0 1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18768 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_12  FILLER_1_196
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19228 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_199
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_0_211
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_208
timestamp 1586364061
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_0_218
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_230
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_220
timestamp 1586364061
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_242
timestamp 1586364061
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_6  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_12  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_258
timestamp 1586364061
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_262
timestamp 1586364061
transform 1 0 25208 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_0_274
timestamp 1586364061
transform 1 0 26312 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_8  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2300 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__230__A
timestamp 1586364061
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2116 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_7
timestamp 1586364061
transform 1 0 1748 0 -1 3808
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_22
timestamp 1586364061
transform 1 0 3128 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_26
timestamp 1586364061
transform 1 0 3496 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_30
timestamp 1586364061
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_3.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5612 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_41
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_8  FILLER_2_52
timestamp 1586364061
transform 1 0 5888 0 -1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  FILLER_2_60
timestamp 1586364061
transform 1 0 6624 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_72
timestamp 1586364061
transform 1 0 7728 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_84
timestamp 1586364061
transform 1 0 8832 0 -1 3808
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9936 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_93
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_99
timestamp 1586364061
transform 1 0 10212 0 -1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11408 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_111
timestamp 1586364061
transform 1 0 11316 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_115
timestamp 1586364061
transform 1 0 11684 0 -1 3808
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 866 592
use scs8hd_fill_1  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_2_135
timestamp 1586364061
transform 1 0 13524 0 -1 3808
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__140__B
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_157
timestamp 1586364061
transform 1 0 15548 0 -1 3808
box -38 -48 774 592
use scs8hd_buf_2  _231_
timestamp 1586364061
transform 1 0 16560 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  FILLER_2_165
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_2_172
timestamp 1586364061
transform 1 0 16928 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_184
timestamp 1586364061
transform 1 0 18032 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_196
timestamp 1586364061
transform 1 0 19136 0 -1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_6  FILLER_2_208
timestamp 1586364061
transform 1 0 20240 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_12  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_227
timestamp 1586364061
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_239
timestamp 1586364061
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_251
timestamp 1586364061
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_263
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_buf_2  _229_
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__191__A
timestamp 1586364061
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_11
timestamp 1586364061
transform 1 0 2116 0 1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_3_16
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_30
timestamp 1586364061
transform 1 0 3864 0 1 3808
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_47
timestamp 1586364061
transform 1 0 5428 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_51
timestamp 1586364061
transform 1 0 5796 0 1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6256 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_54
timestamp 1586364061
transform 1 0 6072 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_58
timestamp 1586364061
transform 1 0 6440 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_71
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_75
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_79
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_84
timestamp 1586364061
transform 1 0 8832 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_88
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 406 592
use scs8hd_inv_1  mux_left_track_11.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9568 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__239__A
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_95
timestamp 1586364061
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_99
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_103
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_107
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_136
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_140
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 406 592
use scs8hd_nor2_4  _140_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14628 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__140__A
timestamp 1586364061
transform 1 0 14444 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_144
timestamp 1586364061
transform 1 0 14352 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_156
timestamp 1586364061
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_160
timestamp 1586364061
transform 1 0 15824 0 1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16284 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16744 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16100 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_168
timestamp 1586364061
transform 1 0 16560 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_172
timestamp 1586364061
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_176
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18216 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_182
timestamp 1586364061
transform 1 0 17848 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_3_188
timestamp 1586364061
transform 1 0 18400 0 1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_199
timestamp 1586364061
transform 1 0 19412 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_3_211
timestamp 1586364061
transform 1 0 20516 0 1 3808
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_221
timestamp 1586364061
transform 1 0 21436 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_3_233
timestamp 1586364061
transform 1 0 22540 0 1 3808
box -38 -48 774 592
use scs8hd_decap_3  FILLER_3_241
timestamp 1586364061
transform 1 0 23276 0 1 3808
box -38 -48 314 592
use scs8hd_decap_12  FILLER_3_245
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_257
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_3_269
timestamp 1586364061
transform 1 0 25852 0 1 3808
box -38 -48 774 592
use scs8hd_inv_8  _191_
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_3.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__229__A
timestamp 1586364061
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_10
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 774 592
use scs8hd_decap_6  FILLER_4_32
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 590 592
use scs8hd_conb_1  _216_
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5888 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5612 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4600 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_40
timestamp 1586364061
transform 1 0 4784 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_44
timestamp 1586364061
transform 1 0 5152 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_48
timestamp 1586364061
transform 1 0 5520 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_51
timestamp 1586364061
transform 1 0 5796 0 -1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_61
timestamp 1586364061
transform 1 0 6716 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_65
timestamp 1586364061
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_78
timestamp 1586364061
transform 1 0 8280 0 -1 4896
box -38 -48 1142 592
use scs8hd_buf_2  _239_
timestamp 1586364061
transform 1 0 10028 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__160__B
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_90
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_4  FILLER_4_101
timestamp 1586364061
transform 1 0 10396 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_107
timestamp 1586364061
transform 1 0 10948 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11132 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12512 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_118
timestamp 1586364061
transform 1 0 11960 0 -1 4896
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12696 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_135
timestamp 1586364061
transform 1 0 13524 0 -1 4896
box -38 -48 590 592
use scs8hd_inv_1  mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_143
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_147
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_8  FILLER_4_157
timestamp 1586364061
transform 1 0 15548 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16652 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_165
timestamp 1586364061
transform 1 0 16284 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_168
timestamp 1586364061
transform 1 0 16560 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_178
timestamp 1586364061
transform 1 0 17480 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_182
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_189
timestamp 1586364061
transform 1 0 18492 0 -1 4896
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_200
timestamp 1586364061
transform 1 0 19504 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_4_212
timestamp 1586364061
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21252 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_4_215
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_222
timestamp 1586364061
transform 1 0 21528 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_234
timestamp 1586364061
transform 1 0 22632 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_246
timestamp 1586364061
transform 1 0 23736 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_258
timestamp 1586364061
transform 1 0 24840 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_270
timestamp 1586364061
transform 1 0 25944 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_buf_2  _228_
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__228__A
timestamp 1586364061
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_11
timestamp 1586364061
transform 1 0 2116 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_15
timestamp 1586364061
transform 1 0 2484 0 1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_3.LATCH_1_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3128 0 1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__198__A
timestamp 1586364061
transform 1 0 4324 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_18
timestamp 1586364061
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_33
timestamp 1586364061
transform 1 0 4140 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _193_
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__193__A
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_37
timestamp 1586364061
transform 1 0 4508 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_41
timestamp 1586364061
transform 1 0 4876 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_5.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _196_
timestamp 1586364061
transform 1 0 8556 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__194__A
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__196__A
timestamp 1586364061
transform 1 0 8372 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_73
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_77
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use scs8hd_nor2_4  _160_
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__160__A
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_90
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_5_95
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_101
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14076 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_133
timestamp 1586364061
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_137
timestamp 1586364061
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15364 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_150
timestamp 1586364061
transform 1 0 14904 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_154
timestamp 1586364061
transform 1 0 15272 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_157
timestamp 1586364061
transform 1 0 15548 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17480 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_161
timestamp 1586364061
transform 1 0 15916 0 1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_5_175
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_180
timestamp 1586364061
transform 1 0 17664 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_193
timestamp 1586364061
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_197
timestamp 1586364061
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_201
timestamp 1586364061
transform 1 0 19596 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_213
timestamp 1586364061
transform 1 0 20700 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_225
timestamp 1586364061
transform 1 0 21804 0 1 4896
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_6  FILLER_5_237
timestamp 1586364061
transform 1 0 22908 0 1 4896
box -38 -48 590 592
use scs8hd_fill_1  FILLER_5_243
timestamp 1586364061
transform 1 0 23460 0 1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_2  _227_
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_decap_3  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_8
timestamp 1586364061
transform 1 0 1840 0 -1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_7.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1564 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_12
timestamp 1586364061
transform 1 0 2208 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_12
timestamp 1586364061
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__227__A
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__225__A
timestamp 1586364061
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_16
timestamp 1586364061
transform 1 0 2576 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _218_
timestamp 1586364061
transform 1 0 2576 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_19
timestamp 1586364061
transform 1 0 2852 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3036 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_3.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2760 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_35
timestamp 1586364061
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_31
timestamp 1586364061
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__226__A
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_3.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2944 0 1 5984
box -38 -48 1050 592
use scs8hd_inv_8  _198_
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_5.LATCH_1_.latch
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4508 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_41
timestamp 1586364061
transform 1 0 4876 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_46
timestamp 1586364061
transform 1 0 5336 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_39
timestamp 1586364061
transform 1 0 4692 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_60
timestamp 1586364061
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_7_69
timestamp 1586364061
transform 1 0 7452 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_65
timestamp 1586364061
transform 1 0 7084 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_64
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _194_
timestamp 1586364061
transform 1 0 7360 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_79
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_75
timestamp 1586364061
transform 1 0 8004 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_77
timestamp 1586364061
transform 1 0 8188 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8188 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_87
timestamp 1586364061
transform 1 0 9108 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_83
timestamp 1586364061
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8556 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8556 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_94
timestamp 1586364061
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_90
timestamp 1586364061
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_96
timestamp 1586364061
transform 1 0 9936 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10120 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_7.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_7_107
timestamp 1586364061
transform 1 0 10948 0 1 5984
box -38 -48 314 592
use scs8hd_decap_4  FILLER_6_100
timestamp 1586364061
transform 1 0 10304 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10856 0 -1 5984
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_3_.latch
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_4_.latch
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_115
timestamp 1586364061
transform 1 0 11684 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_112
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_116
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_134
timestamp 1586364061
transform 1 0 13432 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_134
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_142
timestamp 1586364061
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_151
timestamp 1586364061
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_147
timestamp 1586364061
transform 1 0 14628 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14812 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14352 0 1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_158
timestamp 1586364061
transform 1 0 15640 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_154
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__159__A
timestamp 1586364061
transform 1 0 15456 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 15180 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_4_.latch
timestamp 1586364061
transform 1 0 15732 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15364 0 1 5984
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17480 0 -1 5984
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__159__B
timestamp 1586364061
transform 1 0 16560 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17296 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_170
timestamp 1586364061
transform 1 0 16744 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_166
timestamp 1586364061
transform 1 0 16376 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_170
timestamp 1586364061
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_174
timestamp 1586364061
transform 1 0 17112 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_187
timestamp 1586364061
transform 1 0 18308 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_191
timestamp 1586364061
transform 1 0 18676 0 -1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__139__A
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19044 0 -1 5984
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__139__B
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_204
timestamp 1586364061
transform 1 0 19872 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_6_212
timestamp 1586364061
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_197
timestamp 1586364061
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_201
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_213
timestamp 1586364061
transform 1 0 20700 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_215
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_227
timestamp 1586364061
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_225
timestamp 1586364061
transform 1 0 21804 0 1 5984
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_239
timestamp 1586364061
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_7_237
timestamp 1586364061
transform 1 0 22908 0 1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_7_243
timestamp 1586364061
transform 1 0 23460 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_251
timestamp 1586364061
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_263
timestamp 1586364061
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_9.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__197__A
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__178__B
timestamp 1586364061
transform 1 0 3680 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_30
timestamp 1586364061
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__175__B
timestamp 1586364061
transform 1 0 5428 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_45
timestamp 1586364061
transform 1 0 5244 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__B
timestamp 1586364061
transform 1 0 6624 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_58
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_62
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_70
timestamp 1586364061
transform 1 0 7544 0 -1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_7.LATCH_0_.latch
timestamp 1586364061
transform 1 0 7820 0 -1 7072
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_8_84
timestamp 1586364061
transform 1 0 8832 0 -1 7072
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__158__B
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_2_.latch
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_108
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_121
timestamp 1586364061
transform 1 0 12236 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13156 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_125
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_140
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use scs8hd_nor2_4  _159_
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_144
timestamp 1586364061
transform 1 0 14352 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_152
timestamp 1586364061
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16560 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_163
timestamp 1586364061
transform 1 0 16100 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_167
timestamp 1586364061
transform 1 0 16468 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_170
timestamp 1586364061
transform 1 0 16744 0 -1 7072
box -38 -48 774 592
use scs8hd_nor2_4  _139_
timestamp 1586364061
transform 1 0 19044 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18860 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_187
timestamp 1586364061
transform 1 0 18308 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_191
timestamp 1586364061
transform 1 0 18676 0 -1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_204
timestamp 1586364061
transform 1 0 19872 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_212
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_buf_2  _226_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_7
timestamp 1586364061
transform 1 0 1748 0 1 7072
box -38 -48 406 592
use scs8hd_decap_4  FILLER_9_13
timestamp 1586364061
transform 1 0 2300 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_17
timestamp 1586364061
transform 1 0 2668 0 1 7072
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2944 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_31
timestamp 1586364061
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_35
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__C
timestamp 1586364061
transform 1 0 5888 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_50
timestamp 1586364061
transform 1 0 5704 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_7.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 7544 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__D
timestamp 1586364061
transform 1 0 6256 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__175__A
timestamp 1586364061
transform 1 0 6992 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_54
timestamp 1586364061
transform 1 0 6072 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_58
timestamp 1586364061
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_66
timestamp 1586364061
transform 1 0 7176 0 1 7072
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_7.LATCH_1_.latch
timestamp 1586364061
transform 1 0 7728 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9292 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__195__A
timestamp 1586364061
transform 1 0 8924 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_83
timestamp 1586364061
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_87
timestamp 1586364061
transform 1 0 9108 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9476 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__158__A
timestamp 1586364061
transform 1 0 10856 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_100
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_104
timestamp 1586364061
transform 1 0 10672 0 1 7072
box -38 -48 222 592
use scs8hd_conb_1  _208_
timestamp 1586364061
transform 1 0 11316 0 1 7072
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_108
timestamp 1586364061
transform 1 0 11040 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_114
timestamp 1586364061
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_118
timestamp 1586364061
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__137__A
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_132
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_136
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__096__A
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_149
timestamp 1586364061
transform 1 0 14812 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_153
timestamp 1586364061
transform 1 0 15180 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_160
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_2_.latch
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_179
timestamp 1586364061
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_193
timestamp 1586364061
transform 1 0 18860 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_197
timestamp 1586364061
transform 1 0 19228 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_204
timestamp 1586364061
transform 1 0 19872 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_208
timestamp 1586364061
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_220
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_9_232
timestamp 1586364061
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_inv_8  _197_
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use scs8hd_conb_1  _211_
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_6
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_10
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__179__C
timestamp 1586364061
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__C
timestamp 1586364061
transform 1 0 3680 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_30
timestamp 1586364061
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use scs8hd_nor4_4  _175_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 1602 592
use scs8hd_inv_1  mux_left_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4600 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__179__A
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__A
timestamp 1586364061
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_36
timestamp 1586364061
transform 1 0 4416 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_45
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__C
timestamp 1586364061
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_66
timestamp 1586364061
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_70
timestamp 1586364061
transform 1 0 7544 0 -1 8160
box -38 -48 222 592
use scs8hd_inv_8  _195_
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__177__D
timestamp 1586364061
transform 1 0 7728 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_74
timestamp 1586364061
transform 1 0 7912 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_10_84
timestamp 1586364061
transform 1 0 8832 0 -1 8160
box -38 -48 590 592
use scs8hd_nor2_4  _158_
timestamp 1586364061
transform 1 0 10856 0 -1 8160
box -38 -48 866 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9844 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_98
timestamp 1586364061
transform 1 0 10120 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_5_.latch
timestamp 1586364061
transform 1 0 12420 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_115
timestamp 1586364061
transform 1 0 11684 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_119
timestamp 1586364061
transform 1 0 12052 0 -1 8160
box -38 -48 406 592
use scs8hd_buf_1  _137_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__161__B
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_134
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_138
timestamp 1586364061
transform 1 0 13800 0 -1 8160
box -38 -48 222 592
use scs8hd_buf_1  _096_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15732 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_157
timestamp 1586364061
transform 1 0 15548 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_5_.latch
timestamp 1586364061
transform 1 0 16560 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_161
timestamp 1586364061
transform 1 0 15916 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_167
timestamp 1586364061
transform 1 0 16468 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18308 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_179
timestamp 1586364061
transform 1 0 17572 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_183
timestamp 1586364061
transform 1 0 17940 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_186
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_196
timestamp 1586364061
transform 1 0 19136 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_10_208
timestamp 1586364061
transform 1 0 20240 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_12  FILLER_10_215
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_227
timestamp 1586364061
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_239
timestamp 1586364061
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_251
timestamp 1586364061
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_263
timestamp 1586364061
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_buf_1  _165_
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 314 592
use scs8hd_buf_2  _225_
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__A
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_7
timestamp 1586364061
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_11
timestamp 1586364061
transform 1 0 2116 0 1 8160
box -38 -48 406 592
use scs8hd_nor4_4  _178_
timestamp 1586364061
transform 1 0 3680 0 1 8160
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__165__A
timestamp 1586364061
transform 1 0 3128 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__167__A
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_20
timestamp 1586364061
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_24
timestamp 1586364061
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__174__D
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__179__D
timestamp 1586364061
transform 1 0 5428 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_45
timestamp 1586364061
transform 1 0 5244 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_49
timestamp 1586364061
transform 1 0 5612 0 1 8160
box -38 -48 406 592
use scs8hd_nor4_4  _177_
timestamp 1586364061
transform 1 0 6992 0 1 8160
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__174__C
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_55
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_59
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_62
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 222 592
use scs8hd_conb_1  _217_
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__177__A
timestamp 1586364061
transform 1 0 8740 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__177__B
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_81
timestamp 1586364061
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_85
timestamp 1586364061
transform 1 0 8924 0 1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10580 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_92
timestamp 1586364061
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_96
timestamp 1586364061
transform 1 0 9936 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_100
timestamp 1586364061
transform 1 0 10304 0 1 8160
box -38 -48 130 592
use scs8hd_nor2_4  _157_
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__A
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_114
timestamp 1586364061
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_118
timestamp 1586364061
transform 1 0 11960 0 1 8160
box -38 -48 222 592
use scs8hd_nor2_4  _138_
timestamp 1586364061
transform 1 0 14076 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__138__A
timestamp 1586364061
transform 1 0 13892 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__161__A
timestamp 1586364061
transform 1 0 13432 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_132
timestamp 1586364061
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_136
timestamp 1586364061
transform 1 0 13616 0 1 8160
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_150
timestamp 1586364061
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_154
timestamp 1586364061
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_169
timestamp 1586364061
transform 1 0 16652 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_173
timestamp 1586364061
transform 1 0 17020 0 1 8160
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_179
timestamp 1586364061
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_193
timestamp 1586364061
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use scs8hd_conb_1  _207_
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__156__A
timestamp 1586364061
transform 1 0 20056 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_197
timestamp 1586364061
transform 1 0 19228 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_204
timestamp 1586364061
transform 1 0 19872 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_220
timestamp 1586364061
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_232
timestamp 1586364061
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 866 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__179__B
timestamp 1586364061
transform 1 0 2392 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_12
timestamp 1586364061
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_16
timestamp 1586364061
transform 1 0 2576 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  _167_
timestamp 1586364061
transform 1 0 2944 0 -1 9248
box -38 -48 314 592
use scs8hd_nor4_4  _179_
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__169__B
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__178__D
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__D
timestamp 1586364061
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__D
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_49
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 406 592
use scs8hd_nor4_4  _174_
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_12_55
timestamp 1586364061
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__146__A
timestamp 1586364061
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__A
timestamp 1586364061
transform 1 0 8096 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__A
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9292 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_74
timestamp 1586364061
transform 1 0 7912 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_78
timestamp 1586364061
transform 1 0 8280 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_83
timestamp 1586364061
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_87
timestamp 1586364061
transform 1 0 9108 0 -1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_91
timestamp 1586364061
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 774 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 11684 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11224 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_112
timestamp 1586364061
transform 1 0 11408 0 -1 9248
box -38 -48 314 592
use scs8hd_nor2_4  _161_
timestamp 1586364061
transform 1 0 13432 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__162__B
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__157__B
timestamp 1586364061
transform 1 0 13248 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_126
timestamp 1586364061
transform 1 0 12696 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_130
timestamp 1586364061
transform 1 0 13064 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_1  _086_
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__110__B
timestamp 1586364061
transform 1 0 15732 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__141__B
timestamp 1586364061
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__138__B
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_143
timestamp 1586364061
transform 1 0 14260 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_147
timestamp 1586364061
transform 1 0 14628 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_12_157
timestamp 1586364061
transform 1 0 15548 0 -1 9248
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16284 0 -1 9248
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__141__A
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_161
timestamp 1586364061
transform 1 0 15916 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_12_176
timestamp 1586364061
transform 1 0 17296 0 -1 9248
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_193
timestamp 1586364061
transform 1 0 18860 0 -1 9248
box -38 -48 774 592
use scs8hd_buf_1  _156_
timestamp 1586364061
transform 1 0 19596 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_204
timestamp 1586364061
transform 1 0 19872 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_2  FILLER_12_212
timestamp 1586364061
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_8
timestamp 1586364061
transform 1 0 1840 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__170__A
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_14
timestamp 1586364061
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1564 0 1 9248
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_11.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2116 0 -1 10336
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_14_26
timestamp 1586364061
transform 1 0 3496 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_22
timestamp 1586364061
transform 1 0 3128 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_18
timestamp 1586364061
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__A
timestamp 1586364061
transform 1 0 3312 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__169__C
timestamp 1586364061
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_14_30
timestamp 1586364061
transform 1 0 3864 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__168__C
timestamp 1586364061
transform 1 0 3680 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_nor4_4  _169_
timestamp 1586364061
transform 1 0 3128 0 1 9248
box -38 -48 1602 592
use scs8hd_decap_3  FILLER_14_39
timestamp 1586364061
transform 1 0 4692 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_1  FILLER_14_36
timestamp 1586364061
transform 1 0 4416 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_1  FILLER_13_43
timestamp 1586364061
transform 1 0 5060 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__180__A
timestamp 1586364061
transform 1 0 4508 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__D
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _172_
timestamp 1586364061
transform 1 0 4968 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_49
timestamp 1586364061
transform 1 0 5612 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_45
timestamp 1586364061
transform 1 0 5244 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_53
timestamp 1586364061
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_46
timestamp 1586364061
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__B
timestamp 1586364061
transform 1 0 5796 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__172__A
timestamp 1586364061
transform 1 0 5428 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__181__C
timestamp 1586364061
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _173_
timestamp 1586364061
transform 1 0 5704 0 1 9248
box -38 -48 314 592
use scs8hd_nor4_4  _181_
timestamp 1586364061
transform 1 0 5980 0 -1 10336
box -38 -48 1602 592
use scs8hd_nor4_4  _176_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__181__B
timestamp 1586364061
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__173__A
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_57
timestamp 1586364061
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_70
timestamp 1586364061
transform 1 0 7544 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_79
timestamp 1586364061
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_75
timestamp 1586364061
transform 1 0 8004 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_79
timestamp 1586364061
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__D
timestamp 1586364061
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__171__A
timestamp 1586364061
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_88
timestamp 1586364061
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_84
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_83
timestamp 1586364061
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__A
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__176__C
timestamp 1586364061
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_11.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _146_
timestamp 1586364061
transform 1 0 8556 0 -1 10336
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_11.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9108 0 1 9248
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_14_106
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_102
timestamp 1586364061
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_102
timestamp 1586364061
transform 1 0 10488 0 1 9248
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__200__A
timestamp 1586364061
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use scs8hd_or2_4  _089_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 10948 0 1 9248
box -38 -48 682 592
use scs8hd_ebufn_2  mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_119
timestamp 1586364061
transform 1 0 12052 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__089__B
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_125
timestamp 1586364061
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_132
timestamp 1586364061
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use scs8hd_decap_6  FILLER_14_140
timestamp 1586364061
transform 1 0 13984 0 -1 10336
box -38 -48 590 592
use scs8hd_fill_2  FILLER_14_136
timestamp 1586364061
transform 1 0 13616 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_140
timestamp 1586364061
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_136
timestamp 1586364061
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__B
timestamp 1586364061
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__162__A
timestamp 1586364061
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _162_
timestamp 1586364061
transform 1 0 12788 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_149
timestamp 1586364061
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_146
timestamp 1586364061
transform 1 0 14536 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__142__B
timestamp 1586364061
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_157
timestamp 1586364061
transform 1 0 15548 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_153
timestamp 1586364061
transform 1 0 15180 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__110__C
timestamp 1586364061
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_or3_4  _110_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use scs8hd_inv_8  _085_
timestamp 1586364061
transform 1 0 14352 0 1 9248
box -38 -48 866 592
use scs8hd_decap_3  FILLER_14_168
timestamp 1586364061
transform 1 0 16560 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  FILLER_14_163
timestamp 1586364061
transform 1 0 16100 0 -1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__143__A
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_178
timestamp 1586364061
transform 1 0 17480 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_174
timestamp 1586364061
transform 1 0 17112 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_170
timestamp 1586364061
transform 1 0 16744 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__B
timestamp 1586364061
transform 1 0 17296 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use scs8hd_nor2_4  _141_
timestamp 1586364061
transform 1 0 15916 0 1 9248
box -38 -48 866 592
use scs8hd_or3_4  _107_
timestamp 1586364061
transform 1 0 16836 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_186
timestamp 1586364061
transform 1 0 18216 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_14_180
timestamp 1586364061
transform 1 0 17664 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_13_182
timestamp 1586364061
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__136__B
timestamp 1586364061
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__C
timestamp 1586364061
transform 1 0 17664 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_14_195
timestamp 1586364061
transform 1 0 19044 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_191
timestamp 1586364061
transform 1 0 18676 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_193
timestamp 1586364061
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18860 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use scs8hd_buf_1  _108_
timestamp 1586364061
transform 1 0 18400 0 -1 10336
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use scs8hd_buf_1  _111_
timestamp 1586364061
transform 1 0 19412 0 -1 10336
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_197
timestamp 1586364061
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_204
timestamp 1586364061
transform 1 0 19872 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_inv_8  _199_
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 866 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__170__C
timestamp 1586364061
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_12
timestamp 1586364061
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_16
timestamp 1586364061
transform 1 0 2576 0 1 10336
box -38 -48 314 592
use scs8hd_nor4_4  _168_
timestamp 1586364061
transform 1 0 3036 0 1 10336
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__168__A
timestamp 1586364061
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _135_
timestamp 1586364061
transform 1 0 5704 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__183__D
timestamp 1586364061
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__B
timestamp 1586364061
transform 1 0 5152 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__168__D
timestamp 1586364061
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_38
timestamp 1586364061
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_42
timestamp 1586364061
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_46
timestamp 1586364061
transform 1 0 5336 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_nor4_4  _182_
timestamp 1586364061
transform 1 0 7544 0 1 10336
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__182__B
timestamp 1586364061
transform 1 0 7360 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__C
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__135__A
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__C
timestamp 1586364061
transform 1 0 6992 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_66
timestamp 1586364061
transform 1 0 7176 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__B
timestamp 1586364061
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_87
timestamp 1586364061
transform 1 0 9108 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _200_
timestamp 1586364061
transform 1 0 9844 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__155__A
timestamp 1586364061
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__155__C
timestamp 1586364061
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_91
timestamp 1586364061
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_104
timestamp 1586364061
transform 1 0 10672 0 1 10336
box -38 -48 222 592
use scs8hd_inv_8  _090_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__B
timestamp 1586364061
transform 1 0 12052 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__C
timestamp 1586364061
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_108
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_113
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_117
timestamp 1586364061
transform 1 0 11868 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_121
timestamp 1586364061
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__087__C
timestamp 1586364061
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_15_138
timestamp 1586364061
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_142
timestamp 1586364061
transform 1 0 14168 0 1 10336
box -38 -48 406 592
use scs8hd_nor2_4  _142_
timestamp 1586364061
transform 1 0 14812 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__104__B
timestamp 1586364061
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__C
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_15_146
timestamp 1586364061
transform 1 0 14536 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_158
timestamp 1586364061
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use scs8hd_nor2_4  _143_
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__097__A
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__C
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_162
timestamp 1586364061
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_or2_4  _136_
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__136__A
timestamp 1586364061
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_191
timestamp 1586364061
transform 1 0 18676 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_195
timestamp 1586364061
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use scs8hd_buf_1  _102_
timestamp 1586364061
transform 1 0 19412 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 19872 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__097__B
timestamp 1586364061
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_202
timestamp 1586364061
transform 1 0 19688 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_206
timestamp 1586364061
transform 1 0 20056 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_218
timestamp 1586364061
transform 1 0 21160 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_230
timestamp 1586364061
transform 1 0 22264 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_242
timestamp 1586364061
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_nor4_4  _170_
timestamp 1586364061
transform 1 0 1656 0 -1 11424
box -38 -48 1602 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__168__B
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__D
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use scs8hd_buf_1  _180_
timestamp 1586364061
transform 1 0 4508 0 -1 11424
box -38 -48 314 592
use scs8hd_nor4_4  _183_
timestamp 1586364061
transform 1 0 5520 0 -1 11424
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__188__A
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__183__A
timestamp 1586364061
transform 1 0 4968 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_36
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_40
timestamp 1586364061
transform 1 0 4784 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__182__C
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_65
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_69
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 130 592
use scs8hd_inv_8  _171_
timestamp 1586364061
transform 1 0 7820 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__185__A
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_72
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_16_82
timestamp 1586364061
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_86
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 406 592
use scs8hd_or3_4  _155_
timestamp 1586364061
transform 1 0 10120 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__147__A
timestamp 1586364061
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__B
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_97
timestamp 1586364061
transform 1 0 10028 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_6  FILLER_16_107
timestamp 1586364061
transform 1 0 10948 0 -1 11424
box -38 -48 590 592
use scs8hd_or3_4  _091_
timestamp 1586364061
transform 1 0 11684 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__114__C
timestamp 1586364061
transform 1 0 11500 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_124
timestamp 1586364061
transform 1 0 12512 0 -1 11424
box -38 -48 222 592
use scs8hd_or3_4  _087_
timestamp 1586364061
transform 1 0 13616 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__125__C
timestamp 1586364061
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__A
timestamp 1586364061
transform 1 0 12696 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_128
timestamp 1586364061
transform 1 0 12880 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_134
timestamp 1586364061
transform 1 0 13432 0 -1 11424
box -38 -48 222 592
use scs8hd_or3_4  _104_
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__142__A
timestamp 1586364061
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_145
timestamp 1586364061
transform 1 0 14444 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_151
timestamp 1586364061
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use scs8hd_or3_4  _097_
timestamp 1586364061
transform 1 0 16836 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__143__B
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_16_163
timestamp 1586364061
transform 1 0 16100 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_3  FILLER_16_168
timestamp 1586364061
transform 1 0 16560 0 -1 11424
box -38 -48 314 592
use scs8hd_inv_8  _100_
timestamp 1586364061
transform 1 0 18400 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__C
timestamp 1586364061
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_180
timestamp 1586364061
transform 1 0 17664 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_16_186
timestamp 1586364061
transform 1 0 18216 0 -1 11424
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_197
timestamp 1586364061
transform 1 0 19228 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_201
timestamp 1586364061
transform 1 0 19596 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_213
timestamp 1586364061
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_buf_2  _223_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__170__B
timestamp 1586364061
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__166__B
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_7
timestamp 1586364061
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_11
timestamp 1586364061
transform 1 0 2116 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 130 592
use scs8hd_nor4_4  _166_
timestamp 1586364061
transform 1 0 3128 0 1 11424
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__166__A
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_18
timestamp 1586364061
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _144_
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 5428 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 4876 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_43
timestamp 1586364061
transform 1 0 5060 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_49
timestamp 1586364061
transform 1 0 5612 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _115_
timestamp 1586364061
transform 1 0 7084 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__144__A
timestamp 1586364061
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__188__D
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 7544 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use scs8hd_decap_3  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use scs8hd_fill_2  FILLER_17_68
timestamp 1586364061
transform 1 0 7360 0 1 11424
box -38 -48 222 592
use scs8hd_nor4_4  _185_
timestamp 1586364061
transform 1 0 8096 0 1 11424
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__185__D
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_72
timestamp 1586364061
transform 1 0 7728 0 1 11424
box -38 -48 222 592
use scs8hd_inv_8  _145_
timestamp 1586364061
transform 1 0 10396 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__145__A
timestamp 1586364061
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__147__C
timestamp 1586364061
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_93
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_97
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use scs8hd_or3_4  _134_
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__114__B
timestamp 1586364061
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__134__C
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_114
timestamp 1586364061
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_17_117
timestamp 1586364061
transform 1 0 11868 0 1 11424
box -38 -48 314 592
use scs8hd_inv_8  _084_
timestamp 1586364061
transform 1 0 13984 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__A
timestamp 1586364061
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_132
timestamp 1586364061
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_136
timestamp 1586364061
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use scs8hd_nor2_4  _150_
timestamp 1586364061
transform 1 0 15548 0 1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__116__A
timestamp 1586364061
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_149
timestamp 1586364061
transform 1 0 14812 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_153
timestamp 1586364061
transform 1 0 15180 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_156
timestamp 1586364061
transform 1 0 15456 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__150__B
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_166
timestamp 1586364061
transform 1 0 16376 0 1 11424
box -38 -48 406 592
use scs8hd_fill_2  FILLER_17_172
timestamp 1586364061
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_176
timestamp 1586364061
transform 1 0 17296 0 1 11424
box -38 -48 406 592
use scs8hd_or3_4  _101_
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__101__B
timestamp 1586364061
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_180
timestamp 1586364061
transform 1 0 17664 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_193
timestamp 1586364061
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use scs8hd_buf_1  _088_
timestamp 1586364061
transform 1 0 19596 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 20056 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 19412 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_197
timestamp 1586364061
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_204
timestamp 1586364061
transform 1 0 19872 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_inv_8  _201_
timestamp 1586364061
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_13.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__170__D
timestamp 1586364061
transform 1 0 1840 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__199__A
timestamp 1586364061
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_6
timestamp 1586364061
transform 1 0 1656 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_10
timestamp 1586364061
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__166__C
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__201__A
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4232 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_23
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 314 592
use scs8hd_inv_1  mux_left_track_13.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5428 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__184__B
timestamp 1586364061
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__223__A
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_39
timestamp 1586364061
transform 1 0 4692 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_43
timestamp 1586364061
transform 1 0 5060 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_18_50
timestamp 1586364061
transform 1 0 5704 0 -1 12512
box -38 -48 222 592
use scs8hd_nor4_4  _188_
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__188__B
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_54
timestamp 1586364061
transform 1 0 6072 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__D
timestamp 1586364061
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__C
timestamp 1586364061
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__185__B
timestamp 1586364061
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_75
timestamp 1586364061
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_79
timestamp 1586364061
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_83
timestamp 1586364061
transform 1 0 8740 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_3  FILLER_18_89
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use scs8hd_or3_4  _147_
timestamp 1586364061
transform 1 0 9844 0 -1 12512
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__203__A
timestamp 1586364061
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_104
timestamp 1586364061
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use scs8hd_or3_4  _114_
timestamp 1586364061
transform 1 0 11684 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_108
timestamp 1586364061
transform 1 0 11040 0 -1 12512
box -38 -48 406 592
use scs8hd_fill_1  FILLER_18_112
timestamp 1586364061
transform 1 0 11408 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_124
timestamp 1586364061
transform 1 0 12512 0 -1 12512
box -38 -48 222 592
use scs8hd_or3_4  _125_
timestamp 1586364061
transform 1 0 13248 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__134__B
timestamp 1586364061
transform 1 0 12696 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__125__B
timestamp 1586364061
transform 1 0 13064 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_128
timestamp 1586364061
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 222 592
use scs8hd_or2_4  _116_
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 682 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__116__B
timestamp 1586364061
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__B
timestamp 1586364061
transform 1 0 14260 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_18_145
timestamp 1586364061
transform 1 0 14444 0 -1 12512
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_4_.latch
timestamp 1586364061
transform 1 0 16744 0 -1 12512
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__150__A
timestamp 1586364061
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16468 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_161
timestamp 1586364061
transform 1 0 15916 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_165
timestamp 1586364061
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_169
timestamp 1586364061
transform 1 0 16652 0 -1 12512
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18492 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 18032 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_18_181
timestamp 1586364061
transform 1 0 17756 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_18_186
timestamp 1586364061
transform 1 0 18216 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_198
timestamp 1586364061
transform 1 0 19320 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_18_210
timestamp 1586364061
transform 1 0 20424 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_6
timestamp 1586364061
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_7
timestamp 1586364061
transform 1 0 1748 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_buf_2  _224_
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use scs8hd_conb_1  _212_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_20_10
timestamp 1586364061
transform 1 0 2024 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_16
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_12
timestamp 1586364061
transform 1 0 2208 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__224__A
timestamp 1586364061
transform 1 0 2208 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2024 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_35
timestamp 1586364061
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_31
timestamp 1586364061
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4140 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_13.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2944 0 1 12512
box -38 -48 1050 592
use scs8hd_decap_6  FILLER_20_41
timestamp 1586364061
transform 1 0 4876 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_42
timestamp 1586364061
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__148__A
timestamp 1586364061
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__D
timestamp 1586364061
transform 1 0 5152 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _148_
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_53
timestamp 1586364061
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_46
timestamp 1586364061
transform 1 0 5336 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__A
timestamp 1586364061
transform 1 0 5428 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__184__C
timestamp 1586364061
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _092_
timestamp 1586364061
transform 1 0 5704 0 1 12512
box -38 -48 314 592
use scs8hd_nor4_4  _184_
timestamp 1586364061
transform 1 0 5612 0 -1 13600
box -38 -48 1602 592
use scs8hd_nor4_4  _187_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__187__D
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__092__A
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__B
timestamp 1586364061
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_57
timestamp 1586364061
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_66
timestamp 1586364061
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_70
timestamp 1586364061
transform 1 0 7544 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_74
timestamp 1586364061
transform 1 0 7912 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_79
timestamp 1586364061
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__C
timestamp 1586364061
transform 1 0 7728 0 -1 13600
box -38 -48 222 592
use scs8hd_or2_4  _093_
timestamp 1586364061
transform 1 0 8188 0 -1 13600
box -38 -48 682 592
use scs8hd_decap_3  FILLER_20_89
timestamp 1586364061
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  FILLER_20_84
timestamp 1586364061
transform 1 0 8832 0 -1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_19_83
timestamp 1586364061
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__C
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__B
timestamp 1586364061
transform 1 0 8924 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__093__A
timestamp 1586364061
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use scs8hd_nor4_4  _186_
timestamp 1586364061
transform 1 0 9108 0 1 12512
box -38 -48 1602 592
use scs8hd_inv_8  _203_
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__099__B
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__B
timestamp 1586364061
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_104
timestamp 1586364061
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_102
timestamp 1586364061
transform 1 0 10488 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_4  FILLER_20_107
timestamp 1586364061
transform 1 0 10948 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_111
timestamp 1586364061
transform 1 0 11316 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_112
timestamp 1586364061
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_108
timestamp 1586364061
transform 1 0 11040 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__186__A
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__B
timestamp 1586364061
transform 1 0 11408 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__124__A
timestamp 1586364061
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use scs8hd_decap_6  FILLER_20_123
timestamp 1586364061
transform 1 0 12420 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_4  FILLER_19_116
timestamp 1586364061
transform 1 0 11776 0 1 12512
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_inv_8  _124_
timestamp 1586364061
transform 1 0 11592 0 -1 13600
box -38 -48 866 592
use scs8hd_inv_8  _113_
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use scs8hd_or2_4  _126_
timestamp 1586364061
transform 1 0 13984 0 1 12512
box -38 -48 682 592
use scs8hd_nor2_4  _151_
timestamp 1586364061
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__151__A
timestamp 1586364061
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__151__B
timestamp 1586364061
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_19_132
timestamp 1586364061
transform 1 0 13248 0 1 12512
box -38 -48 406 592
use scs8hd_fill_2  FILLER_19_138
timestamp 1586364061
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use scs8hd_decap_3  FILLER_20_131
timestamp 1586364061
transform 1 0 13156 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_6  FILLER_20_145
timestamp 1586364061
transform 1 0 14444 0 -1 13600
box -38 -48 590 592
use scs8hd_fill_2  FILLER_19_151
timestamp 1586364061
transform 1 0 14996 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__126__A
timestamp 1586364061
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_157
timestamp 1586364061
transform 1 0 15548 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 15732 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__149__A
timestamp 1586364061
transform 1 0 15180 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_1  _098_
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use scs8hd_nor2_4  _149_
timestamp 1586364061
transform 1 0 15364 0 1 12512
box -38 -48 866 592
use scs8hd_fill_2  FILLER_20_165
timestamp 1586364061
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_161
timestamp 1586364061
transform 1 0 15916 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_19_169
timestamp 1586364061
transform 1 0 16652 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  FILLER_19_164
timestamp 1586364061
transform 1 0 16192 0 1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__149__B
timestamp 1586364061
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 16468 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_178
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_175
timestamp 1586364061
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use scs8hd_buf_1  _105_
timestamp 1586364061
transform 1 0 16928 0 1 12512
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_3_.latch
timestamp 1586364061
transform 1 0 16468 0 -1 13600
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_20_182
timestamp 1586364061
transform 1 0 17848 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_179
timestamp 1586364061
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_20_195
timestamp 1586364061
transform 1 0 19044 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_193
timestamp 1586364061
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 866 592
use scs8hd_fill_2  FILLER_19_204
timestamp 1586364061
transform 1 0 19872 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_197
timestamp 1586364061
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 12512
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 -1 13600
box -38 -48 314 592
use scs8hd_buf_1  _164_
timestamp 1586364061
transform 1 0 19596 0 1 12512
box -38 -48 314 592
use scs8hd_decap_8  FILLER_20_206
timestamp 1586364061
transform 1 0 20056 0 -1 13600
box -38 -48 774 592
use scs8hd_fill_2  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__164__A
timestamp 1586364061
transform 1 0 20424 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_212
timestamp 1586364061
transform 1 0 20608 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_224
timestamp 1586364061
transform 1 0 21712 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_236
timestamp 1586364061
transform 1 0 22816 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_263
timestamp 1586364061
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_2  _222_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_11
timestamp 1586364061
transform 1 0 2116 0 1 13600
box -38 -48 314 592
use scs8hd_fill_2  FILLER_21_16
timestamp 1586364061
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 2944 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_31
timestamp 1586364061
transform 1 0 3956 0 1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_21_35
timestamp 1586364061
transform 1 0 4324 0 1 13600
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_13.LATCH_0_.latch
timestamp 1586364061
transform 1 0 4968 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__094__A
timestamp 1586364061
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_38
timestamp 1586364061
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_53
timestamp 1586364061
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use scs8hd_inv_8  _202_
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__187__A
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_57
timestamp 1586364061
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_71
timestamp 1586364061
transform 1 0 7636 0 1 13600
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_15.LATCH_1_.latch
timestamp 1586364061
transform 1 0 8648 0 1 13600
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_77
timestamp 1586364061
transform 1 0 8188 0 1 13600
box -38 -48 314 592
use scs8hd_nor2_4  _099_
timestamp 1586364061
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_93
timestamp 1586364061
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_97
timestamp 1586364061
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_101
timestamp 1586364061
transform 1 0 10396 0 1 13600
box -38 -48 222 592
use scs8hd_nor2_4  _153_
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__153__A
timestamp 1586364061
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__154__A
timestamp 1586364061
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_114
timestamp 1586364061
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_118
timestamp 1586364061
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14076 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_132
timestamp 1586364061
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use scs8hd_decap_3  FILLER_21_136
timestamp 1586364061
transform 1 0 13616 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_150
timestamp 1586364061
transform 1 0 14904 0 1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_21_156
timestamp 1586364061
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use scs8hd_decap_4  FILLER_21_160
timestamp 1586364061
transform 1 0 15824 0 1 13600
box -38 -48 406 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16376 0 1 13600
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17388 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16192 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_175
timestamp 1586364061
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__152__A
timestamp 1586364061
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_179
timestamp 1586364061
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_193
timestamp 1586364061
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__152__B
timestamp 1586364061
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_197
timestamp 1586364061
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_204
timestamp 1586364061
transform 1 0 19872 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_15.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1472 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_3
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_7
timestamp 1586364061
transform 1 0 1748 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_11
timestamp 1586364061
transform 1 0 2116 0 -1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_22_16
timestamp 1586364061
transform 1 0 2576 0 -1 14688
box -38 -48 222 592
use scs8hd_conb_1  _213_
timestamp 1586364061
transform 1 0 2944 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2760 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__222__A
timestamp 1586364061
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_23
timestamp 1586364061
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_27
timestamp 1586364061
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use scs8hd_decap_4  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use scs8hd_buf_1  _094_
timestamp 1586364061
transform 1 0 4508 0 -1 14688
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5520 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_13.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 4968 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5336 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_22_36
timestamp 1586364061
transform 1 0 4416 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_22_40
timestamp 1586364061
transform 1 0 4784 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6532 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__202__A
timestamp 1586364061
transform 1 0 6900 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_57
timestamp 1586364061
transform 1 0 6348 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_61
timestamp 1586364061
transform 1 0 6716 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_65
timestamp 1586364061
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_69
timestamp 1586364061
transform 1 0 7452 0 -1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__205__A
timestamp 1586364061
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_84
timestamp 1586364061
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_88
timestamp 1586364061
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_102
timestamp 1586364061
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_6  FILLER_22_106
timestamp 1586364061
transform 1 0 10856 0 -1 14688
box -38 -48 590 592
use scs8hd_nor2_4  _154_
timestamp 1586364061
transform 1 0 11408 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__153__B
timestamp 1586364061
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_121
timestamp 1586364061
transform 1 0 12236 0 -1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_0_.latch
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_22_125
timestamp 1586364061
transform 1 0 12604 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_2  FILLER_22_140
timestamp 1586364061
transform 1 0 13984 0 -1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_8  FILLER_22_144
timestamp 1586364061
transform 1 0 14352 0 -1 14688
box -38 -48 774 592
use scs8hd_fill_1  FILLER_22_152
timestamp 1586364061
transform 1 0 15088 0 -1 14688
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17112 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16284 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16652 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_163
timestamp 1586364061
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_167
timestamp 1586364061
transform 1 0 16468 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_22_171
timestamp 1586364061
transform 1 0 16836 0 -1 14688
box -38 -48 314 592
use scs8hd_nor2_4  _152_
timestamp 1586364061
transform 1 0 18676 0 -1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18124 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_183
timestamp 1586364061
transform 1 0 17940 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_187
timestamp 1586364061
transform 1 0 18308 0 -1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_200
timestamp 1586364061
transform 1 0 19504 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_22_212
timestamp 1586364061
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_263
timestamp 1586364061
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_17.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1472 0 1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 2668 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2300 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use scs8hd_fill_1  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use scs8hd_fill_2  FILLER_23_7
timestamp 1586364061
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_11
timestamp 1586364061
transform 1 0 2116 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 2852 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__189__A
timestamp 1586364061
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_30
timestamp 1586364061
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_34
timestamp 1586364061
transform 1 0 4232 0 1 14688
box -38 -48 406 592
use scs8hd_ebufn_2  mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_40
timestamp 1586364061
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_53
timestamp 1586364061
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_57
timestamp 1586364061
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_15.LATCH_0_.latch
timestamp 1586364061
transform 1 0 8556 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 8372 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_15.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8004 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_73
timestamp 1586364061
transform 1 0 7820 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_77
timestamp 1586364061
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10304 0 1 14688
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9752 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_92
timestamp 1586364061
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_96
timestamp 1586364061
transform 1 0 9936 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__B
timestamp 1586364061
transform 1 0 11684 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_109
timestamp 1586364061
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_113
timestamp 1586364061
transform 1 0 11500 0 1 14688
box -38 -48 222 592
use scs8hd_decap_4  FILLER_23_117
timestamp 1586364061
transform 1 0 11868 0 1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_23_121
timestamp 1586364061
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13340 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13156 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12788 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_129
timestamp 1586364061
transform 1 0 12972 0 1 14688
box -38 -48 222 592
use scs8hd_buf_1  _127_
timestamp 1586364061
transform 1 0 15088 0 1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__127__A
timestamp 1586364061
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_144
timestamp 1586364061
transform 1 0 14352 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_148
timestamp 1586364061
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use scs8hd_decap_3  FILLER_23_155
timestamp 1586364061
transform 1 0 15364 0 1 14688
box -38 -48 314 592
use scs8hd_fill_2  FILLER_23_160
timestamp 1586364061
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_2_.latch
timestamp 1586364061
transform 1 0 16192 0 1 14688
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_175
timestamp 1586364061
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_179
timestamp 1586364061
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_23_193
timestamp 1586364061
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use scs8hd_conb_1  _209_
timestamp 1586364061
transform 1 0 19596 0 1 14688
box -38 -48 314 592
use scs8hd_decap_4  FILLER_23_197
timestamp 1586364061
transform 1 0 19228 0 1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_23_204
timestamp 1586364061
transform 1 0 19872 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_216
timestamp 1586364061
transform 1 0 20976 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_228
timestamp 1586364061
transform 1 0 22080 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_23_240
timestamp 1586364061
transform 1 0 23184 0 1 14688
box -38 -48 406 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2024 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_6
timestamp 1586364061
transform 1 0 1656 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_24_12
timestamp 1586364061
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_8  _189_
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_23
timestamp 1586364061
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 5060 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_41
timestamp 1586364061
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_45
timestamp 1586364061
transform 1 0 5244 0 -1 15776
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6348 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_66
timestamp 1586364061
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_24_70
timestamp 1586364061
transform 1 0 7544 0 -1 15776
box -38 -48 222 592
use scs8hd_inv_8  _205_
timestamp 1586364061
transform 1 0 7912 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7728 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_83
timestamp 1586364061
transform 1 0 8740 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_91
timestamp 1586364061
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_24_102
timestamp 1586364061
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_24_106
timestamp 1586364061
transform 1 0 10856 0 -1 15776
box -38 -48 406 592
use scs8hd_nor2_4  _106_
timestamp 1586364061
transform 1 0 11224 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_8  FILLER_24_119
timestamp 1586364061
transform 1 0 12052 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__B
timestamp 1586364061
transform 1 0 12880 0 -1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13340 0 -1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_24_127
timestamp 1586364061
transform 1 0 12788 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  FILLER_24_130
timestamp 1586364061
transform 1 0 13064 0 -1 15776
box -38 -48 314 592
use scs8hd_fill_1  FILLER_24_135
timestamp 1586364061
transform 1 0 13524 0 -1 15776
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__131__A
timestamp 1586364061
transform 1 0 15732 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_8  FILLER_24_145
timestamp 1586364061
transform 1 0 14444 0 -1 15776
box -38 -48 774 592
use scs8hd_decap_4  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_24_158
timestamp 1586364061
transform 1 0 15640 0 -1 15776
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_track_9.LATCH_5_.latch
timestamp 1586364061
transform 1 0 16192 0 -1 15776
box -38 -48 1050 592
use scs8hd_decap_3  FILLER_24_161
timestamp 1586364061
transform 1 0 15916 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_24_175
timestamp 1586364061
transform 1 0 17204 0 -1 15776
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17940 0 -1 15776
box -38 -48 866 592
use scs8hd_decap_12  FILLER_24_192
timestamp 1586364061
transform 1 0 18768 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_8  FILLER_24_204
timestamp 1586364061
transform 1 0 19872 0 -1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_24_212
timestamp 1586364061
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1748 0 1 15776
box -38 -48 314 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2576 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 1564 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_10
timestamp 1586364061
transform 1 0 2024 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_14
timestamp 1586364061
transform 1 0 2392 0 1 15776
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4324 0 1 15776
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2760 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4048 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_31
timestamp 1586364061
transform 1 0 3956 0 1 15776
box -38 -48 130 592
use scs8hd_fill_1  FILLER_25_34
timestamp 1586364061
transform 1 0 4232 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5336 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_44
timestamp 1586364061
transform 1 0 5152 0 1 15776
box -38 -48 222 592
use scs8hd_decap_6  FILLER_25_48
timestamp 1586364061
transform 1 0 5520 0 1 15776
box -38 -48 590 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6900 0 1 15776
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_54
timestamp 1586364061
transform 1 0 6072 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_57
timestamp 1586364061
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 130 592
use scs8hd_inv_8  _204_
timestamp 1586364061
transform 1 0 8740 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__204__A
timestamp 1586364061
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_72
timestamp 1586364061
transform 1 0 7728 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_76
timestamp 1586364061
transform 1 0 8096 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_80
timestamp 1586364061
transform 1 0 8464 0 1 15776
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_92
timestamp 1586364061
transform 1 0 9568 0 1 15776
box -38 -48 406 592
use scs8hd_fill_2  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__119__A
timestamp 1586364061
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_111
timestamp 1586364061
transform 1 0 11316 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_115
timestamp 1586364061
transform 1 0 11684 0 1 15776
box -38 -48 406 592
use scs8hd_fill_1  FILLER_25_119
timestamp 1586364061
transform 1 0 12052 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _119_
timestamp 1586364061
transform 1 0 12604 0 1 15776
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14168 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__121__A
timestamp 1586364061
transform 1 0 13616 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_134
timestamp 1586364061
transform 1 0 13432 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_138
timestamp 1586364061
transform 1 0 13800 0 1 15776
box -38 -48 222 592
use scs8hd_nor2_4  _131_
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__129__A
timestamp 1586364061
transform 1 0 15548 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__131__B
timestamp 1586364061
transform 1 0 15180 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_151
timestamp 1586364061
transform 1 0 14996 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_155
timestamp 1586364061
transform 1 0 15364 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17296 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__129__B
timestamp 1586364061
transform 1 0 16744 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_168
timestamp 1586364061
transform 1 0 16560 0 1 15776
box -38 -48 222 592
use scs8hd_decap_4  FILLER_25_172
timestamp 1586364061
transform 1 0 16928 0 1 15776
box -38 -48 406 592
use scs8hd_decap_4  FILLER_25_178
timestamp 1586364061
transform 1 0 17480 0 1 15776
box -38 -48 406 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19044 0 1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18492 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use scs8hd_fill_1  FILLER_25_182
timestamp 1586364061
transform 1 0 17848 0 1 15776
box -38 -48 130 592
use scs8hd_fill_2  FILLER_25_187
timestamp 1586364061
transform 1 0 18308 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_191
timestamp 1586364061
transform 1 0 18676 0 1 15776
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19504 0 1 15776
box -38 -48 222 592
use scs8hd_fill_2  FILLER_25_198
timestamp 1586364061
transform 1 0 19320 0 1 15776
box -38 -48 222 592
use scs8hd_decap_12  FILLER_25_202
timestamp 1586364061
transform 1 0 19688 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_214
timestamp 1586364061
transform 1 0 20792 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_226
timestamp 1586364061
transform 1 0 21896 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_6  FILLER_25_238
timestamp 1586364061
transform 1 0 23000 0 1 15776
box -38 -48 590 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1564 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_conb_1  _210_
timestamp 1586364061
transform 1 0 1748 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_14
timestamp 1586364061
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_10
timestamp 1586364061
transform 1 0 2024 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_9
timestamp 1586364061
transform 1 0 1932 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__190__A
timestamp 1586364061
transform 1 0 2208 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2024 0 -1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 2760 0 1 16864
box -38 -48 866 592
use scs8hd_ebufn_2  mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3036 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_19
timestamp 1586364061
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_23
timestamp 1586364061
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_41
timestamp 1586364061
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_53
timestamp 1586364061
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_27_49
timestamp 1586364061
transform 1 0 5612 0 1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_51
timestamp 1586364061
transform 1 0 5796 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_6  FILLER_26_45
timestamp 1586364061
transform 1 0 5244 0 -1 16864
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__163__A
timestamp 1586364061
transform 1 0 5428 0 1 16864
box -38 -48 222 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5704 0 1 16864
box -38 -48 314 592
use scs8hd_conb_1  _214_
timestamp 1586364061
transform 1 0 5888 0 -1 16864
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_left_track_17.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6900 0 -1 16864
box -38 -48 1050 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7360 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7176 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_55
timestamp 1586364061
transform 1 0 6164 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_57
timestamp 1586364061
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 406 592
use scs8hd_inv_8  _206_
timestamp 1586364061
transform 1 0 8924 0 1 16864
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__206__A
timestamp 1586364061
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8096 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_74
timestamp 1586364061
transform 1 0 7912 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_12  FILLER_26_78
timestamp 1586364061
transform 1 0 8280 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_27_77
timestamp 1586364061
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_81
timestamp 1586364061
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_94
timestamp 1586364061
transform 1 0 9752 0 1 16864
box -38 -48 314 592
use scs8hd_decap_8  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_26_90
timestamp 1586364061
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_2  FILLER_27_99
timestamp 1586364061
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_101
timestamp 1586364061
transform 1 0 10396 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 10580 0 1 16864
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 10580 0 -1 16864
box -38 -48 1050 592
use scs8hd_fill_2  FILLER_27_118
timestamp 1586364061
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_114
timestamp 1586364061
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_26_118
timestamp 1586364061
transform 1 0 11960 0 -1 16864
box -38 -48 590 592
use scs8hd_fill_2  FILLER_26_114
timestamp 1586364061
transform 1 0 11592 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11776 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__117__A
timestamp 1586364061
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_124
timestamp 1586364061
transform 1 0 12512 0 -1 16864
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_buf_1  _117_
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use scs8hd_fill_2  FILLER_27_131
timestamp 1586364061
transform 1 0 13156 0 1 16864
box -38 -48 222 592
use scs8hd_decap_3  FILLER_27_126
timestamp 1586364061
transform 1 0 12696 0 1 16864
box -38 -48 314 592
use scs8hd_fill_1  FILLER_26_127
timestamp 1586364061
transform 1 0 12788 0 -1 16864
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__119__B
timestamp 1586364061
transform 1 0 12604 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 12972 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 13340 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_137
timestamp 1586364061
transform 1 0 13708 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13892 0 -1 16864
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_2_.latch
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 1050 592
use scs8hd_nor2_4  _121_
timestamp 1586364061
transform 1 0 12880 0 -1 16864
box -38 -48 866 592
use scs8hd_decap_4  FILLER_27_150
timestamp 1586364061
transform 1 0 14904 0 1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_146
timestamp 1586364061
transform 1 0 14536 0 1 16864
box -38 -48 222 592
use scs8hd_decap_8  FILLER_26_145
timestamp 1586364061
transform 1 0 14444 0 -1 16864
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14260 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14720 0 1 16864
box -38 -48 222 592
use scs8hd_decap_6  FILLER_27_156
timestamp 1586364061
transform 1 0 15456 0 1 16864
box -38 -48 590 592
use scs8hd_fill_1  FILLER_26_158
timestamp 1586364061
transform 1 0 15640 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15272 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_nor2_4  _129_
timestamp 1586364061
transform 1 0 15732 0 -1 16864
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_2_.latch
timestamp 1586364061
transform 1 0 16192 0 1 16864
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 17296 0 -1 16864
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16744 0 -1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_26_168
timestamp 1586364061
transform 1 0 16560 0 -1 16864
box -38 -48 222 592
use scs8hd_decap_4  FILLER_26_172
timestamp 1586364061
transform 1 0 16928 0 -1 16864
box -38 -48 406 592
use scs8hd_fill_2  FILLER_27_175
timestamp 1586364061
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use scs8hd_fill_2  FILLER_27_179
timestamp 1586364061
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use scs8hd_fill_1  FILLER_26_186
timestamp 1586364061
transform 1 0 18216 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_183
timestamp 1586364061
transform 1 0 17940 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_179
timestamp 1586364061
transform 1 0 17572 0 -1 16864
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18308 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_193
timestamp 1586364061
transform 1 0 18860 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_205
timestamp 1586364061
transform 1 0 19964 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_217
timestamp 1586364061
transform 1 0 21068 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_229
timestamp 1586364061
transform 1 0 22172 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_27_241
timestamp 1586364061
transform 1 0 23276 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_inv_8  _190_
timestamp 1586364061
transform 1 0 2392 0 -1 17952
box -38 -48 866 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_6
timestamp 1586364061
transform 1 0 1656 0 -1 17952
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_23
timestamp 1586364061
transform 1 0 3220 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_buf_1  _163_
timestamp 1586364061
transform 1 0 5428 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_28_50
timestamp 1586364061
transform 1 0 5704 0 -1 17952
box -38 -48 774 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6440 0 -1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_6  FILLER_28_61
timestamp 1586364061
transform 1 0 6716 0 -1 17952
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__095__A
timestamp 1586364061
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_8  FILLER_28_78
timestamp 1586364061
transform 1 0 8280 0 -1 17952
box -38 -48 774 592
use scs8hd_decap_4  FILLER_28_88
timestamp 1586364061
transform 1 0 9200 0 -1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10028 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10580 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_100
timestamp 1586364061
transform 1 0 10304 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11040 0 -1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_121
timestamp 1586364061
transform 1 0 12236 0 -1 17952
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_4_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__118__A
timestamp 1586364061
transform 1 0 12696 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13248 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_1  FILLER_28_125
timestamp 1586364061
transform 1 0 12604 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_128
timestamp 1586364061
transform 1 0 12880 0 -1 17952
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__128__B
timestamp 1586364061
transform 1 0 15732 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_28_145
timestamp 1586364061
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_4  FILLER_28_149
timestamp 1586364061
transform 1 0 14812 0 -1 17952
box -38 -48 406 592
use scs8hd_fill_2  FILLER_28_157
timestamp 1586364061
transform 1 0 15548 0 -1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_4_.latch
timestamp 1586364061
transform 1 0 16744 0 -1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16192 0 -1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16560 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_161
timestamp 1586364061
transform 1 0 15916 0 -1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 222 592
use scs8hd_conb_1  _220_
timestamp 1586364061
transform 1 0 18492 0 -1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18032 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_28_181
timestamp 1586364061
transform 1 0 17756 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_28_186
timestamp 1586364061
transform 1 0 18216 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_192
timestamp 1586364061
transform 1 0 18768 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_8  FILLER_28_204
timestamp 1586364061
transform 1 0 19872 0 -1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_28_212
timestamp 1586364061
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_inv_1  mux_left_track_11.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_6
timestamp 1586364061
transform 1 0 1656 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_10
timestamp 1586364061
transform 1 0 2024 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_22
timestamp 1586364061
transform 1 0 3128 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_34
timestamp 1586364061
transform 1 0 4232 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_46
timestamp 1586364061
transform 1 0 5336 0 1 17952
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6992 0 1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7452 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_58
timestamp 1586364061
transform 1 0 6440 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_67
timestamp 1586364061
transform 1 0 7268 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_71
timestamp 1586364061
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use scs8hd_nor2_4  _095_
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 866 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8004 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8464 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_78
timestamp 1586364061
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_82
timestamp 1586364061
transform 1 0 8648 0 1 17952
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 10580 0 1 17952
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_95
timestamp 1586364061
transform 1 0 9844 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_99
timestamp 1586364061
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__118__B
timestamp 1586364061
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_114
timestamp 1586364061
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_118
timestamp 1586364061
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use scs8hd_nor2_4  _118_
timestamp 1586364061
transform 1 0 12696 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 13708 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14076 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_139
timestamp 1586364061
transform 1 0 13892 0 1 17952
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 17952
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 17952
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__128__A
timestamp 1586364061
transform 1 0 15364 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_152
timestamp 1586364061
transform 1 0 15088 0 1 17952
box -38 -48 314 592
use scs8hd_decap_3  FILLER_29_157
timestamp 1586364061
transform 1 0 15548 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17296 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_169
timestamp 1586364061
transform 1 0 16652 0 1 17952
box -38 -48 314 592
use scs8hd_fill_2  FILLER_29_174
timestamp 1586364061
transform 1 0 17112 0 1 17952
box -38 -48 222 592
use scs8hd_decap_3  FILLER_29_178
timestamp 1586364061
transform 1 0 17480 0 1 17952
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_193
timestamp 1586364061
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 17952
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 17952
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_197
timestamp 1586364061
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use scs8hd_fill_2  FILLER_29_204
timestamp 1586364061
transform 1 0 19872 0 1 17952
box -38 -48 222 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7544 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__095__B
timestamp 1586364061
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_30_73
timestamp 1586364061
transform 1 0 7820 0 -1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_30_84
timestamp 1586364061
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_88
timestamp 1586364061
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10120 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9936 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_30_107
timestamp 1586364061
transform 1 0 10948 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11684 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_111
timestamp 1586364061
transform 1 0 11316 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_2  FILLER_30_124
timestamp 1586364061
transform 1 0 12512 0 -1 19040
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_5_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__123__A
timestamp 1586364061
transform 1 0 12696 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13248 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_128
timestamp 1586364061
transform 1 0 12880 0 -1 19040
box -38 -48 406 592
use scs8hd_nor2_4  _128_
timestamp 1586364061
transform 1 0 15364 0 -1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14628 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_145
timestamp 1586364061
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_30_149
timestamp 1586364061
transform 1 0 14812 0 -1 19040
box -38 -48 406 592
use scs8hd_fill_1  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_5_.latch
timestamp 1586364061
transform 1 0 16928 0 -1 19040
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_164
timestamp 1586364061
transform 1 0 16192 0 -1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_30_168
timestamp 1586364061
transform 1 0 16560 0 -1 19040
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 -1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18216 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_30_183
timestamp 1586364061
transform 1 0 17940 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_30_188
timestamp 1586364061
transform 1 0 18400 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_200
timestamp 1586364061
transform 1 0 19504 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_30_212
timestamp 1586364061
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_decap_8  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  FILLER_31_70
timestamp 1586364061
transform 1 0 7544 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8004 0 1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8556 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_78
timestamp 1586364061
transform 1 0 8280 0 1 19040
box -38 -48 314 592
use scs8hd_decap_3  FILLER_31_83
timestamp 1586364061
transform 1 0 8740 0 1 19040
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10580 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_95
timestamp 1586364061
transform 1 0 9844 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_99
timestamp 1586364061
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__122__A
timestamp 1586364061
transform 1 0 12052 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__123__B
timestamp 1586364061
transform 1 0 11684 0 1 19040
box -38 -48 222 592
use scs8hd_decap_3  FILLER_31_112
timestamp 1586364061
transform 1 0 11408 0 1 19040
box -38 -48 314 592
use scs8hd_fill_2  FILLER_31_117
timestamp 1586364061
transform 1 0 11868 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_121
timestamp 1586364061
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use scs8hd_fill_2  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 222 592
use scs8hd_nor2_4  _123_
timestamp 1586364061
transform 1 0 12604 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__122__B
timestamp 1586364061
transform 1 0 13616 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13984 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_134
timestamp 1586364061
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_138
timestamp 1586364061
transform 1 0 13800 0 1 19040
box -38 -48 222 592
use scs8hd_fill_1  FILLER_31_142
timestamp 1586364061
transform 1 0 14168 0 1 19040
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15824 0 1 19040
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14260 0 1 19040
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 15640 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_152
timestamp 1586364061
transform 1 0 15088 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_156
timestamp 1586364061
transform 1 0 15456 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_169
timestamp 1586364061
transform 1 0 16652 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_173
timestamp 1586364061
transform 1 0 17020 0 1 19040
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18216 0 1 19040
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_179
timestamp 1586364061
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_195
timestamp 1586364061
transform 1 0 19044 0 1 19040
box -38 -48 222 592
use scs8hd_conb_1  _221_
timestamp 1586364061
transform 1 0 20792 0 1 19040
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19780 0 1 19040
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19228 0 1 19040
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19596 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_199
timestamp 1586364061
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use scs8hd_fill_2  FILLER_31_206
timestamp 1586364061
transform 1 0 20056 0 1 19040
box -38 -48 222 592
use scs8hd_decap_4  FILLER_31_210
timestamp 1586364061
transform 1 0 20424 0 1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_31_217
timestamp 1586364061
transform 1 0 21068 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_229
timestamp 1586364061
transform 1 0 22172 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_3  FILLER_31_241
timestamp 1586364061
transform 1 0 23276 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_conb_1  _219_
timestamp 1586364061
transform 1 0 7544 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 -1 20128
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__112__B
timestamp 1586364061
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_32_73
timestamp 1586364061
transform 1 0 7820 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_32_84
timestamp 1586364061
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_88
timestamp 1586364061
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10396 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10212 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9844 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_97
timestamp 1586364061
transform 1 0 10028 0 -1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _122_
timestamp 1586364061
transform 1 0 12052 0 -1 20128
box -38 -48 866 592
use scs8hd_decap_8  FILLER_32_110
timestamp 1586364061
transform 1 0 11224 0 -1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_32_118
timestamp 1586364061
transform 1 0 11960 0 -1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13616 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13156 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_3  FILLER_32_128
timestamp 1586364061
transform 1 0 12880 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_3  FILLER_32_133
timestamp 1586364061
transform 1 0 13340 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_145
timestamp 1586364061
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_149
timestamp 1586364061
transform 1 0 14812 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_6  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 590 592
use scs8hd_fill_1  FILLER_32_160
timestamp 1586364061
transform 1 0 15824 0 -1 20128
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 16100 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17112 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 15916 0 -1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_172
timestamp 1586364061
transform 1 0 16928 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_176
timestamp 1586364061
transform 1 0 17296 0 -1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17664 0 -1 20128
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18676 0 -1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_32_189
timestamp 1586364061
transform 1 0 18492 0 -1 20128
box -38 -48 222 592
use scs8hd_decap_4  FILLER_32_193
timestamp 1586364061
transform 1 0 18860 0 -1 20128
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_8  FILLER_32_206
timestamp 1586364061
transform 1 0 20056 0 -1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_34_74
timestamp 1586364061
transform 1 0 7912 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_77
timestamp 1586364061
transform 1 0 8188 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__109__B
timestamp 1586364061
transform 1 0 8372 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 8004 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_84
timestamp 1586364061
transform 1 0 8832 0 -1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_81
timestamp 1586364061
transform 1 0 8556 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 8740 0 1 20128
box -38 -48 222 592
use scs8hd_nor2_4  _112_
timestamp 1586364061
transform 1 0 8924 0 1 20128
box -38 -48 866 592
use scs8hd_nor2_4  _109_
timestamp 1586364061
transform 1 0 8004 0 -1 21216
box -38 -48 866 592
use scs8hd_decap_3  FILLER_34_98
timestamp 1586364061
transform 1 0 10120 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_3  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_94
timestamp 1586364061
transform 1 0 9752 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9936 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 9936 0 -1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 10304 0 1 20128
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10488 0 1 20128
box -38 -48 866 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 10396 0 -1 21216
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_34_112
timestamp 1586364061
transform 1 0 11408 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_4  FILLER_33_115
timestamp 1586364061
transform 1 0 11684 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_111
timestamp 1586364061
transform 1 0 11316 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 11500 0 1 20128
box -38 -48 222 592
use scs8hd_decap_8  FILLER_34_123
timestamp 1586364061
transform 1 0 12420 0 -1 21216
box -38 -48 774 592
use scs8hd_decap_4  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 406 592
use scs8hd_fill_1  FILLER_33_119
timestamp 1586364061
transform 1 0 12052 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_6_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12144 0 -1 21216
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_0_.latch
timestamp 1586364061
transform 1 0 13156 0 -1 21216
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_1_.latch
timestamp 1586364061
transform 1 0 13340 0 1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 13156 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 12788 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_129
timestamp 1586364061
transform 1 0 12972 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_142
timestamp 1586364061
transform 1 0 14168 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_34_146
timestamp 1586364061
transform 1 0 14536 0 -1 21216
box -38 -48 590 592
use scs8hd_decap_4  FILLER_33_148
timestamp 1586364061
transform 1 0 14720 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_144
timestamp 1586364061
transform 1 0 14352 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14536 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14352 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_152
timestamp 1586364061
transform 1 0 15088 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_33_156
timestamp 1586364061
transform 1 0 15456 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_33_152
timestamp 1586364061
transform 1 0 15088 0 1 20128
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15456 0 -1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15180 0 1 20128
box -38 -48 314 592
use scs8hd_decap_4  FILLER_34_159
timestamp 1586364061
transform 1 0 15732 0 -1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_160
timestamp 1586364061
transform 1 0 15824 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15640 0 1 20128
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_0_.latch
timestamp 1586364061
transform 1 0 16468 0 -1 21216
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_1_.latch
timestamp 1586364061
transform 1 0 16192 0 1 20128
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16008 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 16192 0 -1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_175
timestamp 1586364061
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use scs8hd_fill_1  FILLER_34_163
timestamp 1586364061
transform 1 0 16100 0 -1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_6  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 590 592
use scs8hd_nor2_4  _133_
timestamp 1586364061
transform 1 0 18216 0 -1 21216
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__133__A
timestamp 1586364061
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__133__B
timestamp 1586364061
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18032 0 -1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_179
timestamp 1586364061
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_33_193
timestamp 1586364061
transform 1 0 18860 0 1 20128
box -38 -48 222 592
use scs8hd_fill_2  FILLER_34_195
timestamp 1586364061
transform 1 0 19044 0 -1 21216
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19596 0 1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 20128
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19228 0 -1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_33_197
timestamp 1586364061
transform 1 0 19228 0 1 20128
box -38 -48 406 592
use scs8hd_fill_2  FILLER_33_204
timestamp 1586364061
transform 1 0 19872 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_199
timestamp 1586364061
transform 1 0 19412 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_34_211
timestamp 1586364061
transform 1 0 20516 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_nor2_4  _103_
timestamp 1586364061
transform 1 0 8372 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 314 592
use scs8hd_decap_6  FILLER_35_88
timestamp 1586364061
transform 1 0 9200 0 1 21216
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 9936 0 1 21216
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 9752 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_107
timestamp 1586364061
transform 1 0 10948 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11132 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11500 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_111
timestamp 1586364061
transform 1 0 11316 0 1 21216
box -38 -48 222 592
use scs8hd_decap_6  FILLER_35_115
timestamp 1586364061
transform 1 0 11684 0 1 21216
box -38 -48 590 592
use scs8hd_fill_1  FILLER_35_121
timestamp 1586364061
transform 1 0 12236 0 1 21216
box -38 -48 130 592
use scs8hd_decap_3  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_7_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12880 0 1 21216
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13892 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13340 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13708 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12696 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_131
timestamp 1586364061
transform 1 0 13156 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__130__A
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__A
timestamp 1586364061
transform 1 0 15364 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__132__B
timestamp 1586364061
transform 1 0 14996 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_148
timestamp 1586364061
transform 1 0 14720 0 1 21216
box -38 -48 314 592
use scs8hd_fill_2  FILLER_35_153
timestamp 1586364061
transform 1 0 15180 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_157
timestamp 1586364061
transform 1 0 15548 0 1 21216
box -38 -48 222 592
use scs8hd_nor2_4  _130_
timestamp 1586364061
transform 1 0 15916 0 1 21216
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 17112 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 17480 0 1 21216
box -38 -48 222 592
use scs8hd_decap_4  FILLER_35_170
timestamp 1586364061
transform 1 0 16744 0 1 21216
box -38 -48 406 592
use scs8hd_fill_2  FILLER_35_176
timestamp 1586364061
transform 1 0 17296 0 1 21216
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 1 21216
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18400 0 1 21216
box -38 -48 222 592
use scs8hd_decap_3  FILLER_35_180
timestamp 1586364061
transform 1 0 17664 0 1 21216
box -38 -48 314 592
use scs8hd_decap_4  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19596 0 1 21216
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19964 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_199
timestamp 1586364061
transform 1 0 19412 0 1 21216
box -38 -48 222 592
use scs8hd_fill_2  FILLER_35_203
timestamp 1586364061
transform 1 0 19780 0 1 21216
box -38 -48 222 592
use scs8hd_decap_12  FILLER_35_207
timestamp 1586364061
transform 1 0 20148 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_219
timestamp 1586364061
transform 1 0 21252 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_231
timestamp 1586364061
transform 1 0 22356 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_fill_1  FILLER_35_243
timestamp 1586364061
transform 1 0 23460 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__103__B
timestamp 1586364061
transform 1 0 8372 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_3  FILLER_36_76
timestamp 1586364061
transform 1 0 8096 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_36_81
timestamp 1586364061
transform 1 0 8556 0 -1 22304
box -38 -48 774 592
use scs8hd_decap_3  FILLER_36_89
timestamp 1586364061
transform 1 0 9292 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 10580 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_8  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_36_101
timestamp 1586364061
transform 1 0 10396 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11132 0 -1 22304
box -38 -48 866 592
use scs8hd_decap_8  FILLER_36_118
timestamp 1586364061
transform 1 0 11960 0 -1 22304
box -38 -48 774 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13524 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12788 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_36_126
timestamp 1586364061
transform 1 0 12696 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_6  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 590 592
use scs8hd_nor2_4  _132_
timestamp 1586364061
transform 1 0 15456 0 -1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14536 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_144
timestamp 1586364061
transform 1 0 14352 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_148
timestamp 1586364061
transform 1 0 14720 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_152
timestamp 1586364061
transform 1 0 15088 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_16.LATCH_3_.latch
timestamp 1586364061
transform 1 0 17112 0 -1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__130__B
timestamp 1586364061
transform 1 0 16468 0 -1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_36_165
timestamp 1586364061
transform 1 0 16284 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_36_169
timestamp 1586364061
transform 1 0 16652 0 -1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_36_173
timestamp 1586364061
transform 1 0 17020 0 -1 22304
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18860 0 -1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18676 0 -1 22304
box -38 -48 222 592
use scs8hd_decap_6  FILLER_36_185
timestamp 1586364061
transform 1 0 18124 0 -1 22304
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 590 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 10580 0 1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_track_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 10396 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9660 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10028 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_92
timestamp 1586364061
transform 1 0 9568 0 1 22304
box -38 -48 130 592
use scs8hd_fill_2  FILLER_37_95
timestamp 1586364061
transform 1 0 9844 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_99
timestamp 1586364061
transform 1 0 10212 0 1 22304
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_114
timestamp 1586364061
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_118
timestamp 1586364061
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_track_8.LATCH_3_.latch
timestamp 1586364061
transform 1 0 13616 0 1 22304
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 13432 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_126
timestamp 1586364061
transform 1 0 12696 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_130
timestamp 1586364061
transform 1 0 13064 0 1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15364 0 1 22304
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15180 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_151
timestamp 1586364061
transform 1 0 14996 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16376 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16744 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17112 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_164
timestamp 1586364061
transform 1 0 16192 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_168
timestamp 1586364061
transform 1 0 16560 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_172
timestamp 1586364061
transform 1 0 16928 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_176
timestamp 1586364061
transform 1 0 17296 0 1 22304
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18676 0 1 22304
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 18492 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use scs8hd_fill_1  FILLER_37_180
timestamp 1586364061
transform 1 0 17664 0 1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 406 592
use scs8hd_fill_1  FILLER_37_188
timestamp 1586364061
transform 1 0 18400 0 1 22304
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20056 0 1 22304
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_200
timestamp 1586364061
transform 1 0 19504 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_204
timestamp 1586364061
transform 1 0 19872 0 1 22304
box -38 -48 222 592
use scs8hd_decap_4  FILLER_37_211
timestamp 1586364061
transform 1 0 20516 0 1 22304
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20884 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_217
timestamp 1586364061
transform 1 0 21068 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_229
timestamp 1586364061
transform 1 0 22172 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_3  FILLER_37_241
timestamp 1586364061
transform 1 0 23276 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24564 0 1 22304
box -38 -48 222 592
use scs8hd_fill_2  FILLER_37_253
timestamp 1586364061
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_38_102
timestamp 1586364061
transform 1 0 10488 0 -1 23392
box -38 -48 590 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 11224 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__120__A
timestamp 1586364061
transform 1 0 12512 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11040 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_119
timestamp 1586364061
transform 1 0 12052 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_123
timestamp 1586364061
transform 1 0 12420 0 -1 23392
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12788 0 -1 23392
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13800 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14168 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_38_126
timestamp 1586364061
transform 1 0 12696 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_38_136
timestamp 1586364061
transform 1 0 13616 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_140
timestamp 1586364061
transform 1 0 13984 0 -1 23392
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__244__A
timestamp 1586364061
transform 1 0 14536 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_144
timestamp 1586364061
transform 1 0 14352 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_38_148
timestamp 1586364061
transform 1 0 14720 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_8.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16836 0 -1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 16284 0 -1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_38_163
timestamp 1586364061
transform 1 0 16100 0 -1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_38_167
timestamp 1586364061
transform 1 0 16468 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_174
timestamp 1586364061
transform 1 0 17112 0 -1 23392
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 866 592
use scs8hd_decap_4  FILLER_38_186
timestamp 1586364061
transform 1 0 18216 0 -1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_199
timestamp 1586364061
transform 1 0 19412 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_38_211
timestamp 1586364061
transform 1 0 20516 0 -1 23392
box -38 -48 314 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_218
timestamp 1586364061
transform 1 0 21160 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_230
timestamp 1586364061
transform 1 0 22264 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_242
timestamp 1586364061
transform 1 0 23368 0 -1 23392
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_16.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24564 0 -1 23392
box -38 -48 314 592
use scs8hd_fill_1  FILLER_38_254
timestamp 1586364061
transform 1 0 24472 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_258
timestamp 1586364061
transform 1 0 24840 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_270
timestamp 1586364061
transform 1 0 25944 0 -1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_38_274
timestamp 1586364061
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_6
timestamp 1586364061
transform 1 0 1656 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_10
timestamp 1586364061
transform 1 0 2024 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3036 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3496 0 1 23392
box -38 -48 222 592
use scs8hd_decap_3  FILLER_39_18
timestamp 1586364061
transform 1 0 2760 0 1 23392
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_24
timestamp 1586364061
transform 1 0 3312 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_28
timestamp 1586364061
transform 1 0 3680 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_40
timestamp 1586364061
transform 1 0 4784 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_52
timestamp 1586364061
transform 1 0 5888 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_17.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 7360 0 1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_39_60
timestamp 1586364061
transform 1 0 6624 0 1 23392
box -38 -48 130 592
use scs8hd_decap_6  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_71
timestamp 1586364061
transform 1 0 7636 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_left_track_15.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8556 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7820 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 222 592
use scs8hd_decap_6  FILLER_39_75
timestamp 1586364061
transform 1 0 8004 0 1 23392
box -38 -48 590 592
use scs8hd_fill_2  FILLER_39_84
timestamp 1586364061
transform 1 0 8832 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_39_88
timestamp 1586364061
transform 1 0 9200 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _247_
timestamp 1586364061
transform 1 0 9936 0 -1 24480
box -38 -48 406 592
use scs8hd_buf_2  _248_
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__247__A
timestamp 1586364061
transform 1 0 9936 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__248__A
timestamp 1586364061
transform 1 0 10672 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_102
timestamp 1586364061
transform 1 0 10488 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_106
timestamp 1586364061
transform 1 0 10856 0 1 23392
box -38 -48 406 592
use scs8hd_decap_3  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_100
timestamp 1586364061
transform 1 0 10304 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_40_112
timestamp 1586364061
transform 1 0 11408 0 -1 24480
box -38 -48 314 592
use scs8hd_fill_2  FILLER_39_114
timestamp 1586364061
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 23392
box -38 -48 314 592
use scs8hd_buf_2  _246_
timestamp 1586364061
transform 1 0 11684 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_123
timestamp 1586364061
transform 1 0 12420 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_40_119
timestamp 1586364061
transform 1 0 12052 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_118
timestamp 1586364061
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__120__B
timestamp 1586364061
transform 1 0 12512 0 -1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__246__A
timestamp 1586364061
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_nor2_4  _120_
timestamp 1586364061
transform 1 0 12512 0 1 23392
box -38 -48 866 592
use scs8hd_decap_8  FILLER_40_131
timestamp 1586364061
transform 1 0 13156 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_126
timestamp 1586364061
transform 1 0 12696 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_133
timestamp 1586364061
transform 1 0 13340 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _245_
timestamp 1586364061
transform 1 0 12788 0 -1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_40_139
timestamp 1586364061
transform 1 0 13892 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_137
timestamp 1586364061
transform 1 0 13708 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13892 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__245__A
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 222 592
use scs8hd_buf_2  _244_
timestamp 1586364061
transform 1 0 13984 0 -1 24480
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14076 0 1 23392
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15640 0 1 23392
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15272 0 1 23392
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_150
timestamp 1586364061
transform 1 0 14904 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_156
timestamp 1586364061
transform 1 0 15456 0 1 23392
box -38 -48 222 592
use scs8hd_decap_8  FILLER_40_144
timestamp 1586364061
transform 1 0 14352 0 -1 24480
box -38 -48 774 592
use scs8hd_fill_1  FILLER_40_152
timestamp 1586364061
transform 1 0 15088 0 -1 24480
box -38 -48 130 592
use scs8hd_buf_2  _241_
timestamp 1586364061
transform 1 0 16836 0 -1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__241__A
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 16284 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_39_167
timestamp 1586364061
transform 1 0 16468 0 1 23392
box -38 -48 406 592
use scs8hd_decap_8  FILLER_39_173
timestamp 1586364061
transform 1 0 17020 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_40_163
timestamp 1586364061
transform 1 0 16100 0 -1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_40_167
timestamp 1586364061
transform 1 0 16468 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_8  FILLER_40_175
timestamp 1586364061
transform 1 0 17204 0 -1 24480
box -38 -48 774 592
use scs8hd_decap_3  FILLER_40_183
timestamp 1586364061
transform 1 0 17940 0 -1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__240__A
timestamp 1586364061
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18216 0 -1 24480
box -38 -48 314 592
use scs8hd_buf_2  _240_
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 406 592
use scs8hd_decap_4  FILLER_39_192
timestamp 1586364061
transform 1 0 18768 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_188
timestamp 1586364061
transform 1 0 18400 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 18584 0 1 23392
box -38 -48 222 592
use scs8hd_inv_1  mux_top_track_16.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_189
timestamp 1586364061
transform 1 0 18492 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_39_203
timestamp 1586364061
transform 1 0 19780 0 1 23392
box -38 -48 406 592
use scs8hd_fill_2  FILLER_39_199
timestamp 1586364061
transform 1 0 19412 0 1 23392
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19596 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_40_213
timestamp 1586364061
transform 1 0 20700 0 -1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_39_211
timestamp 1586364061
transform 1 0 20516 0 1 23392
box -38 -48 222 592
use scs8hd_fill_1  FILLER_39_207
timestamp 1586364061
transform 1 0 20148 0 1 23392
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20700 0 1 23392
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_inv_1  mux_top_track_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_40_201
timestamp 1586364061
transform 1 0 19596 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_215
timestamp 1586364061
transform 1 0 20884 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_227
timestamp 1586364061
transform 1 0 21988 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_239
timestamp 1586364061
transform 1 0 23092 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_243
timestamp 1586364061
transform 1 0 23460 0 1 23392
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 24380 0 1 23392
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 24840 0 1 23392
box -38 -48 222 592
use scs8hd_fill_2  FILLER_39_256
timestamp 1586364061
transform 1 0 24656 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_39_260
timestamp 1586364061
transform 1 0 25024 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_4  FILLER_39_272
timestamp 1586364061
transform 1 0 26128 0 1 23392
box -38 -48 406 592
use scs8hd_fill_1  FILLER_39_276
timestamp 1586364061
transform 1 0 26496 0 1 23392
box -38 -48 130 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_inv_1  mux_top_track_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 10580 0 1 24480
box -38 -48 314 592
use scs8hd_decap_4  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 406 592
use scs8hd_fill_1  FILLER_41_102
timestamp 1586364061
transform 1 0 10488 0 1 24480
box -38 -48 130 592
use scs8hd_fill_2  FILLER_41_106
timestamp 1586364061
transform 1 0 10856 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11040 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_buf_2  _243_
timestamp 1586364061
transform 1 0 13892 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 13708 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 222 592
use scs8hd_buf_2  _242_
timestamp 1586364061
transform 1 0 14996 0 1 24480
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__243__A
timestamp 1586364061
transform 1 0 14444 0 1 24480
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__242__A
timestamp 1586364061
transform 1 0 15548 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_143
timestamp 1586364061
transform 1 0 14260 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 406 592
use scs8hd_fill_2  FILLER_41_155
timestamp 1586364061
transform 1 0 15364 0 1 24480
box -38 -48 222 592
use scs8hd_decap_4  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 406 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16100 0 1 24480
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 16560 0 1 24480
box -38 -48 222 592
use scs8hd_fill_2  FILLER_41_166
timestamp 1586364061
transform 1 0 16376 0 1 24480
box -38 -48 222 592
use scs8hd_decap_12  FILLER_41_170
timestamp 1586364061
transform 1 0 16744 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_fill_1  FILLER_41_182
timestamp 1586364061
transform 1 0 17848 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_inv_1  mux_top_track_8.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 13800 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_141
timestamp 1586364061
transform 1 0 14076 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_fill_2  FILLER_42_153
timestamp 1586364061
transform 1 0 15180 0 -1 25568
box -38 -48 222 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal3 s 27520 4496 28000 4616 6 address[0]
port 0 nsew default input
rlabel metal3 s 27520 7624 28000 7744 6 address[1]
port 1 nsew default input
rlabel metal3 s 27520 10752 28000 10872 6 address[2]
port 2 nsew default input
rlabel metal3 s 27520 13880 28000 14000 6 address[3]
port 3 nsew default input
rlabel metal3 s 27520 17008 28000 17128 6 address[4]
port 4 nsew default input
rlabel metal3 s 27520 20136 28000 20256 6 address[5]
port 5 nsew default input
rlabel metal3 s 27520 23264 28000 23384 6 address[6]
port 6 nsew default input
rlabel metal2 s 478 0 534 480 6 bottom_left_grid_pin_13_
port 7 nsew default input
rlabel metal2 s 25318 0 25374 480 6 bottom_right_grid_pin_11_
port 8 nsew default input
rlabel metal2 s 26330 0 26386 480 6 bottom_right_grid_pin_13_
port 9 nsew default input
rlabel metal2 s 27342 0 27398 480 6 bottom_right_grid_pin_15_
port 10 nsew default input
rlabel metal2 s 20074 0 20130 480 6 bottom_right_grid_pin_1_
port 11 nsew default input
rlabel metal2 s 21178 0 21234 480 6 bottom_right_grid_pin_3_
port 12 nsew default input
rlabel metal2 s 22190 0 22246 480 6 bottom_right_grid_pin_5_
port 13 nsew default input
rlabel metal2 s 23202 0 23258 480 6 bottom_right_grid_pin_7_
port 14 nsew default input
rlabel metal2 s 24214 0 24270 480 6 bottom_right_grid_pin_9_
port 15 nsew default input
rlabel metal3 s 0 14696 480 14816 6 chanx_left_in[0]
port 16 nsew default input
rlabel metal3 s 0 16056 480 16176 6 chanx_left_in[1]
port 17 nsew default input
rlabel metal3 s 0 17416 480 17536 6 chanx_left_in[2]
port 18 nsew default input
rlabel metal3 s 0 18776 480 18896 6 chanx_left_in[3]
port 19 nsew default input
rlabel metal3 s 0 20272 480 20392 6 chanx_left_in[4]
port 20 nsew default input
rlabel metal3 s 0 21632 480 21752 6 chanx_left_in[5]
port 21 nsew default input
rlabel metal3 s 0 22992 480 23112 6 chanx_left_in[6]
port 22 nsew default input
rlabel metal3 s 0 24488 480 24608 6 chanx_left_in[7]
port 23 nsew default input
rlabel metal3 s 0 25848 480 25968 6 chanx_left_in[8]
port 24 nsew default input
rlabel metal3 s 0 2048 480 2168 6 chanx_left_out[0]
port 25 nsew default tristate
rlabel metal3 s 0 3408 480 3528 6 chanx_left_out[1]
port 26 nsew default tristate
rlabel metal3 s 0 4768 480 4888 6 chanx_left_out[2]
port 27 nsew default tristate
rlabel metal3 s 0 6264 480 6384 6 chanx_left_out[3]
port 28 nsew default tristate
rlabel metal3 s 0 7624 480 7744 6 chanx_left_out[4]
port 29 nsew default tristate
rlabel metal3 s 0 8984 480 9104 6 chanx_left_out[5]
port 30 nsew default tristate
rlabel metal3 s 0 10480 480 10600 6 chanx_left_out[6]
port 31 nsew default tristate
rlabel metal3 s 0 11840 480 11960 6 chanx_left_out[7]
port 32 nsew default tristate
rlabel metal3 s 0 13200 480 13320 6 chanx_left_out[8]
port 33 nsew default tristate
rlabel metal2 s 1490 0 1546 480 6 chany_bottom_in[0]
port 34 nsew default input
rlabel metal2 s 2502 0 2558 480 6 chany_bottom_in[1]
port 35 nsew default input
rlabel metal2 s 3514 0 3570 480 6 chany_bottom_in[2]
port 36 nsew default input
rlabel metal2 s 4618 0 4674 480 6 chany_bottom_in[3]
port 37 nsew default input
rlabel metal2 s 5630 0 5686 480 6 chany_bottom_in[4]
port 38 nsew default input
rlabel metal2 s 6642 0 6698 480 6 chany_bottom_in[5]
port 39 nsew default input
rlabel metal2 s 7654 0 7710 480 6 chany_bottom_in[6]
port 40 nsew default input
rlabel metal2 s 8758 0 8814 480 6 chany_bottom_in[7]
port 41 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[8]
port 42 nsew default input
rlabel metal2 s 10782 0 10838 480 6 chany_bottom_out[0]
port 43 nsew default tristate
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_out[1]
port 44 nsew default tristate
rlabel metal2 s 12898 0 12954 480 6 chany_bottom_out[2]
port 45 nsew default tristate
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_out[3]
port 46 nsew default tristate
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_out[4]
port 47 nsew default tristate
rlabel metal2 s 15934 0 15990 480 6 chany_bottom_out[5]
port 48 nsew default tristate
rlabel metal2 s 17038 0 17094 480 6 chany_bottom_out[6]
port 49 nsew default tristate
rlabel metal2 s 18050 0 18106 480 6 chany_bottom_out[7]
port 50 nsew default tristate
rlabel metal2 s 19062 0 19118 480 6 chany_bottom_out[8]
port 51 nsew default tristate
rlabel metal2 s 1490 27520 1546 28000 6 chany_top_in[0]
port 52 nsew default input
rlabel metal2 s 2502 27520 2558 28000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 3514 27520 3570 28000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 4618 27520 4674 28000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 5630 27520 5686 28000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 6642 27520 6698 28000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 7654 27520 7710 28000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 8758 27520 8814 28000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 9770 27520 9826 28000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 10782 27520 10838 28000 6 chany_top_out[0]
port 61 nsew default tristate
rlabel metal2 s 11794 27520 11850 28000 6 chany_top_out[1]
port 62 nsew default tristate
rlabel metal2 s 12898 27520 12954 28000 6 chany_top_out[2]
port 63 nsew default tristate
rlabel metal2 s 13910 27520 13966 28000 6 chany_top_out[3]
port 64 nsew default tristate
rlabel metal2 s 14922 27520 14978 28000 6 chany_top_out[4]
port 65 nsew default tristate
rlabel metal2 s 15934 27520 15990 28000 6 chany_top_out[5]
port 66 nsew default tristate
rlabel metal2 s 17038 27520 17094 28000 6 chany_top_out[6]
port 67 nsew default tristate
rlabel metal2 s 18050 27520 18106 28000 6 chany_top_out[7]
port 68 nsew default tristate
rlabel metal2 s 19062 27520 19118 28000 6 chany_top_out[8]
port 69 nsew default tristate
rlabel metal3 s 27520 26392 28000 26512 6 data_in
port 70 nsew default input
rlabel metal3 s 27520 1504 28000 1624 6 enable
port 71 nsew default input
rlabel metal3 s 0 688 480 808 6 left_bottom_grid_pin_12_
port 72 nsew default input
rlabel metal3 s 0 27208 480 27328 6 left_top_grid_pin_10_
port 73 nsew default input
rlabel metal2 s 478 27520 534 28000 6 top_left_grid_pin_13_
port 74 nsew default input
rlabel metal2 s 25318 27520 25374 28000 6 top_right_grid_pin_11_
port 75 nsew default input
rlabel metal2 s 26330 27520 26386 28000 6 top_right_grid_pin_13_
port 76 nsew default input
rlabel metal2 s 27342 27520 27398 28000 6 top_right_grid_pin_15_
port 77 nsew default input
rlabel metal2 s 20074 27520 20130 28000 6 top_right_grid_pin_1_
port 78 nsew default input
rlabel metal2 s 21178 27520 21234 28000 6 top_right_grid_pin_3_
port 79 nsew default input
rlabel metal2 s 22190 27520 22246 28000 6 top_right_grid_pin_5_
port 80 nsew default input
rlabel metal2 s 23202 27520 23258 28000 6 top_right_grid_pin_7_
port 81 nsew default input
rlabel metal2 s 24214 27520 24270 28000 6 top_right_grid_pin_9_
port 82 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 83 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 84 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
