magic
tech sky130A
magscale 1 2
timestamp 1605120744
<< locali >>
rect 14933 9707 14967 19261
rect 14933 595 14967 3349
<< viali >>
rect 1593 31977 1627 32011
rect 5365 31977 5399 32011
rect 1409 31841 1443 31875
rect 4077 31841 4111 31875
rect 5181 31841 5215 31875
rect 4261 31637 4295 31671
rect 1593 31433 1627 31467
rect 8769 31433 8803 31467
rect 12633 31433 12667 31467
rect 1409 31229 1443 31263
rect 8585 31229 8619 31263
rect 12449 31229 12483 31263
rect 13001 31229 13035 31263
rect 2053 31093 2087 31127
rect 4169 31093 4203 31127
rect 5181 31093 5215 31127
rect 9229 31093 9263 31127
rect 9689 30685 9723 30719
rect 1685 30549 1719 30583
rect 9321 30549 9355 30583
rect 9873 30209 9907 30243
rect 9689 30141 9723 30175
rect 9781 30073 9815 30107
rect 9137 30005 9171 30039
rect 9321 30005 9355 30039
rect 9413 29801 9447 29835
rect 7553 29665 7587 29699
rect 7297 29597 7331 29631
rect 8677 29461 8711 29495
rect 2237 29257 2271 29291
rect 2421 29053 2455 29087
rect 2677 29053 2711 29087
rect 7297 28985 7331 29019
rect 7665 28985 7699 29019
rect 3801 28917 3835 28951
rect 2421 28441 2455 28475
rect 4537 27965 4571 27999
rect 4782 27897 4816 27931
rect 4445 27829 4479 27863
rect 5917 27829 5951 27863
rect 4629 27285 4663 27319
rect 1593 25993 1627 26027
rect 1409 25789 1443 25823
rect 1961 25653 1995 25687
rect 4077 25313 4111 25347
rect 4261 25177 4295 25211
rect 4077 24905 4111 24939
rect 6285 24361 6319 24395
rect 12081 24361 12115 24395
rect 6469 24225 6503 24259
rect 11897 24225 11931 24259
rect 6377 23477 6411 23511
rect 11989 23477 12023 23511
rect 10057 23273 10091 23307
rect 9505 23205 9539 23239
rect 10149 23069 10183 23103
rect 10241 23069 10275 23103
rect 9689 22933 9723 22967
rect 10425 22729 10459 22763
rect 10793 22729 10827 22763
rect 9413 22661 9447 22695
rect 9873 22593 9907 22627
rect 10057 22593 10091 22627
rect 7481 22457 7515 22491
rect 7573 22457 7607 22491
rect 8861 22389 8895 22423
rect 9781 22389 9815 22423
rect 10241 22185 10275 22219
rect 9965 22117 9999 22151
rect 6009 22049 6043 22083
rect 6101 21981 6135 22015
rect 6285 21981 6319 22015
rect 9413 21913 9447 21947
rect 5641 21845 5675 21879
rect 6009 21641 6043 21675
rect 6377 21641 6411 21675
rect 5733 21301 5767 21335
rect 7021 21097 7055 21131
rect 7481 20417 7515 20451
rect 7665 20417 7699 20451
rect 8769 20349 8803 20383
rect 9045 20349 9079 20383
rect 6653 20281 6687 20315
rect 7021 20213 7055 20247
rect 7389 20213 7423 20247
rect 8585 20213 8619 20247
rect 7113 20009 7147 20043
rect 12357 19873 12391 19907
rect 12541 19669 12575 19703
rect 12633 19329 12667 19363
rect 14933 19261 14967 19295
rect 4445 16745 4479 16779
rect 12909 16745 12943 16779
rect 11529 16609 11563 16643
rect 11785 16609 11819 16643
rect 11897 16201 11931 16235
rect 4997 16065 5031 16099
rect 4813 15997 4847 16031
rect 4353 15929 4387 15963
rect 4445 15861 4479 15895
rect 4905 15861 4939 15895
rect 11529 15861 11563 15895
rect 5641 15657 5675 15691
rect 7297 15657 7331 15691
rect 4537 15589 4571 15623
rect 5549 15521 5583 15555
rect 5733 15453 5767 15487
rect 5181 15317 5215 15351
rect 1593 15113 1627 15147
rect 2053 15113 2087 15147
rect 5549 15113 5583 15147
rect 5825 15113 5859 15147
rect 8953 15113 8987 15147
rect 3985 14977 4019 15011
rect 4997 14977 5031 15011
rect 7205 14977 7239 15011
rect 7941 14977 7975 15011
rect 9505 14977 9539 15011
rect 1409 14909 1443 14943
rect 4813 14909 4847 14943
rect 7665 14909 7699 14943
rect 9413 14909 9447 14943
rect 9761 14909 9795 14943
rect 4353 14841 4387 14875
rect 7757 14841 7791 14875
rect 4445 14773 4479 14807
rect 4905 14773 4939 14807
rect 7297 14773 7331 14807
rect 10885 14773 10919 14807
rect 5273 14569 5307 14603
rect 7297 14569 7331 14603
rect 8033 14569 8067 14603
rect 4537 14501 4571 14535
rect 7849 13889 7883 13923
rect 8493 13889 8527 13923
rect 2053 13821 2087 13855
rect 2605 13821 2639 13855
rect 8401 13753 8435 13787
rect 2237 13685 2271 13719
rect 7941 13685 7975 13719
rect 8309 13685 8343 13719
rect 7941 13481 7975 13515
rect 1409 12257 1443 12291
rect 1593 12189 1627 12223
rect 1593 11849 1627 11883
rect 1961 11169 1995 11203
rect 2145 11033 2179 11067
rect 2053 10761 2087 10795
rect 13093 10761 13127 10795
rect 12449 10557 12483 10591
rect 12633 10421 12667 10455
rect 14933 9673 14967 9707
rect 2881 9605 2915 9639
rect 2697 9469 2731 9503
rect 3341 9401 3375 9435
rect 10609 9129 10643 9163
rect 12541 9129 12575 9163
rect 10425 8993 10459 9027
rect 12357 8993 12391 9027
rect 12265 8381 12299 8415
rect 12449 8381 12483 8415
rect 10517 8313 10551 8347
rect 13093 8313 13127 8347
rect 12633 8245 12667 8279
rect 4905 8041 4939 8075
rect 4721 7905 4755 7939
rect 7481 7497 7515 7531
rect 6837 7293 6871 7327
rect 4813 7157 4847 7191
rect 7021 7157 7055 7191
rect 1593 6817 1627 6851
rect 6009 6817 6043 6851
rect 10425 6817 10459 6851
rect 6193 6681 6227 6715
rect 1777 6613 1811 6647
rect 10609 6613 10643 6647
rect 1593 6409 1627 6443
rect 8217 6409 8251 6443
rect 10517 6409 10551 6443
rect 11253 6409 11287 6443
rect 8861 6341 8895 6375
rect 4169 6205 4203 6239
rect 4813 6205 4847 6239
rect 7573 6205 7607 6239
rect 8677 6205 8711 6239
rect 10333 6205 10367 6239
rect 4353 6069 4387 6103
rect 6101 6069 6135 6103
rect 7757 6069 7791 6103
rect 9321 6069 9355 6103
rect 10977 6069 11011 6103
rect 1593 3689 1627 3723
rect 4721 3689 4755 3723
rect 1409 3553 1443 3587
rect 4537 3553 4571 3587
rect 14933 3349 14967 3383
rect 1685 3145 1719 3179
rect 2421 3145 2455 3179
rect 4629 3145 4663 3179
rect 5641 3145 5675 3179
rect 9965 3145 9999 3179
rect 10425 3145 10459 3179
rect 13093 3145 13127 3179
rect 2053 3077 2087 3111
rect 5181 3077 5215 3111
rect 11437 3077 11471 3111
rect 1869 2941 1903 2975
rect 4997 2941 5031 2975
rect 8677 2941 8711 2975
rect 9229 2941 9263 2975
rect 9781 2941 9815 2975
rect 11253 2941 11287 2975
rect 12449 2941 12483 2975
rect 11897 2873 11931 2907
rect 8861 2805 8895 2839
rect 12633 2805 12667 2839
rect 2329 2601 2363 2635
rect 3065 2601 3099 2635
rect 5825 2601 5859 2635
rect 7113 2601 7147 2635
rect 11621 2601 11655 2635
rect 13277 2601 13311 2635
rect 6193 2533 6227 2567
rect 1777 2465 1811 2499
rect 2881 2465 2915 2499
rect 4537 2465 4571 2499
rect 5089 2465 5123 2499
rect 5641 2465 5675 2499
rect 6929 2465 6963 2499
rect 8585 2465 8619 2499
rect 9781 2465 9815 2499
rect 10425 2465 10459 2499
rect 11437 2465 11471 2499
rect 12633 2465 12667 2499
rect 12817 2329 12851 2363
rect 1961 2261 1995 2295
rect 3525 2261 3559 2295
rect 4721 2261 4755 2295
rect 7573 2261 7607 2295
rect 8769 2261 8803 2295
rect 9229 2261 9263 2295
rect 9965 2261 9999 2295
rect 12081 2261 12115 2295
rect 14933 561 14967 595
<< metal1 >>
rect 1104 37562 14812 37584
rect 1104 37510 6315 37562
rect 6367 37510 6379 37562
rect 6431 37510 6443 37562
rect 6495 37510 6507 37562
rect 6559 37510 11648 37562
rect 11700 37510 11712 37562
rect 11764 37510 11776 37562
rect 11828 37510 11840 37562
rect 11892 37510 14812 37562
rect 1104 37488 14812 37510
rect 8386 37136 8392 37188
rect 8444 37176 8450 37188
rect 8938 37176 8944 37188
rect 8444 37148 8944 37176
rect 8444 37136 8450 37148
rect 8938 37136 8944 37148
rect 8996 37136 9002 37188
rect 1104 37018 14812 37040
rect 1104 36966 3648 37018
rect 3700 36966 3712 37018
rect 3764 36966 3776 37018
rect 3828 36966 3840 37018
rect 3892 36966 8982 37018
rect 9034 36966 9046 37018
rect 9098 36966 9110 37018
rect 9162 36966 9174 37018
rect 9226 36966 14315 37018
rect 14367 36966 14379 37018
rect 14431 36966 14443 37018
rect 14495 36966 14507 37018
rect 14559 36966 14812 37018
rect 1104 36944 14812 36966
rect 1104 36474 14812 36496
rect 1104 36422 6315 36474
rect 6367 36422 6379 36474
rect 6431 36422 6443 36474
rect 6495 36422 6507 36474
rect 6559 36422 11648 36474
rect 11700 36422 11712 36474
rect 11764 36422 11776 36474
rect 11828 36422 11840 36474
rect 11892 36422 14812 36474
rect 1104 36400 14812 36422
rect 1104 35930 14812 35952
rect 1104 35878 3648 35930
rect 3700 35878 3712 35930
rect 3764 35878 3776 35930
rect 3828 35878 3840 35930
rect 3892 35878 8982 35930
rect 9034 35878 9046 35930
rect 9098 35878 9110 35930
rect 9162 35878 9174 35930
rect 9226 35878 14315 35930
rect 14367 35878 14379 35930
rect 14431 35878 14443 35930
rect 14495 35878 14507 35930
rect 14559 35878 14812 35930
rect 1104 35856 14812 35878
rect 4522 35708 4528 35760
rect 4580 35748 4586 35760
rect 5442 35748 5448 35760
rect 4580 35720 5448 35748
rect 4580 35708 4586 35720
rect 5442 35708 5448 35720
rect 5500 35708 5506 35760
rect 5718 35708 5724 35760
rect 5776 35748 5782 35760
rect 6730 35748 6736 35760
rect 5776 35720 6736 35748
rect 5776 35708 5782 35720
rect 6730 35708 6736 35720
rect 6788 35708 6794 35760
rect 6178 35640 6184 35692
rect 6236 35680 6242 35692
rect 6638 35680 6644 35692
rect 6236 35652 6644 35680
rect 6236 35640 6242 35652
rect 6638 35640 6644 35652
rect 6696 35640 6702 35692
rect 7190 35640 7196 35692
rect 7248 35680 7254 35692
rect 8202 35680 8208 35692
rect 7248 35652 8208 35680
rect 7248 35640 7254 35652
rect 8202 35640 8208 35652
rect 8260 35640 8266 35692
rect 5074 35572 5080 35624
rect 5132 35612 5138 35624
rect 5350 35612 5356 35624
rect 5132 35584 5356 35612
rect 5132 35572 5138 35584
rect 5350 35572 5356 35584
rect 5408 35572 5414 35624
rect 1104 35386 14812 35408
rect 1104 35334 6315 35386
rect 6367 35334 6379 35386
rect 6431 35334 6443 35386
rect 6495 35334 6507 35386
rect 6559 35334 11648 35386
rect 11700 35334 11712 35386
rect 11764 35334 11776 35386
rect 11828 35334 11840 35386
rect 11892 35334 14812 35386
rect 1104 35312 14812 35334
rect 7374 35232 7380 35284
rect 7432 35272 7438 35284
rect 8202 35272 8208 35284
rect 7432 35244 8208 35272
rect 7432 35232 7438 35244
rect 8202 35232 8208 35244
rect 8260 35232 8266 35284
rect 6914 35096 6920 35148
rect 6972 35136 6978 35148
rect 8018 35136 8024 35148
rect 6972 35108 8024 35136
rect 6972 35096 6978 35108
rect 8018 35096 8024 35108
rect 8076 35096 8082 35148
rect 1394 34892 1400 34944
rect 1452 34932 1458 34944
rect 2498 34932 2504 34944
rect 1452 34904 2504 34932
rect 1452 34892 1458 34904
rect 2498 34892 2504 34904
rect 2556 34892 2562 34944
rect 1104 34842 14812 34864
rect 1104 34790 3648 34842
rect 3700 34790 3712 34842
rect 3764 34790 3776 34842
rect 3828 34790 3840 34842
rect 3892 34790 8982 34842
rect 9034 34790 9046 34842
rect 9098 34790 9110 34842
rect 9162 34790 9174 34842
rect 9226 34790 14315 34842
rect 14367 34790 14379 34842
rect 14431 34790 14443 34842
rect 14495 34790 14507 34842
rect 14559 34790 14812 34842
rect 1104 34768 14812 34790
rect 198 34552 204 34604
rect 256 34592 262 34604
rect 1302 34592 1308 34604
rect 256 34564 1308 34592
rect 256 34552 262 34564
rect 1302 34552 1308 34564
rect 1360 34552 1366 34604
rect 566 34484 572 34536
rect 624 34524 630 34536
rect 1118 34524 1124 34536
rect 624 34496 1124 34524
rect 624 34484 630 34496
rect 1118 34484 1124 34496
rect 1176 34484 1182 34536
rect 2130 34484 2136 34536
rect 2188 34524 2194 34536
rect 2590 34524 2596 34536
rect 2188 34496 2596 34524
rect 2188 34484 2194 34496
rect 2590 34484 2596 34496
rect 2648 34484 2654 34536
rect 1104 34298 14812 34320
rect 1104 34246 6315 34298
rect 6367 34246 6379 34298
rect 6431 34246 6443 34298
rect 6495 34246 6507 34298
rect 6559 34246 11648 34298
rect 11700 34246 11712 34298
rect 11764 34246 11776 34298
rect 11828 34246 11840 34298
rect 11892 34246 14812 34298
rect 1104 34224 14812 34246
rect 1104 33754 14812 33776
rect 1104 33702 3648 33754
rect 3700 33702 3712 33754
rect 3764 33702 3776 33754
rect 3828 33702 3840 33754
rect 3892 33702 8982 33754
rect 9034 33702 9046 33754
rect 9098 33702 9110 33754
rect 9162 33702 9174 33754
rect 9226 33702 14315 33754
rect 14367 33702 14379 33754
rect 14431 33702 14443 33754
rect 14495 33702 14507 33754
rect 14559 33702 14812 33754
rect 1104 33680 14812 33702
rect 1104 33210 14812 33232
rect 1104 33158 6315 33210
rect 6367 33158 6379 33210
rect 6431 33158 6443 33210
rect 6495 33158 6507 33210
rect 6559 33158 11648 33210
rect 11700 33158 11712 33210
rect 11764 33158 11776 33210
rect 11828 33158 11840 33210
rect 11892 33158 14812 33210
rect 1104 33136 14812 33158
rect 1104 32666 14812 32688
rect 1104 32614 3648 32666
rect 3700 32614 3712 32666
rect 3764 32614 3776 32666
rect 3828 32614 3840 32666
rect 3892 32614 8982 32666
rect 9034 32614 9046 32666
rect 9098 32614 9110 32666
rect 9162 32614 9174 32666
rect 9226 32614 14315 32666
rect 14367 32614 14379 32666
rect 14431 32614 14443 32666
rect 14495 32614 14507 32666
rect 14559 32614 14812 32666
rect 1104 32592 14812 32614
rect 1104 32122 14812 32144
rect 1104 32070 6315 32122
rect 6367 32070 6379 32122
rect 6431 32070 6443 32122
rect 6495 32070 6507 32122
rect 6559 32070 11648 32122
rect 11700 32070 11712 32122
rect 11764 32070 11776 32122
rect 11828 32070 11840 32122
rect 11892 32070 14812 32122
rect 1104 32048 14812 32070
rect 1394 31968 1400 32020
rect 1452 32008 1458 32020
rect 1581 32011 1639 32017
rect 1581 32008 1593 32011
rect 1452 31980 1593 32008
rect 1452 31968 1458 31980
rect 1581 31977 1593 31980
rect 1627 31977 1639 32011
rect 1581 31971 1639 31977
rect 4154 31968 4160 32020
rect 4212 32008 4218 32020
rect 5353 32011 5411 32017
rect 5353 32008 5365 32011
rect 4212 31980 5365 32008
rect 4212 31968 4218 31980
rect 5353 31977 5365 31980
rect 5399 31977 5411 32011
rect 5353 31971 5411 31977
rect 1397 31875 1455 31881
rect 1397 31841 1409 31875
rect 1443 31872 1455 31875
rect 2222 31872 2228 31884
rect 1443 31844 2228 31872
rect 1443 31841 1455 31844
rect 1397 31835 1455 31841
rect 2222 31832 2228 31844
rect 2280 31832 2286 31884
rect 4062 31872 4068 31884
rect 4023 31844 4068 31872
rect 4062 31832 4068 31844
rect 4120 31832 4126 31884
rect 5166 31872 5172 31884
rect 5127 31844 5172 31872
rect 5166 31832 5172 31844
rect 5224 31832 5230 31884
rect 1762 31628 1768 31680
rect 1820 31668 1826 31680
rect 4249 31671 4307 31677
rect 4249 31668 4261 31671
rect 1820 31640 4261 31668
rect 1820 31628 1826 31640
rect 4249 31637 4261 31640
rect 4295 31637 4307 31671
rect 4249 31631 4307 31637
rect 1104 31578 14812 31600
rect 1104 31526 3648 31578
rect 3700 31526 3712 31578
rect 3764 31526 3776 31578
rect 3828 31526 3840 31578
rect 3892 31526 8982 31578
rect 9034 31526 9046 31578
rect 9098 31526 9110 31578
rect 9162 31526 9174 31578
rect 9226 31526 14315 31578
rect 14367 31526 14379 31578
rect 14431 31526 14443 31578
rect 14495 31526 14507 31578
rect 14559 31526 14812 31578
rect 1104 31504 14812 31526
rect 934 31424 940 31476
rect 992 31464 998 31476
rect 1581 31467 1639 31473
rect 1581 31464 1593 31467
rect 992 31436 1593 31464
rect 992 31424 998 31436
rect 1581 31433 1593 31436
rect 1627 31433 1639 31467
rect 8754 31464 8760 31476
rect 8715 31436 8760 31464
rect 1581 31427 1639 31433
rect 8754 31424 8760 31436
rect 8812 31424 8818 31476
rect 12434 31424 12440 31476
rect 12492 31464 12498 31476
rect 12621 31467 12679 31473
rect 12621 31464 12633 31467
rect 12492 31436 12633 31464
rect 12492 31424 12498 31436
rect 12621 31433 12633 31436
rect 12667 31433 12679 31467
rect 12621 31427 12679 31433
rect 1397 31263 1455 31269
rect 1397 31229 1409 31263
rect 1443 31260 1455 31263
rect 1670 31260 1676 31272
rect 1443 31232 1676 31260
rect 1443 31229 1455 31232
rect 1397 31223 1455 31229
rect 1670 31220 1676 31232
rect 1728 31220 1734 31272
rect 8573 31263 8631 31269
rect 8573 31229 8585 31263
rect 8619 31260 8631 31263
rect 8619 31232 9260 31260
rect 8619 31229 8631 31232
rect 8573 31223 8631 31229
rect 2041 31127 2099 31133
rect 2041 31093 2053 31127
rect 2087 31124 2099 31127
rect 2222 31124 2228 31136
rect 2087 31096 2228 31124
rect 2087 31093 2099 31096
rect 2041 31087 2099 31093
rect 2222 31084 2228 31096
rect 2280 31084 2286 31136
rect 4154 31124 4160 31136
rect 4115 31096 4160 31124
rect 4154 31084 4160 31096
rect 4212 31084 4218 31136
rect 5166 31124 5172 31136
rect 5127 31096 5172 31124
rect 5166 31084 5172 31096
rect 5224 31084 5230 31136
rect 9232 31133 9260 31232
rect 12434 31220 12440 31272
rect 12492 31260 12498 31272
rect 12989 31263 13047 31269
rect 12989 31260 13001 31263
rect 12492 31232 13001 31260
rect 12492 31220 12498 31232
rect 12989 31229 13001 31232
rect 13035 31229 13047 31263
rect 12989 31223 13047 31229
rect 9217 31127 9275 31133
rect 9217 31093 9229 31127
rect 9263 31124 9275 31127
rect 9398 31124 9404 31136
rect 9263 31096 9404 31124
rect 9263 31093 9275 31096
rect 9217 31087 9275 31093
rect 9398 31084 9404 31096
rect 9456 31084 9462 31136
rect 1104 31034 14812 31056
rect 1104 30982 6315 31034
rect 6367 30982 6379 31034
rect 6431 30982 6443 31034
rect 6495 30982 6507 31034
rect 6559 30982 11648 31034
rect 11700 30982 11712 31034
rect 11764 30982 11776 31034
rect 11828 30982 11840 31034
rect 11892 30982 14812 31034
rect 1104 30960 14812 30982
rect 9674 30716 9680 30728
rect 9635 30688 9680 30716
rect 9674 30676 9680 30688
rect 9732 30676 9738 30728
rect 1670 30580 1676 30592
rect 1631 30552 1676 30580
rect 1670 30540 1676 30552
rect 1728 30540 1734 30592
rect 9306 30580 9312 30592
rect 9267 30552 9312 30580
rect 9306 30540 9312 30552
rect 9364 30540 9370 30592
rect 1104 30490 14812 30512
rect 1104 30438 3648 30490
rect 3700 30438 3712 30490
rect 3764 30438 3776 30490
rect 3828 30438 3840 30490
rect 3892 30438 8982 30490
rect 9034 30438 9046 30490
rect 9098 30438 9110 30490
rect 9162 30438 9174 30490
rect 9226 30438 14315 30490
rect 14367 30438 14379 30490
rect 14431 30438 14443 30490
rect 14495 30438 14507 30490
rect 14559 30438 14812 30490
rect 1104 30416 14812 30438
rect 9766 30336 9772 30388
rect 9824 30376 9830 30388
rect 9950 30376 9956 30388
rect 9824 30348 9956 30376
rect 9824 30336 9830 30348
rect 9950 30336 9956 30348
rect 10008 30336 10014 30388
rect 9306 30200 9312 30252
rect 9364 30240 9370 30252
rect 9861 30243 9919 30249
rect 9861 30240 9873 30243
rect 9364 30212 9873 30240
rect 9364 30200 9370 30212
rect 9861 30209 9873 30212
rect 9907 30209 9919 30243
rect 9861 30203 9919 30209
rect 9674 30172 9680 30184
rect 9635 30144 9680 30172
rect 9674 30132 9680 30144
rect 9732 30132 9738 30184
rect 9766 30104 9772 30116
rect 9140 30076 9772 30104
rect 8478 29996 8484 30048
rect 8536 30036 8542 30048
rect 9140 30045 9168 30076
rect 9766 30064 9772 30076
rect 9824 30064 9830 30116
rect 9125 30039 9183 30045
rect 9125 30036 9137 30039
rect 8536 30008 9137 30036
rect 8536 29996 8542 30008
rect 9125 30005 9137 30008
rect 9171 30005 9183 30039
rect 9125 29999 9183 30005
rect 9309 30039 9367 30045
rect 9309 30005 9321 30039
rect 9355 30036 9367 30039
rect 9582 30036 9588 30048
rect 9355 30008 9588 30036
rect 9355 30005 9367 30008
rect 9309 29999 9367 30005
rect 9582 29996 9588 30008
rect 9640 29996 9646 30048
rect 1104 29946 14812 29968
rect 1104 29894 6315 29946
rect 6367 29894 6379 29946
rect 6431 29894 6443 29946
rect 6495 29894 6507 29946
rect 6559 29894 11648 29946
rect 11700 29894 11712 29946
rect 11764 29894 11776 29946
rect 11828 29894 11840 29946
rect 11892 29894 14812 29946
rect 1104 29872 14812 29894
rect 9401 29835 9459 29841
rect 9401 29801 9413 29835
rect 9447 29832 9459 29835
rect 9674 29832 9680 29844
rect 9447 29804 9680 29832
rect 9447 29801 9459 29804
rect 9401 29795 9459 29801
rect 9674 29792 9680 29804
rect 9732 29792 9738 29844
rect 7374 29656 7380 29708
rect 7432 29696 7438 29708
rect 7541 29699 7599 29705
rect 7541 29696 7553 29699
rect 7432 29668 7553 29696
rect 7432 29656 7438 29668
rect 7541 29665 7553 29668
rect 7587 29696 7599 29699
rect 9306 29696 9312 29708
rect 7587 29668 9312 29696
rect 7587 29665 7599 29668
rect 7541 29659 7599 29665
rect 9306 29656 9312 29668
rect 9364 29656 9370 29708
rect 7285 29631 7343 29637
rect 7285 29597 7297 29631
rect 7331 29597 7343 29631
rect 7285 29591 7343 29597
rect 7300 29492 7328 29591
rect 7650 29492 7656 29504
rect 7300 29464 7656 29492
rect 7650 29452 7656 29464
rect 7708 29452 7714 29504
rect 8665 29495 8723 29501
rect 8665 29461 8677 29495
rect 8711 29492 8723 29495
rect 9490 29492 9496 29504
rect 8711 29464 9496 29492
rect 8711 29461 8723 29464
rect 8665 29455 8723 29461
rect 9490 29452 9496 29464
rect 9548 29452 9554 29504
rect 1104 29402 14812 29424
rect 1104 29350 3648 29402
rect 3700 29350 3712 29402
rect 3764 29350 3776 29402
rect 3828 29350 3840 29402
rect 3892 29350 8982 29402
rect 9034 29350 9046 29402
rect 9098 29350 9110 29402
rect 9162 29350 9174 29402
rect 9226 29350 14315 29402
rect 14367 29350 14379 29402
rect 14431 29350 14443 29402
rect 14495 29350 14507 29402
rect 14559 29350 14812 29402
rect 1104 29328 14812 29350
rect 1946 29248 1952 29300
rect 2004 29288 2010 29300
rect 2225 29291 2283 29297
rect 2225 29288 2237 29291
rect 2004 29260 2237 29288
rect 2004 29248 2010 29260
rect 2225 29257 2237 29260
rect 2271 29257 2283 29291
rect 2225 29251 2283 29257
rect 2240 29152 2268 29251
rect 2240 29124 2544 29152
rect 2406 29084 2412 29096
rect 2367 29056 2412 29084
rect 2406 29044 2412 29056
rect 2464 29044 2470 29096
rect 2516 29084 2544 29124
rect 2665 29087 2723 29093
rect 2665 29084 2677 29087
rect 2516 29056 2677 29084
rect 2665 29053 2677 29056
rect 2711 29053 2723 29087
rect 2665 29047 2723 29053
rect 7285 29019 7343 29025
rect 7285 29016 7297 29019
rect 6840 28988 7297 29016
rect 3789 28951 3847 28957
rect 3789 28917 3801 28951
rect 3835 28948 3847 28951
rect 4430 28948 4436 28960
rect 3835 28920 4436 28948
rect 3835 28917 3847 28920
rect 3789 28911 3847 28917
rect 4430 28908 4436 28920
rect 4488 28908 4494 28960
rect 5718 28908 5724 28960
rect 5776 28948 5782 28960
rect 6840 28948 6868 28988
rect 7285 28985 7297 28988
rect 7331 29016 7343 29019
rect 7374 29016 7380 29028
rect 7331 28988 7380 29016
rect 7331 28985 7343 28988
rect 7285 28979 7343 28985
rect 7374 28976 7380 28988
rect 7432 28976 7438 29028
rect 7650 29016 7656 29028
rect 7611 28988 7656 29016
rect 7650 28976 7656 28988
rect 7708 28976 7714 29028
rect 5776 28920 6868 28948
rect 5776 28908 5782 28920
rect 10318 28908 10324 28960
rect 10376 28948 10382 28960
rect 10594 28948 10600 28960
rect 10376 28920 10600 28948
rect 10376 28908 10382 28920
rect 10594 28908 10600 28920
rect 10652 28908 10658 28960
rect 12710 28908 12716 28960
rect 12768 28948 12774 28960
rect 12894 28948 12900 28960
rect 12768 28920 12900 28948
rect 12768 28908 12774 28920
rect 12894 28908 12900 28920
rect 12952 28908 12958 28960
rect 1104 28858 14812 28880
rect 1104 28806 6315 28858
rect 6367 28806 6379 28858
rect 6431 28806 6443 28858
rect 6495 28806 6507 28858
rect 6559 28806 11648 28858
rect 11700 28806 11712 28858
rect 11764 28806 11776 28858
rect 11828 28806 11840 28858
rect 11892 28806 14812 28858
rect 1104 28784 14812 28806
rect 2406 28472 2412 28484
rect 2367 28444 2412 28472
rect 2406 28432 2412 28444
rect 2464 28432 2470 28484
rect 1104 28314 14812 28336
rect 1104 28262 3648 28314
rect 3700 28262 3712 28314
rect 3764 28262 3776 28314
rect 3828 28262 3840 28314
rect 3892 28262 8982 28314
rect 9034 28262 9046 28314
rect 9098 28262 9110 28314
rect 9162 28262 9174 28314
rect 9226 28262 14315 28314
rect 14367 28262 14379 28314
rect 14431 28262 14443 28314
rect 14495 28262 14507 28314
rect 14559 28262 14812 28314
rect 1104 28240 14812 28262
rect 4522 27996 4528 28008
rect 4483 27968 4528 27996
rect 4522 27956 4528 27968
rect 4580 27956 4586 28008
rect 4770 27931 4828 27937
rect 4770 27928 4782 27931
rect 4448 27900 4782 27928
rect 4448 27872 4476 27900
rect 4770 27897 4782 27900
rect 4816 27897 4828 27931
rect 4770 27891 4828 27897
rect 4430 27860 4436 27872
rect 4391 27832 4436 27860
rect 4430 27820 4436 27832
rect 4488 27820 4494 27872
rect 5718 27820 5724 27872
rect 5776 27860 5782 27872
rect 5905 27863 5963 27869
rect 5905 27860 5917 27863
rect 5776 27832 5917 27860
rect 5776 27820 5782 27832
rect 5905 27829 5917 27832
rect 5951 27829 5963 27863
rect 5905 27823 5963 27829
rect 1104 27770 14812 27792
rect 1104 27718 6315 27770
rect 6367 27718 6379 27770
rect 6431 27718 6443 27770
rect 6495 27718 6507 27770
rect 6559 27718 11648 27770
rect 11700 27718 11712 27770
rect 11764 27718 11776 27770
rect 11828 27718 11840 27770
rect 11892 27718 14812 27770
rect 1104 27696 14812 27718
rect 4338 27548 4344 27600
rect 4396 27588 4402 27600
rect 4614 27588 4620 27600
rect 4396 27560 4620 27588
rect 4396 27548 4402 27560
rect 4614 27548 4620 27560
rect 4672 27548 4678 27600
rect 4522 27276 4528 27328
rect 4580 27316 4586 27328
rect 4617 27319 4675 27325
rect 4617 27316 4629 27319
rect 4580 27288 4629 27316
rect 4580 27276 4586 27288
rect 4617 27285 4629 27288
rect 4663 27316 4675 27319
rect 5350 27316 5356 27328
rect 4663 27288 5356 27316
rect 4663 27285 4675 27288
rect 4617 27279 4675 27285
rect 5350 27276 5356 27288
rect 5408 27276 5414 27328
rect 1104 27226 14812 27248
rect 1104 27174 3648 27226
rect 3700 27174 3712 27226
rect 3764 27174 3776 27226
rect 3828 27174 3840 27226
rect 3892 27174 8982 27226
rect 9034 27174 9046 27226
rect 9098 27174 9110 27226
rect 9162 27174 9174 27226
rect 9226 27174 14315 27226
rect 14367 27174 14379 27226
rect 14431 27174 14443 27226
rect 14495 27174 14507 27226
rect 14559 27174 14812 27226
rect 1104 27152 14812 27174
rect 14090 27004 14096 27056
rect 14148 27044 14154 27056
rect 14826 27044 14832 27056
rect 14148 27016 14832 27044
rect 14148 27004 14154 27016
rect 14826 27004 14832 27016
rect 14884 27004 14890 27056
rect 12526 26936 12532 26988
rect 12584 26976 12590 26988
rect 13170 26976 13176 26988
rect 12584 26948 13176 26976
rect 12584 26936 12590 26948
rect 13170 26936 13176 26948
rect 13228 26936 13234 26988
rect 13906 26936 13912 26988
rect 13964 26976 13970 26988
rect 15378 26976 15384 26988
rect 13964 26948 15384 26976
rect 13964 26936 13970 26948
rect 15378 26936 15384 26948
rect 15436 26936 15442 26988
rect 8570 26868 8576 26920
rect 8628 26908 8634 26920
rect 9306 26908 9312 26920
rect 8628 26880 9312 26908
rect 8628 26868 8634 26880
rect 9306 26868 9312 26880
rect 9364 26868 9370 26920
rect 12802 26868 12808 26920
rect 12860 26908 12866 26920
rect 13722 26908 13728 26920
rect 12860 26880 13728 26908
rect 12860 26868 12866 26880
rect 13722 26868 13728 26880
rect 13780 26868 13786 26920
rect 13998 26868 14004 26920
rect 14056 26908 14062 26920
rect 14918 26908 14924 26920
rect 14056 26880 14924 26908
rect 14056 26868 14062 26880
rect 14918 26868 14924 26880
rect 14976 26868 14982 26920
rect 14090 26732 14096 26784
rect 14148 26772 14154 26784
rect 15746 26772 15752 26784
rect 14148 26744 15752 26772
rect 14148 26732 14154 26744
rect 15746 26732 15752 26744
rect 15804 26732 15810 26784
rect 1104 26682 14812 26704
rect 1104 26630 6315 26682
rect 6367 26630 6379 26682
rect 6431 26630 6443 26682
rect 6495 26630 6507 26682
rect 6559 26630 11648 26682
rect 11700 26630 11712 26682
rect 11764 26630 11776 26682
rect 11828 26630 11840 26682
rect 11892 26630 14812 26682
rect 1104 26608 14812 26630
rect 1104 26138 14812 26160
rect 1104 26086 3648 26138
rect 3700 26086 3712 26138
rect 3764 26086 3776 26138
rect 3828 26086 3840 26138
rect 3892 26086 8982 26138
rect 9034 26086 9046 26138
rect 9098 26086 9110 26138
rect 9162 26086 9174 26138
rect 9226 26086 14315 26138
rect 14367 26086 14379 26138
rect 14431 26086 14443 26138
rect 14495 26086 14507 26138
rect 14559 26086 14812 26138
rect 1104 26064 14812 26086
rect 1578 26024 1584 26036
rect 1539 25996 1584 26024
rect 1578 25984 1584 25996
rect 1636 25984 1642 26036
rect 1397 25823 1455 25829
rect 1397 25789 1409 25823
rect 1443 25820 1455 25823
rect 1443 25792 1808 25820
rect 1443 25789 1455 25792
rect 1397 25783 1455 25789
rect 1780 25696 1808 25792
rect 1762 25644 1768 25696
rect 1820 25684 1826 25696
rect 1949 25687 2007 25693
rect 1949 25684 1961 25687
rect 1820 25656 1961 25684
rect 1820 25644 1826 25656
rect 1949 25653 1961 25656
rect 1995 25653 2007 25687
rect 1949 25647 2007 25653
rect 1104 25594 14812 25616
rect 1104 25542 6315 25594
rect 6367 25542 6379 25594
rect 6431 25542 6443 25594
rect 6495 25542 6507 25594
rect 6559 25542 11648 25594
rect 11700 25542 11712 25594
rect 11764 25542 11776 25594
rect 11828 25542 11840 25594
rect 11892 25542 14812 25594
rect 1104 25520 14812 25542
rect 4062 25344 4068 25356
rect 4023 25316 4068 25344
rect 4062 25304 4068 25316
rect 4120 25304 4126 25356
rect 4246 25208 4252 25220
rect 4207 25180 4252 25208
rect 4246 25168 4252 25180
rect 4304 25168 4310 25220
rect 1104 25050 14812 25072
rect 1104 24998 3648 25050
rect 3700 24998 3712 25050
rect 3764 24998 3776 25050
rect 3828 24998 3840 25050
rect 3892 24998 8982 25050
rect 9034 24998 9046 25050
rect 9098 24998 9110 25050
rect 9162 24998 9174 25050
rect 9226 24998 14315 25050
rect 14367 24998 14379 25050
rect 14431 24998 14443 25050
rect 14495 24998 14507 25050
rect 14559 24998 14812 25050
rect 1104 24976 14812 24998
rect 4062 24936 4068 24948
rect 4023 24908 4068 24936
rect 4062 24896 4068 24908
rect 4120 24896 4126 24948
rect 1104 24506 14812 24528
rect 1104 24454 6315 24506
rect 6367 24454 6379 24506
rect 6431 24454 6443 24506
rect 6495 24454 6507 24506
rect 6559 24454 11648 24506
rect 11700 24454 11712 24506
rect 11764 24454 11776 24506
rect 11828 24454 11840 24506
rect 11892 24454 14812 24506
rect 1104 24432 14812 24454
rect 5350 24352 5356 24404
rect 5408 24392 5414 24404
rect 6273 24395 6331 24401
rect 6273 24392 6285 24395
rect 5408 24364 6285 24392
rect 5408 24352 5414 24364
rect 6273 24361 6285 24364
rect 6319 24361 6331 24395
rect 12066 24392 12072 24404
rect 12027 24364 12072 24392
rect 6273 24355 6331 24361
rect 12066 24352 12072 24364
rect 12124 24352 12130 24404
rect 6457 24259 6515 24265
rect 6457 24225 6469 24259
rect 6503 24256 6515 24259
rect 6822 24256 6828 24268
rect 6503 24228 6828 24256
rect 6503 24225 6515 24228
rect 6457 24219 6515 24225
rect 6822 24216 6828 24228
rect 6880 24216 6886 24268
rect 11885 24259 11943 24265
rect 11885 24225 11897 24259
rect 11931 24256 11943 24259
rect 12066 24256 12072 24268
rect 11931 24228 12072 24256
rect 11931 24225 11943 24228
rect 11885 24219 11943 24225
rect 12066 24216 12072 24228
rect 12124 24216 12130 24268
rect 1104 23962 14812 23984
rect 1104 23910 3648 23962
rect 3700 23910 3712 23962
rect 3764 23910 3776 23962
rect 3828 23910 3840 23962
rect 3892 23910 8982 23962
rect 9034 23910 9046 23962
rect 9098 23910 9110 23962
rect 9162 23910 9174 23962
rect 9226 23910 14315 23962
rect 14367 23910 14379 23962
rect 14431 23910 14443 23962
rect 14495 23910 14507 23962
rect 14559 23910 14812 23962
rect 1104 23888 14812 23910
rect 6365 23511 6423 23517
rect 6365 23477 6377 23511
rect 6411 23508 6423 23511
rect 6822 23508 6828 23520
rect 6411 23480 6828 23508
rect 6411 23477 6423 23480
rect 6365 23471 6423 23477
rect 6822 23468 6828 23480
rect 6880 23468 6886 23520
rect 11977 23511 12035 23517
rect 11977 23477 11989 23511
rect 12023 23508 12035 23511
rect 12066 23508 12072 23520
rect 12023 23480 12072 23508
rect 12023 23477 12035 23480
rect 11977 23471 12035 23477
rect 12066 23468 12072 23480
rect 12124 23468 12130 23520
rect 1104 23418 14812 23440
rect 1104 23366 6315 23418
rect 6367 23366 6379 23418
rect 6431 23366 6443 23418
rect 6495 23366 6507 23418
rect 6559 23366 11648 23418
rect 11700 23366 11712 23418
rect 11764 23366 11776 23418
rect 11828 23366 11840 23418
rect 11892 23366 14812 23418
rect 1104 23344 14812 23366
rect 9674 23264 9680 23316
rect 9732 23304 9738 23316
rect 10045 23307 10103 23313
rect 10045 23304 10057 23307
rect 9732 23276 10057 23304
rect 9732 23264 9738 23276
rect 10045 23273 10057 23276
rect 10091 23304 10103 23307
rect 10778 23304 10784 23316
rect 10091 23276 10784 23304
rect 10091 23273 10103 23276
rect 10045 23267 10103 23273
rect 10778 23264 10784 23276
rect 10836 23264 10842 23316
rect 9493 23239 9551 23245
rect 9493 23205 9505 23239
rect 9539 23236 9551 23239
rect 9858 23236 9864 23248
rect 9539 23208 9864 23236
rect 9539 23205 9551 23208
rect 9493 23199 9551 23205
rect 9858 23196 9864 23208
rect 9916 23236 9922 23248
rect 11974 23236 11980 23248
rect 9916 23208 11980 23236
rect 9916 23196 9922 23208
rect 11974 23196 11980 23208
rect 12032 23196 12038 23248
rect 9674 23128 9680 23180
rect 9732 23168 9738 23180
rect 9732 23140 10272 23168
rect 9732 23128 9738 23140
rect 10134 23100 10140 23112
rect 10095 23072 10140 23100
rect 10134 23060 10140 23072
rect 10192 23060 10198 23112
rect 10244 23109 10272 23140
rect 10229 23103 10287 23109
rect 10229 23069 10241 23103
rect 10275 23100 10287 23103
rect 10318 23100 10324 23112
rect 10275 23072 10324 23100
rect 10275 23069 10287 23072
rect 10229 23063 10287 23069
rect 10318 23060 10324 23072
rect 10376 23060 10382 23112
rect 9674 22964 9680 22976
rect 9635 22936 9680 22964
rect 9674 22924 9680 22936
rect 9732 22924 9738 22976
rect 1104 22874 14812 22896
rect 1104 22822 3648 22874
rect 3700 22822 3712 22874
rect 3764 22822 3776 22874
rect 3828 22822 3840 22874
rect 3892 22822 8982 22874
rect 9034 22822 9046 22874
rect 9098 22822 9110 22874
rect 9162 22822 9174 22874
rect 9226 22822 14315 22874
rect 14367 22822 14379 22874
rect 14431 22822 14443 22874
rect 14495 22822 14507 22874
rect 14559 22822 14812 22874
rect 1104 22800 14812 22822
rect 10318 22720 10324 22772
rect 10376 22760 10382 22772
rect 10413 22763 10471 22769
rect 10413 22760 10425 22763
rect 10376 22732 10425 22760
rect 10376 22720 10382 22732
rect 10413 22729 10425 22732
rect 10459 22729 10471 22763
rect 10778 22760 10784 22772
rect 10739 22732 10784 22760
rect 10413 22723 10471 22729
rect 10778 22720 10784 22732
rect 10836 22720 10842 22772
rect 9401 22695 9459 22701
rect 9401 22661 9413 22695
rect 9447 22692 9459 22695
rect 10134 22692 10140 22704
rect 9447 22664 10140 22692
rect 9447 22661 9459 22664
rect 9401 22655 9459 22661
rect 10134 22652 10140 22664
rect 10192 22652 10198 22704
rect 9858 22624 9864 22636
rect 9819 22596 9864 22624
rect 9858 22584 9864 22596
rect 9916 22584 9922 22636
rect 10042 22624 10048 22636
rect 10003 22596 10048 22624
rect 10042 22584 10048 22596
rect 10100 22584 10106 22636
rect 7469 22491 7527 22497
rect 7469 22457 7481 22491
rect 7515 22488 7527 22491
rect 7558 22488 7564 22500
rect 7515 22460 7564 22488
rect 7515 22457 7527 22460
rect 7469 22451 7527 22457
rect 7558 22448 7564 22460
rect 7616 22448 7622 22500
rect 8754 22380 8760 22432
rect 8812 22420 8818 22432
rect 8849 22423 8907 22429
rect 8849 22420 8861 22423
rect 8812 22392 8861 22420
rect 8812 22380 8818 22392
rect 8849 22389 8861 22392
rect 8895 22389 8907 22423
rect 9766 22420 9772 22432
rect 9727 22392 9772 22420
rect 8849 22383 8907 22389
rect 9766 22380 9772 22392
rect 9824 22380 9830 22432
rect 1104 22330 14812 22352
rect 1104 22278 6315 22330
rect 6367 22278 6379 22330
rect 6431 22278 6443 22330
rect 6495 22278 6507 22330
rect 6559 22278 11648 22330
rect 11700 22278 11712 22330
rect 11764 22278 11776 22330
rect 11828 22278 11840 22330
rect 11892 22278 14812 22330
rect 1104 22256 14812 22278
rect 10134 22176 10140 22228
rect 10192 22216 10198 22228
rect 10229 22219 10287 22225
rect 10229 22216 10241 22219
rect 10192 22188 10241 22216
rect 10192 22176 10198 22188
rect 10229 22185 10241 22188
rect 10275 22185 10287 22219
rect 10229 22179 10287 22185
rect 9953 22151 10011 22157
rect 9953 22117 9965 22151
rect 9999 22148 10011 22151
rect 10042 22148 10048 22160
rect 9999 22120 10048 22148
rect 9999 22117 10011 22120
rect 9953 22111 10011 22117
rect 10042 22108 10048 22120
rect 10100 22108 10106 22160
rect 5994 22080 6000 22092
rect 5955 22052 6000 22080
rect 5994 22040 6000 22052
rect 6052 22040 6058 22092
rect 6086 22012 6092 22024
rect 6047 21984 6092 22012
rect 6086 21972 6092 21984
rect 6144 21972 6150 22024
rect 6270 22012 6276 22024
rect 6231 21984 6276 22012
rect 6270 21972 6276 21984
rect 6328 21972 6334 22024
rect 9398 21944 9404 21956
rect 9359 21916 9404 21944
rect 9398 21904 9404 21916
rect 9456 21904 9462 21956
rect 5626 21876 5632 21888
rect 5587 21848 5632 21876
rect 5626 21836 5632 21848
rect 5684 21836 5690 21888
rect 1104 21786 14812 21808
rect 1104 21734 3648 21786
rect 3700 21734 3712 21786
rect 3764 21734 3776 21786
rect 3828 21734 3840 21786
rect 3892 21734 8982 21786
rect 9034 21734 9046 21786
rect 9098 21734 9110 21786
rect 9162 21734 9174 21786
rect 9226 21734 14315 21786
rect 14367 21734 14379 21786
rect 14431 21734 14443 21786
rect 14495 21734 14507 21786
rect 14559 21734 14812 21786
rect 1104 21712 14812 21734
rect 5994 21672 6000 21684
rect 5955 21644 6000 21672
rect 5994 21632 6000 21644
rect 6052 21632 6058 21684
rect 6270 21632 6276 21684
rect 6328 21672 6334 21684
rect 6365 21675 6423 21681
rect 6365 21672 6377 21675
rect 6328 21644 6377 21672
rect 6328 21632 6334 21644
rect 6365 21641 6377 21644
rect 6411 21641 6423 21675
rect 6365 21635 6423 21641
rect 5721 21335 5779 21341
rect 5721 21301 5733 21335
rect 5767 21332 5779 21335
rect 5994 21332 6000 21344
rect 5767 21304 6000 21332
rect 5767 21301 5779 21304
rect 5721 21295 5779 21301
rect 5994 21292 6000 21304
rect 6052 21292 6058 21344
rect 1104 21242 14812 21264
rect 1104 21190 6315 21242
rect 6367 21190 6379 21242
rect 6431 21190 6443 21242
rect 6495 21190 6507 21242
rect 6559 21190 11648 21242
rect 11700 21190 11712 21242
rect 11764 21190 11776 21242
rect 11828 21190 11840 21242
rect 11892 21190 14812 21242
rect 1104 21168 14812 21190
rect 5626 21088 5632 21140
rect 5684 21128 5690 21140
rect 7006 21128 7012 21140
rect 5684 21100 7012 21128
rect 5684 21088 5690 21100
rect 7006 21088 7012 21100
rect 7064 21088 7070 21140
rect 1104 20698 14812 20720
rect 1104 20646 3648 20698
rect 3700 20646 3712 20698
rect 3764 20646 3776 20698
rect 3828 20646 3840 20698
rect 3892 20646 8982 20698
rect 9034 20646 9046 20698
rect 9098 20646 9110 20698
rect 9162 20646 9174 20698
rect 9226 20646 14315 20698
rect 14367 20646 14379 20698
rect 14431 20646 14443 20698
rect 14495 20646 14507 20698
rect 14559 20646 14812 20698
rect 1104 20624 14812 20646
rect 7006 20408 7012 20460
rect 7064 20448 7070 20460
rect 7469 20451 7527 20457
rect 7469 20448 7481 20451
rect 7064 20420 7481 20448
rect 7064 20408 7070 20420
rect 7469 20417 7481 20420
rect 7515 20417 7527 20451
rect 7650 20448 7656 20460
rect 7611 20420 7656 20448
rect 7469 20411 7527 20417
rect 7650 20408 7656 20420
rect 7708 20408 7714 20460
rect 8754 20380 8760 20392
rect 8715 20352 8760 20380
rect 8754 20340 8760 20352
rect 8812 20380 8818 20392
rect 9033 20383 9091 20389
rect 9033 20380 9045 20383
rect 8812 20352 9045 20380
rect 8812 20340 8818 20352
rect 9033 20349 9045 20352
rect 9079 20349 9091 20383
rect 9033 20343 9091 20349
rect 5166 20272 5172 20324
rect 5224 20312 5230 20324
rect 6641 20315 6699 20321
rect 6641 20312 6653 20315
rect 5224 20284 6653 20312
rect 5224 20272 5230 20284
rect 6641 20281 6653 20284
rect 6687 20312 6699 20315
rect 6687 20284 7420 20312
rect 6687 20281 6699 20284
rect 6641 20275 6699 20281
rect 7392 20256 7420 20284
rect 7006 20244 7012 20256
rect 6967 20216 7012 20244
rect 7006 20204 7012 20216
rect 7064 20204 7070 20256
rect 7374 20244 7380 20256
rect 7335 20216 7380 20244
rect 7374 20204 7380 20216
rect 7432 20204 7438 20256
rect 8570 20244 8576 20256
rect 8531 20216 8576 20244
rect 8570 20204 8576 20216
rect 8628 20204 8634 20256
rect 1104 20154 14812 20176
rect 1104 20102 6315 20154
rect 6367 20102 6379 20154
rect 6431 20102 6443 20154
rect 6495 20102 6507 20154
rect 6559 20102 11648 20154
rect 11700 20102 11712 20154
rect 11764 20102 11776 20154
rect 11828 20102 11840 20154
rect 11892 20102 14812 20154
rect 1104 20080 14812 20102
rect 7101 20043 7159 20049
rect 7101 20009 7113 20043
rect 7147 20040 7159 20043
rect 7650 20040 7656 20052
rect 7147 20012 7656 20040
rect 7147 20009 7159 20012
rect 7101 20003 7159 20009
rect 7650 20000 7656 20012
rect 7708 20000 7714 20052
rect 12342 19904 12348 19916
rect 12303 19876 12348 19904
rect 12342 19864 12348 19876
rect 12400 19864 12406 19916
rect 12434 19660 12440 19712
rect 12492 19700 12498 19712
rect 12529 19703 12587 19709
rect 12529 19700 12541 19703
rect 12492 19672 12541 19700
rect 12492 19660 12498 19672
rect 12529 19669 12541 19672
rect 12575 19669 12587 19703
rect 12529 19663 12587 19669
rect 1104 19610 14812 19632
rect 1104 19558 3648 19610
rect 3700 19558 3712 19610
rect 3764 19558 3776 19610
rect 3828 19558 3840 19610
rect 3892 19558 8982 19610
rect 9034 19558 9046 19610
rect 9098 19558 9110 19610
rect 9162 19558 9174 19610
rect 9226 19558 14315 19610
rect 14367 19558 14379 19610
rect 14431 19558 14443 19610
rect 14495 19558 14507 19610
rect 14559 19558 14812 19610
rect 1104 19536 14812 19558
rect 10410 19320 10416 19372
rect 10468 19360 10474 19372
rect 10594 19360 10600 19372
rect 10468 19332 10600 19360
rect 10468 19320 10474 19332
rect 10594 19320 10600 19332
rect 10652 19320 10658 19372
rect 12342 19320 12348 19372
rect 12400 19360 12406 19372
rect 12621 19363 12679 19369
rect 12621 19360 12633 19363
rect 12400 19332 12633 19360
rect 12400 19320 12406 19332
rect 12621 19329 12633 19332
rect 12667 19329 12679 19363
rect 12621 19323 12679 19329
rect 12710 19320 12716 19372
rect 12768 19360 12774 19372
rect 12986 19360 12992 19372
rect 12768 19332 12992 19360
rect 12768 19320 12774 19332
rect 12986 19320 12992 19332
rect 13044 19320 13050 19372
rect 3142 19252 3148 19304
rect 3200 19292 3206 19304
rect 3418 19292 3424 19304
rect 3200 19264 3424 19292
rect 3200 19252 3206 19264
rect 3418 19252 3424 19264
rect 3476 19252 3482 19304
rect 14182 19252 14188 19304
rect 14240 19292 14246 19304
rect 14921 19295 14979 19301
rect 14921 19292 14933 19295
rect 14240 19264 14933 19292
rect 14240 19252 14246 19264
rect 14921 19261 14933 19264
rect 14967 19261 14979 19295
rect 14921 19255 14979 19261
rect 4338 19184 4344 19236
rect 4396 19224 4402 19236
rect 4522 19224 4528 19236
rect 4396 19196 4528 19224
rect 4396 19184 4402 19196
rect 4522 19184 4528 19196
rect 4580 19184 4586 19236
rect 1104 19066 14812 19088
rect 1104 19014 6315 19066
rect 6367 19014 6379 19066
rect 6431 19014 6443 19066
rect 6495 19014 6507 19066
rect 6559 19014 11648 19066
rect 11700 19014 11712 19066
rect 11764 19014 11776 19066
rect 11828 19014 11840 19066
rect 11892 19014 14812 19066
rect 1104 18992 14812 19014
rect 1104 18522 14812 18544
rect 1104 18470 3648 18522
rect 3700 18470 3712 18522
rect 3764 18470 3776 18522
rect 3828 18470 3840 18522
rect 3892 18470 8982 18522
rect 9034 18470 9046 18522
rect 9098 18470 9110 18522
rect 9162 18470 9174 18522
rect 9226 18470 14315 18522
rect 14367 18470 14379 18522
rect 14431 18470 14443 18522
rect 14495 18470 14507 18522
rect 14559 18470 14812 18522
rect 1104 18448 14812 18470
rect 1104 17978 14812 18000
rect 1104 17926 6315 17978
rect 6367 17926 6379 17978
rect 6431 17926 6443 17978
rect 6495 17926 6507 17978
rect 6559 17926 11648 17978
rect 11700 17926 11712 17978
rect 11764 17926 11776 17978
rect 11828 17926 11840 17978
rect 11892 17926 14812 17978
rect 1104 17904 14812 17926
rect 1104 17434 14812 17456
rect 1104 17382 3648 17434
rect 3700 17382 3712 17434
rect 3764 17382 3776 17434
rect 3828 17382 3840 17434
rect 3892 17382 8982 17434
rect 9034 17382 9046 17434
rect 9098 17382 9110 17434
rect 9162 17382 9174 17434
rect 9226 17382 14315 17434
rect 14367 17382 14379 17434
rect 14431 17382 14443 17434
rect 14495 17382 14507 17434
rect 14559 17382 14812 17434
rect 1104 17360 14812 17382
rect 1104 16890 14812 16912
rect 1104 16838 6315 16890
rect 6367 16838 6379 16890
rect 6431 16838 6443 16890
rect 6495 16838 6507 16890
rect 6559 16838 11648 16890
rect 11700 16838 11712 16890
rect 11764 16838 11776 16890
rect 11828 16838 11840 16890
rect 11892 16838 14812 16890
rect 1104 16816 14812 16838
rect 4430 16776 4436 16788
rect 4391 16748 4436 16776
rect 4430 16736 4436 16748
rect 4488 16736 4494 16788
rect 12250 16736 12256 16788
rect 12308 16776 12314 16788
rect 12897 16779 12955 16785
rect 12897 16776 12909 16779
rect 12308 16748 12909 16776
rect 12308 16736 12314 16748
rect 12897 16745 12909 16748
rect 12943 16745 12955 16779
rect 12897 16739 12955 16745
rect 1946 16600 1952 16652
rect 2004 16640 2010 16652
rect 2222 16640 2228 16652
rect 2004 16612 2228 16640
rect 2004 16600 2010 16612
rect 2222 16600 2228 16612
rect 2280 16600 2286 16652
rect 11514 16640 11520 16652
rect 11475 16612 11520 16640
rect 11514 16600 11520 16612
rect 11572 16600 11578 16652
rect 11606 16600 11612 16652
rect 11664 16640 11670 16652
rect 11773 16643 11831 16649
rect 11773 16640 11785 16643
rect 11664 16612 11785 16640
rect 11664 16600 11670 16612
rect 11773 16609 11785 16612
rect 11819 16609 11831 16643
rect 11773 16603 11831 16609
rect 1104 16346 14812 16368
rect 1104 16294 3648 16346
rect 3700 16294 3712 16346
rect 3764 16294 3776 16346
rect 3828 16294 3840 16346
rect 3892 16294 8982 16346
rect 9034 16294 9046 16346
rect 9098 16294 9110 16346
rect 9162 16294 9174 16346
rect 9226 16294 14315 16346
rect 14367 16294 14379 16346
rect 14431 16294 14443 16346
rect 14495 16294 14507 16346
rect 14559 16294 14812 16346
rect 1104 16272 14812 16294
rect 11514 16192 11520 16244
rect 11572 16232 11578 16244
rect 11885 16235 11943 16241
rect 11885 16232 11897 16235
rect 11572 16204 11897 16232
rect 11572 16192 11578 16204
rect 11885 16201 11897 16204
rect 11931 16201 11943 16235
rect 11885 16195 11943 16201
rect 4430 16056 4436 16108
rect 4488 16096 4494 16108
rect 4982 16096 4988 16108
rect 4488 16068 4988 16096
rect 4488 16056 4494 16068
rect 4982 16056 4988 16068
rect 5040 16056 5046 16108
rect 4798 16028 4804 16040
rect 4759 16000 4804 16028
rect 4798 15988 4804 16000
rect 4856 15988 4862 16040
rect 4338 15960 4344 15972
rect 4251 15932 4344 15960
rect 4338 15920 4344 15932
rect 4396 15960 4402 15972
rect 11606 15960 11612 15972
rect 4396 15932 4936 15960
rect 4396 15920 4402 15932
rect 4908 15904 4936 15932
rect 11532 15932 11612 15960
rect 4430 15892 4436 15904
rect 4391 15864 4436 15892
rect 4430 15852 4436 15864
rect 4488 15852 4494 15904
rect 4890 15852 4896 15904
rect 4948 15892 4954 15904
rect 4948 15864 4993 15892
rect 4948 15852 4954 15864
rect 11054 15852 11060 15904
rect 11112 15892 11118 15904
rect 11532 15901 11560 15932
rect 11606 15920 11612 15932
rect 11664 15920 11670 15972
rect 11517 15895 11575 15901
rect 11517 15892 11529 15895
rect 11112 15864 11529 15892
rect 11112 15852 11118 15864
rect 11517 15861 11529 15864
rect 11563 15861 11575 15895
rect 11517 15855 11575 15861
rect 1104 15802 14812 15824
rect 1104 15750 6315 15802
rect 6367 15750 6379 15802
rect 6431 15750 6443 15802
rect 6495 15750 6507 15802
rect 6559 15750 11648 15802
rect 11700 15750 11712 15802
rect 11764 15750 11776 15802
rect 11828 15750 11840 15802
rect 11892 15750 14812 15802
rect 1104 15728 14812 15750
rect 4430 15648 4436 15700
rect 4488 15688 4494 15700
rect 5629 15691 5687 15697
rect 5629 15688 5641 15691
rect 4488 15660 5641 15688
rect 4488 15648 4494 15660
rect 5629 15657 5641 15660
rect 5675 15688 5687 15691
rect 5718 15688 5724 15700
rect 5675 15660 5724 15688
rect 5675 15657 5687 15660
rect 5629 15651 5687 15657
rect 5718 15648 5724 15660
rect 5776 15648 5782 15700
rect 7006 15648 7012 15700
rect 7064 15688 7070 15700
rect 7285 15691 7343 15697
rect 7285 15688 7297 15691
rect 7064 15660 7297 15688
rect 7064 15648 7070 15660
rect 7285 15657 7297 15660
rect 7331 15657 7343 15691
rect 7285 15651 7343 15657
rect 4525 15623 4583 15629
rect 4525 15589 4537 15623
rect 4571 15620 4583 15623
rect 4798 15620 4804 15632
rect 4571 15592 4804 15620
rect 4571 15589 4583 15592
rect 4525 15583 4583 15589
rect 4798 15580 4804 15592
rect 4856 15580 4862 15632
rect 5534 15552 5540 15564
rect 5495 15524 5540 15552
rect 5534 15512 5540 15524
rect 5592 15512 5598 15564
rect 5626 15444 5632 15496
rect 5684 15484 5690 15496
rect 5721 15487 5779 15493
rect 5721 15484 5733 15487
rect 5684 15456 5733 15484
rect 5684 15444 5690 15456
rect 5721 15453 5733 15456
rect 5767 15453 5779 15487
rect 5721 15447 5779 15453
rect 5166 15348 5172 15360
rect 5127 15320 5172 15348
rect 5166 15308 5172 15320
rect 5224 15308 5230 15360
rect 1104 15258 14812 15280
rect 1104 15206 3648 15258
rect 3700 15206 3712 15258
rect 3764 15206 3776 15258
rect 3828 15206 3840 15258
rect 3892 15206 8982 15258
rect 9034 15206 9046 15258
rect 9098 15206 9110 15258
rect 9162 15206 9174 15258
rect 9226 15206 14315 15258
rect 14367 15206 14379 15258
rect 14431 15206 14443 15258
rect 14495 15206 14507 15258
rect 14559 15206 14812 15258
rect 1104 15184 14812 15206
rect 1578 15144 1584 15156
rect 1539 15116 1584 15144
rect 1578 15104 1584 15116
rect 1636 15104 1642 15156
rect 2038 15144 2044 15156
rect 1999 15116 2044 15144
rect 2038 15104 2044 15116
rect 2096 15104 2102 15156
rect 5537 15147 5595 15153
rect 5537 15113 5549 15147
rect 5583 15144 5595 15147
rect 5626 15144 5632 15156
rect 5583 15116 5632 15144
rect 5583 15113 5595 15116
rect 5537 15107 5595 15113
rect 5626 15104 5632 15116
rect 5684 15104 5690 15156
rect 5718 15104 5724 15156
rect 5776 15144 5782 15156
rect 5813 15147 5871 15153
rect 5813 15144 5825 15147
rect 5776 15116 5825 15144
rect 5776 15104 5782 15116
rect 5813 15113 5825 15116
rect 5859 15113 5871 15147
rect 5813 15107 5871 15113
rect 8570 15104 8576 15156
rect 8628 15144 8634 15156
rect 8941 15147 8999 15153
rect 8941 15144 8953 15147
rect 8628 15116 8953 15144
rect 8628 15104 8634 15116
rect 8941 15113 8953 15116
rect 8987 15113 8999 15147
rect 8941 15107 8999 15113
rect 3973 15011 4031 15017
rect 3973 14977 3985 15011
rect 4019 15008 4031 15011
rect 4982 15008 4988 15020
rect 4019 14980 4988 15008
rect 4019 14977 4031 14980
rect 3973 14971 4031 14977
rect 4982 14968 4988 14980
rect 5040 14968 5046 15020
rect 7193 15011 7251 15017
rect 7193 14977 7205 15011
rect 7239 15008 7251 15011
rect 7929 15011 7987 15017
rect 7929 15008 7941 15011
rect 7239 14980 7941 15008
rect 7239 14977 7251 14980
rect 7193 14971 7251 14977
rect 7929 14977 7941 14980
rect 7975 14977 7987 15011
rect 8956 15008 8984 15107
rect 9493 15011 9551 15017
rect 9493 15008 9505 15011
rect 8956 14980 9505 15008
rect 7929 14971 7987 14977
rect 9493 14977 9505 14980
rect 9539 14977 9551 15011
rect 9493 14971 9551 14977
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14940 1455 14943
rect 2038 14940 2044 14952
rect 1443 14912 2044 14940
rect 1443 14909 1455 14912
rect 1397 14903 1455 14909
rect 2038 14900 2044 14912
rect 2096 14900 2102 14952
rect 4798 14940 4804 14952
rect 4759 14912 4804 14940
rect 4798 14900 4804 14912
rect 4856 14900 4862 14952
rect 7006 14900 7012 14952
rect 7064 14940 7070 14952
rect 7653 14943 7711 14949
rect 7653 14940 7665 14943
rect 7064 14912 7665 14940
rect 7064 14900 7070 14912
rect 7653 14909 7665 14912
rect 7699 14909 7711 14943
rect 7944 14940 7972 14971
rect 9401 14943 9459 14949
rect 9401 14940 9413 14943
rect 7944 14912 9413 14940
rect 7653 14903 7711 14909
rect 9401 14909 9413 14912
rect 9447 14940 9459 14943
rect 9582 14940 9588 14952
rect 9447 14912 9588 14940
rect 9447 14909 9459 14912
rect 9401 14903 9459 14909
rect 9582 14900 9588 14912
rect 9640 14940 9646 14952
rect 9749 14943 9807 14949
rect 9749 14940 9761 14943
rect 9640 14912 9761 14940
rect 9640 14900 9646 14912
rect 9749 14909 9761 14912
rect 9795 14909 9807 14943
rect 9749 14903 9807 14909
rect 4338 14872 4344 14884
rect 4251 14844 4344 14872
rect 4338 14832 4344 14844
rect 4396 14872 4402 14884
rect 4396 14844 4936 14872
rect 4396 14832 4402 14844
rect 4908 14816 4936 14844
rect 7190 14832 7196 14884
rect 7248 14872 7254 14884
rect 7745 14875 7803 14881
rect 7745 14872 7757 14875
rect 7248 14844 7757 14872
rect 7248 14832 7254 14844
rect 7745 14841 7757 14844
rect 7791 14841 7803 14875
rect 7745 14835 7803 14841
rect 4430 14804 4436 14816
rect 4391 14776 4436 14804
rect 4430 14764 4436 14776
rect 4488 14764 4494 14816
rect 4890 14764 4896 14816
rect 4948 14804 4954 14816
rect 7282 14804 7288 14816
rect 4948 14776 4993 14804
rect 7243 14776 7288 14804
rect 4948 14764 4954 14776
rect 7282 14764 7288 14776
rect 7340 14764 7346 14816
rect 10870 14804 10876 14816
rect 10831 14776 10876 14804
rect 10870 14764 10876 14776
rect 10928 14764 10934 14816
rect 1104 14714 14812 14736
rect 1104 14662 6315 14714
rect 6367 14662 6379 14714
rect 6431 14662 6443 14714
rect 6495 14662 6507 14714
rect 6559 14662 11648 14714
rect 11700 14662 11712 14714
rect 11764 14662 11776 14714
rect 11828 14662 11840 14714
rect 11892 14662 14812 14714
rect 1104 14640 14812 14662
rect 4430 14560 4436 14612
rect 4488 14600 4494 14612
rect 5261 14603 5319 14609
rect 5261 14600 5273 14603
rect 4488 14572 5273 14600
rect 4488 14560 4494 14572
rect 5261 14569 5273 14572
rect 5307 14600 5319 14603
rect 5534 14600 5540 14612
rect 5307 14572 5540 14600
rect 5307 14569 5319 14572
rect 5261 14563 5319 14569
rect 5534 14560 5540 14572
rect 5592 14560 5598 14612
rect 7190 14560 7196 14612
rect 7248 14600 7254 14612
rect 7285 14603 7343 14609
rect 7285 14600 7297 14603
rect 7248 14572 7297 14600
rect 7248 14560 7254 14572
rect 7285 14569 7297 14572
rect 7331 14569 7343 14603
rect 8018 14600 8024 14612
rect 7979 14572 8024 14600
rect 7285 14563 7343 14569
rect 8018 14560 8024 14572
rect 8076 14560 8082 14612
rect 4525 14535 4583 14541
rect 4525 14501 4537 14535
rect 4571 14532 4583 14535
rect 4798 14532 4804 14544
rect 4571 14504 4804 14532
rect 4571 14501 4583 14504
rect 4525 14495 4583 14501
rect 4798 14492 4804 14504
rect 4856 14492 4862 14544
rect 1104 14170 14812 14192
rect 1104 14118 3648 14170
rect 3700 14118 3712 14170
rect 3764 14118 3776 14170
rect 3828 14118 3840 14170
rect 3892 14118 8982 14170
rect 9034 14118 9046 14170
rect 9098 14118 9110 14170
rect 9162 14118 9174 14170
rect 9226 14118 14315 14170
rect 14367 14118 14379 14170
rect 14431 14118 14443 14170
rect 14495 14118 14507 14170
rect 14559 14118 14812 14170
rect 1104 14096 14812 14118
rect 7837 13923 7895 13929
rect 7837 13889 7849 13923
rect 7883 13920 7895 13923
rect 8481 13923 8539 13929
rect 8481 13920 8493 13923
rect 7883 13892 8493 13920
rect 7883 13889 7895 13892
rect 7837 13883 7895 13889
rect 8481 13889 8493 13892
rect 8527 13920 8539 13923
rect 10870 13920 10876 13932
rect 8527 13892 10876 13920
rect 8527 13889 8539 13892
rect 8481 13883 8539 13889
rect 10870 13880 10876 13892
rect 10928 13880 10934 13932
rect 1854 13812 1860 13864
rect 1912 13852 1918 13864
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 1912 13824 2053 13852
rect 1912 13812 1918 13824
rect 2041 13821 2053 13824
rect 2087 13852 2099 13855
rect 2593 13855 2651 13861
rect 2593 13852 2605 13855
rect 2087 13824 2605 13852
rect 2087 13821 2099 13824
rect 2041 13815 2099 13821
rect 2593 13821 2605 13824
rect 2639 13821 2651 13855
rect 2593 13815 2651 13821
rect 8018 13744 8024 13796
rect 8076 13784 8082 13796
rect 8389 13787 8447 13793
rect 8389 13784 8401 13787
rect 8076 13756 8401 13784
rect 8076 13744 8082 13756
rect 8389 13753 8401 13756
rect 8435 13753 8447 13787
rect 8389 13747 8447 13753
rect 2222 13716 2228 13728
rect 2183 13688 2228 13716
rect 2222 13676 2228 13688
rect 2280 13676 2286 13728
rect 7926 13716 7932 13728
rect 7887 13688 7932 13716
rect 7926 13676 7932 13688
rect 7984 13676 7990 13728
rect 8294 13716 8300 13728
rect 8255 13688 8300 13716
rect 8294 13676 8300 13688
rect 8352 13676 8358 13728
rect 1104 13626 14812 13648
rect 1104 13574 6315 13626
rect 6367 13574 6379 13626
rect 6431 13574 6443 13626
rect 6495 13574 6507 13626
rect 6559 13574 11648 13626
rect 11700 13574 11712 13626
rect 11764 13574 11776 13626
rect 11828 13574 11840 13626
rect 11892 13574 14812 13626
rect 1104 13552 14812 13574
rect 7282 13472 7288 13524
rect 7340 13512 7346 13524
rect 7929 13515 7987 13521
rect 7929 13512 7941 13515
rect 7340 13484 7941 13512
rect 7340 13472 7346 13484
rect 7929 13481 7941 13484
rect 7975 13512 7987 13515
rect 8018 13512 8024 13524
rect 7975 13484 8024 13512
rect 7975 13481 7987 13484
rect 7929 13475 7987 13481
rect 8018 13472 8024 13484
rect 8076 13472 8082 13524
rect 1104 13082 14812 13104
rect 1104 13030 3648 13082
rect 3700 13030 3712 13082
rect 3764 13030 3776 13082
rect 3828 13030 3840 13082
rect 3892 13030 8982 13082
rect 9034 13030 9046 13082
rect 9098 13030 9110 13082
rect 9162 13030 9174 13082
rect 9226 13030 14315 13082
rect 14367 13030 14379 13082
rect 14431 13030 14443 13082
rect 14495 13030 14507 13082
rect 14559 13030 14812 13082
rect 1104 13008 14812 13030
rect 8938 12860 8944 12912
rect 8996 12900 9002 12912
rect 9398 12900 9404 12912
rect 8996 12872 9404 12900
rect 8996 12860 9002 12872
rect 9398 12860 9404 12872
rect 9456 12860 9462 12912
rect 1104 12538 14812 12560
rect 1104 12486 6315 12538
rect 6367 12486 6379 12538
rect 6431 12486 6443 12538
rect 6495 12486 6507 12538
rect 6559 12486 11648 12538
rect 11700 12486 11712 12538
rect 11764 12486 11776 12538
rect 11828 12486 11840 12538
rect 11892 12486 14812 12538
rect 1104 12464 14812 12486
rect 1394 12288 1400 12300
rect 1355 12260 1400 12288
rect 1394 12248 1400 12260
rect 1452 12248 1458 12300
rect 1578 12220 1584 12232
rect 1539 12192 1584 12220
rect 1578 12180 1584 12192
rect 1636 12180 1642 12232
rect 1104 11994 14812 12016
rect 1104 11942 3648 11994
rect 3700 11942 3712 11994
rect 3764 11942 3776 11994
rect 3828 11942 3840 11994
rect 3892 11942 8982 11994
rect 9034 11942 9046 11994
rect 9098 11942 9110 11994
rect 9162 11942 9174 11994
rect 9226 11942 14315 11994
rect 14367 11942 14379 11994
rect 14431 11942 14443 11994
rect 14495 11942 14507 11994
rect 14559 11942 14812 11994
rect 1104 11920 14812 11942
rect 1394 11840 1400 11892
rect 1452 11880 1458 11892
rect 1581 11883 1639 11889
rect 1581 11880 1593 11883
rect 1452 11852 1593 11880
rect 1452 11840 1458 11852
rect 1581 11849 1593 11852
rect 1627 11849 1639 11883
rect 1581 11843 1639 11849
rect 1104 11450 14812 11472
rect 1104 11398 6315 11450
rect 6367 11398 6379 11450
rect 6431 11398 6443 11450
rect 6495 11398 6507 11450
rect 6559 11398 11648 11450
rect 11700 11398 11712 11450
rect 11764 11398 11776 11450
rect 11828 11398 11840 11450
rect 11892 11398 14812 11450
rect 1104 11376 14812 11398
rect 1949 11203 2007 11209
rect 1949 11169 1961 11203
rect 1995 11200 2007 11203
rect 2314 11200 2320 11212
rect 1995 11172 2320 11200
rect 1995 11169 2007 11172
rect 1949 11163 2007 11169
rect 2314 11160 2320 11172
rect 2372 11160 2378 11212
rect 1210 11024 1216 11076
rect 1268 11064 1274 11076
rect 2133 11067 2191 11073
rect 2133 11064 2145 11067
rect 1268 11036 2145 11064
rect 1268 11024 1274 11036
rect 2133 11033 2145 11036
rect 2179 11033 2191 11067
rect 2133 11027 2191 11033
rect 1104 10906 14812 10928
rect 1104 10854 3648 10906
rect 3700 10854 3712 10906
rect 3764 10854 3776 10906
rect 3828 10854 3840 10906
rect 3892 10854 8982 10906
rect 9034 10854 9046 10906
rect 9098 10854 9110 10906
rect 9162 10854 9174 10906
rect 9226 10854 14315 10906
rect 14367 10854 14379 10906
rect 14431 10854 14443 10906
rect 14495 10854 14507 10906
rect 14559 10854 14812 10906
rect 1104 10832 14812 10854
rect 2041 10795 2099 10801
rect 2041 10761 2053 10795
rect 2087 10792 2099 10795
rect 2314 10792 2320 10804
rect 2087 10764 2320 10792
rect 2087 10761 2099 10764
rect 2041 10755 2099 10761
rect 2314 10752 2320 10764
rect 2372 10752 2378 10804
rect 13081 10795 13139 10801
rect 13081 10761 13093 10795
rect 13127 10792 13139 10795
rect 14090 10792 14096 10804
rect 13127 10764 14096 10792
rect 13127 10761 13139 10764
rect 13081 10755 13139 10761
rect 2038 10616 2044 10668
rect 2096 10656 2102 10668
rect 2314 10656 2320 10668
rect 2096 10628 2320 10656
rect 2096 10616 2102 10628
rect 2314 10616 2320 10628
rect 2372 10616 2378 10668
rect 12437 10591 12495 10597
rect 12437 10557 12449 10591
rect 12483 10588 12495 10591
rect 13096 10588 13124 10755
rect 14090 10752 14096 10764
rect 14148 10752 14154 10804
rect 12483 10560 13124 10588
rect 12483 10557 12495 10560
rect 12437 10551 12495 10557
rect 6914 10412 6920 10464
rect 6972 10452 6978 10464
rect 8202 10452 8208 10464
rect 6972 10424 8208 10452
rect 6972 10412 6978 10424
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12621 10455 12679 10461
rect 12621 10452 12633 10455
rect 12492 10424 12633 10452
rect 12492 10412 12498 10424
rect 12621 10421 12633 10424
rect 12667 10421 12679 10455
rect 12621 10415 12679 10421
rect 1104 10362 14812 10384
rect 1104 10310 6315 10362
rect 6367 10310 6379 10362
rect 6431 10310 6443 10362
rect 6495 10310 6507 10362
rect 6559 10310 11648 10362
rect 11700 10310 11712 10362
rect 11764 10310 11776 10362
rect 11828 10310 11840 10362
rect 11892 10310 14812 10362
rect 1104 10288 14812 10310
rect 1104 9818 14812 9840
rect 1104 9766 3648 9818
rect 3700 9766 3712 9818
rect 3764 9766 3776 9818
rect 3828 9766 3840 9818
rect 3892 9766 8982 9818
rect 9034 9766 9046 9818
rect 9098 9766 9110 9818
rect 9162 9766 9174 9818
rect 9226 9766 14315 9818
rect 14367 9766 14379 9818
rect 14431 9766 14443 9818
rect 14495 9766 14507 9818
rect 14559 9766 14812 9818
rect 1104 9744 14812 9766
rect 3142 9664 3148 9716
rect 3200 9704 3206 9716
rect 3418 9704 3424 9716
rect 3200 9676 3424 9704
rect 3200 9664 3206 9676
rect 3418 9664 3424 9676
rect 3476 9664 3482 9716
rect 14734 9664 14740 9716
rect 14792 9704 14798 9716
rect 14921 9707 14979 9713
rect 14921 9704 14933 9707
rect 14792 9676 14933 9704
rect 14792 9664 14798 9676
rect 14921 9673 14933 9676
rect 14967 9673 14979 9707
rect 14921 9667 14979 9673
rect 2590 9596 2596 9648
rect 2648 9636 2654 9648
rect 2869 9639 2927 9645
rect 2869 9636 2881 9639
rect 2648 9608 2881 9636
rect 2648 9596 2654 9608
rect 2869 9605 2881 9608
rect 2915 9605 2927 9639
rect 2869 9599 2927 9605
rect 2685 9503 2743 9509
rect 2685 9469 2697 9503
rect 2731 9469 2743 9503
rect 2685 9463 2743 9469
rect 2700 9432 2728 9463
rect 3329 9435 3387 9441
rect 3329 9432 3341 9435
rect 2700 9404 3341 9432
rect 3329 9401 3341 9404
rect 3375 9432 3387 9435
rect 3510 9432 3516 9444
rect 3375 9404 3516 9432
rect 3375 9401 3387 9404
rect 3329 9395 3387 9401
rect 3510 9392 3516 9404
rect 3568 9392 3574 9444
rect 1104 9274 14812 9296
rect 1104 9222 6315 9274
rect 6367 9222 6379 9274
rect 6431 9222 6443 9274
rect 6495 9222 6507 9274
rect 6559 9222 11648 9274
rect 11700 9222 11712 9274
rect 11764 9222 11776 9274
rect 11828 9222 11840 9274
rect 11892 9222 14812 9274
rect 1104 9200 14812 9222
rect 10594 9160 10600 9172
rect 10555 9132 10600 9160
rect 10594 9120 10600 9132
rect 10652 9120 10658 9172
rect 12526 9160 12532 9172
rect 12487 9132 12532 9160
rect 12526 9120 12532 9132
rect 12584 9120 12590 9172
rect 10413 9027 10471 9033
rect 10413 8993 10425 9027
rect 10459 9024 10471 9027
rect 10502 9024 10508 9036
rect 10459 8996 10508 9024
rect 10459 8993 10471 8996
rect 10413 8987 10471 8993
rect 10502 8984 10508 8996
rect 10560 8984 10566 9036
rect 12345 9027 12403 9033
rect 12345 8993 12357 9027
rect 12391 9024 12403 9027
rect 13078 9024 13084 9036
rect 12391 8996 13084 9024
rect 12391 8993 12403 8996
rect 12345 8987 12403 8993
rect 13078 8984 13084 8996
rect 13136 8984 13142 9036
rect 1104 8730 14812 8752
rect 1104 8678 3648 8730
rect 3700 8678 3712 8730
rect 3764 8678 3776 8730
rect 3828 8678 3840 8730
rect 3892 8678 8982 8730
rect 9034 8678 9046 8730
rect 9098 8678 9110 8730
rect 9162 8678 9174 8730
rect 9226 8678 14315 8730
rect 14367 8678 14379 8730
rect 14431 8678 14443 8730
rect 14495 8678 14507 8730
rect 14559 8678 14812 8730
rect 1104 8656 14812 8678
rect 12253 8415 12311 8421
rect 12253 8381 12265 8415
rect 12299 8412 12311 8415
rect 12437 8415 12495 8421
rect 12437 8412 12449 8415
rect 12299 8384 12449 8412
rect 12299 8381 12311 8384
rect 12253 8375 12311 8381
rect 12437 8381 12449 8384
rect 12483 8412 12495 8415
rect 13998 8412 14004 8424
rect 12483 8384 14004 8412
rect 12483 8381 12495 8384
rect 12437 8375 12495 8381
rect 13998 8372 14004 8384
rect 14056 8372 14062 8424
rect 10502 8344 10508 8356
rect 10463 8316 10508 8344
rect 10502 8304 10508 8316
rect 10560 8304 10566 8356
rect 13078 8344 13084 8356
rect 13039 8316 13084 8344
rect 13078 8304 13084 8316
rect 13136 8304 13142 8356
rect 12618 8276 12624 8288
rect 12579 8248 12624 8276
rect 12618 8236 12624 8248
rect 12676 8236 12682 8288
rect 1104 8186 14812 8208
rect 1104 8134 6315 8186
rect 6367 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 11648 8186
rect 11700 8134 11712 8186
rect 11764 8134 11776 8186
rect 11828 8134 11840 8186
rect 11892 8134 14812 8186
rect 1104 8112 14812 8134
rect 3418 8032 3424 8084
rect 3476 8072 3482 8084
rect 4893 8075 4951 8081
rect 4893 8072 4905 8075
rect 3476 8044 4905 8072
rect 3476 8032 3482 8044
rect 4893 8041 4905 8044
rect 4939 8041 4951 8075
rect 4893 8035 4951 8041
rect 4709 7939 4767 7945
rect 4709 7905 4721 7939
rect 4755 7936 4767 7939
rect 4890 7936 4896 7948
rect 4755 7908 4896 7936
rect 4755 7905 4767 7908
rect 4709 7899 4767 7905
rect 4890 7896 4896 7908
rect 4948 7896 4954 7948
rect 1104 7642 14812 7664
rect 1104 7590 3648 7642
rect 3700 7590 3712 7642
rect 3764 7590 3776 7642
rect 3828 7590 3840 7642
rect 3892 7590 8982 7642
rect 9034 7590 9046 7642
rect 9098 7590 9110 7642
rect 9162 7590 9174 7642
rect 9226 7590 14315 7642
rect 14367 7590 14379 7642
rect 14431 7590 14443 7642
rect 14495 7590 14507 7642
rect 14559 7590 14812 7642
rect 1104 7568 14812 7590
rect 7466 7528 7472 7540
rect 7427 7500 7472 7528
rect 7466 7488 7472 7500
rect 7524 7488 7530 7540
rect 6825 7327 6883 7333
rect 6825 7293 6837 7327
rect 6871 7324 6883 7327
rect 7466 7324 7472 7336
rect 6871 7296 7472 7324
rect 6871 7293 6883 7296
rect 6825 7287 6883 7293
rect 7466 7284 7472 7296
rect 7524 7284 7530 7336
rect 4801 7191 4859 7197
rect 4801 7157 4813 7191
rect 4847 7188 4859 7191
rect 4890 7188 4896 7200
rect 4847 7160 4896 7188
rect 4847 7157 4859 7160
rect 4801 7151 4859 7157
rect 4890 7148 4896 7160
rect 4948 7148 4954 7200
rect 7006 7188 7012 7200
rect 6967 7160 7012 7188
rect 7006 7148 7012 7160
rect 7064 7148 7070 7200
rect 1104 7098 14812 7120
rect 1104 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 11648 7098
rect 11700 7046 11712 7098
rect 11764 7046 11776 7098
rect 11828 7046 11840 7098
rect 11892 7046 14812 7098
rect 1104 7024 14812 7046
rect 1578 6848 1584 6860
rect 1539 6820 1584 6848
rect 1578 6808 1584 6820
rect 1636 6808 1642 6860
rect 5997 6851 6055 6857
rect 5997 6817 6009 6851
rect 6043 6848 6055 6851
rect 6270 6848 6276 6860
rect 6043 6820 6276 6848
rect 6043 6817 6055 6820
rect 5997 6811 6055 6817
rect 6270 6808 6276 6820
rect 6328 6808 6334 6860
rect 10413 6851 10471 6857
rect 10413 6817 10425 6851
rect 10459 6848 10471 6851
rect 11238 6848 11244 6860
rect 10459 6820 11244 6848
rect 10459 6817 10471 6820
rect 10413 6811 10471 6817
rect 11238 6808 11244 6820
rect 11296 6808 11302 6860
rect 6178 6712 6184 6724
rect 6139 6684 6184 6712
rect 6178 6672 6184 6684
rect 6236 6672 6242 6724
rect 566 6604 572 6656
rect 624 6644 630 6656
rect 1765 6647 1823 6653
rect 1765 6644 1777 6647
rect 624 6616 1777 6644
rect 624 6604 630 6616
rect 1765 6613 1777 6616
rect 1811 6613 1823 6647
rect 10594 6644 10600 6656
rect 10555 6616 10600 6644
rect 1765 6607 1823 6613
rect 10594 6604 10600 6616
rect 10652 6604 10658 6656
rect 1104 6554 14812 6576
rect 1104 6502 3648 6554
rect 3700 6502 3712 6554
rect 3764 6502 3776 6554
rect 3828 6502 3840 6554
rect 3892 6502 8982 6554
rect 9034 6502 9046 6554
rect 9098 6502 9110 6554
rect 9162 6502 9174 6554
rect 9226 6502 14315 6554
rect 14367 6502 14379 6554
rect 14431 6502 14443 6554
rect 14495 6502 14507 6554
rect 14559 6502 14812 6554
rect 1104 6480 14812 6502
rect 1578 6440 1584 6452
rect 1539 6412 1584 6440
rect 1578 6400 1584 6412
rect 1636 6400 1642 6452
rect 8205 6443 8263 6449
rect 8205 6409 8217 6443
rect 8251 6440 8263 6443
rect 8478 6440 8484 6452
rect 8251 6412 8484 6440
rect 8251 6409 8263 6412
rect 8205 6403 8263 6409
rect 4157 6239 4215 6245
rect 4157 6205 4169 6239
rect 4203 6236 4215 6239
rect 4798 6236 4804 6248
rect 4203 6208 4804 6236
rect 4203 6205 4215 6208
rect 4157 6199 4215 6205
rect 4798 6196 4804 6208
rect 4856 6196 4862 6248
rect 7561 6239 7619 6245
rect 7561 6205 7573 6239
rect 7607 6236 7619 6239
rect 8220 6236 8248 6403
rect 8478 6400 8484 6412
rect 8536 6400 8542 6452
rect 10410 6400 10416 6452
rect 10468 6440 10474 6452
rect 10505 6443 10563 6449
rect 10505 6440 10517 6443
rect 10468 6412 10517 6440
rect 10468 6400 10474 6412
rect 10505 6409 10517 6412
rect 10551 6409 10563 6443
rect 11238 6440 11244 6452
rect 11199 6412 11244 6440
rect 10505 6403 10563 6409
rect 11238 6400 11244 6412
rect 11296 6440 11302 6452
rect 12802 6440 12808 6452
rect 11296 6412 12808 6440
rect 11296 6400 11302 6412
rect 12802 6400 12808 6412
rect 12860 6400 12866 6452
rect 8846 6372 8852 6384
rect 8807 6344 8852 6372
rect 8846 6332 8852 6344
rect 8904 6332 8910 6384
rect 7607 6208 8248 6236
rect 8665 6239 8723 6245
rect 7607 6205 7619 6208
rect 7561 6199 7619 6205
rect 8665 6205 8677 6239
rect 8711 6236 8723 6239
rect 10321 6239 10379 6245
rect 8711 6208 9352 6236
rect 8711 6205 8723 6208
rect 8665 6199 8723 6205
rect 6270 6128 6276 6180
rect 6328 6128 6334 6180
rect 4338 6100 4344 6112
rect 4299 6072 4344 6100
rect 4338 6060 4344 6072
rect 4396 6060 4402 6112
rect 6086 6100 6092 6112
rect 6047 6072 6092 6100
rect 6086 6060 6092 6072
rect 6144 6100 6150 6112
rect 6288 6100 6316 6128
rect 6144 6072 6316 6100
rect 6144 6060 6150 6072
rect 6638 6060 6644 6112
rect 6696 6100 6702 6112
rect 9324 6109 9352 6208
rect 10321 6205 10333 6239
rect 10367 6236 10379 6239
rect 10367 6208 11008 6236
rect 10367 6205 10379 6208
rect 10321 6199 10379 6205
rect 10980 6112 11008 6208
rect 7745 6103 7803 6109
rect 7745 6100 7757 6103
rect 6696 6072 7757 6100
rect 6696 6060 6702 6072
rect 7745 6069 7757 6072
rect 7791 6069 7803 6103
rect 7745 6063 7803 6069
rect 9309 6103 9367 6109
rect 9309 6069 9321 6103
rect 9355 6100 9367 6103
rect 9398 6100 9404 6112
rect 9355 6072 9404 6100
rect 9355 6069 9367 6072
rect 9309 6063 9367 6069
rect 9398 6060 9404 6072
rect 9456 6060 9462 6112
rect 10962 6100 10968 6112
rect 10923 6072 10968 6100
rect 10962 6060 10968 6072
rect 11020 6060 11026 6112
rect 1104 6010 14812 6032
rect 1104 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 11648 6010
rect 11700 5958 11712 6010
rect 11764 5958 11776 6010
rect 11828 5958 11840 6010
rect 11892 5958 14812 6010
rect 1104 5936 14812 5958
rect 1104 5466 14812 5488
rect 1104 5414 3648 5466
rect 3700 5414 3712 5466
rect 3764 5414 3776 5466
rect 3828 5414 3840 5466
rect 3892 5414 8982 5466
rect 9034 5414 9046 5466
rect 9098 5414 9110 5466
rect 9162 5414 9174 5466
rect 9226 5414 14315 5466
rect 14367 5414 14379 5466
rect 14431 5414 14443 5466
rect 14495 5414 14507 5466
rect 14559 5414 14812 5466
rect 1104 5392 14812 5414
rect 1104 4922 14812 4944
rect 1104 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 11648 4922
rect 11700 4870 11712 4922
rect 11764 4870 11776 4922
rect 11828 4870 11840 4922
rect 11892 4870 14812 4922
rect 1104 4848 14812 4870
rect 1104 4378 14812 4400
rect 1104 4326 3648 4378
rect 3700 4326 3712 4378
rect 3764 4326 3776 4378
rect 3828 4326 3840 4378
rect 3892 4326 8982 4378
rect 9034 4326 9046 4378
rect 9098 4326 9110 4378
rect 9162 4326 9174 4378
rect 9226 4326 14315 4378
rect 14367 4326 14379 4378
rect 14431 4326 14443 4378
rect 14495 4326 14507 4378
rect 14559 4326 14812 4378
rect 1104 4304 14812 4326
rect 198 4088 204 4140
rect 256 4128 262 4140
rect 1210 4128 1216 4140
rect 256 4100 1216 4128
rect 256 4088 262 4100
rect 1210 4088 1216 4100
rect 1268 4088 1274 4140
rect 1104 3834 14812 3856
rect 1104 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 11648 3834
rect 11700 3782 11712 3834
rect 11764 3782 11776 3834
rect 11828 3782 11840 3834
rect 11892 3782 14812 3834
rect 1104 3760 14812 3782
rect 1118 3680 1124 3732
rect 1176 3720 1182 3732
rect 1581 3723 1639 3729
rect 1581 3720 1593 3723
rect 1176 3692 1593 3720
rect 1176 3680 1182 3692
rect 1581 3689 1593 3692
rect 1627 3689 1639 3723
rect 1581 3683 1639 3689
rect 4154 3680 4160 3732
rect 4212 3720 4218 3732
rect 4709 3723 4767 3729
rect 4709 3720 4721 3723
rect 4212 3692 4721 3720
rect 4212 3680 4218 3692
rect 4709 3689 4721 3692
rect 4755 3689 4767 3723
rect 4709 3683 4767 3689
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3584 1455 3587
rect 1670 3584 1676 3596
rect 1443 3556 1676 3584
rect 1443 3553 1455 3556
rect 1397 3547 1455 3553
rect 1670 3544 1676 3556
rect 1728 3544 1734 3596
rect 4525 3587 4583 3593
rect 4525 3553 4537 3587
rect 4571 3584 4583 3587
rect 4706 3584 4712 3596
rect 4571 3556 4712 3584
rect 4571 3553 4583 3556
rect 4525 3547 4583 3553
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 14642 3340 14648 3392
rect 14700 3380 14706 3392
rect 14921 3383 14979 3389
rect 14921 3380 14933 3383
rect 14700 3352 14933 3380
rect 14700 3340 14706 3352
rect 14921 3349 14933 3352
rect 14967 3349 14979 3383
rect 14921 3343 14979 3349
rect 1104 3290 14812 3312
rect 1104 3238 3648 3290
rect 3700 3238 3712 3290
rect 3764 3238 3776 3290
rect 3828 3238 3840 3290
rect 3892 3238 8982 3290
rect 9034 3238 9046 3290
rect 9098 3238 9110 3290
rect 9162 3238 9174 3290
rect 9226 3238 14315 3290
rect 14367 3238 14379 3290
rect 14431 3238 14443 3290
rect 14495 3238 14507 3290
rect 14559 3238 14812 3290
rect 1104 3216 14812 3238
rect 1670 3176 1676 3188
rect 1631 3148 1676 3176
rect 1670 3136 1676 3148
rect 1728 3136 1734 3188
rect 1762 3136 1768 3188
rect 1820 3176 1826 3188
rect 2222 3176 2228 3188
rect 1820 3148 2228 3176
rect 1820 3136 1826 3148
rect 2222 3136 2228 3148
rect 2280 3136 2286 3188
rect 2406 3176 2412 3188
rect 2367 3148 2412 3176
rect 2406 3136 2412 3148
rect 2464 3136 2470 3188
rect 4617 3179 4675 3185
rect 4617 3145 4629 3179
rect 4663 3176 4675 3179
rect 4706 3176 4712 3188
rect 4663 3148 4712 3176
rect 4663 3145 4675 3148
rect 4617 3139 4675 3145
rect 4706 3136 4712 3148
rect 4764 3136 4770 3188
rect 5629 3179 5687 3185
rect 5629 3145 5641 3179
rect 5675 3176 5687 3179
rect 5810 3176 5816 3188
rect 5675 3148 5816 3176
rect 5675 3145 5687 3148
rect 5629 3139 5687 3145
rect 1394 3068 1400 3120
rect 1452 3108 1458 3120
rect 2041 3111 2099 3117
rect 2041 3108 2053 3111
rect 1452 3080 2053 3108
rect 1452 3068 1458 3080
rect 2041 3077 2053 3080
rect 2087 3077 2099 3111
rect 2041 3071 2099 3077
rect 3326 3068 3332 3120
rect 3384 3108 3390 3120
rect 5169 3111 5227 3117
rect 5169 3108 5181 3111
rect 3384 3080 5181 3108
rect 3384 3068 3390 3080
rect 5169 3077 5181 3080
rect 5215 3077 5227 3111
rect 5169 3071 5227 3077
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2972 1915 2975
rect 2406 2972 2412 2984
rect 1903 2944 2412 2972
rect 1903 2941 1915 2944
rect 1857 2935 1915 2941
rect 2406 2932 2412 2944
rect 2464 2932 2470 2984
rect 4985 2975 5043 2981
rect 4985 2941 4997 2975
rect 5031 2972 5043 2975
rect 5644 2972 5672 3139
rect 5810 3136 5816 3148
rect 5868 3136 5874 3188
rect 9950 3176 9956 3188
rect 9911 3148 9956 3176
rect 9950 3136 9956 3148
rect 10008 3136 10014 3188
rect 10410 3176 10416 3188
rect 10371 3148 10416 3176
rect 10410 3136 10416 3148
rect 10468 3136 10474 3188
rect 13081 3179 13139 3185
rect 13081 3145 13093 3179
rect 13127 3176 13139 3179
rect 13906 3176 13912 3188
rect 13127 3148 13912 3176
rect 13127 3145 13139 3148
rect 13081 3139 13139 3145
rect 11422 3108 11428 3120
rect 11383 3080 11428 3108
rect 11422 3068 11428 3080
rect 11480 3068 11486 3120
rect 8662 2972 8668 2984
rect 5031 2944 5672 2972
rect 8623 2944 8668 2972
rect 5031 2941 5043 2944
rect 4985 2935 5043 2941
rect 8662 2932 8668 2944
rect 8720 2972 8726 2984
rect 9217 2975 9275 2981
rect 9217 2972 9229 2975
rect 8720 2944 9229 2972
rect 8720 2932 8726 2944
rect 9217 2941 9229 2944
rect 9263 2941 9275 2975
rect 9217 2935 9275 2941
rect 9769 2975 9827 2981
rect 9769 2941 9781 2975
rect 9815 2972 9827 2975
rect 10410 2972 10416 2984
rect 9815 2944 10416 2972
rect 9815 2941 9827 2944
rect 9769 2935 9827 2941
rect 10410 2932 10416 2944
rect 10468 2932 10474 2984
rect 11241 2975 11299 2981
rect 11241 2941 11253 2975
rect 11287 2941 11299 2975
rect 11241 2935 11299 2941
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2972 12495 2975
rect 13096 2972 13124 3139
rect 13906 3136 13912 3148
rect 13964 3136 13970 3188
rect 12483 2944 13124 2972
rect 12483 2941 12495 2944
rect 12437 2935 12495 2941
rect 11256 2904 11284 2935
rect 11885 2907 11943 2913
rect 11885 2904 11897 2907
rect 11256 2876 11897 2904
rect 11885 2873 11897 2876
rect 11931 2904 11943 2907
rect 14826 2904 14832 2916
rect 11931 2876 14832 2904
rect 11931 2873 11943 2876
rect 11885 2867 11943 2873
rect 14826 2864 14832 2876
rect 14884 2864 14890 2916
rect 8846 2836 8852 2848
rect 8807 2808 8852 2836
rect 8846 2796 8852 2808
rect 8904 2796 8910 2848
rect 12618 2836 12624 2848
rect 12579 2808 12624 2836
rect 12618 2796 12624 2808
rect 12676 2796 12682 2848
rect 1104 2746 14812 2768
rect 1104 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 11648 2746
rect 11700 2694 11712 2746
rect 11764 2694 11776 2746
rect 11828 2694 11840 2746
rect 11892 2694 14812 2746
rect 1104 2672 14812 2694
rect 2314 2632 2320 2644
rect 2275 2604 2320 2632
rect 2314 2592 2320 2604
rect 2372 2592 2378 2644
rect 2774 2592 2780 2644
rect 2832 2632 2838 2644
rect 3053 2635 3111 2641
rect 3053 2632 3065 2635
rect 2832 2604 3065 2632
rect 2832 2592 2838 2604
rect 3053 2601 3065 2604
rect 3099 2601 3111 2635
rect 5810 2632 5816 2644
rect 5771 2604 5816 2632
rect 3053 2595 3111 2601
rect 5810 2592 5816 2604
rect 5868 2592 5874 2644
rect 7098 2632 7104 2644
rect 7059 2604 7104 2632
rect 7098 2592 7104 2604
rect 7156 2592 7162 2644
rect 11422 2592 11428 2644
rect 11480 2632 11486 2644
rect 11609 2635 11667 2641
rect 11609 2632 11621 2635
rect 11480 2604 11621 2632
rect 11480 2592 11486 2604
rect 11609 2601 11621 2604
rect 11655 2601 11667 2635
rect 13262 2632 13268 2644
rect 13223 2604 13268 2632
rect 11609 2595 11667 2601
rect 13262 2592 13268 2604
rect 13320 2592 13326 2644
rect 1765 2499 1823 2505
rect 1765 2465 1777 2499
rect 1811 2496 1823 2499
rect 2332 2496 2360 2592
rect 6178 2564 6184 2576
rect 5644 2536 6184 2564
rect 1811 2468 2360 2496
rect 2869 2499 2927 2505
rect 1811 2465 1823 2468
rect 1765 2459 1823 2465
rect 2869 2465 2881 2499
rect 2915 2496 2927 2499
rect 3510 2496 3516 2508
rect 2915 2468 3516 2496
rect 2915 2465 2927 2468
rect 2869 2459 2927 2465
rect 3510 2456 3516 2468
rect 3568 2456 3574 2508
rect 4522 2496 4528 2508
rect 4483 2468 4528 2496
rect 4522 2456 4528 2468
rect 4580 2496 4586 2508
rect 5644 2505 5672 2536
rect 6178 2524 6184 2536
rect 6236 2524 6242 2576
rect 5077 2499 5135 2505
rect 5077 2496 5089 2499
rect 4580 2468 5089 2496
rect 4580 2456 4586 2468
rect 5077 2465 5089 2468
rect 5123 2465 5135 2499
rect 5077 2459 5135 2465
rect 5629 2499 5687 2505
rect 5629 2465 5641 2499
rect 5675 2465 5687 2499
rect 5629 2459 5687 2465
rect 6917 2499 6975 2505
rect 6917 2465 6929 2499
rect 6963 2496 6975 2499
rect 7558 2496 7564 2508
rect 6963 2468 7564 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 7558 2456 7564 2468
rect 7616 2456 7622 2508
rect 8573 2499 8631 2505
rect 8573 2465 8585 2499
rect 8619 2496 8631 2499
rect 9769 2499 9827 2505
rect 8619 2468 9260 2496
rect 8619 2465 8631 2468
rect 8573 2459 8631 2465
rect 934 2252 940 2304
rect 992 2292 998 2304
rect 1949 2295 2007 2301
rect 1949 2292 1961 2295
rect 992 2264 1961 2292
rect 992 2252 998 2264
rect 1949 2261 1961 2264
rect 1995 2261 2007 2295
rect 3510 2292 3516 2304
rect 3471 2264 3516 2292
rect 1949 2255 2007 2261
rect 3510 2252 3516 2264
rect 3568 2252 3574 2304
rect 3970 2252 3976 2304
rect 4028 2292 4034 2304
rect 4709 2295 4767 2301
rect 4709 2292 4721 2295
rect 4028 2264 4721 2292
rect 4028 2252 4034 2264
rect 4709 2261 4721 2264
rect 4755 2261 4767 2295
rect 7558 2292 7564 2304
rect 7519 2264 7564 2292
rect 4709 2255 4767 2261
rect 7558 2252 7564 2264
rect 7616 2252 7622 2304
rect 8754 2292 8760 2304
rect 8715 2264 8760 2292
rect 8754 2252 8760 2264
rect 8812 2252 8818 2304
rect 9232 2301 9260 2468
rect 9769 2465 9781 2499
rect 9815 2496 9827 2499
rect 10410 2496 10416 2508
rect 9815 2468 10416 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 10410 2456 10416 2468
rect 10468 2456 10474 2508
rect 11425 2499 11483 2505
rect 11425 2465 11437 2499
rect 11471 2496 11483 2499
rect 12066 2496 12072 2508
rect 11471 2468 12072 2496
rect 11471 2465 11483 2468
rect 11425 2459 11483 2465
rect 12066 2456 12072 2468
rect 12124 2456 12130 2508
rect 12621 2499 12679 2505
rect 12621 2465 12633 2499
rect 12667 2496 12679 2499
rect 13280 2496 13308 2592
rect 12667 2468 13308 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 12802 2360 12808 2372
rect 12763 2332 12808 2360
rect 12802 2320 12808 2332
rect 12860 2320 12866 2372
rect 9217 2295 9275 2301
rect 9217 2261 9229 2295
rect 9263 2292 9275 2295
rect 9398 2292 9404 2304
rect 9263 2264 9404 2292
rect 9263 2261 9275 2264
rect 9217 2255 9275 2261
rect 9398 2252 9404 2264
rect 9456 2252 9462 2304
rect 9950 2292 9956 2304
rect 9911 2264 9956 2292
rect 9950 2252 9956 2264
rect 10008 2252 10014 2304
rect 12066 2292 12072 2304
rect 12027 2264 12072 2292
rect 12066 2252 12072 2264
rect 12124 2252 12130 2304
rect 1104 2202 14812 2224
rect 1104 2150 3648 2202
rect 3700 2150 3712 2202
rect 3764 2150 3776 2202
rect 3828 2150 3840 2202
rect 3892 2150 8982 2202
rect 9034 2150 9046 2202
rect 9098 2150 9110 2202
rect 9162 2150 9174 2202
rect 9226 2150 14315 2202
rect 14367 2150 14379 2202
rect 14431 2150 14443 2202
rect 14495 2150 14507 2202
rect 14559 2150 14812 2202
rect 1104 2128 14812 2150
rect 12066 1844 12072 1896
rect 12124 1884 12130 1896
rect 14090 1884 14096 1896
rect 12124 1856 14096 1884
rect 12124 1844 12130 1856
rect 14090 1844 14096 1856
rect 14148 1844 14154 1896
rect 11054 1368 11060 1420
rect 11112 1408 11118 1420
rect 12158 1408 12164 1420
rect 11112 1380 12164 1408
rect 11112 1368 11118 1380
rect 12158 1368 12164 1380
rect 12216 1368 12222 1420
rect 13814 1368 13820 1420
rect 13872 1408 13878 1420
rect 14550 1408 14556 1420
rect 13872 1380 14556 1408
rect 13872 1368 13878 1380
rect 14550 1368 14556 1380
rect 14608 1368 14614 1420
rect 14918 592 14924 604
rect 14879 564 14924 592
rect 14918 552 14924 564
rect 14976 552 14982 604
<< via1 >>
rect 6315 37510 6367 37562
rect 6379 37510 6431 37562
rect 6443 37510 6495 37562
rect 6507 37510 6559 37562
rect 11648 37510 11700 37562
rect 11712 37510 11764 37562
rect 11776 37510 11828 37562
rect 11840 37510 11892 37562
rect 8392 37136 8444 37188
rect 8944 37136 8996 37188
rect 3648 36966 3700 37018
rect 3712 36966 3764 37018
rect 3776 36966 3828 37018
rect 3840 36966 3892 37018
rect 8982 36966 9034 37018
rect 9046 36966 9098 37018
rect 9110 36966 9162 37018
rect 9174 36966 9226 37018
rect 14315 36966 14367 37018
rect 14379 36966 14431 37018
rect 14443 36966 14495 37018
rect 14507 36966 14559 37018
rect 6315 36422 6367 36474
rect 6379 36422 6431 36474
rect 6443 36422 6495 36474
rect 6507 36422 6559 36474
rect 11648 36422 11700 36474
rect 11712 36422 11764 36474
rect 11776 36422 11828 36474
rect 11840 36422 11892 36474
rect 3648 35878 3700 35930
rect 3712 35878 3764 35930
rect 3776 35878 3828 35930
rect 3840 35878 3892 35930
rect 8982 35878 9034 35930
rect 9046 35878 9098 35930
rect 9110 35878 9162 35930
rect 9174 35878 9226 35930
rect 14315 35878 14367 35930
rect 14379 35878 14431 35930
rect 14443 35878 14495 35930
rect 14507 35878 14559 35930
rect 4528 35708 4580 35760
rect 5448 35708 5500 35760
rect 5724 35708 5776 35760
rect 6736 35708 6788 35760
rect 6184 35640 6236 35692
rect 6644 35640 6696 35692
rect 7196 35640 7248 35692
rect 8208 35640 8260 35692
rect 5080 35572 5132 35624
rect 5356 35572 5408 35624
rect 6315 35334 6367 35386
rect 6379 35334 6431 35386
rect 6443 35334 6495 35386
rect 6507 35334 6559 35386
rect 11648 35334 11700 35386
rect 11712 35334 11764 35386
rect 11776 35334 11828 35386
rect 11840 35334 11892 35386
rect 7380 35232 7432 35284
rect 8208 35232 8260 35284
rect 6920 35096 6972 35148
rect 8024 35096 8076 35148
rect 1400 34892 1452 34944
rect 2504 34892 2556 34944
rect 3648 34790 3700 34842
rect 3712 34790 3764 34842
rect 3776 34790 3828 34842
rect 3840 34790 3892 34842
rect 8982 34790 9034 34842
rect 9046 34790 9098 34842
rect 9110 34790 9162 34842
rect 9174 34790 9226 34842
rect 14315 34790 14367 34842
rect 14379 34790 14431 34842
rect 14443 34790 14495 34842
rect 14507 34790 14559 34842
rect 204 34552 256 34604
rect 1308 34552 1360 34604
rect 572 34484 624 34536
rect 1124 34484 1176 34536
rect 2136 34484 2188 34536
rect 2596 34484 2648 34536
rect 6315 34246 6367 34298
rect 6379 34246 6431 34298
rect 6443 34246 6495 34298
rect 6507 34246 6559 34298
rect 11648 34246 11700 34298
rect 11712 34246 11764 34298
rect 11776 34246 11828 34298
rect 11840 34246 11892 34298
rect 3648 33702 3700 33754
rect 3712 33702 3764 33754
rect 3776 33702 3828 33754
rect 3840 33702 3892 33754
rect 8982 33702 9034 33754
rect 9046 33702 9098 33754
rect 9110 33702 9162 33754
rect 9174 33702 9226 33754
rect 14315 33702 14367 33754
rect 14379 33702 14431 33754
rect 14443 33702 14495 33754
rect 14507 33702 14559 33754
rect 6315 33158 6367 33210
rect 6379 33158 6431 33210
rect 6443 33158 6495 33210
rect 6507 33158 6559 33210
rect 11648 33158 11700 33210
rect 11712 33158 11764 33210
rect 11776 33158 11828 33210
rect 11840 33158 11892 33210
rect 3648 32614 3700 32666
rect 3712 32614 3764 32666
rect 3776 32614 3828 32666
rect 3840 32614 3892 32666
rect 8982 32614 9034 32666
rect 9046 32614 9098 32666
rect 9110 32614 9162 32666
rect 9174 32614 9226 32666
rect 14315 32614 14367 32666
rect 14379 32614 14431 32666
rect 14443 32614 14495 32666
rect 14507 32614 14559 32666
rect 6315 32070 6367 32122
rect 6379 32070 6431 32122
rect 6443 32070 6495 32122
rect 6507 32070 6559 32122
rect 11648 32070 11700 32122
rect 11712 32070 11764 32122
rect 11776 32070 11828 32122
rect 11840 32070 11892 32122
rect 1400 31968 1452 32020
rect 4160 31968 4212 32020
rect 2228 31832 2280 31884
rect 4068 31875 4120 31884
rect 4068 31841 4077 31875
rect 4077 31841 4111 31875
rect 4111 31841 4120 31875
rect 4068 31832 4120 31841
rect 5172 31875 5224 31884
rect 5172 31841 5181 31875
rect 5181 31841 5215 31875
rect 5215 31841 5224 31875
rect 5172 31832 5224 31841
rect 1768 31628 1820 31680
rect 3648 31526 3700 31578
rect 3712 31526 3764 31578
rect 3776 31526 3828 31578
rect 3840 31526 3892 31578
rect 8982 31526 9034 31578
rect 9046 31526 9098 31578
rect 9110 31526 9162 31578
rect 9174 31526 9226 31578
rect 14315 31526 14367 31578
rect 14379 31526 14431 31578
rect 14443 31526 14495 31578
rect 14507 31526 14559 31578
rect 940 31424 992 31476
rect 8760 31467 8812 31476
rect 8760 31433 8769 31467
rect 8769 31433 8803 31467
rect 8803 31433 8812 31467
rect 8760 31424 8812 31433
rect 12440 31424 12492 31476
rect 1676 31220 1728 31272
rect 2228 31084 2280 31136
rect 4160 31127 4212 31136
rect 4160 31093 4169 31127
rect 4169 31093 4203 31127
rect 4203 31093 4212 31127
rect 4160 31084 4212 31093
rect 5172 31127 5224 31136
rect 5172 31093 5181 31127
rect 5181 31093 5215 31127
rect 5215 31093 5224 31127
rect 5172 31084 5224 31093
rect 12440 31263 12492 31272
rect 12440 31229 12449 31263
rect 12449 31229 12483 31263
rect 12483 31229 12492 31263
rect 12440 31220 12492 31229
rect 9404 31084 9456 31136
rect 6315 30982 6367 31034
rect 6379 30982 6431 31034
rect 6443 30982 6495 31034
rect 6507 30982 6559 31034
rect 11648 30982 11700 31034
rect 11712 30982 11764 31034
rect 11776 30982 11828 31034
rect 11840 30982 11892 31034
rect 9680 30719 9732 30728
rect 9680 30685 9689 30719
rect 9689 30685 9723 30719
rect 9723 30685 9732 30719
rect 9680 30676 9732 30685
rect 1676 30583 1728 30592
rect 1676 30549 1685 30583
rect 1685 30549 1719 30583
rect 1719 30549 1728 30583
rect 1676 30540 1728 30549
rect 9312 30583 9364 30592
rect 9312 30549 9321 30583
rect 9321 30549 9355 30583
rect 9355 30549 9364 30583
rect 9312 30540 9364 30549
rect 3648 30438 3700 30490
rect 3712 30438 3764 30490
rect 3776 30438 3828 30490
rect 3840 30438 3892 30490
rect 8982 30438 9034 30490
rect 9046 30438 9098 30490
rect 9110 30438 9162 30490
rect 9174 30438 9226 30490
rect 14315 30438 14367 30490
rect 14379 30438 14431 30490
rect 14443 30438 14495 30490
rect 14507 30438 14559 30490
rect 9772 30336 9824 30388
rect 9956 30336 10008 30388
rect 9312 30200 9364 30252
rect 9680 30175 9732 30184
rect 9680 30141 9689 30175
rect 9689 30141 9723 30175
rect 9723 30141 9732 30175
rect 9680 30132 9732 30141
rect 9772 30107 9824 30116
rect 8484 29996 8536 30048
rect 9772 30073 9781 30107
rect 9781 30073 9815 30107
rect 9815 30073 9824 30107
rect 9772 30064 9824 30073
rect 9588 29996 9640 30048
rect 6315 29894 6367 29946
rect 6379 29894 6431 29946
rect 6443 29894 6495 29946
rect 6507 29894 6559 29946
rect 11648 29894 11700 29946
rect 11712 29894 11764 29946
rect 11776 29894 11828 29946
rect 11840 29894 11892 29946
rect 9680 29792 9732 29844
rect 7380 29656 7432 29708
rect 9312 29656 9364 29708
rect 7656 29452 7708 29504
rect 9496 29452 9548 29504
rect 3648 29350 3700 29402
rect 3712 29350 3764 29402
rect 3776 29350 3828 29402
rect 3840 29350 3892 29402
rect 8982 29350 9034 29402
rect 9046 29350 9098 29402
rect 9110 29350 9162 29402
rect 9174 29350 9226 29402
rect 14315 29350 14367 29402
rect 14379 29350 14431 29402
rect 14443 29350 14495 29402
rect 14507 29350 14559 29402
rect 1952 29248 2004 29300
rect 2412 29087 2464 29096
rect 2412 29053 2421 29087
rect 2421 29053 2455 29087
rect 2455 29053 2464 29087
rect 2412 29044 2464 29053
rect 4436 28908 4488 28960
rect 5724 28908 5776 28960
rect 7380 28976 7432 29028
rect 7656 29019 7708 29028
rect 7656 28985 7665 29019
rect 7665 28985 7699 29019
rect 7699 28985 7708 29019
rect 7656 28976 7708 28985
rect 10324 28908 10376 28960
rect 10600 28908 10652 28960
rect 12716 28908 12768 28960
rect 12900 28908 12952 28960
rect 6315 28806 6367 28858
rect 6379 28806 6431 28858
rect 6443 28806 6495 28858
rect 6507 28806 6559 28858
rect 11648 28806 11700 28858
rect 11712 28806 11764 28858
rect 11776 28806 11828 28858
rect 11840 28806 11892 28858
rect 2412 28475 2464 28484
rect 2412 28441 2421 28475
rect 2421 28441 2455 28475
rect 2455 28441 2464 28475
rect 2412 28432 2464 28441
rect 3648 28262 3700 28314
rect 3712 28262 3764 28314
rect 3776 28262 3828 28314
rect 3840 28262 3892 28314
rect 8982 28262 9034 28314
rect 9046 28262 9098 28314
rect 9110 28262 9162 28314
rect 9174 28262 9226 28314
rect 14315 28262 14367 28314
rect 14379 28262 14431 28314
rect 14443 28262 14495 28314
rect 14507 28262 14559 28314
rect 4528 27999 4580 28008
rect 4528 27965 4537 27999
rect 4537 27965 4571 27999
rect 4571 27965 4580 27999
rect 4528 27956 4580 27965
rect 4436 27863 4488 27872
rect 4436 27829 4445 27863
rect 4445 27829 4479 27863
rect 4479 27829 4488 27863
rect 4436 27820 4488 27829
rect 5724 27820 5776 27872
rect 6315 27718 6367 27770
rect 6379 27718 6431 27770
rect 6443 27718 6495 27770
rect 6507 27718 6559 27770
rect 11648 27718 11700 27770
rect 11712 27718 11764 27770
rect 11776 27718 11828 27770
rect 11840 27718 11892 27770
rect 4344 27548 4396 27600
rect 4620 27548 4672 27600
rect 4528 27276 4580 27328
rect 5356 27276 5408 27328
rect 3648 27174 3700 27226
rect 3712 27174 3764 27226
rect 3776 27174 3828 27226
rect 3840 27174 3892 27226
rect 8982 27174 9034 27226
rect 9046 27174 9098 27226
rect 9110 27174 9162 27226
rect 9174 27174 9226 27226
rect 14315 27174 14367 27226
rect 14379 27174 14431 27226
rect 14443 27174 14495 27226
rect 14507 27174 14559 27226
rect 14096 27004 14148 27056
rect 14832 27004 14884 27056
rect 12532 26936 12584 26988
rect 13176 26936 13228 26988
rect 13912 26936 13964 26988
rect 15384 26936 15436 26988
rect 8576 26868 8628 26920
rect 9312 26868 9364 26920
rect 12808 26868 12860 26920
rect 13728 26868 13780 26920
rect 14004 26868 14056 26920
rect 14924 26868 14976 26920
rect 14096 26732 14148 26784
rect 15752 26732 15804 26784
rect 6315 26630 6367 26682
rect 6379 26630 6431 26682
rect 6443 26630 6495 26682
rect 6507 26630 6559 26682
rect 11648 26630 11700 26682
rect 11712 26630 11764 26682
rect 11776 26630 11828 26682
rect 11840 26630 11892 26682
rect 3648 26086 3700 26138
rect 3712 26086 3764 26138
rect 3776 26086 3828 26138
rect 3840 26086 3892 26138
rect 8982 26086 9034 26138
rect 9046 26086 9098 26138
rect 9110 26086 9162 26138
rect 9174 26086 9226 26138
rect 14315 26086 14367 26138
rect 14379 26086 14431 26138
rect 14443 26086 14495 26138
rect 14507 26086 14559 26138
rect 1584 26027 1636 26036
rect 1584 25993 1593 26027
rect 1593 25993 1627 26027
rect 1627 25993 1636 26027
rect 1584 25984 1636 25993
rect 1768 25644 1820 25696
rect 6315 25542 6367 25594
rect 6379 25542 6431 25594
rect 6443 25542 6495 25594
rect 6507 25542 6559 25594
rect 11648 25542 11700 25594
rect 11712 25542 11764 25594
rect 11776 25542 11828 25594
rect 11840 25542 11892 25594
rect 4068 25347 4120 25356
rect 4068 25313 4077 25347
rect 4077 25313 4111 25347
rect 4111 25313 4120 25347
rect 4068 25304 4120 25313
rect 4252 25211 4304 25220
rect 4252 25177 4261 25211
rect 4261 25177 4295 25211
rect 4295 25177 4304 25211
rect 4252 25168 4304 25177
rect 3648 24998 3700 25050
rect 3712 24998 3764 25050
rect 3776 24998 3828 25050
rect 3840 24998 3892 25050
rect 8982 24998 9034 25050
rect 9046 24998 9098 25050
rect 9110 24998 9162 25050
rect 9174 24998 9226 25050
rect 14315 24998 14367 25050
rect 14379 24998 14431 25050
rect 14443 24998 14495 25050
rect 14507 24998 14559 25050
rect 4068 24939 4120 24948
rect 4068 24905 4077 24939
rect 4077 24905 4111 24939
rect 4111 24905 4120 24939
rect 4068 24896 4120 24905
rect 6315 24454 6367 24506
rect 6379 24454 6431 24506
rect 6443 24454 6495 24506
rect 6507 24454 6559 24506
rect 11648 24454 11700 24506
rect 11712 24454 11764 24506
rect 11776 24454 11828 24506
rect 11840 24454 11892 24506
rect 5356 24352 5408 24404
rect 12072 24395 12124 24404
rect 12072 24361 12081 24395
rect 12081 24361 12115 24395
rect 12115 24361 12124 24395
rect 12072 24352 12124 24361
rect 6828 24216 6880 24268
rect 12072 24216 12124 24268
rect 3648 23910 3700 23962
rect 3712 23910 3764 23962
rect 3776 23910 3828 23962
rect 3840 23910 3892 23962
rect 8982 23910 9034 23962
rect 9046 23910 9098 23962
rect 9110 23910 9162 23962
rect 9174 23910 9226 23962
rect 14315 23910 14367 23962
rect 14379 23910 14431 23962
rect 14443 23910 14495 23962
rect 14507 23910 14559 23962
rect 6828 23468 6880 23520
rect 12072 23468 12124 23520
rect 6315 23366 6367 23418
rect 6379 23366 6431 23418
rect 6443 23366 6495 23418
rect 6507 23366 6559 23418
rect 11648 23366 11700 23418
rect 11712 23366 11764 23418
rect 11776 23366 11828 23418
rect 11840 23366 11892 23418
rect 9680 23264 9732 23316
rect 10784 23264 10836 23316
rect 9864 23196 9916 23248
rect 11980 23196 12032 23248
rect 9680 23128 9732 23180
rect 10140 23103 10192 23112
rect 10140 23069 10149 23103
rect 10149 23069 10183 23103
rect 10183 23069 10192 23103
rect 10140 23060 10192 23069
rect 10324 23060 10376 23112
rect 9680 22967 9732 22976
rect 9680 22933 9689 22967
rect 9689 22933 9723 22967
rect 9723 22933 9732 22967
rect 9680 22924 9732 22933
rect 3648 22822 3700 22874
rect 3712 22822 3764 22874
rect 3776 22822 3828 22874
rect 3840 22822 3892 22874
rect 8982 22822 9034 22874
rect 9046 22822 9098 22874
rect 9110 22822 9162 22874
rect 9174 22822 9226 22874
rect 14315 22822 14367 22874
rect 14379 22822 14431 22874
rect 14443 22822 14495 22874
rect 14507 22822 14559 22874
rect 10324 22720 10376 22772
rect 10784 22763 10836 22772
rect 10784 22729 10793 22763
rect 10793 22729 10827 22763
rect 10827 22729 10836 22763
rect 10784 22720 10836 22729
rect 10140 22652 10192 22704
rect 9864 22627 9916 22636
rect 9864 22593 9873 22627
rect 9873 22593 9907 22627
rect 9907 22593 9916 22627
rect 9864 22584 9916 22593
rect 10048 22627 10100 22636
rect 10048 22593 10057 22627
rect 10057 22593 10091 22627
rect 10091 22593 10100 22627
rect 10048 22584 10100 22593
rect 7564 22491 7616 22500
rect 7564 22457 7573 22491
rect 7573 22457 7607 22491
rect 7607 22457 7616 22491
rect 7564 22448 7616 22457
rect 8760 22380 8812 22432
rect 9772 22423 9824 22432
rect 9772 22389 9781 22423
rect 9781 22389 9815 22423
rect 9815 22389 9824 22423
rect 9772 22380 9824 22389
rect 6315 22278 6367 22330
rect 6379 22278 6431 22330
rect 6443 22278 6495 22330
rect 6507 22278 6559 22330
rect 11648 22278 11700 22330
rect 11712 22278 11764 22330
rect 11776 22278 11828 22330
rect 11840 22278 11892 22330
rect 10140 22176 10192 22228
rect 10048 22108 10100 22160
rect 6000 22083 6052 22092
rect 6000 22049 6009 22083
rect 6009 22049 6043 22083
rect 6043 22049 6052 22083
rect 6000 22040 6052 22049
rect 6092 22015 6144 22024
rect 6092 21981 6101 22015
rect 6101 21981 6135 22015
rect 6135 21981 6144 22015
rect 6092 21972 6144 21981
rect 6276 22015 6328 22024
rect 6276 21981 6285 22015
rect 6285 21981 6319 22015
rect 6319 21981 6328 22015
rect 6276 21972 6328 21981
rect 9404 21947 9456 21956
rect 9404 21913 9413 21947
rect 9413 21913 9447 21947
rect 9447 21913 9456 21947
rect 9404 21904 9456 21913
rect 5632 21879 5684 21888
rect 5632 21845 5641 21879
rect 5641 21845 5675 21879
rect 5675 21845 5684 21879
rect 5632 21836 5684 21845
rect 3648 21734 3700 21786
rect 3712 21734 3764 21786
rect 3776 21734 3828 21786
rect 3840 21734 3892 21786
rect 8982 21734 9034 21786
rect 9046 21734 9098 21786
rect 9110 21734 9162 21786
rect 9174 21734 9226 21786
rect 14315 21734 14367 21786
rect 14379 21734 14431 21786
rect 14443 21734 14495 21786
rect 14507 21734 14559 21786
rect 6000 21675 6052 21684
rect 6000 21641 6009 21675
rect 6009 21641 6043 21675
rect 6043 21641 6052 21675
rect 6000 21632 6052 21641
rect 6276 21632 6328 21684
rect 6000 21292 6052 21344
rect 6315 21190 6367 21242
rect 6379 21190 6431 21242
rect 6443 21190 6495 21242
rect 6507 21190 6559 21242
rect 11648 21190 11700 21242
rect 11712 21190 11764 21242
rect 11776 21190 11828 21242
rect 11840 21190 11892 21242
rect 5632 21088 5684 21140
rect 7012 21131 7064 21140
rect 7012 21097 7021 21131
rect 7021 21097 7055 21131
rect 7055 21097 7064 21131
rect 7012 21088 7064 21097
rect 3648 20646 3700 20698
rect 3712 20646 3764 20698
rect 3776 20646 3828 20698
rect 3840 20646 3892 20698
rect 8982 20646 9034 20698
rect 9046 20646 9098 20698
rect 9110 20646 9162 20698
rect 9174 20646 9226 20698
rect 14315 20646 14367 20698
rect 14379 20646 14431 20698
rect 14443 20646 14495 20698
rect 14507 20646 14559 20698
rect 7012 20408 7064 20460
rect 7656 20451 7708 20460
rect 7656 20417 7665 20451
rect 7665 20417 7699 20451
rect 7699 20417 7708 20451
rect 7656 20408 7708 20417
rect 8760 20383 8812 20392
rect 8760 20349 8769 20383
rect 8769 20349 8803 20383
rect 8803 20349 8812 20383
rect 8760 20340 8812 20349
rect 5172 20272 5224 20324
rect 7012 20247 7064 20256
rect 7012 20213 7021 20247
rect 7021 20213 7055 20247
rect 7055 20213 7064 20247
rect 7012 20204 7064 20213
rect 7380 20247 7432 20256
rect 7380 20213 7389 20247
rect 7389 20213 7423 20247
rect 7423 20213 7432 20247
rect 7380 20204 7432 20213
rect 8576 20247 8628 20256
rect 8576 20213 8585 20247
rect 8585 20213 8619 20247
rect 8619 20213 8628 20247
rect 8576 20204 8628 20213
rect 6315 20102 6367 20154
rect 6379 20102 6431 20154
rect 6443 20102 6495 20154
rect 6507 20102 6559 20154
rect 11648 20102 11700 20154
rect 11712 20102 11764 20154
rect 11776 20102 11828 20154
rect 11840 20102 11892 20154
rect 7656 20000 7708 20052
rect 12348 19907 12400 19916
rect 12348 19873 12357 19907
rect 12357 19873 12391 19907
rect 12391 19873 12400 19907
rect 12348 19864 12400 19873
rect 12440 19660 12492 19712
rect 3648 19558 3700 19610
rect 3712 19558 3764 19610
rect 3776 19558 3828 19610
rect 3840 19558 3892 19610
rect 8982 19558 9034 19610
rect 9046 19558 9098 19610
rect 9110 19558 9162 19610
rect 9174 19558 9226 19610
rect 14315 19558 14367 19610
rect 14379 19558 14431 19610
rect 14443 19558 14495 19610
rect 14507 19558 14559 19610
rect 10416 19320 10468 19372
rect 10600 19320 10652 19372
rect 12348 19320 12400 19372
rect 12716 19320 12768 19372
rect 12992 19320 13044 19372
rect 3148 19252 3200 19304
rect 3424 19252 3476 19304
rect 14188 19252 14240 19304
rect 4344 19184 4396 19236
rect 4528 19184 4580 19236
rect 6315 19014 6367 19066
rect 6379 19014 6431 19066
rect 6443 19014 6495 19066
rect 6507 19014 6559 19066
rect 11648 19014 11700 19066
rect 11712 19014 11764 19066
rect 11776 19014 11828 19066
rect 11840 19014 11892 19066
rect 3648 18470 3700 18522
rect 3712 18470 3764 18522
rect 3776 18470 3828 18522
rect 3840 18470 3892 18522
rect 8982 18470 9034 18522
rect 9046 18470 9098 18522
rect 9110 18470 9162 18522
rect 9174 18470 9226 18522
rect 14315 18470 14367 18522
rect 14379 18470 14431 18522
rect 14443 18470 14495 18522
rect 14507 18470 14559 18522
rect 6315 17926 6367 17978
rect 6379 17926 6431 17978
rect 6443 17926 6495 17978
rect 6507 17926 6559 17978
rect 11648 17926 11700 17978
rect 11712 17926 11764 17978
rect 11776 17926 11828 17978
rect 11840 17926 11892 17978
rect 3648 17382 3700 17434
rect 3712 17382 3764 17434
rect 3776 17382 3828 17434
rect 3840 17382 3892 17434
rect 8982 17382 9034 17434
rect 9046 17382 9098 17434
rect 9110 17382 9162 17434
rect 9174 17382 9226 17434
rect 14315 17382 14367 17434
rect 14379 17382 14431 17434
rect 14443 17382 14495 17434
rect 14507 17382 14559 17434
rect 6315 16838 6367 16890
rect 6379 16838 6431 16890
rect 6443 16838 6495 16890
rect 6507 16838 6559 16890
rect 11648 16838 11700 16890
rect 11712 16838 11764 16890
rect 11776 16838 11828 16890
rect 11840 16838 11892 16890
rect 4436 16779 4488 16788
rect 4436 16745 4445 16779
rect 4445 16745 4479 16779
rect 4479 16745 4488 16779
rect 4436 16736 4488 16745
rect 12256 16736 12308 16788
rect 1952 16600 2004 16652
rect 2228 16600 2280 16652
rect 11520 16643 11572 16652
rect 11520 16609 11529 16643
rect 11529 16609 11563 16643
rect 11563 16609 11572 16643
rect 11520 16600 11572 16609
rect 11612 16600 11664 16652
rect 3648 16294 3700 16346
rect 3712 16294 3764 16346
rect 3776 16294 3828 16346
rect 3840 16294 3892 16346
rect 8982 16294 9034 16346
rect 9046 16294 9098 16346
rect 9110 16294 9162 16346
rect 9174 16294 9226 16346
rect 14315 16294 14367 16346
rect 14379 16294 14431 16346
rect 14443 16294 14495 16346
rect 14507 16294 14559 16346
rect 11520 16192 11572 16244
rect 4436 16056 4488 16108
rect 4988 16099 5040 16108
rect 4988 16065 4997 16099
rect 4997 16065 5031 16099
rect 5031 16065 5040 16099
rect 4988 16056 5040 16065
rect 4804 16031 4856 16040
rect 4804 15997 4813 16031
rect 4813 15997 4847 16031
rect 4847 15997 4856 16031
rect 4804 15988 4856 15997
rect 4344 15963 4396 15972
rect 4344 15929 4353 15963
rect 4353 15929 4387 15963
rect 4387 15929 4396 15963
rect 4344 15920 4396 15929
rect 4436 15895 4488 15904
rect 4436 15861 4445 15895
rect 4445 15861 4479 15895
rect 4479 15861 4488 15895
rect 4436 15852 4488 15861
rect 4896 15895 4948 15904
rect 4896 15861 4905 15895
rect 4905 15861 4939 15895
rect 4939 15861 4948 15895
rect 4896 15852 4948 15861
rect 11060 15852 11112 15904
rect 11612 15920 11664 15972
rect 6315 15750 6367 15802
rect 6379 15750 6431 15802
rect 6443 15750 6495 15802
rect 6507 15750 6559 15802
rect 11648 15750 11700 15802
rect 11712 15750 11764 15802
rect 11776 15750 11828 15802
rect 11840 15750 11892 15802
rect 4436 15648 4488 15700
rect 5724 15648 5776 15700
rect 7012 15648 7064 15700
rect 4804 15580 4856 15632
rect 5540 15555 5592 15564
rect 5540 15521 5549 15555
rect 5549 15521 5583 15555
rect 5583 15521 5592 15555
rect 5540 15512 5592 15521
rect 5632 15444 5684 15496
rect 5172 15351 5224 15360
rect 5172 15317 5181 15351
rect 5181 15317 5215 15351
rect 5215 15317 5224 15351
rect 5172 15308 5224 15317
rect 3648 15206 3700 15258
rect 3712 15206 3764 15258
rect 3776 15206 3828 15258
rect 3840 15206 3892 15258
rect 8982 15206 9034 15258
rect 9046 15206 9098 15258
rect 9110 15206 9162 15258
rect 9174 15206 9226 15258
rect 14315 15206 14367 15258
rect 14379 15206 14431 15258
rect 14443 15206 14495 15258
rect 14507 15206 14559 15258
rect 1584 15147 1636 15156
rect 1584 15113 1593 15147
rect 1593 15113 1627 15147
rect 1627 15113 1636 15147
rect 1584 15104 1636 15113
rect 2044 15147 2096 15156
rect 2044 15113 2053 15147
rect 2053 15113 2087 15147
rect 2087 15113 2096 15147
rect 2044 15104 2096 15113
rect 5632 15104 5684 15156
rect 5724 15104 5776 15156
rect 8576 15104 8628 15156
rect 4988 15011 5040 15020
rect 4988 14977 4997 15011
rect 4997 14977 5031 15011
rect 5031 14977 5040 15011
rect 4988 14968 5040 14977
rect 2044 14900 2096 14952
rect 4804 14943 4856 14952
rect 4804 14909 4813 14943
rect 4813 14909 4847 14943
rect 4847 14909 4856 14943
rect 4804 14900 4856 14909
rect 7012 14900 7064 14952
rect 9588 14900 9640 14952
rect 4344 14875 4396 14884
rect 4344 14841 4353 14875
rect 4353 14841 4387 14875
rect 4387 14841 4396 14875
rect 4344 14832 4396 14841
rect 7196 14832 7248 14884
rect 4436 14807 4488 14816
rect 4436 14773 4445 14807
rect 4445 14773 4479 14807
rect 4479 14773 4488 14807
rect 4436 14764 4488 14773
rect 4896 14807 4948 14816
rect 4896 14773 4905 14807
rect 4905 14773 4939 14807
rect 4939 14773 4948 14807
rect 7288 14807 7340 14816
rect 4896 14764 4948 14773
rect 7288 14773 7297 14807
rect 7297 14773 7331 14807
rect 7331 14773 7340 14807
rect 7288 14764 7340 14773
rect 10876 14807 10928 14816
rect 10876 14773 10885 14807
rect 10885 14773 10919 14807
rect 10919 14773 10928 14807
rect 10876 14764 10928 14773
rect 6315 14662 6367 14714
rect 6379 14662 6431 14714
rect 6443 14662 6495 14714
rect 6507 14662 6559 14714
rect 11648 14662 11700 14714
rect 11712 14662 11764 14714
rect 11776 14662 11828 14714
rect 11840 14662 11892 14714
rect 4436 14560 4488 14612
rect 5540 14560 5592 14612
rect 7196 14560 7248 14612
rect 8024 14603 8076 14612
rect 8024 14569 8033 14603
rect 8033 14569 8067 14603
rect 8067 14569 8076 14603
rect 8024 14560 8076 14569
rect 4804 14492 4856 14544
rect 3648 14118 3700 14170
rect 3712 14118 3764 14170
rect 3776 14118 3828 14170
rect 3840 14118 3892 14170
rect 8982 14118 9034 14170
rect 9046 14118 9098 14170
rect 9110 14118 9162 14170
rect 9174 14118 9226 14170
rect 14315 14118 14367 14170
rect 14379 14118 14431 14170
rect 14443 14118 14495 14170
rect 14507 14118 14559 14170
rect 10876 13880 10928 13932
rect 1860 13812 1912 13864
rect 8024 13744 8076 13796
rect 2228 13719 2280 13728
rect 2228 13685 2237 13719
rect 2237 13685 2271 13719
rect 2271 13685 2280 13719
rect 2228 13676 2280 13685
rect 7932 13719 7984 13728
rect 7932 13685 7941 13719
rect 7941 13685 7975 13719
rect 7975 13685 7984 13719
rect 7932 13676 7984 13685
rect 8300 13719 8352 13728
rect 8300 13685 8309 13719
rect 8309 13685 8343 13719
rect 8343 13685 8352 13719
rect 8300 13676 8352 13685
rect 6315 13574 6367 13626
rect 6379 13574 6431 13626
rect 6443 13574 6495 13626
rect 6507 13574 6559 13626
rect 11648 13574 11700 13626
rect 11712 13574 11764 13626
rect 11776 13574 11828 13626
rect 11840 13574 11892 13626
rect 7288 13472 7340 13524
rect 8024 13472 8076 13524
rect 3648 13030 3700 13082
rect 3712 13030 3764 13082
rect 3776 13030 3828 13082
rect 3840 13030 3892 13082
rect 8982 13030 9034 13082
rect 9046 13030 9098 13082
rect 9110 13030 9162 13082
rect 9174 13030 9226 13082
rect 14315 13030 14367 13082
rect 14379 13030 14431 13082
rect 14443 13030 14495 13082
rect 14507 13030 14559 13082
rect 8944 12860 8996 12912
rect 9404 12860 9456 12912
rect 6315 12486 6367 12538
rect 6379 12486 6431 12538
rect 6443 12486 6495 12538
rect 6507 12486 6559 12538
rect 11648 12486 11700 12538
rect 11712 12486 11764 12538
rect 11776 12486 11828 12538
rect 11840 12486 11892 12538
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 1584 12223 1636 12232
rect 1584 12189 1593 12223
rect 1593 12189 1627 12223
rect 1627 12189 1636 12223
rect 1584 12180 1636 12189
rect 3648 11942 3700 11994
rect 3712 11942 3764 11994
rect 3776 11942 3828 11994
rect 3840 11942 3892 11994
rect 8982 11942 9034 11994
rect 9046 11942 9098 11994
rect 9110 11942 9162 11994
rect 9174 11942 9226 11994
rect 14315 11942 14367 11994
rect 14379 11942 14431 11994
rect 14443 11942 14495 11994
rect 14507 11942 14559 11994
rect 1400 11840 1452 11892
rect 6315 11398 6367 11450
rect 6379 11398 6431 11450
rect 6443 11398 6495 11450
rect 6507 11398 6559 11450
rect 11648 11398 11700 11450
rect 11712 11398 11764 11450
rect 11776 11398 11828 11450
rect 11840 11398 11892 11450
rect 2320 11160 2372 11212
rect 1216 11024 1268 11076
rect 3648 10854 3700 10906
rect 3712 10854 3764 10906
rect 3776 10854 3828 10906
rect 3840 10854 3892 10906
rect 8982 10854 9034 10906
rect 9046 10854 9098 10906
rect 9110 10854 9162 10906
rect 9174 10854 9226 10906
rect 14315 10854 14367 10906
rect 14379 10854 14431 10906
rect 14443 10854 14495 10906
rect 14507 10854 14559 10906
rect 2320 10752 2372 10804
rect 2044 10616 2096 10668
rect 2320 10616 2372 10668
rect 14096 10752 14148 10804
rect 6920 10412 6972 10464
rect 8208 10412 8260 10464
rect 12440 10412 12492 10464
rect 6315 10310 6367 10362
rect 6379 10310 6431 10362
rect 6443 10310 6495 10362
rect 6507 10310 6559 10362
rect 11648 10310 11700 10362
rect 11712 10310 11764 10362
rect 11776 10310 11828 10362
rect 11840 10310 11892 10362
rect 3648 9766 3700 9818
rect 3712 9766 3764 9818
rect 3776 9766 3828 9818
rect 3840 9766 3892 9818
rect 8982 9766 9034 9818
rect 9046 9766 9098 9818
rect 9110 9766 9162 9818
rect 9174 9766 9226 9818
rect 14315 9766 14367 9818
rect 14379 9766 14431 9818
rect 14443 9766 14495 9818
rect 14507 9766 14559 9818
rect 3148 9664 3200 9716
rect 3424 9664 3476 9716
rect 14740 9664 14792 9716
rect 2596 9596 2648 9648
rect 3516 9392 3568 9444
rect 6315 9222 6367 9274
rect 6379 9222 6431 9274
rect 6443 9222 6495 9274
rect 6507 9222 6559 9274
rect 11648 9222 11700 9274
rect 11712 9222 11764 9274
rect 11776 9222 11828 9274
rect 11840 9222 11892 9274
rect 10600 9163 10652 9172
rect 10600 9129 10609 9163
rect 10609 9129 10643 9163
rect 10643 9129 10652 9163
rect 10600 9120 10652 9129
rect 12532 9163 12584 9172
rect 12532 9129 12541 9163
rect 12541 9129 12575 9163
rect 12575 9129 12584 9163
rect 12532 9120 12584 9129
rect 10508 8984 10560 9036
rect 13084 8984 13136 9036
rect 3648 8678 3700 8730
rect 3712 8678 3764 8730
rect 3776 8678 3828 8730
rect 3840 8678 3892 8730
rect 8982 8678 9034 8730
rect 9046 8678 9098 8730
rect 9110 8678 9162 8730
rect 9174 8678 9226 8730
rect 14315 8678 14367 8730
rect 14379 8678 14431 8730
rect 14443 8678 14495 8730
rect 14507 8678 14559 8730
rect 14004 8372 14056 8424
rect 10508 8347 10560 8356
rect 10508 8313 10517 8347
rect 10517 8313 10551 8347
rect 10551 8313 10560 8347
rect 10508 8304 10560 8313
rect 13084 8347 13136 8356
rect 13084 8313 13093 8347
rect 13093 8313 13127 8347
rect 13127 8313 13136 8347
rect 13084 8304 13136 8313
rect 12624 8279 12676 8288
rect 12624 8245 12633 8279
rect 12633 8245 12667 8279
rect 12667 8245 12676 8279
rect 12624 8236 12676 8245
rect 6315 8134 6367 8186
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 11648 8134 11700 8186
rect 11712 8134 11764 8186
rect 11776 8134 11828 8186
rect 11840 8134 11892 8186
rect 3424 8032 3476 8084
rect 4896 7896 4948 7948
rect 3648 7590 3700 7642
rect 3712 7590 3764 7642
rect 3776 7590 3828 7642
rect 3840 7590 3892 7642
rect 8982 7590 9034 7642
rect 9046 7590 9098 7642
rect 9110 7590 9162 7642
rect 9174 7590 9226 7642
rect 14315 7590 14367 7642
rect 14379 7590 14431 7642
rect 14443 7590 14495 7642
rect 14507 7590 14559 7642
rect 7472 7531 7524 7540
rect 7472 7497 7481 7531
rect 7481 7497 7515 7531
rect 7515 7497 7524 7531
rect 7472 7488 7524 7497
rect 7472 7284 7524 7336
rect 4896 7148 4948 7200
rect 7012 7191 7064 7200
rect 7012 7157 7021 7191
rect 7021 7157 7055 7191
rect 7055 7157 7064 7191
rect 7012 7148 7064 7157
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 11648 7046 11700 7098
rect 11712 7046 11764 7098
rect 11776 7046 11828 7098
rect 11840 7046 11892 7098
rect 1584 6851 1636 6860
rect 1584 6817 1593 6851
rect 1593 6817 1627 6851
rect 1627 6817 1636 6851
rect 1584 6808 1636 6817
rect 6276 6808 6328 6860
rect 11244 6808 11296 6860
rect 6184 6715 6236 6724
rect 6184 6681 6193 6715
rect 6193 6681 6227 6715
rect 6227 6681 6236 6715
rect 6184 6672 6236 6681
rect 572 6604 624 6656
rect 10600 6647 10652 6656
rect 10600 6613 10609 6647
rect 10609 6613 10643 6647
rect 10643 6613 10652 6647
rect 10600 6604 10652 6613
rect 3648 6502 3700 6554
rect 3712 6502 3764 6554
rect 3776 6502 3828 6554
rect 3840 6502 3892 6554
rect 8982 6502 9034 6554
rect 9046 6502 9098 6554
rect 9110 6502 9162 6554
rect 9174 6502 9226 6554
rect 14315 6502 14367 6554
rect 14379 6502 14431 6554
rect 14443 6502 14495 6554
rect 14507 6502 14559 6554
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 4804 6239 4856 6248
rect 4804 6205 4813 6239
rect 4813 6205 4847 6239
rect 4847 6205 4856 6239
rect 4804 6196 4856 6205
rect 8484 6400 8536 6452
rect 10416 6400 10468 6452
rect 11244 6443 11296 6452
rect 11244 6409 11253 6443
rect 11253 6409 11287 6443
rect 11287 6409 11296 6443
rect 11244 6400 11296 6409
rect 12808 6400 12860 6452
rect 8852 6375 8904 6384
rect 8852 6341 8861 6375
rect 8861 6341 8895 6375
rect 8895 6341 8904 6375
rect 8852 6332 8904 6341
rect 6276 6128 6328 6180
rect 4344 6103 4396 6112
rect 4344 6069 4353 6103
rect 4353 6069 4387 6103
rect 4387 6069 4396 6103
rect 4344 6060 4396 6069
rect 6092 6103 6144 6112
rect 6092 6069 6101 6103
rect 6101 6069 6135 6103
rect 6135 6069 6144 6103
rect 6092 6060 6144 6069
rect 6644 6060 6696 6112
rect 9404 6060 9456 6112
rect 10968 6103 11020 6112
rect 10968 6069 10977 6103
rect 10977 6069 11011 6103
rect 11011 6069 11020 6103
rect 10968 6060 11020 6069
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 11648 5958 11700 6010
rect 11712 5958 11764 6010
rect 11776 5958 11828 6010
rect 11840 5958 11892 6010
rect 3648 5414 3700 5466
rect 3712 5414 3764 5466
rect 3776 5414 3828 5466
rect 3840 5414 3892 5466
rect 8982 5414 9034 5466
rect 9046 5414 9098 5466
rect 9110 5414 9162 5466
rect 9174 5414 9226 5466
rect 14315 5414 14367 5466
rect 14379 5414 14431 5466
rect 14443 5414 14495 5466
rect 14507 5414 14559 5466
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 11648 4870 11700 4922
rect 11712 4870 11764 4922
rect 11776 4870 11828 4922
rect 11840 4870 11892 4922
rect 3648 4326 3700 4378
rect 3712 4326 3764 4378
rect 3776 4326 3828 4378
rect 3840 4326 3892 4378
rect 8982 4326 9034 4378
rect 9046 4326 9098 4378
rect 9110 4326 9162 4378
rect 9174 4326 9226 4378
rect 14315 4326 14367 4378
rect 14379 4326 14431 4378
rect 14443 4326 14495 4378
rect 14507 4326 14559 4378
rect 204 4088 256 4140
rect 1216 4088 1268 4140
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 11648 3782 11700 3834
rect 11712 3782 11764 3834
rect 11776 3782 11828 3834
rect 11840 3782 11892 3834
rect 1124 3680 1176 3732
rect 4160 3680 4212 3732
rect 1676 3544 1728 3596
rect 4712 3544 4764 3596
rect 14648 3340 14700 3392
rect 3648 3238 3700 3290
rect 3712 3238 3764 3290
rect 3776 3238 3828 3290
rect 3840 3238 3892 3290
rect 8982 3238 9034 3290
rect 9046 3238 9098 3290
rect 9110 3238 9162 3290
rect 9174 3238 9226 3290
rect 14315 3238 14367 3290
rect 14379 3238 14431 3290
rect 14443 3238 14495 3290
rect 14507 3238 14559 3290
rect 1676 3179 1728 3188
rect 1676 3145 1685 3179
rect 1685 3145 1719 3179
rect 1719 3145 1728 3179
rect 1676 3136 1728 3145
rect 1768 3136 1820 3188
rect 2228 3136 2280 3188
rect 2412 3179 2464 3188
rect 2412 3145 2421 3179
rect 2421 3145 2455 3179
rect 2455 3145 2464 3179
rect 2412 3136 2464 3145
rect 4712 3136 4764 3188
rect 1400 3068 1452 3120
rect 3332 3068 3384 3120
rect 2412 2932 2464 2984
rect 5816 3136 5868 3188
rect 9956 3179 10008 3188
rect 9956 3145 9965 3179
rect 9965 3145 9999 3179
rect 9999 3145 10008 3179
rect 9956 3136 10008 3145
rect 10416 3179 10468 3188
rect 10416 3145 10425 3179
rect 10425 3145 10459 3179
rect 10459 3145 10468 3179
rect 10416 3136 10468 3145
rect 11428 3111 11480 3120
rect 11428 3077 11437 3111
rect 11437 3077 11471 3111
rect 11471 3077 11480 3111
rect 11428 3068 11480 3077
rect 8668 2975 8720 2984
rect 8668 2941 8677 2975
rect 8677 2941 8711 2975
rect 8711 2941 8720 2975
rect 8668 2932 8720 2941
rect 10416 2932 10468 2984
rect 13912 3136 13964 3188
rect 14832 2864 14884 2916
rect 8852 2839 8904 2848
rect 8852 2805 8861 2839
rect 8861 2805 8895 2839
rect 8895 2805 8904 2839
rect 8852 2796 8904 2805
rect 12624 2839 12676 2848
rect 12624 2805 12633 2839
rect 12633 2805 12667 2839
rect 12667 2805 12676 2839
rect 12624 2796 12676 2805
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 11648 2694 11700 2746
rect 11712 2694 11764 2746
rect 11776 2694 11828 2746
rect 11840 2694 11892 2746
rect 2320 2635 2372 2644
rect 2320 2601 2329 2635
rect 2329 2601 2363 2635
rect 2363 2601 2372 2635
rect 2320 2592 2372 2601
rect 2780 2592 2832 2644
rect 5816 2635 5868 2644
rect 5816 2601 5825 2635
rect 5825 2601 5859 2635
rect 5859 2601 5868 2635
rect 5816 2592 5868 2601
rect 7104 2635 7156 2644
rect 7104 2601 7113 2635
rect 7113 2601 7147 2635
rect 7147 2601 7156 2635
rect 7104 2592 7156 2601
rect 11428 2592 11480 2644
rect 13268 2635 13320 2644
rect 13268 2601 13277 2635
rect 13277 2601 13311 2635
rect 13311 2601 13320 2635
rect 13268 2592 13320 2601
rect 6184 2567 6236 2576
rect 3516 2456 3568 2508
rect 4528 2499 4580 2508
rect 4528 2465 4537 2499
rect 4537 2465 4571 2499
rect 4571 2465 4580 2499
rect 6184 2533 6193 2567
rect 6193 2533 6227 2567
rect 6227 2533 6236 2567
rect 6184 2524 6236 2533
rect 4528 2456 4580 2465
rect 7564 2456 7616 2508
rect 940 2252 992 2304
rect 3516 2295 3568 2304
rect 3516 2261 3525 2295
rect 3525 2261 3559 2295
rect 3559 2261 3568 2295
rect 3516 2252 3568 2261
rect 3976 2252 4028 2304
rect 7564 2295 7616 2304
rect 7564 2261 7573 2295
rect 7573 2261 7607 2295
rect 7607 2261 7616 2295
rect 7564 2252 7616 2261
rect 8760 2295 8812 2304
rect 8760 2261 8769 2295
rect 8769 2261 8803 2295
rect 8803 2261 8812 2295
rect 8760 2252 8812 2261
rect 10416 2499 10468 2508
rect 10416 2465 10425 2499
rect 10425 2465 10459 2499
rect 10459 2465 10468 2499
rect 10416 2456 10468 2465
rect 12072 2456 12124 2508
rect 12808 2363 12860 2372
rect 12808 2329 12817 2363
rect 12817 2329 12851 2363
rect 12851 2329 12860 2363
rect 12808 2320 12860 2329
rect 9404 2252 9456 2304
rect 9956 2295 10008 2304
rect 9956 2261 9965 2295
rect 9965 2261 9999 2295
rect 9999 2261 10008 2295
rect 9956 2252 10008 2261
rect 12072 2295 12124 2304
rect 12072 2261 12081 2295
rect 12081 2261 12115 2295
rect 12115 2261 12124 2295
rect 12072 2252 12124 2261
rect 3648 2150 3700 2202
rect 3712 2150 3764 2202
rect 3776 2150 3828 2202
rect 3840 2150 3892 2202
rect 8982 2150 9034 2202
rect 9046 2150 9098 2202
rect 9110 2150 9162 2202
rect 9174 2150 9226 2202
rect 14315 2150 14367 2202
rect 14379 2150 14431 2202
rect 14443 2150 14495 2202
rect 14507 2150 14559 2202
rect 12072 1844 12124 1896
rect 14096 1844 14148 1896
rect 11060 1368 11112 1420
rect 12164 1368 12216 1420
rect 13820 1368 13872 1420
rect 14556 1368 14608 1420
rect 14924 595 14976 604
rect 14924 561 14933 595
rect 14933 561 14967 595
rect 14967 561 14976 595
rect 14924 552 14976 561
<< metal2 >>
rect 202 39520 258 40000
rect 570 39520 626 40000
rect 938 39520 994 40000
rect 1398 39520 1454 40000
rect 1766 39520 1822 40000
rect 2134 39520 2190 40000
rect 2594 39520 2650 40000
rect 2962 39522 3018 40000
rect 2962 39520 3096 39522
rect 3330 39520 3386 40000
rect 3790 39520 3846 40000
rect 4158 39520 4214 40000
rect 4526 39520 4582 40000
rect 4986 39520 5042 40000
rect 5354 39520 5410 40000
rect 5722 39520 5778 40000
rect 6182 39520 6238 40000
rect 6550 39520 6606 40000
rect 6918 39520 6974 40000
rect 7378 39520 7434 40000
rect 7746 39520 7802 40000
rect 8206 39520 8262 40000
rect 8574 39520 8630 40000
rect 8942 39520 8998 40000
rect 9402 39520 9458 40000
rect 9770 39520 9826 40000
rect 10138 39522 10194 40000
rect 10598 39522 10654 40000
rect 9876 39520 10194 39522
rect 10336 39520 10654 39522
rect 10966 39520 11022 40000
rect 11334 39520 11390 40000
rect 11794 39520 11850 40000
rect 12162 39522 12218 40000
rect 11992 39520 12218 39522
rect 12530 39520 12586 40000
rect 12990 39520 13046 40000
rect 13358 39520 13414 40000
rect 13726 39520 13782 40000
rect 14186 39522 14242 40000
rect 14108 39520 14242 39522
rect 14554 39520 14610 40000
rect 14922 39520 14978 40000
rect 15382 39520 15438 40000
rect 15750 39520 15806 40000
rect 216 34610 244 39520
rect 204 34604 256 34610
rect 204 34546 256 34552
rect 584 34542 612 39520
rect 572 34536 624 34542
rect 572 34478 624 34484
rect 952 31482 980 39520
rect 1412 34950 1440 39520
rect 1400 34944 1452 34950
rect 1400 34886 1452 34892
rect 1308 34604 1360 34610
rect 1308 34546 1360 34552
rect 1124 34536 1176 34542
rect 1124 34478 1176 34484
rect 940 31476 992 31482
rect 940 31418 992 31424
rect 572 6656 624 6662
rect 572 6598 624 6604
rect 204 4140 256 4146
rect 204 4082 256 4088
rect 216 480 244 4082
rect 584 480 612 6598
rect 1136 3738 1164 34478
rect 1320 33266 1348 34546
rect 1320 33238 1440 33266
rect 1412 32026 1440 33238
rect 1400 32020 1452 32026
rect 1400 31962 1452 31968
rect 1780 31686 1808 39520
rect 1950 36680 2006 36689
rect 1950 36615 2006 36624
rect 1768 31680 1820 31686
rect 1768 31622 1820 31628
rect 1676 31272 1728 31278
rect 1676 31214 1728 31220
rect 1688 30598 1716 31214
rect 1676 30592 1728 30598
rect 1676 30534 1728 30540
rect 1582 30016 1638 30025
rect 1582 29951 1638 29960
rect 1596 26042 1624 29951
rect 1584 26036 1636 26042
rect 1584 25978 1636 25984
rect 1582 16688 1638 16697
rect 1582 16623 1638 16632
rect 1596 15162 1624 16623
rect 1584 15156 1636 15162
rect 1584 15098 1636 15104
rect 1688 15065 1716 30534
rect 1964 29306 1992 36615
rect 2148 34542 2176 39520
rect 2318 35592 2374 35601
rect 2318 35527 2374 35536
rect 2136 34536 2188 34542
rect 2136 34478 2188 34484
rect 2228 31884 2280 31890
rect 2228 31826 2280 31832
rect 2240 31142 2268 31826
rect 2228 31136 2280 31142
rect 2228 31078 2280 31084
rect 1952 29300 2004 29306
rect 1952 29242 2004 29248
rect 1768 25696 1820 25702
rect 1768 25638 1820 25644
rect 1674 15056 1730 15065
rect 1674 14991 1730 15000
rect 1398 12744 1454 12753
rect 1398 12679 1454 12688
rect 1412 12306 1440 12679
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 1412 11898 1440 12242
rect 1584 12232 1636 12238
rect 1584 12174 1636 12180
rect 1400 11892 1452 11898
rect 1400 11834 1452 11840
rect 1216 11076 1268 11082
rect 1216 11018 1268 11024
rect 1228 4146 1256 11018
rect 1596 10033 1624 12174
rect 1582 10024 1638 10033
rect 1582 9959 1638 9968
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 1596 6769 1624 6802
rect 1582 6760 1638 6769
rect 1582 6695 1638 6704
rect 1596 6458 1624 6695
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 1216 4140 1268 4146
rect 1216 4082 1268 4088
rect 1124 3732 1176 3738
rect 1124 3674 1176 3680
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1688 3505 1716 3538
rect 1674 3496 1730 3505
rect 1674 3431 1730 3440
rect 1688 3194 1716 3431
rect 1780 3369 1808 25638
rect 2134 25256 2190 25265
rect 2134 25191 2190 25200
rect 1858 22128 1914 22137
rect 1858 22063 1914 22072
rect 1872 13870 1900 22063
rect 2042 17232 2098 17241
rect 2042 17167 2098 17176
rect 1952 16652 2004 16658
rect 1952 16594 2004 16600
rect 1964 16017 1992 16594
rect 1950 16008 2006 16017
rect 1950 15943 2006 15952
rect 2056 15162 2084 17167
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 2056 14958 2084 15098
rect 2044 14952 2096 14958
rect 2044 14894 2096 14900
rect 2042 13968 2098 13977
rect 2042 13903 2098 13912
rect 1860 13864 1912 13870
rect 1860 13806 1912 13812
rect 2056 10674 2084 13903
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 1766 3360 1822 3369
rect 1766 3295 1822 3304
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 1400 3120 1452 3126
rect 1400 3062 1452 3068
rect 940 2304 992 2310
rect 940 2246 992 2252
rect 952 480 980 2246
rect 1412 480 1440 3062
rect 1780 480 1808 3130
rect 2148 480 2176 25191
rect 2240 16658 2268 31078
rect 2332 28370 2360 35527
rect 2504 34944 2556 34950
rect 2504 34886 2556 34892
rect 2412 29096 2464 29102
rect 2412 29038 2464 29044
rect 2424 28529 2452 29038
rect 2410 28520 2466 28529
rect 2410 28455 2412 28464
rect 2464 28455 2466 28464
rect 2412 28426 2464 28432
rect 2332 28342 2452 28370
rect 2228 16652 2280 16658
rect 2228 16594 2280 16600
rect 2318 16144 2374 16153
rect 2318 16079 2374 16088
rect 2228 13728 2280 13734
rect 2228 13670 2280 13676
rect 2240 3194 2268 13670
rect 2332 11218 2360 16079
rect 2320 11212 2372 11218
rect 2320 11154 2372 11160
rect 2332 10810 2360 11154
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2332 2650 2360 10610
rect 2424 3194 2452 28342
rect 2516 5794 2544 34886
rect 2608 34626 2636 39520
rect 2976 39494 3096 39520
rect 2608 34598 2728 34626
rect 2596 34536 2648 34542
rect 2596 34478 2648 34484
rect 2608 9654 2636 34478
rect 2596 9648 2648 9654
rect 2596 9590 2648 9596
rect 2700 6905 2728 34598
rect 3068 26738 3096 39494
rect 3344 26874 3372 39520
rect 3804 37210 3832 39520
rect 3804 37182 4016 37210
rect 3622 37020 3918 37040
rect 3678 37018 3702 37020
rect 3758 37018 3782 37020
rect 3838 37018 3862 37020
rect 3700 36966 3702 37018
rect 3764 36966 3776 37018
rect 3838 36966 3840 37018
rect 3678 36964 3702 36966
rect 3758 36964 3782 36966
rect 3838 36964 3862 36966
rect 3622 36944 3918 36964
rect 3622 35932 3918 35952
rect 3678 35930 3702 35932
rect 3758 35930 3782 35932
rect 3838 35930 3862 35932
rect 3700 35878 3702 35930
rect 3764 35878 3776 35930
rect 3838 35878 3840 35930
rect 3678 35876 3702 35878
rect 3758 35876 3782 35878
rect 3838 35876 3862 35878
rect 3622 35856 3918 35876
rect 3622 34844 3918 34864
rect 3678 34842 3702 34844
rect 3758 34842 3782 34844
rect 3838 34842 3862 34844
rect 3700 34790 3702 34842
rect 3764 34790 3776 34842
rect 3838 34790 3840 34842
rect 3678 34788 3702 34790
rect 3758 34788 3782 34790
rect 3838 34788 3862 34790
rect 3622 34768 3918 34788
rect 3622 33756 3918 33776
rect 3678 33754 3702 33756
rect 3758 33754 3782 33756
rect 3838 33754 3862 33756
rect 3700 33702 3702 33754
rect 3764 33702 3776 33754
rect 3838 33702 3840 33754
rect 3678 33700 3702 33702
rect 3758 33700 3782 33702
rect 3838 33700 3862 33702
rect 3622 33680 3918 33700
rect 3622 32668 3918 32688
rect 3678 32666 3702 32668
rect 3758 32666 3782 32668
rect 3838 32666 3862 32668
rect 3700 32614 3702 32666
rect 3764 32614 3776 32666
rect 3838 32614 3840 32666
rect 3678 32612 3702 32614
rect 3758 32612 3782 32614
rect 3838 32612 3862 32614
rect 3622 32592 3918 32612
rect 3622 31580 3918 31600
rect 3678 31578 3702 31580
rect 3758 31578 3782 31580
rect 3838 31578 3862 31580
rect 3700 31526 3702 31578
rect 3764 31526 3776 31578
rect 3838 31526 3840 31578
rect 3678 31524 3702 31526
rect 3758 31524 3782 31526
rect 3838 31524 3862 31526
rect 3622 31504 3918 31524
rect 3622 30492 3918 30512
rect 3678 30490 3702 30492
rect 3758 30490 3782 30492
rect 3838 30490 3862 30492
rect 3700 30438 3702 30490
rect 3764 30438 3776 30490
rect 3838 30438 3840 30490
rect 3678 30436 3702 30438
rect 3758 30436 3782 30438
rect 3838 30436 3862 30438
rect 3622 30416 3918 30436
rect 3622 29404 3918 29424
rect 3678 29402 3702 29404
rect 3758 29402 3782 29404
rect 3838 29402 3862 29404
rect 3700 29350 3702 29402
rect 3764 29350 3776 29402
rect 3838 29350 3840 29402
rect 3678 29348 3702 29350
rect 3758 29348 3782 29350
rect 3838 29348 3862 29350
rect 3622 29328 3918 29348
rect 3622 28316 3918 28336
rect 3678 28314 3702 28316
rect 3758 28314 3782 28316
rect 3838 28314 3862 28316
rect 3700 28262 3702 28314
rect 3764 28262 3776 28314
rect 3838 28262 3840 28314
rect 3678 28260 3702 28262
rect 3758 28260 3782 28262
rect 3838 28260 3862 28262
rect 3622 28240 3918 28260
rect 3622 27228 3918 27248
rect 3678 27226 3702 27228
rect 3758 27226 3782 27228
rect 3838 27226 3862 27228
rect 3700 27174 3702 27226
rect 3764 27174 3776 27226
rect 3838 27174 3840 27226
rect 3678 27172 3702 27174
rect 3758 27172 3782 27174
rect 3838 27172 3862 27174
rect 3622 27152 3918 27172
rect 3344 26846 3464 26874
rect 3068 26710 3372 26738
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 3160 9722 3188 19246
rect 3148 9716 3200 9722
rect 3148 9658 3200 9664
rect 2686 6896 2742 6905
rect 2686 6831 2742 6840
rect 3344 6361 3372 26710
rect 3436 19310 3464 26846
rect 3622 26140 3918 26160
rect 3678 26138 3702 26140
rect 3758 26138 3782 26140
rect 3838 26138 3862 26140
rect 3700 26086 3702 26138
rect 3764 26086 3776 26138
rect 3838 26086 3840 26138
rect 3678 26084 3702 26086
rect 3758 26084 3782 26086
rect 3838 26084 3862 26086
rect 3622 26064 3918 26084
rect 3622 25052 3918 25072
rect 3678 25050 3702 25052
rect 3758 25050 3782 25052
rect 3838 25050 3862 25052
rect 3700 24998 3702 25050
rect 3764 24998 3776 25050
rect 3838 24998 3840 25050
rect 3678 24996 3702 24998
rect 3758 24996 3782 24998
rect 3838 24996 3862 24998
rect 3622 24976 3918 24996
rect 3622 23964 3918 23984
rect 3678 23962 3702 23964
rect 3758 23962 3782 23964
rect 3838 23962 3862 23964
rect 3700 23910 3702 23962
rect 3764 23910 3776 23962
rect 3838 23910 3840 23962
rect 3678 23908 3702 23910
rect 3758 23908 3782 23910
rect 3838 23908 3862 23910
rect 3622 23888 3918 23908
rect 3622 22876 3918 22896
rect 3678 22874 3702 22876
rect 3758 22874 3782 22876
rect 3838 22874 3862 22876
rect 3700 22822 3702 22874
rect 3764 22822 3776 22874
rect 3838 22822 3840 22874
rect 3678 22820 3702 22822
rect 3758 22820 3782 22822
rect 3838 22820 3862 22822
rect 3622 22800 3918 22820
rect 3622 21788 3918 21808
rect 3678 21786 3702 21788
rect 3758 21786 3782 21788
rect 3838 21786 3862 21788
rect 3700 21734 3702 21786
rect 3764 21734 3776 21786
rect 3838 21734 3840 21786
rect 3678 21732 3702 21734
rect 3758 21732 3782 21734
rect 3838 21732 3862 21734
rect 3622 21712 3918 21732
rect 3622 20700 3918 20720
rect 3678 20698 3702 20700
rect 3758 20698 3782 20700
rect 3838 20698 3862 20700
rect 3700 20646 3702 20698
rect 3764 20646 3776 20698
rect 3838 20646 3840 20698
rect 3678 20644 3702 20646
rect 3758 20644 3782 20646
rect 3838 20644 3862 20646
rect 3622 20624 3918 20644
rect 3622 19612 3918 19632
rect 3678 19610 3702 19612
rect 3758 19610 3782 19612
rect 3838 19610 3862 19612
rect 3700 19558 3702 19610
rect 3764 19558 3776 19610
rect 3838 19558 3840 19610
rect 3678 19556 3702 19558
rect 3758 19556 3782 19558
rect 3838 19556 3862 19558
rect 3622 19536 3918 19556
rect 3424 19304 3476 19310
rect 3424 19246 3476 19252
rect 3622 18524 3918 18544
rect 3678 18522 3702 18524
rect 3758 18522 3782 18524
rect 3838 18522 3862 18524
rect 3700 18470 3702 18522
rect 3764 18470 3776 18522
rect 3838 18470 3840 18522
rect 3678 18468 3702 18470
rect 3758 18468 3782 18470
rect 3838 18468 3862 18470
rect 3622 18448 3918 18468
rect 3622 17436 3918 17456
rect 3678 17434 3702 17436
rect 3758 17434 3782 17436
rect 3838 17434 3862 17436
rect 3700 17382 3702 17434
rect 3764 17382 3776 17434
rect 3838 17382 3840 17434
rect 3678 17380 3702 17382
rect 3758 17380 3782 17382
rect 3838 17380 3862 17382
rect 3622 17360 3918 17380
rect 3622 16348 3918 16368
rect 3678 16346 3702 16348
rect 3758 16346 3782 16348
rect 3838 16346 3862 16348
rect 3700 16294 3702 16346
rect 3764 16294 3776 16346
rect 3838 16294 3840 16346
rect 3678 16292 3702 16294
rect 3758 16292 3782 16294
rect 3838 16292 3862 16294
rect 3622 16272 3918 16292
rect 3622 15260 3918 15280
rect 3678 15258 3702 15260
rect 3758 15258 3782 15260
rect 3838 15258 3862 15260
rect 3700 15206 3702 15258
rect 3764 15206 3776 15258
rect 3838 15206 3840 15258
rect 3678 15204 3702 15206
rect 3758 15204 3782 15206
rect 3838 15204 3862 15206
rect 3622 15184 3918 15204
rect 3622 14172 3918 14192
rect 3678 14170 3702 14172
rect 3758 14170 3782 14172
rect 3838 14170 3862 14172
rect 3700 14118 3702 14170
rect 3764 14118 3776 14170
rect 3838 14118 3840 14170
rect 3678 14116 3702 14118
rect 3758 14116 3782 14118
rect 3838 14116 3862 14118
rect 3622 14096 3918 14116
rect 3622 13084 3918 13104
rect 3678 13082 3702 13084
rect 3758 13082 3782 13084
rect 3838 13082 3862 13084
rect 3700 13030 3702 13082
rect 3764 13030 3776 13082
rect 3838 13030 3840 13082
rect 3678 13028 3702 13030
rect 3758 13028 3782 13030
rect 3838 13028 3862 13030
rect 3622 13008 3918 13028
rect 3622 11996 3918 12016
rect 3678 11994 3702 11996
rect 3758 11994 3782 11996
rect 3838 11994 3862 11996
rect 3700 11942 3702 11994
rect 3764 11942 3776 11994
rect 3838 11942 3840 11994
rect 3678 11940 3702 11942
rect 3758 11940 3782 11942
rect 3838 11940 3862 11942
rect 3622 11920 3918 11940
rect 3622 10908 3918 10928
rect 3678 10906 3702 10908
rect 3758 10906 3782 10908
rect 3838 10906 3862 10908
rect 3700 10854 3702 10906
rect 3764 10854 3776 10906
rect 3838 10854 3840 10906
rect 3678 10852 3702 10854
rect 3758 10852 3782 10854
rect 3838 10852 3862 10854
rect 3622 10832 3918 10852
rect 3622 9820 3918 9840
rect 3678 9818 3702 9820
rect 3758 9818 3782 9820
rect 3838 9818 3862 9820
rect 3700 9766 3702 9818
rect 3764 9766 3776 9818
rect 3838 9766 3840 9818
rect 3678 9764 3702 9766
rect 3758 9764 3782 9766
rect 3838 9764 3862 9766
rect 3622 9744 3918 9764
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 3436 8090 3464 9658
rect 3516 9444 3568 9450
rect 3516 9386 3568 9392
rect 3528 9081 3556 9386
rect 3514 9072 3570 9081
rect 3514 9007 3570 9016
rect 3622 8732 3918 8752
rect 3678 8730 3702 8732
rect 3758 8730 3782 8732
rect 3838 8730 3862 8732
rect 3700 8678 3702 8730
rect 3764 8678 3776 8730
rect 3838 8678 3840 8730
rect 3678 8676 3702 8678
rect 3758 8676 3782 8678
rect 3838 8676 3862 8678
rect 3622 8656 3918 8676
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3622 7644 3918 7664
rect 3678 7642 3702 7644
rect 3758 7642 3782 7644
rect 3838 7642 3862 7644
rect 3700 7590 3702 7642
rect 3764 7590 3776 7642
rect 3838 7590 3840 7642
rect 3678 7588 3702 7590
rect 3758 7588 3782 7590
rect 3838 7588 3862 7590
rect 3622 7568 3918 7588
rect 3622 6556 3918 6576
rect 3678 6554 3702 6556
rect 3758 6554 3782 6556
rect 3838 6554 3862 6556
rect 3700 6502 3702 6554
rect 3764 6502 3776 6554
rect 3838 6502 3840 6554
rect 3678 6500 3702 6502
rect 3758 6500 3782 6502
rect 3838 6500 3862 6502
rect 3622 6480 3918 6500
rect 3330 6352 3386 6361
rect 3330 6287 3386 6296
rect 2516 5766 2728 5794
rect 2594 5672 2650 5681
rect 2594 5607 2650 5616
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 2424 2990 2452 3130
rect 2412 2984 2464 2990
rect 2412 2926 2464 2932
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 2608 480 2636 5607
rect 2700 2666 2728 5766
rect 3622 5468 3918 5488
rect 3678 5466 3702 5468
rect 3758 5466 3782 5468
rect 3838 5466 3862 5468
rect 3700 5414 3702 5466
rect 3764 5414 3776 5466
rect 3838 5414 3840 5466
rect 3678 5412 3702 5414
rect 3758 5412 3782 5414
rect 3838 5412 3862 5414
rect 3622 5392 3918 5412
rect 3622 4380 3918 4400
rect 3678 4378 3702 4380
rect 3758 4378 3782 4380
rect 3838 4378 3862 4380
rect 3700 4326 3702 4378
rect 3764 4326 3776 4378
rect 3838 4326 3840 4378
rect 3678 4324 3702 4326
rect 3758 4324 3782 4326
rect 3838 4324 3862 4326
rect 3622 4304 3918 4324
rect 3988 3890 4016 37182
rect 4172 32026 4200 39520
rect 4540 35766 4568 39520
rect 4528 35760 4580 35766
rect 4528 35702 4580 35708
rect 5000 35714 5028 39520
rect 5000 35686 5304 35714
rect 5080 35624 5132 35630
rect 5080 35566 5132 35572
rect 4434 34640 4490 34649
rect 4434 34575 4490 34584
rect 4160 32020 4212 32026
rect 4160 31962 4212 31968
rect 4068 31884 4120 31890
rect 4068 31826 4120 31832
rect 4080 31226 4108 31826
rect 4080 31198 4200 31226
rect 4172 31142 4200 31198
rect 4160 31136 4212 31142
rect 4160 31078 4212 31084
rect 4066 25392 4122 25401
rect 4066 25327 4068 25336
rect 4120 25327 4122 25336
rect 4068 25298 4120 25304
rect 4080 24954 4108 25298
rect 4068 24948 4120 24954
rect 4068 24890 4120 24896
rect 4172 21865 4200 31078
rect 4448 29073 4476 34575
rect 4434 29064 4490 29073
rect 4434 28999 4490 29008
rect 4618 29030 4674 29039
rect 4436 28960 4488 28966
rect 4618 28965 4674 28974
rect 4436 28902 4488 28908
rect 4448 27878 4476 28902
rect 4526 28520 4582 28529
rect 4526 28455 4582 28464
rect 4540 28014 4568 28455
rect 4528 28008 4580 28014
rect 4528 27950 4580 27956
rect 4436 27872 4488 27878
rect 4436 27814 4488 27820
rect 4344 27600 4396 27606
rect 4344 27542 4396 27548
rect 4250 25256 4306 25265
rect 4250 25191 4252 25200
rect 4304 25191 4306 25200
rect 4252 25162 4304 25168
rect 4158 21856 4214 21865
rect 4158 21791 4214 21800
rect 4356 19242 4384 27542
rect 4448 22001 4476 27814
rect 4540 27334 4568 27950
rect 4632 27606 4660 28965
rect 4620 27600 4672 27606
rect 4620 27542 4672 27548
rect 4528 27328 4580 27334
rect 4528 27270 4580 27276
rect 4434 21992 4490 22001
rect 4434 21927 4490 21936
rect 4344 19236 4396 19242
rect 4344 19178 4396 19184
rect 4448 16794 4476 21927
rect 4528 19236 4580 19242
rect 4528 19178 4580 19184
rect 4436 16788 4488 16794
rect 4436 16730 4488 16736
rect 4448 16114 4476 16730
rect 4436 16108 4488 16114
rect 4436 16050 4488 16056
rect 4342 16008 4398 16017
rect 4342 15943 4344 15952
rect 4396 15943 4398 15952
rect 4344 15914 4396 15920
rect 4436 15904 4488 15910
rect 4436 15846 4488 15852
rect 4448 15706 4476 15846
rect 4436 15700 4488 15706
rect 4436 15642 4488 15648
rect 4342 15056 4398 15065
rect 4342 14991 4398 15000
rect 4356 14890 4384 14991
rect 4344 14884 4396 14890
rect 4344 14826 4396 14832
rect 4436 14816 4488 14822
rect 4436 14758 4488 14764
rect 4448 14618 4476 14758
rect 4436 14612 4488 14618
rect 4436 14554 4488 14560
rect 4540 12594 4568 19178
rect 4802 16144 4858 16153
rect 4802 16079 4858 16088
rect 4988 16108 5040 16114
rect 4816 16046 4844 16079
rect 4988 16050 5040 16056
rect 4804 16040 4856 16046
rect 4804 15982 4856 15988
rect 4816 15638 4844 15982
rect 4896 15904 4948 15910
rect 4896 15846 4948 15852
rect 4804 15632 4856 15638
rect 4908 15609 4936 15846
rect 4804 15574 4856 15580
rect 4894 15600 4950 15609
rect 4894 15535 4950 15544
rect 4802 15056 4858 15065
rect 5000 15026 5028 16050
rect 4802 14991 4858 15000
rect 4988 15020 5040 15026
rect 4816 14958 4844 14991
rect 4988 14962 5040 14968
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 4816 14550 4844 14894
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 4804 14544 4856 14550
rect 4908 14521 4936 14758
rect 4804 14486 4856 14492
rect 4894 14512 4950 14521
rect 4816 13977 4844 14486
rect 4894 14447 4950 14456
rect 4802 13968 4858 13977
rect 4802 13903 4858 13912
rect 4356 12566 4568 12594
rect 4356 12322 4384 12566
rect 4356 12294 4568 12322
rect 4250 7304 4306 7313
rect 4250 7239 4306 7248
rect 3988 3862 4200 3890
rect 4172 3738 4200 3862
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4264 3618 4292 7239
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4356 5681 4384 6054
rect 4342 5672 4398 5681
rect 4342 5607 4398 5616
rect 4172 3590 4292 3618
rect 3622 3292 3918 3312
rect 3678 3290 3702 3292
rect 3758 3290 3782 3292
rect 3838 3290 3862 3292
rect 3700 3238 3702 3290
rect 3764 3238 3776 3290
rect 3838 3238 3840 3290
rect 3678 3236 3702 3238
rect 3758 3236 3782 3238
rect 3838 3236 3862 3238
rect 3622 3216 3918 3236
rect 3332 3120 3384 3126
rect 3332 3062 3384 3068
rect 2962 2816 3018 2825
rect 2962 2751 3018 2760
rect 2700 2650 2820 2666
rect 2700 2644 2832 2650
rect 2700 2638 2780 2644
rect 2780 2586 2832 2592
rect 2976 480 3004 2751
rect 3344 480 3372 3062
rect 3516 2508 3568 2514
rect 3516 2450 3568 2456
rect 3528 2310 3556 2450
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 3528 1873 3556 2246
rect 3622 2204 3918 2224
rect 3678 2202 3702 2204
rect 3758 2202 3782 2204
rect 3838 2202 3862 2204
rect 3700 2150 3702 2202
rect 3764 2150 3776 2202
rect 3838 2150 3840 2202
rect 3678 2148 3702 2150
rect 3758 2148 3782 2150
rect 3838 2148 3862 2150
rect 3622 2128 3918 2148
rect 3514 1864 3570 1873
rect 3514 1799 3570 1808
rect 3988 1170 4016 2246
rect 3804 1142 4016 1170
rect 3804 480 3832 1142
rect 4172 480 4200 3590
rect 4434 3496 4490 3505
rect 4434 3431 4490 3440
rect 4448 1034 4476 3431
rect 4540 2514 4568 12294
rect 5092 9489 5120 35566
rect 5172 31884 5224 31890
rect 5172 31826 5224 31832
rect 5184 31142 5212 31826
rect 5172 31136 5224 31142
rect 5172 31078 5224 31084
rect 5184 20330 5212 31078
rect 5172 20324 5224 20330
rect 5172 20266 5224 20272
rect 5172 15360 5224 15366
rect 5170 15328 5172 15337
rect 5224 15328 5226 15337
rect 5170 15263 5226 15272
rect 5078 9480 5134 9489
rect 5078 9415 5134 9424
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 4908 7206 4936 7890
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4804 6248 4856 6254
rect 4802 6216 4804 6225
rect 4856 6216 4858 6225
rect 4802 6151 4858 6160
rect 4908 5817 4936 7142
rect 4894 5808 4950 5817
rect 4894 5743 4950 5752
rect 4710 3632 4766 3641
rect 4710 3567 4712 3576
rect 4764 3567 4766 3576
rect 4712 3538 4764 3544
rect 4724 3194 4752 3538
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 5276 2553 5304 35686
rect 5368 35630 5396 39520
rect 5736 35766 5764 39520
rect 5448 35760 5500 35766
rect 5448 35702 5500 35708
rect 5724 35760 5776 35766
rect 5724 35702 5776 35708
rect 5356 35624 5408 35630
rect 5356 35566 5408 35572
rect 5354 28656 5410 28665
rect 5354 28591 5410 28600
rect 5368 27334 5396 28591
rect 5356 27328 5408 27334
rect 5356 27270 5408 27276
rect 5368 24410 5396 27270
rect 5356 24404 5408 24410
rect 5356 24346 5408 24352
rect 5354 2952 5410 2961
rect 5354 2887 5410 2896
rect 5262 2544 5318 2553
rect 4528 2508 4580 2514
rect 5262 2479 5318 2488
rect 4528 2450 4580 2456
rect 4986 1456 5042 1465
rect 4986 1391 5042 1400
rect 4448 1006 4568 1034
rect 4540 480 4568 1006
rect 5000 480 5028 1391
rect 5368 480 5396 2887
rect 5460 2281 5488 35702
rect 6196 35698 6224 39520
rect 6564 37754 6592 39520
rect 6564 37726 6868 37754
rect 6289 37564 6585 37584
rect 6345 37562 6369 37564
rect 6425 37562 6449 37564
rect 6505 37562 6529 37564
rect 6367 37510 6369 37562
rect 6431 37510 6443 37562
rect 6505 37510 6507 37562
rect 6345 37508 6369 37510
rect 6425 37508 6449 37510
rect 6505 37508 6529 37510
rect 6289 37488 6585 37508
rect 6289 36476 6585 36496
rect 6345 36474 6369 36476
rect 6425 36474 6449 36476
rect 6505 36474 6529 36476
rect 6367 36422 6369 36474
rect 6431 36422 6443 36474
rect 6505 36422 6507 36474
rect 6345 36420 6369 36422
rect 6425 36420 6449 36422
rect 6505 36420 6529 36422
rect 6289 36400 6585 36420
rect 6736 35760 6788 35766
rect 6736 35702 6788 35708
rect 6184 35692 6236 35698
rect 6184 35634 6236 35640
rect 6644 35692 6696 35698
rect 6644 35634 6696 35640
rect 6289 35388 6585 35408
rect 6345 35386 6369 35388
rect 6425 35386 6449 35388
rect 6505 35386 6529 35388
rect 6367 35334 6369 35386
rect 6431 35334 6443 35386
rect 6505 35334 6507 35386
rect 6345 35332 6369 35334
rect 6425 35332 6449 35334
rect 6505 35332 6529 35334
rect 6289 35312 6585 35332
rect 5998 35184 6054 35193
rect 5998 35119 6054 35128
rect 5814 35048 5870 35057
rect 5814 34983 5870 34992
rect 5724 28960 5776 28966
rect 5724 28902 5776 28908
rect 5736 27878 5764 28902
rect 5724 27872 5776 27878
rect 5724 27814 5776 27820
rect 5632 21888 5684 21894
rect 5632 21830 5684 21836
rect 5644 21146 5672 21830
rect 5632 21140 5684 21146
rect 5632 21082 5684 21088
rect 5736 20505 5764 27814
rect 5722 20496 5778 20505
rect 5644 20454 5722 20482
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5552 14618 5580 15506
rect 5644 15502 5672 20454
rect 5722 20431 5778 20440
rect 5724 15700 5776 15706
rect 5724 15642 5776 15648
rect 5632 15496 5684 15502
rect 5632 15438 5684 15444
rect 5644 15162 5672 15438
rect 5736 15162 5764 15642
rect 5632 15156 5684 15162
rect 5632 15098 5684 15104
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5540 14612 5592 14618
rect 5540 14554 5592 14560
rect 5722 4720 5778 4729
rect 5722 4655 5778 4664
rect 5446 2272 5502 2281
rect 5446 2207 5502 2216
rect 5736 480 5764 4655
rect 5828 3194 5856 34983
rect 6012 26874 6040 35119
rect 6289 34300 6585 34320
rect 6345 34298 6369 34300
rect 6425 34298 6449 34300
rect 6505 34298 6529 34300
rect 6367 34246 6369 34298
rect 6431 34246 6443 34298
rect 6505 34246 6507 34298
rect 6345 34244 6369 34246
rect 6425 34244 6449 34246
rect 6505 34244 6529 34246
rect 6289 34224 6585 34244
rect 6289 33212 6585 33232
rect 6345 33210 6369 33212
rect 6425 33210 6449 33212
rect 6505 33210 6529 33212
rect 6367 33158 6369 33210
rect 6431 33158 6443 33210
rect 6505 33158 6507 33210
rect 6345 33156 6369 33158
rect 6425 33156 6449 33158
rect 6505 33156 6529 33158
rect 6289 33136 6585 33156
rect 6289 32124 6585 32144
rect 6345 32122 6369 32124
rect 6425 32122 6449 32124
rect 6505 32122 6529 32124
rect 6367 32070 6369 32122
rect 6431 32070 6443 32122
rect 6505 32070 6507 32122
rect 6345 32068 6369 32070
rect 6425 32068 6449 32070
rect 6505 32068 6529 32070
rect 6289 32048 6585 32068
rect 6289 31036 6585 31056
rect 6345 31034 6369 31036
rect 6425 31034 6449 31036
rect 6505 31034 6529 31036
rect 6367 30982 6369 31034
rect 6431 30982 6443 31034
rect 6505 30982 6507 31034
rect 6345 30980 6369 30982
rect 6425 30980 6449 30982
rect 6505 30980 6529 30982
rect 6289 30960 6585 30980
rect 6289 29948 6585 29968
rect 6345 29946 6369 29948
rect 6425 29946 6449 29948
rect 6505 29946 6529 29948
rect 6367 29894 6369 29946
rect 6431 29894 6443 29946
rect 6505 29894 6507 29946
rect 6345 29892 6369 29894
rect 6425 29892 6449 29894
rect 6505 29892 6529 29894
rect 6289 29872 6585 29892
rect 6289 28860 6585 28880
rect 6345 28858 6369 28860
rect 6425 28858 6449 28860
rect 6505 28858 6529 28860
rect 6367 28806 6369 28858
rect 6431 28806 6443 28858
rect 6505 28806 6507 28858
rect 6345 28804 6369 28806
rect 6425 28804 6449 28806
rect 6505 28804 6529 28806
rect 6289 28784 6585 28804
rect 6289 27772 6585 27792
rect 6345 27770 6369 27772
rect 6425 27770 6449 27772
rect 6505 27770 6529 27772
rect 6367 27718 6369 27770
rect 6431 27718 6443 27770
rect 6505 27718 6507 27770
rect 6345 27716 6369 27718
rect 6425 27716 6449 27718
rect 6505 27716 6529 27718
rect 6289 27696 6585 27716
rect 5920 26846 6040 26874
rect 5920 6610 5948 26846
rect 6289 26684 6585 26704
rect 6345 26682 6369 26684
rect 6425 26682 6449 26684
rect 6505 26682 6529 26684
rect 6367 26630 6369 26682
rect 6431 26630 6443 26682
rect 6505 26630 6507 26682
rect 6345 26628 6369 26630
rect 6425 26628 6449 26630
rect 6505 26628 6529 26630
rect 6289 26608 6585 26628
rect 6289 25596 6585 25616
rect 6345 25594 6369 25596
rect 6425 25594 6449 25596
rect 6505 25594 6529 25596
rect 6367 25542 6369 25594
rect 6431 25542 6443 25594
rect 6505 25542 6507 25594
rect 6345 25540 6369 25542
rect 6425 25540 6449 25542
rect 6505 25540 6529 25542
rect 6289 25520 6585 25540
rect 6289 24508 6585 24528
rect 6345 24506 6369 24508
rect 6425 24506 6449 24508
rect 6505 24506 6529 24508
rect 6367 24454 6369 24506
rect 6431 24454 6443 24506
rect 6505 24454 6507 24506
rect 6345 24452 6369 24454
rect 6425 24452 6449 24454
rect 6505 24452 6529 24454
rect 6289 24432 6585 24452
rect 6289 23420 6585 23440
rect 6345 23418 6369 23420
rect 6425 23418 6449 23420
rect 6505 23418 6529 23420
rect 6367 23366 6369 23418
rect 6431 23366 6443 23418
rect 6505 23366 6507 23418
rect 6345 23364 6369 23366
rect 6425 23364 6449 23366
rect 6505 23364 6529 23366
rect 6289 23344 6585 23364
rect 5998 23080 6054 23089
rect 5998 23015 6054 23024
rect 6012 22137 6040 23015
rect 6289 22332 6585 22352
rect 6345 22330 6369 22332
rect 6425 22330 6449 22332
rect 6505 22330 6529 22332
rect 6367 22278 6369 22330
rect 6431 22278 6443 22330
rect 6505 22278 6507 22330
rect 6345 22276 6369 22278
rect 6425 22276 6449 22278
rect 6505 22276 6529 22278
rect 6289 22256 6585 22276
rect 5998 22128 6054 22137
rect 5998 22063 6000 22072
rect 6052 22063 6054 22072
rect 6000 22034 6052 22040
rect 6012 21690 6040 22034
rect 6092 22024 6144 22030
rect 6276 22024 6328 22030
rect 6092 21966 6144 21972
rect 6274 21992 6276 22001
rect 6328 21992 6330 22001
rect 6104 21865 6132 21966
rect 6274 21927 6330 21936
rect 6090 21856 6146 21865
rect 6090 21791 6146 21800
rect 6000 21684 6052 21690
rect 6000 21626 6052 21632
rect 6104 21434 6132 21791
rect 6288 21690 6316 21927
rect 6276 21684 6328 21690
rect 6276 21626 6328 21632
rect 6012 21406 6132 21434
rect 6012 21350 6040 21406
rect 6000 21344 6052 21350
rect 6000 21286 6052 21292
rect 6012 21049 6040 21286
rect 6289 21244 6585 21264
rect 6345 21242 6369 21244
rect 6425 21242 6449 21244
rect 6505 21242 6529 21244
rect 6367 21190 6369 21242
rect 6431 21190 6443 21242
rect 6505 21190 6507 21242
rect 6345 21188 6369 21190
rect 6425 21188 6449 21190
rect 6505 21188 6529 21190
rect 6289 21168 6585 21188
rect 5998 21040 6054 21049
rect 5998 20975 6054 20984
rect 6289 20156 6585 20176
rect 6345 20154 6369 20156
rect 6425 20154 6449 20156
rect 6505 20154 6529 20156
rect 6367 20102 6369 20154
rect 6431 20102 6443 20154
rect 6505 20102 6507 20154
rect 6345 20100 6369 20102
rect 6425 20100 6449 20102
rect 6505 20100 6529 20102
rect 6289 20080 6585 20100
rect 6289 19068 6585 19088
rect 6345 19066 6369 19068
rect 6425 19066 6449 19068
rect 6505 19066 6529 19068
rect 6367 19014 6369 19066
rect 6431 19014 6443 19066
rect 6505 19014 6507 19066
rect 6345 19012 6369 19014
rect 6425 19012 6449 19014
rect 6505 19012 6529 19014
rect 6289 18992 6585 19012
rect 6289 17980 6585 18000
rect 6345 17978 6369 17980
rect 6425 17978 6449 17980
rect 6505 17978 6529 17980
rect 6367 17926 6369 17978
rect 6431 17926 6443 17978
rect 6505 17926 6507 17978
rect 6345 17924 6369 17926
rect 6425 17924 6449 17926
rect 6505 17924 6529 17926
rect 6289 17904 6585 17924
rect 6289 16892 6585 16912
rect 6345 16890 6369 16892
rect 6425 16890 6449 16892
rect 6505 16890 6529 16892
rect 6367 16838 6369 16890
rect 6431 16838 6443 16890
rect 6505 16838 6507 16890
rect 6345 16836 6369 16838
rect 6425 16836 6449 16838
rect 6505 16836 6529 16838
rect 6289 16816 6585 16836
rect 6289 15804 6585 15824
rect 6345 15802 6369 15804
rect 6425 15802 6449 15804
rect 6505 15802 6529 15804
rect 6367 15750 6369 15802
rect 6431 15750 6443 15802
rect 6505 15750 6507 15802
rect 6345 15748 6369 15750
rect 6425 15748 6449 15750
rect 6505 15748 6529 15750
rect 6289 15728 6585 15748
rect 6289 14716 6585 14736
rect 6345 14714 6369 14716
rect 6425 14714 6449 14716
rect 6505 14714 6529 14716
rect 6367 14662 6369 14714
rect 6431 14662 6443 14714
rect 6505 14662 6507 14714
rect 6345 14660 6369 14662
rect 6425 14660 6449 14662
rect 6505 14660 6529 14662
rect 6289 14640 6585 14660
rect 6289 13628 6585 13648
rect 6345 13626 6369 13628
rect 6425 13626 6449 13628
rect 6505 13626 6529 13628
rect 6367 13574 6369 13626
rect 6431 13574 6443 13626
rect 6505 13574 6507 13626
rect 6345 13572 6369 13574
rect 6425 13572 6449 13574
rect 6505 13572 6529 13574
rect 6289 13552 6585 13572
rect 6289 12540 6585 12560
rect 6345 12538 6369 12540
rect 6425 12538 6449 12540
rect 6505 12538 6529 12540
rect 6367 12486 6369 12538
rect 6431 12486 6443 12538
rect 6505 12486 6507 12538
rect 6345 12484 6369 12486
rect 6425 12484 6449 12486
rect 6505 12484 6529 12486
rect 6289 12464 6585 12484
rect 6289 11452 6585 11472
rect 6345 11450 6369 11452
rect 6425 11450 6449 11452
rect 6505 11450 6529 11452
rect 6367 11398 6369 11450
rect 6431 11398 6443 11450
rect 6505 11398 6507 11450
rect 6345 11396 6369 11398
rect 6425 11396 6449 11398
rect 6505 11396 6529 11398
rect 6289 11376 6585 11396
rect 6289 10364 6585 10384
rect 6345 10362 6369 10364
rect 6425 10362 6449 10364
rect 6505 10362 6529 10364
rect 6367 10310 6369 10362
rect 6431 10310 6443 10362
rect 6505 10310 6507 10362
rect 6345 10308 6369 10310
rect 6425 10308 6449 10310
rect 6505 10308 6529 10310
rect 6289 10288 6585 10308
rect 6289 9276 6585 9296
rect 6345 9274 6369 9276
rect 6425 9274 6449 9276
rect 6505 9274 6529 9276
rect 6367 9222 6369 9274
rect 6431 9222 6443 9274
rect 6505 9222 6507 9274
rect 6345 9220 6369 9222
rect 6425 9220 6449 9222
rect 6505 9220 6529 9222
rect 6289 9200 6585 9220
rect 6289 8188 6585 8208
rect 6345 8186 6369 8188
rect 6425 8186 6449 8188
rect 6505 8186 6529 8188
rect 6367 8134 6369 8186
rect 6431 8134 6443 8186
rect 6505 8134 6507 8186
rect 6345 8132 6369 8134
rect 6425 8132 6449 8134
rect 6505 8132 6529 8134
rect 6289 8112 6585 8132
rect 6656 7562 6684 35634
rect 6748 7698 6776 35702
rect 6840 33153 6868 37726
rect 6932 35154 6960 39520
rect 7196 35692 7248 35698
rect 7196 35634 7248 35640
rect 6920 35148 6972 35154
rect 6920 35090 6972 35096
rect 6826 33144 6882 33153
rect 6826 33079 6882 33088
rect 6828 24268 6880 24274
rect 6828 24210 6880 24216
rect 6840 23526 6868 24210
rect 6828 23520 6880 23526
rect 6826 23488 6828 23497
rect 6880 23488 6882 23497
rect 6826 23423 6882 23432
rect 7012 21140 7064 21146
rect 7012 21082 7064 21088
rect 7024 20466 7052 21082
rect 7012 20460 7064 20466
rect 7012 20402 7064 20408
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 7024 15706 7052 20198
rect 7208 16153 7236 35634
rect 7392 35290 7420 39520
rect 7760 35714 7788 39520
rect 7760 35686 8156 35714
rect 8220 35698 8248 39520
rect 8392 37188 8444 37194
rect 8392 37130 8444 37136
rect 7380 35284 7432 35290
rect 7380 35226 7432 35232
rect 8024 35148 8076 35154
rect 8024 35090 8076 35096
rect 7380 29708 7432 29714
rect 7380 29650 7432 29656
rect 7392 29034 7420 29650
rect 7656 29504 7708 29510
rect 7656 29446 7708 29452
rect 7668 29034 7696 29446
rect 7380 29028 7432 29034
rect 7380 28970 7432 28976
rect 7656 29028 7708 29034
rect 7656 28970 7708 28976
rect 7668 28665 7696 28970
rect 7654 28656 7710 28665
rect 7654 28591 7710 28600
rect 8036 24721 8064 35090
rect 8022 24712 8078 24721
rect 8022 24647 8078 24656
rect 8128 24562 8156 35686
rect 8208 35692 8260 35698
rect 8208 35634 8260 35640
rect 8208 35284 8260 35290
rect 8208 35226 8260 35232
rect 7852 24534 8156 24562
rect 7470 22536 7526 22545
rect 7470 22471 7526 22480
rect 7564 22500 7616 22506
rect 7380 20256 7432 20262
rect 7378 20224 7380 20233
rect 7432 20224 7434 20233
rect 7378 20159 7434 20168
rect 7194 16144 7250 16153
rect 7194 16079 7250 16088
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 6918 15600 6974 15609
rect 6918 15535 6974 15544
rect 6932 10470 6960 15535
rect 7024 14958 7052 15642
rect 7194 15328 7250 15337
rect 7194 15263 7250 15272
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 7208 14890 7236 15263
rect 7196 14884 7248 14890
rect 7196 14826 7248 14832
rect 7208 14618 7236 14826
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7196 14612 7248 14618
rect 7196 14554 7248 14560
rect 7300 13530 7328 14758
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6748 7670 6868 7698
rect 6656 7534 6776 7562
rect 6289 7100 6585 7120
rect 6345 7098 6369 7100
rect 6425 7098 6449 7100
rect 6505 7098 6529 7100
rect 6367 7046 6369 7098
rect 6431 7046 6443 7098
rect 6505 7046 6507 7098
rect 6345 7044 6369 7046
rect 6425 7044 6449 7046
rect 6505 7044 6529 7046
rect 6289 7024 6585 7044
rect 6182 6896 6238 6905
rect 6182 6831 6238 6840
rect 6276 6860 6328 6866
rect 6196 6730 6224 6831
rect 6276 6802 6328 6808
rect 6184 6724 6236 6730
rect 6184 6666 6236 6672
rect 5920 6582 6224 6610
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 6104 4049 6132 6054
rect 6090 4040 6146 4049
rect 6090 3975 6146 3984
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 6090 3088 6146 3097
rect 6090 3023 6146 3032
rect 5814 2816 5870 2825
rect 5814 2751 5870 2760
rect 5828 2650 5856 2751
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 6104 1034 6132 3023
rect 6196 2582 6224 6582
rect 6288 6186 6316 6802
rect 6276 6180 6328 6186
rect 6276 6122 6328 6128
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6289 6012 6585 6032
rect 6345 6010 6369 6012
rect 6425 6010 6449 6012
rect 6505 6010 6529 6012
rect 6367 5958 6369 6010
rect 6431 5958 6443 6010
rect 6505 5958 6507 6010
rect 6345 5956 6369 5958
rect 6425 5956 6449 5958
rect 6505 5956 6529 5958
rect 6289 5936 6585 5956
rect 6289 4924 6585 4944
rect 6345 4922 6369 4924
rect 6425 4922 6449 4924
rect 6505 4922 6529 4924
rect 6367 4870 6369 4922
rect 6431 4870 6443 4922
rect 6505 4870 6507 4922
rect 6345 4868 6369 4870
rect 6425 4868 6449 4870
rect 6505 4868 6529 4870
rect 6289 4848 6585 4868
rect 6289 3836 6585 3856
rect 6345 3834 6369 3836
rect 6425 3834 6449 3836
rect 6505 3834 6529 3836
rect 6367 3782 6369 3834
rect 6431 3782 6443 3834
rect 6505 3782 6507 3834
rect 6345 3780 6369 3782
rect 6425 3780 6449 3782
rect 6505 3780 6529 3782
rect 6289 3760 6585 3780
rect 6289 2748 6585 2768
rect 6345 2746 6369 2748
rect 6425 2746 6449 2748
rect 6505 2746 6529 2748
rect 6367 2694 6369 2746
rect 6431 2694 6443 2746
rect 6505 2694 6507 2746
rect 6345 2692 6369 2694
rect 6425 2692 6449 2694
rect 6505 2692 6529 2694
rect 6289 2672 6585 2692
rect 6184 2576 6236 2582
rect 6184 2518 6236 2524
rect 6656 1034 6684 6054
rect 6748 2689 6776 7534
rect 6840 6769 6868 7670
rect 7484 7546 7512 22471
rect 7564 22442 7616 22448
rect 7576 14929 7604 22442
rect 7654 20496 7710 20505
rect 7654 20431 7656 20440
rect 7708 20431 7710 20440
rect 7656 20402 7708 20408
rect 7668 20058 7696 20402
rect 7656 20052 7708 20058
rect 7656 19994 7708 20000
rect 7562 14920 7618 14929
rect 7562 14855 7618 14864
rect 7852 9625 7880 24534
rect 8022 14648 8078 14657
rect 8022 14583 8024 14592
rect 8076 14583 8078 14592
rect 8024 14554 8076 14560
rect 8024 13796 8076 13802
rect 8024 13738 8076 13744
rect 7932 13728 7984 13734
rect 7932 13670 7984 13676
rect 7944 12753 7972 13670
rect 8036 13530 8064 13738
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 7930 12744 7986 12753
rect 7930 12679 7986 12688
rect 8220 10554 8248 35226
rect 8404 15065 8432 37130
rect 8484 30048 8536 30054
rect 8484 29990 8536 29996
rect 8390 15056 8446 15065
rect 8390 14991 8446 15000
rect 8298 14648 8354 14657
rect 8298 14583 8354 14592
rect 8312 13734 8340 14583
rect 8300 13728 8352 13734
rect 8300 13670 8352 13676
rect 8128 10526 8248 10554
rect 7838 9616 7894 9625
rect 7838 9551 7894 9560
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7484 7342 7512 7482
rect 7472 7336 7524 7342
rect 7010 7304 7066 7313
rect 7472 7278 7524 7284
rect 7010 7239 7066 7248
rect 7024 7206 7052 7239
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 6826 6760 6882 6769
rect 6826 6695 6882 6704
rect 6918 3768 6974 3777
rect 6918 3703 6974 3712
rect 6734 2680 6790 2689
rect 6734 2615 6790 2624
rect 6104 1006 6224 1034
rect 6196 480 6224 1006
rect 6564 1006 6684 1034
rect 6564 480 6592 1006
rect 6932 480 6960 3703
rect 7746 3632 7802 3641
rect 7746 3567 7802 3576
rect 7378 2816 7434 2825
rect 7378 2751 7434 2760
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7116 2553 7144 2586
rect 7102 2544 7158 2553
rect 7102 2479 7158 2488
rect 7392 480 7420 2751
rect 7564 2508 7616 2514
rect 7564 2450 7616 2456
rect 7576 2310 7604 2450
rect 7564 2304 7616 2310
rect 7564 2246 7616 2252
rect 7576 2009 7604 2246
rect 7562 2000 7618 2009
rect 7562 1935 7618 1944
rect 7760 480 7788 3567
rect 8128 2417 8156 10526
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8114 2408 8170 2417
rect 8114 2343 8170 2352
rect 8220 480 8248 10406
rect 8496 6458 8524 29990
rect 8588 26926 8616 39520
rect 8956 37194 8984 39520
rect 8944 37188 8996 37194
rect 8944 37130 8996 37136
rect 8956 37020 9252 37040
rect 9012 37018 9036 37020
rect 9092 37018 9116 37020
rect 9172 37018 9196 37020
rect 9034 36966 9036 37018
rect 9098 36966 9110 37018
rect 9172 36966 9174 37018
rect 9012 36964 9036 36966
rect 9092 36964 9116 36966
rect 9172 36964 9196 36966
rect 8956 36944 9252 36964
rect 8956 35932 9252 35952
rect 9012 35930 9036 35932
rect 9092 35930 9116 35932
rect 9172 35930 9196 35932
rect 9034 35878 9036 35930
rect 9098 35878 9110 35930
rect 9172 35878 9174 35930
rect 9012 35876 9036 35878
rect 9092 35876 9116 35878
rect 9172 35876 9196 35878
rect 8956 35856 9252 35876
rect 9416 35737 9444 39520
rect 9402 35728 9458 35737
rect 9402 35663 9458 35672
rect 8666 35592 8722 35601
rect 8666 35527 8722 35536
rect 8576 26920 8628 26926
rect 8576 26862 8628 26868
rect 8576 20256 8628 20262
rect 8576 20198 8628 20204
rect 8588 16697 8616 20198
rect 8574 16688 8630 16697
rect 8574 16623 8630 16632
rect 8588 15162 8616 16623
rect 8576 15156 8628 15162
rect 8576 15098 8628 15104
rect 8484 6452 8536 6458
rect 8484 6394 8536 6400
rect 8574 3360 8630 3369
rect 8574 3295 8630 3304
rect 8588 480 8616 3295
rect 8680 2990 8708 35527
rect 8956 34844 9252 34864
rect 9012 34842 9036 34844
rect 9092 34842 9116 34844
rect 9172 34842 9196 34844
rect 9034 34790 9036 34842
rect 9098 34790 9110 34842
rect 9172 34790 9174 34842
rect 9012 34788 9036 34790
rect 9092 34788 9116 34790
rect 9172 34788 9196 34790
rect 8956 34768 9252 34788
rect 8956 33756 9252 33776
rect 9012 33754 9036 33756
rect 9092 33754 9116 33756
rect 9172 33754 9196 33756
rect 9034 33702 9036 33754
rect 9098 33702 9110 33754
rect 9172 33702 9174 33754
rect 9012 33700 9036 33702
rect 9092 33700 9116 33702
rect 9172 33700 9196 33702
rect 8956 33680 9252 33700
rect 8758 33144 8814 33153
rect 8758 33079 8814 33088
rect 8772 31482 8800 33079
rect 8956 32668 9252 32688
rect 9012 32666 9036 32668
rect 9092 32666 9116 32668
rect 9172 32666 9196 32668
rect 9034 32614 9036 32666
rect 9098 32614 9110 32666
rect 9172 32614 9174 32666
rect 9012 32612 9036 32614
rect 9092 32612 9116 32614
rect 9172 32612 9196 32614
rect 8956 32592 9252 32612
rect 8956 31580 9252 31600
rect 9012 31578 9036 31580
rect 9092 31578 9116 31580
rect 9172 31578 9196 31580
rect 9034 31526 9036 31578
rect 9098 31526 9110 31578
rect 9172 31526 9174 31578
rect 9012 31524 9036 31526
rect 9092 31524 9116 31526
rect 9172 31524 9196 31526
rect 8956 31504 9252 31524
rect 8760 31476 8812 31482
rect 8760 31418 8812 31424
rect 9404 31136 9456 31142
rect 9404 31078 9456 31084
rect 9312 30592 9364 30598
rect 9312 30534 9364 30540
rect 8956 30492 9252 30512
rect 9012 30490 9036 30492
rect 9092 30490 9116 30492
rect 9172 30490 9196 30492
rect 9034 30438 9036 30490
rect 9098 30438 9110 30490
rect 9172 30438 9174 30490
rect 9012 30436 9036 30438
rect 9092 30436 9116 30438
rect 9172 30436 9196 30438
rect 8956 30416 9252 30436
rect 9324 30258 9352 30534
rect 9312 30252 9364 30258
rect 9312 30194 9364 30200
rect 9324 29714 9352 30194
rect 9312 29708 9364 29714
rect 9312 29650 9364 29656
rect 8956 29404 9252 29424
rect 9012 29402 9036 29404
rect 9092 29402 9116 29404
rect 9172 29402 9196 29404
rect 9034 29350 9036 29402
rect 9098 29350 9110 29402
rect 9172 29350 9174 29402
rect 9012 29348 9036 29350
rect 9092 29348 9116 29350
rect 9172 29348 9196 29350
rect 8956 29328 9252 29348
rect 8956 28316 9252 28336
rect 9012 28314 9036 28316
rect 9092 28314 9116 28316
rect 9172 28314 9196 28316
rect 9034 28262 9036 28314
rect 9098 28262 9110 28314
rect 9172 28262 9174 28314
rect 9012 28260 9036 28262
rect 9092 28260 9116 28262
rect 9172 28260 9196 28262
rect 8956 28240 9252 28260
rect 8956 27228 9252 27248
rect 9012 27226 9036 27228
rect 9092 27226 9116 27228
rect 9172 27226 9196 27228
rect 9034 27174 9036 27226
rect 9098 27174 9110 27226
rect 9172 27174 9174 27226
rect 9012 27172 9036 27174
rect 9092 27172 9116 27174
rect 9172 27172 9196 27174
rect 8956 27152 9252 27172
rect 9312 26920 9364 26926
rect 9312 26862 9364 26868
rect 8956 26140 9252 26160
rect 9012 26138 9036 26140
rect 9092 26138 9116 26140
rect 9172 26138 9196 26140
rect 9034 26086 9036 26138
rect 9098 26086 9110 26138
rect 9172 26086 9174 26138
rect 9012 26084 9036 26086
rect 9092 26084 9116 26086
rect 9172 26084 9196 26086
rect 8956 26064 9252 26084
rect 8956 25052 9252 25072
rect 9012 25050 9036 25052
rect 9092 25050 9116 25052
rect 9172 25050 9196 25052
rect 9034 24998 9036 25050
rect 9098 24998 9110 25050
rect 9172 24998 9174 25050
rect 9012 24996 9036 24998
rect 9092 24996 9116 24998
rect 9172 24996 9196 24998
rect 8956 24976 9252 24996
rect 8956 23964 9252 23984
rect 9012 23962 9036 23964
rect 9092 23962 9116 23964
rect 9172 23962 9196 23964
rect 9034 23910 9036 23962
rect 9098 23910 9110 23962
rect 9172 23910 9174 23962
rect 9012 23908 9036 23910
rect 9092 23908 9116 23910
rect 9172 23908 9196 23910
rect 8956 23888 9252 23908
rect 8758 23488 8814 23497
rect 8758 23423 8814 23432
rect 8772 22438 8800 23423
rect 8956 22876 9252 22896
rect 9012 22874 9036 22876
rect 9092 22874 9116 22876
rect 9172 22874 9196 22876
rect 9034 22822 9036 22874
rect 9098 22822 9110 22874
rect 9172 22822 9174 22874
rect 9012 22820 9036 22822
rect 9092 22820 9116 22822
rect 9172 22820 9196 22822
rect 8956 22800 9252 22820
rect 8760 22432 8812 22438
rect 8760 22374 8812 22380
rect 8772 20398 8800 22374
rect 8956 21788 9252 21808
rect 9012 21786 9036 21788
rect 9092 21786 9116 21788
rect 9172 21786 9196 21788
rect 9034 21734 9036 21786
rect 9098 21734 9110 21786
rect 9172 21734 9174 21786
rect 9012 21732 9036 21734
rect 9092 21732 9116 21734
rect 9172 21732 9196 21734
rect 8956 21712 9252 21732
rect 8956 20700 9252 20720
rect 9012 20698 9036 20700
rect 9092 20698 9116 20700
rect 9172 20698 9196 20700
rect 9034 20646 9036 20698
rect 9098 20646 9110 20698
rect 9172 20646 9174 20698
rect 9012 20644 9036 20646
rect 9092 20644 9116 20646
rect 9172 20644 9196 20646
rect 8956 20624 9252 20644
rect 8760 20392 8812 20398
rect 8760 20334 8812 20340
rect 8956 19612 9252 19632
rect 9012 19610 9036 19612
rect 9092 19610 9116 19612
rect 9172 19610 9196 19612
rect 9034 19558 9036 19610
rect 9098 19558 9110 19610
rect 9172 19558 9174 19610
rect 9012 19556 9036 19558
rect 9092 19556 9116 19558
rect 9172 19556 9196 19558
rect 8956 19536 9252 19556
rect 8956 18524 9252 18544
rect 9012 18522 9036 18524
rect 9092 18522 9116 18524
rect 9172 18522 9196 18524
rect 9034 18470 9036 18522
rect 9098 18470 9110 18522
rect 9172 18470 9174 18522
rect 9012 18468 9036 18470
rect 9092 18468 9116 18470
rect 9172 18468 9196 18470
rect 8956 18448 9252 18468
rect 8956 17436 9252 17456
rect 9012 17434 9036 17436
rect 9092 17434 9116 17436
rect 9172 17434 9196 17436
rect 9034 17382 9036 17434
rect 9098 17382 9110 17434
rect 9172 17382 9174 17434
rect 9012 17380 9036 17382
rect 9092 17380 9116 17382
rect 9172 17380 9196 17382
rect 8956 17360 9252 17380
rect 8956 16348 9252 16368
rect 9012 16346 9036 16348
rect 9092 16346 9116 16348
rect 9172 16346 9196 16348
rect 9034 16294 9036 16346
rect 9098 16294 9110 16346
rect 9172 16294 9174 16346
rect 9012 16292 9036 16294
rect 9092 16292 9116 16294
rect 9172 16292 9196 16294
rect 8956 16272 9252 16292
rect 8956 15260 9252 15280
rect 9012 15258 9036 15260
rect 9092 15258 9116 15260
rect 9172 15258 9196 15260
rect 9034 15206 9036 15258
rect 9098 15206 9110 15258
rect 9172 15206 9174 15258
rect 9012 15204 9036 15206
rect 9092 15204 9116 15206
rect 9172 15204 9196 15206
rect 8956 15184 9252 15204
rect 9324 14634 9352 26862
rect 9416 21962 9444 31078
rect 9680 30728 9732 30734
rect 9680 30670 9732 30676
rect 9692 30190 9720 30670
rect 9784 30394 9812 39520
rect 9876 39494 10180 39520
rect 10336 39494 10640 39520
rect 9772 30388 9824 30394
rect 9772 30330 9824 30336
rect 9770 30288 9826 30297
rect 9770 30223 9826 30232
rect 9680 30184 9732 30190
rect 9680 30126 9732 30132
rect 9588 30048 9640 30054
rect 9588 29990 9640 29996
rect 9496 29504 9548 29510
rect 9496 29446 9548 29452
rect 9508 23202 9536 29446
rect 9600 23338 9628 29990
rect 9692 29850 9720 30126
rect 9784 30122 9812 30223
rect 9772 30116 9824 30122
rect 9772 30058 9824 30064
rect 9680 29844 9732 29850
rect 9680 29786 9732 29792
rect 9876 25401 9904 39494
rect 9956 30388 10008 30394
rect 9956 30330 10008 30336
rect 9862 25392 9918 25401
rect 9862 25327 9918 25336
rect 9600 23322 9720 23338
rect 9600 23316 9732 23322
rect 9600 23310 9680 23316
rect 9680 23258 9732 23264
rect 9864 23248 9916 23254
rect 9508 23186 9720 23202
rect 9864 23190 9916 23196
rect 9508 23180 9732 23186
rect 9508 23174 9680 23180
rect 9404 21956 9456 21962
rect 9404 21898 9456 21904
rect 9416 21865 9444 21898
rect 9402 21856 9458 21865
rect 9402 21791 9458 21800
rect 9600 14958 9628 23174
rect 9680 23122 9732 23128
rect 9680 22976 9732 22982
rect 9680 22918 9732 22924
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 9692 14657 9720 22918
rect 9876 22642 9904 23190
rect 9968 23089 9996 30330
rect 10336 28966 10364 39494
rect 10980 35193 11008 39520
rect 10966 35184 11022 35193
rect 10966 35119 11022 35128
rect 11348 35057 11376 39520
rect 11808 37754 11836 39520
rect 11532 37726 11836 37754
rect 11992 39494 12204 39520
rect 11334 35048 11390 35057
rect 11334 34983 11390 34992
rect 11532 34649 11560 37726
rect 11622 37564 11918 37584
rect 11678 37562 11702 37564
rect 11758 37562 11782 37564
rect 11838 37562 11862 37564
rect 11700 37510 11702 37562
rect 11764 37510 11776 37562
rect 11838 37510 11840 37562
rect 11678 37508 11702 37510
rect 11758 37508 11782 37510
rect 11838 37508 11862 37510
rect 11622 37488 11918 37508
rect 11622 36476 11918 36496
rect 11678 36474 11702 36476
rect 11758 36474 11782 36476
rect 11838 36474 11862 36476
rect 11700 36422 11702 36474
rect 11764 36422 11776 36474
rect 11838 36422 11840 36474
rect 11678 36420 11702 36422
rect 11758 36420 11782 36422
rect 11838 36420 11862 36422
rect 11622 36400 11918 36420
rect 11622 35388 11918 35408
rect 11678 35386 11702 35388
rect 11758 35386 11782 35388
rect 11838 35386 11862 35388
rect 11700 35334 11702 35386
rect 11764 35334 11776 35386
rect 11838 35334 11840 35386
rect 11678 35332 11702 35334
rect 11758 35332 11782 35334
rect 11838 35332 11862 35334
rect 11622 35312 11918 35332
rect 11518 34640 11574 34649
rect 11518 34575 11574 34584
rect 11622 34300 11918 34320
rect 11678 34298 11702 34300
rect 11758 34298 11782 34300
rect 11838 34298 11862 34300
rect 11700 34246 11702 34298
rect 11764 34246 11776 34298
rect 11838 34246 11840 34298
rect 11678 34244 11702 34246
rect 11758 34244 11782 34246
rect 11838 34244 11862 34246
rect 11622 34224 11918 34244
rect 11622 33212 11918 33232
rect 11678 33210 11702 33212
rect 11758 33210 11782 33212
rect 11838 33210 11862 33212
rect 11700 33158 11702 33210
rect 11764 33158 11776 33210
rect 11838 33158 11840 33210
rect 11678 33156 11702 33158
rect 11758 33156 11782 33158
rect 11838 33156 11862 33158
rect 11622 33136 11918 33156
rect 11622 32124 11918 32144
rect 11678 32122 11702 32124
rect 11758 32122 11782 32124
rect 11838 32122 11862 32124
rect 11700 32070 11702 32122
rect 11764 32070 11776 32122
rect 11838 32070 11840 32122
rect 11678 32068 11702 32070
rect 11758 32068 11782 32070
rect 11838 32068 11862 32070
rect 11622 32048 11918 32068
rect 11622 31036 11918 31056
rect 11678 31034 11702 31036
rect 11758 31034 11782 31036
rect 11838 31034 11862 31036
rect 11700 30982 11702 31034
rect 11764 30982 11776 31034
rect 11838 30982 11840 31034
rect 11678 30980 11702 30982
rect 11758 30980 11782 30982
rect 11838 30980 11862 30982
rect 11622 30960 11918 30980
rect 11622 29948 11918 29968
rect 11678 29946 11702 29948
rect 11758 29946 11782 29948
rect 11838 29946 11862 29948
rect 11700 29894 11702 29946
rect 11764 29894 11776 29946
rect 11838 29894 11840 29946
rect 11678 29892 11702 29894
rect 11758 29892 11782 29894
rect 11838 29892 11862 29894
rect 11622 29872 11918 29892
rect 10324 28960 10376 28966
rect 10324 28902 10376 28908
rect 10600 28960 10652 28966
rect 10600 28902 10652 28908
rect 10140 23112 10192 23118
rect 9954 23080 10010 23089
rect 10140 23054 10192 23060
rect 10324 23112 10376 23118
rect 10324 23054 10376 23060
rect 9954 23015 10010 23024
rect 10152 22710 10180 23054
rect 10336 22778 10364 23054
rect 10324 22772 10376 22778
rect 10324 22714 10376 22720
rect 10140 22704 10192 22710
rect 10140 22646 10192 22652
rect 9864 22636 9916 22642
rect 9864 22578 9916 22584
rect 10048 22636 10100 22642
rect 10048 22578 10100 22584
rect 9876 22545 9904 22578
rect 9862 22536 9918 22545
rect 9862 22471 9918 22480
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9784 21865 9812 22374
rect 10060 22166 10088 22578
rect 10152 22234 10180 22646
rect 10140 22228 10192 22234
rect 10140 22170 10192 22176
rect 10048 22160 10100 22166
rect 10048 22102 10100 22108
rect 9770 21856 9826 21865
rect 9770 21791 9826 21800
rect 9770 21040 9826 21049
rect 9770 20975 9826 20984
rect 9678 14648 9734 14657
rect 9324 14606 9444 14634
rect 9310 14512 9366 14521
rect 9310 14447 9366 14456
rect 8956 14172 9252 14192
rect 9012 14170 9036 14172
rect 9092 14170 9116 14172
rect 9172 14170 9196 14172
rect 9034 14118 9036 14170
rect 9098 14118 9110 14170
rect 9172 14118 9174 14170
rect 9012 14116 9036 14118
rect 9092 14116 9116 14118
rect 9172 14116 9196 14118
rect 8956 14096 9252 14116
rect 8956 13084 9252 13104
rect 9012 13082 9036 13084
rect 9092 13082 9116 13084
rect 9172 13082 9196 13084
rect 9034 13030 9036 13082
rect 9098 13030 9110 13082
rect 9172 13030 9174 13082
rect 9012 13028 9036 13030
rect 9092 13028 9116 13030
rect 9172 13028 9196 13030
rect 8956 13008 9252 13028
rect 8944 12912 8996 12918
rect 8944 12854 8996 12860
rect 8956 12186 8984 12854
rect 8864 12158 8984 12186
rect 8864 6905 8892 12158
rect 8956 11996 9252 12016
rect 9012 11994 9036 11996
rect 9092 11994 9116 11996
rect 9172 11994 9196 11996
rect 9034 11942 9036 11994
rect 9098 11942 9110 11994
rect 9172 11942 9174 11994
rect 9012 11940 9036 11942
rect 9092 11940 9116 11942
rect 9172 11940 9196 11942
rect 8956 11920 9252 11940
rect 8956 10908 9252 10928
rect 9012 10906 9036 10908
rect 9092 10906 9116 10908
rect 9172 10906 9196 10908
rect 9034 10854 9036 10906
rect 9098 10854 9110 10906
rect 9172 10854 9174 10906
rect 9012 10852 9036 10854
rect 9092 10852 9116 10854
rect 9172 10852 9196 10854
rect 8956 10832 9252 10852
rect 8956 9820 9252 9840
rect 9012 9818 9036 9820
rect 9092 9818 9116 9820
rect 9172 9818 9196 9820
rect 9034 9766 9036 9818
rect 9098 9766 9110 9818
rect 9172 9766 9174 9818
rect 9012 9764 9036 9766
rect 9092 9764 9116 9766
rect 9172 9764 9196 9766
rect 8956 9744 9252 9764
rect 8956 8732 9252 8752
rect 9012 8730 9036 8732
rect 9092 8730 9116 8732
rect 9172 8730 9196 8732
rect 9034 8678 9036 8730
rect 9098 8678 9110 8730
rect 9172 8678 9174 8730
rect 9012 8676 9036 8678
rect 9092 8676 9116 8678
rect 9172 8676 9196 8678
rect 8956 8656 9252 8676
rect 8956 7644 9252 7664
rect 9012 7642 9036 7644
rect 9092 7642 9116 7644
rect 9172 7642 9196 7644
rect 9034 7590 9036 7642
rect 9098 7590 9110 7642
rect 9172 7590 9174 7642
rect 9012 7588 9036 7590
rect 9092 7588 9116 7590
rect 9172 7588 9196 7590
rect 8956 7568 9252 7588
rect 8850 6896 8906 6905
rect 8850 6831 8906 6840
rect 8956 6556 9252 6576
rect 9012 6554 9036 6556
rect 9092 6554 9116 6556
rect 9172 6554 9196 6556
rect 9034 6502 9036 6554
rect 9098 6502 9110 6554
rect 9172 6502 9174 6554
rect 9012 6500 9036 6502
rect 9092 6500 9116 6502
rect 9172 6500 9196 6502
rect 8956 6480 9252 6500
rect 8852 6384 8904 6390
rect 8850 6352 8852 6361
rect 8904 6352 8906 6361
rect 8850 6287 8906 6296
rect 8956 5468 9252 5488
rect 9012 5466 9036 5468
rect 9092 5466 9116 5468
rect 9172 5466 9196 5468
rect 9034 5414 9036 5466
rect 9098 5414 9110 5466
rect 9172 5414 9174 5466
rect 9012 5412 9036 5414
rect 9092 5412 9116 5414
rect 9172 5412 9196 5414
rect 8956 5392 9252 5412
rect 8956 4380 9252 4400
rect 9012 4378 9036 4380
rect 9092 4378 9116 4380
rect 9172 4378 9196 4380
rect 9034 4326 9036 4378
rect 9098 4326 9110 4378
rect 9172 4326 9174 4378
rect 9012 4324 9036 4326
rect 9092 4324 9116 4326
rect 9172 4324 9196 4326
rect 8956 4304 9252 4324
rect 8956 3292 9252 3312
rect 9012 3290 9036 3292
rect 9092 3290 9116 3292
rect 9172 3290 9196 3292
rect 9034 3238 9036 3290
rect 9098 3238 9110 3290
rect 9172 3238 9174 3290
rect 9012 3236 9036 3238
rect 9092 3236 9116 3238
rect 9172 3236 9196 3238
rect 8956 3216 9252 3236
rect 8668 2984 8720 2990
rect 8668 2926 8720 2932
rect 8850 2952 8906 2961
rect 8850 2887 8906 2896
rect 8864 2854 8892 2887
rect 8852 2848 8904 2854
rect 8852 2790 8904 2796
rect 8760 2304 8812 2310
rect 8758 2272 8760 2281
rect 8812 2272 8814 2281
rect 8758 2207 8814 2216
rect 8956 2204 9252 2224
rect 9012 2202 9036 2204
rect 9092 2202 9116 2204
rect 9172 2202 9196 2204
rect 9034 2150 9036 2202
rect 9098 2150 9110 2202
rect 9172 2150 9174 2202
rect 9012 2148 9036 2150
rect 9092 2148 9116 2150
rect 9172 2148 9196 2150
rect 8956 2128 9252 2148
rect 9324 1442 9352 14447
rect 9416 12918 9444 14606
rect 9678 14583 9734 14592
rect 9404 12912 9456 12918
rect 9404 12854 9456 12860
rect 9404 6112 9456 6118
rect 9404 6054 9456 6060
rect 9416 3369 9444 6054
rect 9402 3360 9458 3369
rect 9402 3295 9458 3304
rect 9404 2304 9456 2310
rect 9402 2272 9404 2281
rect 9456 2272 9458 2281
rect 9402 2207 9458 2216
rect 9402 1864 9458 1873
rect 9402 1799 9458 1808
rect 8956 1414 9352 1442
rect 8956 480 8984 1414
rect 9416 480 9444 1799
rect 9784 480 9812 20975
rect 10060 20505 10088 22102
rect 10046 20496 10102 20505
rect 10046 20431 10102 20440
rect 10612 19378 10640 28902
rect 11622 28860 11918 28880
rect 11678 28858 11702 28860
rect 11758 28858 11782 28860
rect 11838 28858 11862 28860
rect 11700 28806 11702 28858
rect 11764 28806 11776 28858
rect 11838 28806 11840 28858
rect 11678 28804 11702 28806
rect 11758 28804 11782 28806
rect 11838 28804 11862 28806
rect 11622 28784 11918 28804
rect 11622 27772 11918 27792
rect 11678 27770 11702 27772
rect 11758 27770 11782 27772
rect 11838 27770 11862 27772
rect 11700 27718 11702 27770
rect 11764 27718 11776 27770
rect 11838 27718 11840 27770
rect 11678 27716 11702 27718
rect 11758 27716 11782 27718
rect 11838 27716 11862 27718
rect 11622 27696 11918 27716
rect 11622 26684 11918 26704
rect 11678 26682 11702 26684
rect 11758 26682 11782 26684
rect 11838 26682 11862 26684
rect 11700 26630 11702 26682
rect 11764 26630 11776 26682
rect 11838 26630 11840 26682
rect 11678 26628 11702 26630
rect 11758 26628 11782 26630
rect 11838 26628 11862 26630
rect 11622 26608 11918 26628
rect 11622 25596 11918 25616
rect 11678 25594 11702 25596
rect 11758 25594 11782 25596
rect 11838 25594 11862 25596
rect 11700 25542 11702 25594
rect 11764 25542 11776 25594
rect 11838 25542 11840 25594
rect 11678 25540 11702 25542
rect 11758 25540 11782 25542
rect 11838 25540 11862 25542
rect 11622 25520 11918 25540
rect 11622 24508 11918 24528
rect 11678 24506 11702 24508
rect 11758 24506 11782 24508
rect 11838 24506 11862 24508
rect 11700 24454 11702 24506
rect 11764 24454 11776 24506
rect 11838 24454 11840 24506
rect 11678 24452 11702 24454
rect 11758 24452 11782 24454
rect 11838 24452 11862 24454
rect 11622 24432 11918 24452
rect 11622 23420 11918 23440
rect 11678 23418 11702 23420
rect 11758 23418 11782 23420
rect 11838 23418 11862 23420
rect 11700 23366 11702 23418
rect 11764 23366 11776 23418
rect 11838 23366 11840 23418
rect 11678 23364 11702 23366
rect 11758 23364 11782 23366
rect 11838 23364 11862 23366
rect 11622 23344 11918 23364
rect 10784 23316 10836 23322
rect 10784 23258 10836 23264
rect 10796 22778 10824 23258
rect 11992 23254 12020 39494
rect 12346 34640 12402 34649
rect 12346 34575 12402 34584
rect 12360 31498 12388 34575
rect 12360 31482 12480 31498
rect 12360 31476 12492 31482
rect 12360 31470 12440 31476
rect 12440 31418 12492 31424
rect 12440 31272 12492 31278
rect 12440 31214 12492 31220
rect 12254 25256 12310 25265
rect 12254 25191 12310 25200
rect 12070 24712 12126 24721
rect 12070 24647 12126 24656
rect 12084 24410 12112 24647
rect 12072 24404 12124 24410
rect 12072 24346 12124 24352
rect 12072 24268 12124 24274
rect 12072 24210 12124 24216
rect 12084 23526 12112 24210
rect 12072 23520 12124 23526
rect 12070 23488 12072 23497
rect 12124 23488 12126 23497
rect 12070 23423 12126 23432
rect 11980 23248 12032 23254
rect 11058 23216 11114 23225
rect 11980 23190 12032 23196
rect 11058 23151 11114 23160
rect 10784 22772 10836 22778
rect 10784 22714 10836 22720
rect 11072 22137 11100 23151
rect 11622 22332 11918 22352
rect 11678 22330 11702 22332
rect 11758 22330 11782 22332
rect 11838 22330 11862 22332
rect 11700 22278 11702 22330
rect 11764 22278 11776 22330
rect 11838 22278 11840 22330
rect 11678 22276 11702 22278
rect 11758 22276 11782 22278
rect 11838 22276 11862 22278
rect 11622 22256 11918 22276
rect 11058 22128 11114 22137
rect 11058 22063 11114 22072
rect 11622 21244 11918 21264
rect 11678 21242 11702 21244
rect 11758 21242 11782 21244
rect 11838 21242 11862 21244
rect 11700 21190 11702 21242
rect 11764 21190 11776 21242
rect 11838 21190 11840 21242
rect 11678 21188 11702 21190
rect 11758 21188 11782 21190
rect 11838 21188 11862 21190
rect 11622 21168 11918 21188
rect 11150 20224 11206 20233
rect 11150 20159 11206 20168
rect 10416 19372 10468 19378
rect 10416 19314 10468 19320
rect 10600 19372 10652 19378
rect 10600 19314 10652 19320
rect 10138 9072 10194 9081
rect 10138 9007 10194 9016
rect 9954 3496 10010 3505
rect 9954 3431 10010 3440
rect 9968 3194 9996 3431
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 9968 1465 9996 2246
rect 9954 1456 10010 1465
rect 9954 1391 10010 1400
rect 10152 480 10180 9007
rect 10428 6882 10456 19314
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 11072 15178 11100 15846
rect 10888 15150 11100 15178
rect 10888 14822 10916 15150
rect 11164 15042 11192 20159
rect 11622 20156 11918 20176
rect 11678 20154 11702 20156
rect 11758 20154 11782 20156
rect 11838 20154 11862 20156
rect 11700 20102 11702 20154
rect 11764 20102 11776 20154
rect 11838 20102 11840 20154
rect 11678 20100 11702 20102
rect 11758 20100 11782 20102
rect 11838 20100 11862 20102
rect 11622 20080 11918 20100
rect 11622 19068 11918 19088
rect 11678 19066 11702 19068
rect 11758 19066 11782 19068
rect 11838 19066 11862 19068
rect 11700 19014 11702 19066
rect 11764 19014 11776 19066
rect 11838 19014 11840 19066
rect 11678 19012 11702 19014
rect 11758 19012 11782 19014
rect 11838 19012 11862 19014
rect 11622 18992 11918 19012
rect 11622 17980 11918 18000
rect 11678 17978 11702 17980
rect 11758 17978 11782 17980
rect 11838 17978 11862 17980
rect 11700 17926 11702 17978
rect 11764 17926 11776 17978
rect 11838 17926 11840 17978
rect 11678 17924 11702 17926
rect 11758 17924 11782 17926
rect 11838 17924 11862 17926
rect 11622 17904 11918 17924
rect 12268 17241 12296 25191
rect 12452 22137 12480 31214
rect 12544 26994 12572 39520
rect 13004 31770 13032 39520
rect 13372 35601 13400 39520
rect 13358 35592 13414 35601
rect 13358 35527 13414 35536
rect 12912 31742 13032 31770
rect 12912 28966 12940 31742
rect 12716 28960 12768 28966
rect 12716 28902 12768 28908
rect 12900 28960 12952 28966
rect 12900 28902 12952 28908
rect 12532 26988 12584 26994
rect 12532 26930 12584 26936
rect 12438 22128 12494 22137
rect 12438 22063 12494 22072
rect 12452 21842 12480 22063
rect 12360 21814 12480 21842
rect 12360 19922 12388 21814
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12360 19378 12388 19858
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 12452 18170 12480 19654
rect 12728 19378 12756 28902
rect 13176 26988 13228 26994
rect 13176 26930 13228 26936
rect 12808 26920 12860 26926
rect 12808 26862 12860 26868
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12360 18142 12480 18170
rect 12254 17232 12310 17241
rect 12254 17167 12310 17176
rect 11622 16892 11918 16912
rect 11678 16890 11702 16892
rect 11758 16890 11782 16892
rect 11838 16890 11862 16892
rect 11700 16838 11702 16890
rect 11764 16838 11776 16890
rect 11838 16838 11840 16890
rect 11678 16836 11702 16838
rect 11758 16836 11782 16838
rect 11838 16836 11862 16838
rect 11622 16816 11918 16836
rect 12268 16794 12296 17167
rect 12256 16788 12308 16794
rect 12256 16730 12308 16736
rect 11518 16688 11574 16697
rect 11518 16623 11520 16632
rect 11572 16623 11574 16632
rect 11612 16652 11664 16658
rect 11520 16594 11572 16600
rect 11612 16594 11664 16600
rect 11532 16250 11560 16594
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11624 15978 11652 16594
rect 11612 15972 11664 15978
rect 11612 15914 11664 15920
rect 11622 15804 11918 15824
rect 11678 15802 11702 15804
rect 11758 15802 11782 15804
rect 11838 15802 11862 15804
rect 11700 15750 11702 15802
rect 11764 15750 11776 15802
rect 11838 15750 11840 15802
rect 11678 15748 11702 15750
rect 11758 15748 11782 15750
rect 11838 15748 11862 15750
rect 11622 15728 11918 15748
rect 11072 15014 11192 15042
rect 10876 14816 10928 14822
rect 10876 14758 10928 14764
rect 10888 13938 10916 14758
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10598 9480 10654 9489
rect 10598 9415 10654 9424
rect 10612 9178 10640 9415
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10520 8362 10548 8978
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10336 6854 10456 6882
rect 10336 6225 10364 6854
rect 10414 6760 10470 6769
rect 10414 6695 10470 6704
rect 10428 6458 10456 6695
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10322 6216 10378 6225
rect 10322 6151 10378 6160
rect 10520 4185 10548 8298
rect 10600 6656 10652 6662
rect 10600 6598 10652 6604
rect 10612 4729 10640 6598
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10598 4720 10654 4729
rect 10598 4655 10654 4664
rect 10506 4176 10562 4185
rect 10506 4111 10562 4120
rect 10598 4040 10654 4049
rect 10598 3975 10654 3984
rect 10414 3224 10470 3233
rect 10414 3159 10416 3168
rect 10468 3159 10470 3168
rect 10416 3130 10468 3136
rect 10428 2990 10456 3130
rect 10416 2984 10468 2990
rect 10416 2926 10468 2932
rect 10414 2544 10470 2553
rect 10414 2479 10416 2488
rect 10468 2479 10470 2488
rect 10416 2450 10468 2456
rect 10612 480 10640 3975
rect 10980 3505 11008 6054
rect 10966 3496 11022 3505
rect 10966 3431 11022 3440
rect 10966 3360 11022 3369
rect 10966 3295 11022 3304
rect 10980 480 11008 3295
rect 11072 1426 11100 15014
rect 11622 14716 11918 14736
rect 11678 14714 11702 14716
rect 11758 14714 11782 14716
rect 11838 14714 11862 14716
rect 11700 14662 11702 14714
rect 11764 14662 11776 14714
rect 11838 14662 11840 14714
rect 11678 14660 11702 14662
rect 11758 14660 11782 14662
rect 11838 14660 11862 14662
rect 11622 14640 11918 14660
rect 11622 13628 11918 13648
rect 11678 13626 11702 13628
rect 11758 13626 11782 13628
rect 11838 13626 11862 13628
rect 11700 13574 11702 13626
rect 11764 13574 11776 13626
rect 11838 13574 11840 13626
rect 11678 13572 11702 13574
rect 11758 13572 11782 13574
rect 11838 13572 11862 13574
rect 11622 13552 11918 13572
rect 11622 12540 11918 12560
rect 11678 12538 11702 12540
rect 11758 12538 11782 12540
rect 11838 12538 11862 12540
rect 11700 12486 11702 12538
rect 11764 12486 11776 12538
rect 11838 12486 11840 12538
rect 11678 12484 11702 12486
rect 11758 12484 11782 12486
rect 11838 12484 11862 12486
rect 11622 12464 11918 12484
rect 11622 11452 11918 11472
rect 11678 11450 11702 11452
rect 11758 11450 11782 11452
rect 11838 11450 11862 11452
rect 11700 11398 11702 11450
rect 11764 11398 11776 11450
rect 11838 11398 11840 11450
rect 11678 11396 11702 11398
rect 11758 11396 11782 11398
rect 11838 11396 11862 11398
rect 11622 11376 11918 11396
rect 11622 10364 11918 10384
rect 11678 10362 11702 10364
rect 11758 10362 11782 10364
rect 11838 10362 11862 10364
rect 11700 10310 11702 10362
rect 11764 10310 11776 10362
rect 11838 10310 11840 10362
rect 11678 10308 11702 10310
rect 11758 10308 11782 10310
rect 11838 10308 11862 10310
rect 11622 10288 11918 10308
rect 11622 9276 11918 9296
rect 11678 9274 11702 9276
rect 11758 9274 11782 9276
rect 11838 9274 11862 9276
rect 11700 9222 11702 9274
rect 11764 9222 11776 9274
rect 11838 9222 11840 9274
rect 11678 9220 11702 9222
rect 11758 9220 11782 9222
rect 11838 9220 11862 9222
rect 11622 9200 11918 9220
rect 11622 8188 11918 8208
rect 11678 8186 11702 8188
rect 11758 8186 11782 8188
rect 11838 8186 11862 8188
rect 11700 8134 11702 8186
rect 11764 8134 11776 8186
rect 11838 8134 11840 8186
rect 11678 8132 11702 8134
rect 11758 8132 11782 8134
rect 11838 8132 11862 8134
rect 11622 8112 11918 8132
rect 11622 7100 11918 7120
rect 11678 7098 11702 7100
rect 11758 7098 11782 7100
rect 11838 7098 11862 7100
rect 11700 7046 11702 7098
rect 11764 7046 11776 7098
rect 11838 7046 11840 7098
rect 11678 7044 11702 7046
rect 11758 7044 11782 7046
rect 11838 7044 11862 7046
rect 11622 7024 11918 7044
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 11256 6458 11284 6802
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 11622 6012 11918 6032
rect 11678 6010 11702 6012
rect 11758 6010 11782 6012
rect 11838 6010 11862 6012
rect 11700 5958 11702 6010
rect 11764 5958 11776 6010
rect 11838 5958 11840 6010
rect 11678 5956 11702 5958
rect 11758 5956 11782 5958
rect 11838 5956 11862 5958
rect 11622 5936 11918 5956
rect 11334 5808 11390 5817
rect 11334 5743 11390 5752
rect 11150 3768 11206 3777
rect 11150 3703 11206 3712
rect 11164 3369 11192 3703
rect 11150 3360 11206 3369
rect 11150 3295 11206 3304
rect 11060 1420 11112 1426
rect 11060 1362 11112 1368
rect 11348 480 11376 5743
rect 12360 5001 12388 18142
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12346 4992 12402 5001
rect 11622 4924 11918 4944
rect 12346 4927 12402 4936
rect 11678 4922 11702 4924
rect 11758 4922 11782 4924
rect 11838 4922 11862 4924
rect 11700 4870 11702 4922
rect 11764 4870 11776 4922
rect 11838 4870 11840 4922
rect 11678 4868 11702 4870
rect 11758 4868 11782 4870
rect 11838 4868 11862 4870
rect 11622 4848 11918 4868
rect 11426 3904 11482 3913
rect 11482 3862 11560 3890
rect 11426 3839 11482 3848
rect 11428 3120 11480 3126
rect 11426 3088 11428 3097
rect 11480 3088 11482 3097
rect 11426 3023 11482 3032
rect 11426 2680 11482 2689
rect 11426 2615 11428 2624
rect 11480 2615 11482 2624
rect 11428 2586 11480 2592
rect 11532 762 11560 3862
rect 11622 3836 11918 3856
rect 11678 3834 11702 3836
rect 11758 3834 11782 3836
rect 11838 3834 11862 3836
rect 11700 3782 11702 3834
rect 11764 3782 11776 3834
rect 11838 3782 11840 3834
rect 11678 3780 11702 3782
rect 11758 3780 11782 3782
rect 11838 3780 11862 3782
rect 11622 3760 11918 3780
rect 11610 3632 11666 3641
rect 11610 3567 11666 3576
rect 11624 3097 11652 3567
rect 12452 3097 12480 10406
rect 12530 9616 12586 9625
rect 12530 9551 12586 9560
rect 12544 9178 12572 9551
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12636 3369 12664 8230
rect 12820 6458 12848 26862
rect 12992 19372 13044 19378
rect 12992 19314 13044 19320
rect 13004 12458 13032 19314
rect 12912 12430 13032 12458
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 12622 3360 12678 3369
rect 12622 3295 12678 3304
rect 11610 3088 11666 3097
rect 11610 3023 11666 3032
rect 12438 3088 12494 3097
rect 12438 3023 12494 3032
rect 12622 2952 12678 2961
rect 12622 2887 12678 2896
rect 12636 2854 12664 2887
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 11622 2748 11918 2768
rect 11678 2746 11702 2748
rect 11758 2746 11782 2748
rect 11838 2746 11862 2748
rect 11700 2694 11702 2746
rect 11764 2694 11776 2746
rect 11838 2694 11840 2746
rect 11678 2692 11702 2694
rect 11758 2692 11782 2694
rect 11838 2692 11862 2694
rect 11622 2672 11918 2692
rect 12912 2553 12940 12430
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 13096 8401 13124 8978
rect 13082 8392 13138 8401
rect 13082 8327 13084 8336
rect 13136 8327 13138 8336
rect 13084 8298 13136 8304
rect 13188 3233 13216 26930
rect 13740 26926 13768 39520
rect 14108 39494 14228 39520
rect 14108 27062 14136 39494
rect 14568 37210 14596 39520
rect 14568 37182 14688 37210
rect 14289 37020 14585 37040
rect 14345 37018 14369 37020
rect 14425 37018 14449 37020
rect 14505 37018 14529 37020
rect 14367 36966 14369 37018
rect 14431 36966 14443 37018
rect 14505 36966 14507 37018
rect 14345 36964 14369 36966
rect 14425 36964 14449 36966
rect 14505 36964 14529 36966
rect 14289 36944 14585 36964
rect 14289 35932 14585 35952
rect 14345 35930 14369 35932
rect 14425 35930 14449 35932
rect 14505 35930 14529 35932
rect 14367 35878 14369 35930
rect 14431 35878 14443 35930
rect 14505 35878 14507 35930
rect 14345 35876 14369 35878
rect 14425 35876 14449 35878
rect 14505 35876 14529 35878
rect 14289 35856 14585 35876
rect 14289 34844 14585 34864
rect 14345 34842 14369 34844
rect 14425 34842 14449 34844
rect 14505 34842 14529 34844
rect 14367 34790 14369 34842
rect 14431 34790 14443 34842
rect 14505 34790 14507 34842
rect 14345 34788 14369 34790
rect 14425 34788 14449 34790
rect 14505 34788 14529 34790
rect 14289 34768 14585 34788
rect 14289 33756 14585 33776
rect 14345 33754 14369 33756
rect 14425 33754 14449 33756
rect 14505 33754 14529 33756
rect 14367 33702 14369 33754
rect 14431 33702 14443 33754
rect 14505 33702 14507 33754
rect 14345 33700 14369 33702
rect 14425 33700 14449 33702
rect 14505 33700 14529 33702
rect 14289 33680 14585 33700
rect 14289 32668 14585 32688
rect 14345 32666 14369 32668
rect 14425 32666 14449 32668
rect 14505 32666 14529 32668
rect 14367 32614 14369 32666
rect 14431 32614 14443 32666
rect 14505 32614 14507 32666
rect 14345 32612 14369 32614
rect 14425 32612 14449 32614
rect 14505 32612 14529 32614
rect 14289 32592 14585 32612
rect 14289 31580 14585 31600
rect 14345 31578 14369 31580
rect 14425 31578 14449 31580
rect 14505 31578 14529 31580
rect 14367 31526 14369 31578
rect 14431 31526 14443 31578
rect 14505 31526 14507 31578
rect 14345 31524 14369 31526
rect 14425 31524 14449 31526
rect 14505 31524 14529 31526
rect 14289 31504 14585 31524
rect 14289 30492 14585 30512
rect 14345 30490 14369 30492
rect 14425 30490 14449 30492
rect 14505 30490 14529 30492
rect 14367 30438 14369 30490
rect 14431 30438 14443 30490
rect 14505 30438 14507 30490
rect 14345 30436 14369 30438
rect 14425 30436 14449 30438
rect 14505 30436 14529 30438
rect 14289 30416 14585 30436
rect 14660 30297 14688 37182
rect 14646 30288 14702 30297
rect 14646 30223 14702 30232
rect 14289 29404 14585 29424
rect 14345 29402 14369 29404
rect 14425 29402 14449 29404
rect 14505 29402 14529 29404
rect 14367 29350 14369 29402
rect 14431 29350 14443 29402
rect 14505 29350 14507 29402
rect 14345 29348 14369 29350
rect 14425 29348 14449 29350
rect 14505 29348 14529 29350
rect 14289 29328 14585 29348
rect 14289 28316 14585 28336
rect 14345 28314 14369 28316
rect 14425 28314 14449 28316
rect 14505 28314 14529 28316
rect 14367 28262 14369 28314
rect 14431 28262 14443 28314
rect 14505 28262 14507 28314
rect 14345 28260 14369 28262
rect 14425 28260 14449 28262
rect 14505 28260 14529 28262
rect 14289 28240 14585 28260
rect 14289 27228 14585 27248
rect 14345 27226 14369 27228
rect 14425 27226 14449 27228
rect 14505 27226 14529 27228
rect 14367 27174 14369 27226
rect 14431 27174 14443 27226
rect 14505 27174 14507 27226
rect 14345 27172 14369 27174
rect 14425 27172 14449 27174
rect 14505 27172 14529 27174
rect 14289 27152 14585 27172
rect 14096 27056 14148 27062
rect 14096 26998 14148 27004
rect 14832 27056 14884 27062
rect 14832 26998 14884 27004
rect 13912 26988 13964 26994
rect 13912 26930 13964 26936
rect 13728 26920 13780 26926
rect 13728 26862 13780 26868
rect 13818 21856 13874 21865
rect 13818 21791 13874 21800
rect 13358 4176 13414 4185
rect 13358 4111 13414 4120
rect 13174 3224 13230 3233
rect 13174 3159 13230 3168
rect 13266 2816 13322 2825
rect 13266 2751 13322 2760
rect 13280 2650 13308 2751
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 12898 2544 12954 2553
rect 12072 2508 12124 2514
rect 12898 2479 12954 2488
rect 12072 2450 12124 2456
rect 12084 2310 12112 2450
rect 12806 2408 12862 2417
rect 12806 2343 12808 2352
rect 12860 2343 12862 2352
rect 12808 2314 12860 2320
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 12530 2272 12586 2281
rect 12084 1902 12112 2246
rect 12530 2207 12586 2216
rect 12072 1896 12124 1902
rect 12072 1838 12124 1844
rect 12164 1420 12216 1426
rect 12164 1362 12216 1368
rect 11532 734 11836 762
rect 11808 480 11836 734
rect 12176 480 12204 1362
rect 12544 480 12572 2207
rect 12990 2000 13046 2009
rect 12990 1935 13046 1944
rect 13004 480 13032 1935
rect 13372 480 13400 4111
rect 13726 3496 13782 3505
rect 13726 3431 13782 3440
rect 13740 480 13768 3431
rect 13832 1426 13860 21791
rect 13924 3194 13952 26930
rect 14004 26920 14056 26926
rect 14004 26862 14056 26868
rect 14016 8430 14044 26862
rect 14096 26784 14148 26790
rect 14096 26726 14148 26732
rect 14108 10810 14136 26726
rect 14289 26140 14585 26160
rect 14345 26138 14369 26140
rect 14425 26138 14449 26140
rect 14505 26138 14529 26140
rect 14367 26086 14369 26138
rect 14431 26086 14443 26138
rect 14505 26086 14507 26138
rect 14345 26084 14369 26086
rect 14425 26084 14449 26086
rect 14505 26084 14529 26086
rect 14289 26064 14585 26084
rect 14289 25052 14585 25072
rect 14345 25050 14369 25052
rect 14425 25050 14449 25052
rect 14505 25050 14529 25052
rect 14367 24998 14369 25050
rect 14431 24998 14443 25050
rect 14505 24998 14507 25050
rect 14345 24996 14369 24998
rect 14425 24996 14449 24998
rect 14505 24996 14529 24998
rect 14289 24976 14585 24996
rect 14289 23964 14585 23984
rect 14345 23962 14369 23964
rect 14425 23962 14449 23964
rect 14505 23962 14529 23964
rect 14367 23910 14369 23962
rect 14431 23910 14443 23962
rect 14505 23910 14507 23962
rect 14345 23908 14369 23910
rect 14425 23908 14449 23910
rect 14505 23908 14529 23910
rect 14289 23888 14585 23908
rect 14186 23488 14242 23497
rect 14186 23423 14242 23432
rect 14200 19310 14228 23423
rect 14289 22876 14585 22896
rect 14345 22874 14369 22876
rect 14425 22874 14449 22876
rect 14505 22874 14529 22876
rect 14367 22822 14369 22874
rect 14431 22822 14443 22874
rect 14505 22822 14507 22874
rect 14345 22820 14369 22822
rect 14425 22820 14449 22822
rect 14505 22820 14529 22822
rect 14289 22800 14585 22820
rect 14289 21788 14585 21808
rect 14345 21786 14369 21788
rect 14425 21786 14449 21788
rect 14505 21786 14529 21788
rect 14367 21734 14369 21786
rect 14431 21734 14443 21786
rect 14505 21734 14507 21786
rect 14345 21732 14369 21734
rect 14425 21732 14449 21734
rect 14505 21732 14529 21734
rect 14289 21712 14585 21732
rect 14289 20700 14585 20720
rect 14345 20698 14369 20700
rect 14425 20698 14449 20700
rect 14505 20698 14529 20700
rect 14367 20646 14369 20698
rect 14431 20646 14443 20698
rect 14505 20646 14507 20698
rect 14345 20644 14369 20646
rect 14425 20644 14449 20646
rect 14505 20644 14529 20646
rect 14289 20624 14585 20644
rect 14289 19612 14585 19632
rect 14345 19610 14369 19612
rect 14425 19610 14449 19612
rect 14505 19610 14529 19612
rect 14367 19558 14369 19610
rect 14431 19558 14443 19610
rect 14505 19558 14507 19610
rect 14345 19556 14369 19558
rect 14425 19556 14449 19558
rect 14505 19556 14529 19558
rect 14289 19536 14585 19556
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 14289 18524 14585 18544
rect 14345 18522 14369 18524
rect 14425 18522 14449 18524
rect 14505 18522 14529 18524
rect 14367 18470 14369 18522
rect 14431 18470 14443 18522
rect 14505 18470 14507 18522
rect 14345 18468 14369 18470
rect 14425 18468 14449 18470
rect 14505 18468 14529 18470
rect 14289 18448 14585 18468
rect 14289 17436 14585 17456
rect 14345 17434 14369 17436
rect 14425 17434 14449 17436
rect 14505 17434 14529 17436
rect 14367 17382 14369 17434
rect 14431 17382 14443 17434
rect 14505 17382 14507 17434
rect 14345 17380 14369 17382
rect 14425 17380 14449 17382
rect 14505 17380 14529 17382
rect 14289 17360 14585 17380
rect 14289 16348 14585 16368
rect 14345 16346 14369 16348
rect 14425 16346 14449 16348
rect 14505 16346 14529 16348
rect 14367 16294 14369 16346
rect 14431 16294 14443 16346
rect 14505 16294 14507 16346
rect 14345 16292 14369 16294
rect 14425 16292 14449 16294
rect 14505 16292 14529 16294
rect 14289 16272 14585 16292
rect 14289 15260 14585 15280
rect 14345 15258 14369 15260
rect 14425 15258 14449 15260
rect 14505 15258 14529 15260
rect 14367 15206 14369 15258
rect 14431 15206 14443 15258
rect 14505 15206 14507 15258
rect 14345 15204 14369 15206
rect 14425 15204 14449 15206
rect 14505 15204 14529 15206
rect 14289 15184 14585 15204
rect 14289 14172 14585 14192
rect 14345 14170 14369 14172
rect 14425 14170 14449 14172
rect 14505 14170 14529 14172
rect 14367 14118 14369 14170
rect 14431 14118 14443 14170
rect 14505 14118 14507 14170
rect 14345 14116 14369 14118
rect 14425 14116 14449 14118
rect 14505 14116 14529 14118
rect 14289 14096 14585 14116
rect 14289 13084 14585 13104
rect 14345 13082 14369 13084
rect 14425 13082 14449 13084
rect 14505 13082 14529 13084
rect 14367 13030 14369 13082
rect 14431 13030 14443 13082
rect 14505 13030 14507 13082
rect 14345 13028 14369 13030
rect 14425 13028 14449 13030
rect 14505 13028 14529 13030
rect 14289 13008 14585 13028
rect 14289 11996 14585 12016
rect 14345 11994 14369 11996
rect 14425 11994 14449 11996
rect 14505 11994 14529 11996
rect 14367 11942 14369 11994
rect 14431 11942 14443 11994
rect 14505 11942 14507 11994
rect 14345 11940 14369 11942
rect 14425 11940 14449 11942
rect 14505 11940 14529 11942
rect 14289 11920 14585 11940
rect 14289 10908 14585 10928
rect 14345 10906 14369 10908
rect 14425 10906 14449 10908
rect 14505 10906 14529 10908
rect 14367 10854 14369 10906
rect 14431 10854 14443 10906
rect 14505 10854 14507 10906
rect 14345 10852 14369 10854
rect 14425 10852 14449 10854
rect 14505 10852 14529 10854
rect 14289 10832 14585 10852
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 14289 9820 14585 9840
rect 14345 9818 14369 9820
rect 14425 9818 14449 9820
rect 14505 9818 14529 9820
rect 14367 9766 14369 9818
rect 14431 9766 14443 9818
rect 14505 9766 14507 9818
rect 14345 9764 14369 9766
rect 14425 9764 14449 9766
rect 14505 9764 14529 9766
rect 14289 9744 14585 9764
rect 14740 9716 14792 9722
rect 14740 9658 14792 9664
rect 14752 9602 14780 9658
rect 14660 9574 14780 9602
rect 14289 8732 14585 8752
rect 14345 8730 14369 8732
rect 14425 8730 14449 8732
rect 14505 8730 14529 8732
rect 14367 8678 14369 8730
rect 14431 8678 14443 8730
rect 14505 8678 14507 8730
rect 14345 8676 14369 8678
rect 14425 8676 14449 8678
rect 14505 8676 14529 8678
rect 14289 8656 14585 8676
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 14289 7644 14585 7664
rect 14345 7642 14369 7644
rect 14425 7642 14449 7644
rect 14505 7642 14529 7644
rect 14367 7590 14369 7642
rect 14431 7590 14443 7642
rect 14505 7590 14507 7642
rect 14345 7588 14369 7590
rect 14425 7588 14449 7590
rect 14505 7588 14529 7590
rect 14289 7568 14585 7588
rect 14289 6556 14585 6576
rect 14345 6554 14369 6556
rect 14425 6554 14449 6556
rect 14505 6554 14529 6556
rect 14367 6502 14369 6554
rect 14431 6502 14443 6554
rect 14505 6502 14507 6554
rect 14345 6500 14369 6502
rect 14425 6500 14449 6502
rect 14505 6500 14529 6502
rect 14289 6480 14585 6500
rect 14289 5468 14585 5488
rect 14345 5466 14369 5468
rect 14425 5466 14449 5468
rect 14505 5466 14529 5468
rect 14367 5414 14369 5466
rect 14431 5414 14443 5466
rect 14505 5414 14507 5466
rect 14345 5412 14369 5414
rect 14425 5412 14449 5414
rect 14505 5412 14529 5414
rect 14289 5392 14585 5412
rect 14289 4380 14585 4400
rect 14345 4378 14369 4380
rect 14425 4378 14449 4380
rect 14505 4378 14529 4380
rect 14367 4326 14369 4378
rect 14431 4326 14443 4378
rect 14505 4326 14507 4378
rect 14345 4324 14369 4326
rect 14425 4324 14449 4326
rect 14505 4324 14529 4326
rect 14289 4304 14585 4324
rect 14660 3398 14688 9574
rect 14648 3392 14700 3398
rect 14648 3334 14700 3340
rect 14289 3292 14585 3312
rect 14345 3290 14369 3292
rect 14425 3290 14449 3292
rect 14505 3290 14529 3292
rect 14367 3238 14369 3290
rect 14431 3238 14443 3290
rect 14505 3238 14507 3290
rect 14345 3236 14369 3238
rect 14425 3236 14449 3238
rect 14505 3236 14529 3238
rect 14289 3216 14585 3236
rect 13912 3188 13964 3194
rect 13912 3130 13964 3136
rect 14844 2922 14872 26998
rect 14936 26926 14964 39520
rect 15396 26994 15424 39520
rect 15384 26988 15436 26994
rect 15384 26930 15436 26936
rect 14924 26920 14976 26926
rect 14924 26862 14976 26868
rect 15764 26790 15792 39520
rect 15752 26784 15804 26790
rect 15752 26726 15804 26732
rect 15750 8392 15806 8401
rect 15750 8327 15806 8336
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 15382 2816 15438 2825
rect 15382 2751 15438 2760
rect 14289 2204 14585 2224
rect 14345 2202 14369 2204
rect 14425 2202 14449 2204
rect 14505 2202 14529 2204
rect 14367 2150 14369 2202
rect 14431 2150 14443 2202
rect 14505 2150 14507 2202
rect 14345 2148 14369 2150
rect 14425 2148 14449 2150
rect 14505 2148 14529 2150
rect 14289 2128 14585 2148
rect 14096 1896 14148 1902
rect 14096 1838 14148 1844
rect 13820 1420 13872 1426
rect 13820 1362 13872 1368
rect 14108 1306 14136 1838
rect 14556 1420 14608 1426
rect 14556 1362 14608 1368
rect 14108 1278 14228 1306
rect 14200 480 14228 1278
rect 14568 480 14596 1362
rect 14924 604 14976 610
rect 14924 546 14976 552
rect 14936 480 14964 546
rect 15396 480 15424 2751
rect 15764 480 15792 8327
rect 202 0 258 480
rect 570 0 626 480
rect 938 0 994 480
rect 1398 0 1454 480
rect 1766 0 1822 480
rect 2134 0 2190 480
rect 2594 0 2650 480
rect 2962 0 3018 480
rect 3330 0 3386 480
rect 3790 0 3846 480
rect 4158 0 4214 480
rect 4526 0 4582 480
rect 4986 0 5042 480
rect 5354 0 5410 480
rect 5722 0 5778 480
rect 6182 0 6238 480
rect 6550 0 6606 480
rect 6918 0 6974 480
rect 7378 0 7434 480
rect 7746 0 7802 480
rect 8206 0 8262 480
rect 8574 0 8630 480
rect 8942 0 8998 480
rect 9402 0 9458 480
rect 9770 0 9826 480
rect 10138 0 10194 480
rect 10598 0 10654 480
rect 10966 0 11022 480
rect 11334 0 11390 480
rect 11794 0 11850 480
rect 12162 0 12218 480
rect 12530 0 12586 480
rect 12990 0 13046 480
rect 13358 0 13414 480
rect 13726 0 13782 480
rect 14186 0 14242 480
rect 14554 0 14610 480
rect 14922 0 14978 480
rect 15382 0 15438 480
rect 15750 0 15806 480
<< via2 >>
rect 1950 36624 2006 36680
rect 1582 29960 1638 30016
rect 1582 16632 1638 16688
rect 2318 35536 2374 35592
rect 1674 15000 1730 15056
rect 1398 12688 1454 12744
rect 1582 9968 1638 10024
rect 1582 6704 1638 6760
rect 1674 3440 1730 3496
rect 2134 25200 2190 25256
rect 1858 22072 1914 22128
rect 2042 17176 2098 17232
rect 1950 15952 2006 16008
rect 2042 13912 2098 13968
rect 1766 3304 1822 3360
rect 2410 28484 2466 28520
rect 2410 28464 2412 28484
rect 2412 28464 2464 28484
rect 2464 28464 2466 28484
rect 2318 16088 2374 16144
rect 3622 37018 3678 37020
rect 3702 37018 3758 37020
rect 3782 37018 3838 37020
rect 3862 37018 3918 37020
rect 3622 36966 3648 37018
rect 3648 36966 3678 37018
rect 3702 36966 3712 37018
rect 3712 36966 3758 37018
rect 3782 36966 3828 37018
rect 3828 36966 3838 37018
rect 3862 36966 3892 37018
rect 3892 36966 3918 37018
rect 3622 36964 3678 36966
rect 3702 36964 3758 36966
rect 3782 36964 3838 36966
rect 3862 36964 3918 36966
rect 3622 35930 3678 35932
rect 3702 35930 3758 35932
rect 3782 35930 3838 35932
rect 3862 35930 3918 35932
rect 3622 35878 3648 35930
rect 3648 35878 3678 35930
rect 3702 35878 3712 35930
rect 3712 35878 3758 35930
rect 3782 35878 3828 35930
rect 3828 35878 3838 35930
rect 3862 35878 3892 35930
rect 3892 35878 3918 35930
rect 3622 35876 3678 35878
rect 3702 35876 3758 35878
rect 3782 35876 3838 35878
rect 3862 35876 3918 35878
rect 3622 34842 3678 34844
rect 3702 34842 3758 34844
rect 3782 34842 3838 34844
rect 3862 34842 3918 34844
rect 3622 34790 3648 34842
rect 3648 34790 3678 34842
rect 3702 34790 3712 34842
rect 3712 34790 3758 34842
rect 3782 34790 3828 34842
rect 3828 34790 3838 34842
rect 3862 34790 3892 34842
rect 3892 34790 3918 34842
rect 3622 34788 3678 34790
rect 3702 34788 3758 34790
rect 3782 34788 3838 34790
rect 3862 34788 3918 34790
rect 3622 33754 3678 33756
rect 3702 33754 3758 33756
rect 3782 33754 3838 33756
rect 3862 33754 3918 33756
rect 3622 33702 3648 33754
rect 3648 33702 3678 33754
rect 3702 33702 3712 33754
rect 3712 33702 3758 33754
rect 3782 33702 3828 33754
rect 3828 33702 3838 33754
rect 3862 33702 3892 33754
rect 3892 33702 3918 33754
rect 3622 33700 3678 33702
rect 3702 33700 3758 33702
rect 3782 33700 3838 33702
rect 3862 33700 3918 33702
rect 3622 32666 3678 32668
rect 3702 32666 3758 32668
rect 3782 32666 3838 32668
rect 3862 32666 3918 32668
rect 3622 32614 3648 32666
rect 3648 32614 3678 32666
rect 3702 32614 3712 32666
rect 3712 32614 3758 32666
rect 3782 32614 3828 32666
rect 3828 32614 3838 32666
rect 3862 32614 3892 32666
rect 3892 32614 3918 32666
rect 3622 32612 3678 32614
rect 3702 32612 3758 32614
rect 3782 32612 3838 32614
rect 3862 32612 3918 32614
rect 3622 31578 3678 31580
rect 3702 31578 3758 31580
rect 3782 31578 3838 31580
rect 3862 31578 3918 31580
rect 3622 31526 3648 31578
rect 3648 31526 3678 31578
rect 3702 31526 3712 31578
rect 3712 31526 3758 31578
rect 3782 31526 3828 31578
rect 3828 31526 3838 31578
rect 3862 31526 3892 31578
rect 3892 31526 3918 31578
rect 3622 31524 3678 31526
rect 3702 31524 3758 31526
rect 3782 31524 3838 31526
rect 3862 31524 3918 31526
rect 3622 30490 3678 30492
rect 3702 30490 3758 30492
rect 3782 30490 3838 30492
rect 3862 30490 3918 30492
rect 3622 30438 3648 30490
rect 3648 30438 3678 30490
rect 3702 30438 3712 30490
rect 3712 30438 3758 30490
rect 3782 30438 3828 30490
rect 3828 30438 3838 30490
rect 3862 30438 3892 30490
rect 3892 30438 3918 30490
rect 3622 30436 3678 30438
rect 3702 30436 3758 30438
rect 3782 30436 3838 30438
rect 3862 30436 3918 30438
rect 3622 29402 3678 29404
rect 3702 29402 3758 29404
rect 3782 29402 3838 29404
rect 3862 29402 3918 29404
rect 3622 29350 3648 29402
rect 3648 29350 3678 29402
rect 3702 29350 3712 29402
rect 3712 29350 3758 29402
rect 3782 29350 3828 29402
rect 3828 29350 3838 29402
rect 3862 29350 3892 29402
rect 3892 29350 3918 29402
rect 3622 29348 3678 29350
rect 3702 29348 3758 29350
rect 3782 29348 3838 29350
rect 3862 29348 3918 29350
rect 3622 28314 3678 28316
rect 3702 28314 3758 28316
rect 3782 28314 3838 28316
rect 3862 28314 3918 28316
rect 3622 28262 3648 28314
rect 3648 28262 3678 28314
rect 3702 28262 3712 28314
rect 3712 28262 3758 28314
rect 3782 28262 3828 28314
rect 3828 28262 3838 28314
rect 3862 28262 3892 28314
rect 3892 28262 3918 28314
rect 3622 28260 3678 28262
rect 3702 28260 3758 28262
rect 3782 28260 3838 28262
rect 3862 28260 3918 28262
rect 3622 27226 3678 27228
rect 3702 27226 3758 27228
rect 3782 27226 3838 27228
rect 3862 27226 3918 27228
rect 3622 27174 3648 27226
rect 3648 27174 3678 27226
rect 3702 27174 3712 27226
rect 3712 27174 3758 27226
rect 3782 27174 3828 27226
rect 3828 27174 3838 27226
rect 3862 27174 3892 27226
rect 3892 27174 3918 27226
rect 3622 27172 3678 27174
rect 3702 27172 3758 27174
rect 3782 27172 3838 27174
rect 3862 27172 3918 27174
rect 2686 6840 2742 6896
rect 3622 26138 3678 26140
rect 3702 26138 3758 26140
rect 3782 26138 3838 26140
rect 3862 26138 3918 26140
rect 3622 26086 3648 26138
rect 3648 26086 3678 26138
rect 3702 26086 3712 26138
rect 3712 26086 3758 26138
rect 3782 26086 3828 26138
rect 3828 26086 3838 26138
rect 3862 26086 3892 26138
rect 3892 26086 3918 26138
rect 3622 26084 3678 26086
rect 3702 26084 3758 26086
rect 3782 26084 3838 26086
rect 3862 26084 3918 26086
rect 3622 25050 3678 25052
rect 3702 25050 3758 25052
rect 3782 25050 3838 25052
rect 3862 25050 3918 25052
rect 3622 24998 3648 25050
rect 3648 24998 3678 25050
rect 3702 24998 3712 25050
rect 3712 24998 3758 25050
rect 3782 24998 3828 25050
rect 3828 24998 3838 25050
rect 3862 24998 3892 25050
rect 3892 24998 3918 25050
rect 3622 24996 3678 24998
rect 3702 24996 3758 24998
rect 3782 24996 3838 24998
rect 3862 24996 3918 24998
rect 3622 23962 3678 23964
rect 3702 23962 3758 23964
rect 3782 23962 3838 23964
rect 3862 23962 3918 23964
rect 3622 23910 3648 23962
rect 3648 23910 3678 23962
rect 3702 23910 3712 23962
rect 3712 23910 3758 23962
rect 3782 23910 3828 23962
rect 3828 23910 3838 23962
rect 3862 23910 3892 23962
rect 3892 23910 3918 23962
rect 3622 23908 3678 23910
rect 3702 23908 3758 23910
rect 3782 23908 3838 23910
rect 3862 23908 3918 23910
rect 3622 22874 3678 22876
rect 3702 22874 3758 22876
rect 3782 22874 3838 22876
rect 3862 22874 3918 22876
rect 3622 22822 3648 22874
rect 3648 22822 3678 22874
rect 3702 22822 3712 22874
rect 3712 22822 3758 22874
rect 3782 22822 3828 22874
rect 3828 22822 3838 22874
rect 3862 22822 3892 22874
rect 3892 22822 3918 22874
rect 3622 22820 3678 22822
rect 3702 22820 3758 22822
rect 3782 22820 3838 22822
rect 3862 22820 3918 22822
rect 3622 21786 3678 21788
rect 3702 21786 3758 21788
rect 3782 21786 3838 21788
rect 3862 21786 3918 21788
rect 3622 21734 3648 21786
rect 3648 21734 3678 21786
rect 3702 21734 3712 21786
rect 3712 21734 3758 21786
rect 3782 21734 3828 21786
rect 3828 21734 3838 21786
rect 3862 21734 3892 21786
rect 3892 21734 3918 21786
rect 3622 21732 3678 21734
rect 3702 21732 3758 21734
rect 3782 21732 3838 21734
rect 3862 21732 3918 21734
rect 3622 20698 3678 20700
rect 3702 20698 3758 20700
rect 3782 20698 3838 20700
rect 3862 20698 3918 20700
rect 3622 20646 3648 20698
rect 3648 20646 3678 20698
rect 3702 20646 3712 20698
rect 3712 20646 3758 20698
rect 3782 20646 3828 20698
rect 3828 20646 3838 20698
rect 3862 20646 3892 20698
rect 3892 20646 3918 20698
rect 3622 20644 3678 20646
rect 3702 20644 3758 20646
rect 3782 20644 3838 20646
rect 3862 20644 3918 20646
rect 3622 19610 3678 19612
rect 3702 19610 3758 19612
rect 3782 19610 3838 19612
rect 3862 19610 3918 19612
rect 3622 19558 3648 19610
rect 3648 19558 3678 19610
rect 3702 19558 3712 19610
rect 3712 19558 3758 19610
rect 3782 19558 3828 19610
rect 3828 19558 3838 19610
rect 3862 19558 3892 19610
rect 3892 19558 3918 19610
rect 3622 19556 3678 19558
rect 3702 19556 3758 19558
rect 3782 19556 3838 19558
rect 3862 19556 3918 19558
rect 3622 18522 3678 18524
rect 3702 18522 3758 18524
rect 3782 18522 3838 18524
rect 3862 18522 3918 18524
rect 3622 18470 3648 18522
rect 3648 18470 3678 18522
rect 3702 18470 3712 18522
rect 3712 18470 3758 18522
rect 3782 18470 3828 18522
rect 3828 18470 3838 18522
rect 3862 18470 3892 18522
rect 3892 18470 3918 18522
rect 3622 18468 3678 18470
rect 3702 18468 3758 18470
rect 3782 18468 3838 18470
rect 3862 18468 3918 18470
rect 3622 17434 3678 17436
rect 3702 17434 3758 17436
rect 3782 17434 3838 17436
rect 3862 17434 3918 17436
rect 3622 17382 3648 17434
rect 3648 17382 3678 17434
rect 3702 17382 3712 17434
rect 3712 17382 3758 17434
rect 3782 17382 3828 17434
rect 3828 17382 3838 17434
rect 3862 17382 3892 17434
rect 3892 17382 3918 17434
rect 3622 17380 3678 17382
rect 3702 17380 3758 17382
rect 3782 17380 3838 17382
rect 3862 17380 3918 17382
rect 3622 16346 3678 16348
rect 3702 16346 3758 16348
rect 3782 16346 3838 16348
rect 3862 16346 3918 16348
rect 3622 16294 3648 16346
rect 3648 16294 3678 16346
rect 3702 16294 3712 16346
rect 3712 16294 3758 16346
rect 3782 16294 3828 16346
rect 3828 16294 3838 16346
rect 3862 16294 3892 16346
rect 3892 16294 3918 16346
rect 3622 16292 3678 16294
rect 3702 16292 3758 16294
rect 3782 16292 3838 16294
rect 3862 16292 3918 16294
rect 3622 15258 3678 15260
rect 3702 15258 3758 15260
rect 3782 15258 3838 15260
rect 3862 15258 3918 15260
rect 3622 15206 3648 15258
rect 3648 15206 3678 15258
rect 3702 15206 3712 15258
rect 3712 15206 3758 15258
rect 3782 15206 3828 15258
rect 3828 15206 3838 15258
rect 3862 15206 3892 15258
rect 3892 15206 3918 15258
rect 3622 15204 3678 15206
rect 3702 15204 3758 15206
rect 3782 15204 3838 15206
rect 3862 15204 3918 15206
rect 3622 14170 3678 14172
rect 3702 14170 3758 14172
rect 3782 14170 3838 14172
rect 3862 14170 3918 14172
rect 3622 14118 3648 14170
rect 3648 14118 3678 14170
rect 3702 14118 3712 14170
rect 3712 14118 3758 14170
rect 3782 14118 3828 14170
rect 3828 14118 3838 14170
rect 3862 14118 3892 14170
rect 3892 14118 3918 14170
rect 3622 14116 3678 14118
rect 3702 14116 3758 14118
rect 3782 14116 3838 14118
rect 3862 14116 3918 14118
rect 3622 13082 3678 13084
rect 3702 13082 3758 13084
rect 3782 13082 3838 13084
rect 3862 13082 3918 13084
rect 3622 13030 3648 13082
rect 3648 13030 3678 13082
rect 3702 13030 3712 13082
rect 3712 13030 3758 13082
rect 3782 13030 3828 13082
rect 3828 13030 3838 13082
rect 3862 13030 3892 13082
rect 3892 13030 3918 13082
rect 3622 13028 3678 13030
rect 3702 13028 3758 13030
rect 3782 13028 3838 13030
rect 3862 13028 3918 13030
rect 3622 11994 3678 11996
rect 3702 11994 3758 11996
rect 3782 11994 3838 11996
rect 3862 11994 3918 11996
rect 3622 11942 3648 11994
rect 3648 11942 3678 11994
rect 3702 11942 3712 11994
rect 3712 11942 3758 11994
rect 3782 11942 3828 11994
rect 3828 11942 3838 11994
rect 3862 11942 3892 11994
rect 3892 11942 3918 11994
rect 3622 11940 3678 11942
rect 3702 11940 3758 11942
rect 3782 11940 3838 11942
rect 3862 11940 3918 11942
rect 3622 10906 3678 10908
rect 3702 10906 3758 10908
rect 3782 10906 3838 10908
rect 3862 10906 3918 10908
rect 3622 10854 3648 10906
rect 3648 10854 3678 10906
rect 3702 10854 3712 10906
rect 3712 10854 3758 10906
rect 3782 10854 3828 10906
rect 3828 10854 3838 10906
rect 3862 10854 3892 10906
rect 3892 10854 3918 10906
rect 3622 10852 3678 10854
rect 3702 10852 3758 10854
rect 3782 10852 3838 10854
rect 3862 10852 3918 10854
rect 3622 9818 3678 9820
rect 3702 9818 3758 9820
rect 3782 9818 3838 9820
rect 3862 9818 3918 9820
rect 3622 9766 3648 9818
rect 3648 9766 3678 9818
rect 3702 9766 3712 9818
rect 3712 9766 3758 9818
rect 3782 9766 3828 9818
rect 3828 9766 3838 9818
rect 3862 9766 3892 9818
rect 3892 9766 3918 9818
rect 3622 9764 3678 9766
rect 3702 9764 3758 9766
rect 3782 9764 3838 9766
rect 3862 9764 3918 9766
rect 3514 9016 3570 9072
rect 3622 8730 3678 8732
rect 3702 8730 3758 8732
rect 3782 8730 3838 8732
rect 3862 8730 3918 8732
rect 3622 8678 3648 8730
rect 3648 8678 3678 8730
rect 3702 8678 3712 8730
rect 3712 8678 3758 8730
rect 3782 8678 3828 8730
rect 3828 8678 3838 8730
rect 3862 8678 3892 8730
rect 3892 8678 3918 8730
rect 3622 8676 3678 8678
rect 3702 8676 3758 8678
rect 3782 8676 3838 8678
rect 3862 8676 3918 8678
rect 3622 7642 3678 7644
rect 3702 7642 3758 7644
rect 3782 7642 3838 7644
rect 3862 7642 3918 7644
rect 3622 7590 3648 7642
rect 3648 7590 3678 7642
rect 3702 7590 3712 7642
rect 3712 7590 3758 7642
rect 3782 7590 3828 7642
rect 3828 7590 3838 7642
rect 3862 7590 3892 7642
rect 3892 7590 3918 7642
rect 3622 7588 3678 7590
rect 3702 7588 3758 7590
rect 3782 7588 3838 7590
rect 3862 7588 3918 7590
rect 3622 6554 3678 6556
rect 3702 6554 3758 6556
rect 3782 6554 3838 6556
rect 3862 6554 3918 6556
rect 3622 6502 3648 6554
rect 3648 6502 3678 6554
rect 3702 6502 3712 6554
rect 3712 6502 3758 6554
rect 3782 6502 3828 6554
rect 3828 6502 3838 6554
rect 3862 6502 3892 6554
rect 3892 6502 3918 6554
rect 3622 6500 3678 6502
rect 3702 6500 3758 6502
rect 3782 6500 3838 6502
rect 3862 6500 3918 6502
rect 3330 6296 3386 6352
rect 2594 5616 2650 5672
rect 3622 5466 3678 5468
rect 3702 5466 3758 5468
rect 3782 5466 3838 5468
rect 3862 5466 3918 5468
rect 3622 5414 3648 5466
rect 3648 5414 3678 5466
rect 3702 5414 3712 5466
rect 3712 5414 3758 5466
rect 3782 5414 3828 5466
rect 3828 5414 3838 5466
rect 3862 5414 3892 5466
rect 3892 5414 3918 5466
rect 3622 5412 3678 5414
rect 3702 5412 3758 5414
rect 3782 5412 3838 5414
rect 3862 5412 3918 5414
rect 3622 4378 3678 4380
rect 3702 4378 3758 4380
rect 3782 4378 3838 4380
rect 3862 4378 3918 4380
rect 3622 4326 3648 4378
rect 3648 4326 3678 4378
rect 3702 4326 3712 4378
rect 3712 4326 3758 4378
rect 3782 4326 3828 4378
rect 3828 4326 3838 4378
rect 3862 4326 3892 4378
rect 3892 4326 3918 4378
rect 3622 4324 3678 4326
rect 3702 4324 3758 4326
rect 3782 4324 3838 4326
rect 3862 4324 3918 4326
rect 4434 34584 4490 34640
rect 4066 25356 4122 25392
rect 4066 25336 4068 25356
rect 4068 25336 4120 25356
rect 4120 25336 4122 25356
rect 4434 29008 4490 29064
rect 4618 28974 4674 29030
rect 4526 28464 4582 28520
rect 4250 25220 4306 25256
rect 4250 25200 4252 25220
rect 4252 25200 4304 25220
rect 4304 25200 4306 25220
rect 4158 21800 4214 21856
rect 4434 21936 4490 21992
rect 4342 15972 4398 16008
rect 4342 15952 4344 15972
rect 4344 15952 4396 15972
rect 4396 15952 4398 15972
rect 4342 15000 4398 15056
rect 4802 16088 4858 16144
rect 4894 15544 4950 15600
rect 4802 15000 4858 15056
rect 4894 14456 4950 14512
rect 4802 13912 4858 13968
rect 4250 7248 4306 7304
rect 4342 5616 4398 5672
rect 3622 3290 3678 3292
rect 3702 3290 3758 3292
rect 3782 3290 3838 3292
rect 3862 3290 3918 3292
rect 3622 3238 3648 3290
rect 3648 3238 3678 3290
rect 3702 3238 3712 3290
rect 3712 3238 3758 3290
rect 3782 3238 3828 3290
rect 3828 3238 3838 3290
rect 3862 3238 3892 3290
rect 3892 3238 3918 3290
rect 3622 3236 3678 3238
rect 3702 3236 3758 3238
rect 3782 3236 3838 3238
rect 3862 3236 3918 3238
rect 2962 2760 3018 2816
rect 3622 2202 3678 2204
rect 3702 2202 3758 2204
rect 3782 2202 3838 2204
rect 3862 2202 3918 2204
rect 3622 2150 3648 2202
rect 3648 2150 3678 2202
rect 3702 2150 3712 2202
rect 3712 2150 3758 2202
rect 3782 2150 3828 2202
rect 3828 2150 3838 2202
rect 3862 2150 3892 2202
rect 3892 2150 3918 2202
rect 3622 2148 3678 2150
rect 3702 2148 3758 2150
rect 3782 2148 3838 2150
rect 3862 2148 3918 2150
rect 3514 1808 3570 1864
rect 4434 3440 4490 3496
rect 5170 15308 5172 15328
rect 5172 15308 5224 15328
rect 5224 15308 5226 15328
rect 5170 15272 5226 15308
rect 5078 9424 5134 9480
rect 4802 6196 4804 6216
rect 4804 6196 4856 6216
rect 4856 6196 4858 6216
rect 4802 6160 4858 6196
rect 4894 5752 4950 5808
rect 4710 3596 4766 3632
rect 4710 3576 4712 3596
rect 4712 3576 4764 3596
rect 4764 3576 4766 3596
rect 5354 28600 5410 28656
rect 5354 2896 5410 2952
rect 5262 2488 5318 2544
rect 4986 1400 5042 1456
rect 6289 37562 6345 37564
rect 6369 37562 6425 37564
rect 6449 37562 6505 37564
rect 6529 37562 6585 37564
rect 6289 37510 6315 37562
rect 6315 37510 6345 37562
rect 6369 37510 6379 37562
rect 6379 37510 6425 37562
rect 6449 37510 6495 37562
rect 6495 37510 6505 37562
rect 6529 37510 6559 37562
rect 6559 37510 6585 37562
rect 6289 37508 6345 37510
rect 6369 37508 6425 37510
rect 6449 37508 6505 37510
rect 6529 37508 6585 37510
rect 6289 36474 6345 36476
rect 6369 36474 6425 36476
rect 6449 36474 6505 36476
rect 6529 36474 6585 36476
rect 6289 36422 6315 36474
rect 6315 36422 6345 36474
rect 6369 36422 6379 36474
rect 6379 36422 6425 36474
rect 6449 36422 6495 36474
rect 6495 36422 6505 36474
rect 6529 36422 6559 36474
rect 6559 36422 6585 36474
rect 6289 36420 6345 36422
rect 6369 36420 6425 36422
rect 6449 36420 6505 36422
rect 6529 36420 6585 36422
rect 6289 35386 6345 35388
rect 6369 35386 6425 35388
rect 6449 35386 6505 35388
rect 6529 35386 6585 35388
rect 6289 35334 6315 35386
rect 6315 35334 6345 35386
rect 6369 35334 6379 35386
rect 6379 35334 6425 35386
rect 6449 35334 6495 35386
rect 6495 35334 6505 35386
rect 6529 35334 6559 35386
rect 6559 35334 6585 35386
rect 6289 35332 6345 35334
rect 6369 35332 6425 35334
rect 6449 35332 6505 35334
rect 6529 35332 6585 35334
rect 5998 35128 6054 35184
rect 5814 34992 5870 35048
rect 5722 20440 5778 20496
rect 5722 4664 5778 4720
rect 5446 2216 5502 2272
rect 6289 34298 6345 34300
rect 6369 34298 6425 34300
rect 6449 34298 6505 34300
rect 6529 34298 6585 34300
rect 6289 34246 6315 34298
rect 6315 34246 6345 34298
rect 6369 34246 6379 34298
rect 6379 34246 6425 34298
rect 6449 34246 6495 34298
rect 6495 34246 6505 34298
rect 6529 34246 6559 34298
rect 6559 34246 6585 34298
rect 6289 34244 6345 34246
rect 6369 34244 6425 34246
rect 6449 34244 6505 34246
rect 6529 34244 6585 34246
rect 6289 33210 6345 33212
rect 6369 33210 6425 33212
rect 6449 33210 6505 33212
rect 6529 33210 6585 33212
rect 6289 33158 6315 33210
rect 6315 33158 6345 33210
rect 6369 33158 6379 33210
rect 6379 33158 6425 33210
rect 6449 33158 6495 33210
rect 6495 33158 6505 33210
rect 6529 33158 6559 33210
rect 6559 33158 6585 33210
rect 6289 33156 6345 33158
rect 6369 33156 6425 33158
rect 6449 33156 6505 33158
rect 6529 33156 6585 33158
rect 6289 32122 6345 32124
rect 6369 32122 6425 32124
rect 6449 32122 6505 32124
rect 6529 32122 6585 32124
rect 6289 32070 6315 32122
rect 6315 32070 6345 32122
rect 6369 32070 6379 32122
rect 6379 32070 6425 32122
rect 6449 32070 6495 32122
rect 6495 32070 6505 32122
rect 6529 32070 6559 32122
rect 6559 32070 6585 32122
rect 6289 32068 6345 32070
rect 6369 32068 6425 32070
rect 6449 32068 6505 32070
rect 6529 32068 6585 32070
rect 6289 31034 6345 31036
rect 6369 31034 6425 31036
rect 6449 31034 6505 31036
rect 6529 31034 6585 31036
rect 6289 30982 6315 31034
rect 6315 30982 6345 31034
rect 6369 30982 6379 31034
rect 6379 30982 6425 31034
rect 6449 30982 6495 31034
rect 6495 30982 6505 31034
rect 6529 30982 6559 31034
rect 6559 30982 6585 31034
rect 6289 30980 6345 30982
rect 6369 30980 6425 30982
rect 6449 30980 6505 30982
rect 6529 30980 6585 30982
rect 6289 29946 6345 29948
rect 6369 29946 6425 29948
rect 6449 29946 6505 29948
rect 6529 29946 6585 29948
rect 6289 29894 6315 29946
rect 6315 29894 6345 29946
rect 6369 29894 6379 29946
rect 6379 29894 6425 29946
rect 6449 29894 6495 29946
rect 6495 29894 6505 29946
rect 6529 29894 6559 29946
rect 6559 29894 6585 29946
rect 6289 29892 6345 29894
rect 6369 29892 6425 29894
rect 6449 29892 6505 29894
rect 6529 29892 6585 29894
rect 6289 28858 6345 28860
rect 6369 28858 6425 28860
rect 6449 28858 6505 28860
rect 6529 28858 6585 28860
rect 6289 28806 6315 28858
rect 6315 28806 6345 28858
rect 6369 28806 6379 28858
rect 6379 28806 6425 28858
rect 6449 28806 6495 28858
rect 6495 28806 6505 28858
rect 6529 28806 6559 28858
rect 6559 28806 6585 28858
rect 6289 28804 6345 28806
rect 6369 28804 6425 28806
rect 6449 28804 6505 28806
rect 6529 28804 6585 28806
rect 6289 27770 6345 27772
rect 6369 27770 6425 27772
rect 6449 27770 6505 27772
rect 6529 27770 6585 27772
rect 6289 27718 6315 27770
rect 6315 27718 6345 27770
rect 6369 27718 6379 27770
rect 6379 27718 6425 27770
rect 6449 27718 6495 27770
rect 6495 27718 6505 27770
rect 6529 27718 6559 27770
rect 6559 27718 6585 27770
rect 6289 27716 6345 27718
rect 6369 27716 6425 27718
rect 6449 27716 6505 27718
rect 6529 27716 6585 27718
rect 6289 26682 6345 26684
rect 6369 26682 6425 26684
rect 6449 26682 6505 26684
rect 6529 26682 6585 26684
rect 6289 26630 6315 26682
rect 6315 26630 6345 26682
rect 6369 26630 6379 26682
rect 6379 26630 6425 26682
rect 6449 26630 6495 26682
rect 6495 26630 6505 26682
rect 6529 26630 6559 26682
rect 6559 26630 6585 26682
rect 6289 26628 6345 26630
rect 6369 26628 6425 26630
rect 6449 26628 6505 26630
rect 6529 26628 6585 26630
rect 6289 25594 6345 25596
rect 6369 25594 6425 25596
rect 6449 25594 6505 25596
rect 6529 25594 6585 25596
rect 6289 25542 6315 25594
rect 6315 25542 6345 25594
rect 6369 25542 6379 25594
rect 6379 25542 6425 25594
rect 6449 25542 6495 25594
rect 6495 25542 6505 25594
rect 6529 25542 6559 25594
rect 6559 25542 6585 25594
rect 6289 25540 6345 25542
rect 6369 25540 6425 25542
rect 6449 25540 6505 25542
rect 6529 25540 6585 25542
rect 6289 24506 6345 24508
rect 6369 24506 6425 24508
rect 6449 24506 6505 24508
rect 6529 24506 6585 24508
rect 6289 24454 6315 24506
rect 6315 24454 6345 24506
rect 6369 24454 6379 24506
rect 6379 24454 6425 24506
rect 6449 24454 6495 24506
rect 6495 24454 6505 24506
rect 6529 24454 6559 24506
rect 6559 24454 6585 24506
rect 6289 24452 6345 24454
rect 6369 24452 6425 24454
rect 6449 24452 6505 24454
rect 6529 24452 6585 24454
rect 6289 23418 6345 23420
rect 6369 23418 6425 23420
rect 6449 23418 6505 23420
rect 6529 23418 6585 23420
rect 6289 23366 6315 23418
rect 6315 23366 6345 23418
rect 6369 23366 6379 23418
rect 6379 23366 6425 23418
rect 6449 23366 6495 23418
rect 6495 23366 6505 23418
rect 6529 23366 6559 23418
rect 6559 23366 6585 23418
rect 6289 23364 6345 23366
rect 6369 23364 6425 23366
rect 6449 23364 6505 23366
rect 6529 23364 6585 23366
rect 5998 23024 6054 23080
rect 6289 22330 6345 22332
rect 6369 22330 6425 22332
rect 6449 22330 6505 22332
rect 6529 22330 6585 22332
rect 6289 22278 6315 22330
rect 6315 22278 6345 22330
rect 6369 22278 6379 22330
rect 6379 22278 6425 22330
rect 6449 22278 6495 22330
rect 6495 22278 6505 22330
rect 6529 22278 6559 22330
rect 6559 22278 6585 22330
rect 6289 22276 6345 22278
rect 6369 22276 6425 22278
rect 6449 22276 6505 22278
rect 6529 22276 6585 22278
rect 5998 22092 6054 22128
rect 5998 22072 6000 22092
rect 6000 22072 6052 22092
rect 6052 22072 6054 22092
rect 6274 21972 6276 21992
rect 6276 21972 6328 21992
rect 6328 21972 6330 21992
rect 6274 21936 6330 21972
rect 6090 21800 6146 21856
rect 6289 21242 6345 21244
rect 6369 21242 6425 21244
rect 6449 21242 6505 21244
rect 6529 21242 6585 21244
rect 6289 21190 6315 21242
rect 6315 21190 6345 21242
rect 6369 21190 6379 21242
rect 6379 21190 6425 21242
rect 6449 21190 6495 21242
rect 6495 21190 6505 21242
rect 6529 21190 6559 21242
rect 6559 21190 6585 21242
rect 6289 21188 6345 21190
rect 6369 21188 6425 21190
rect 6449 21188 6505 21190
rect 6529 21188 6585 21190
rect 5998 20984 6054 21040
rect 6289 20154 6345 20156
rect 6369 20154 6425 20156
rect 6449 20154 6505 20156
rect 6529 20154 6585 20156
rect 6289 20102 6315 20154
rect 6315 20102 6345 20154
rect 6369 20102 6379 20154
rect 6379 20102 6425 20154
rect 6449 20102 6495 20154
rect 6495 20102 6505 20154
rect 6529 20102 6559 20154
rect 6559 20102 6585 20154
rect 6289 20100 6345 20102
rect 6369 20100 6425 20102
rect 6449 20100 6505 20102
rect 6529 20100 6585 20102
rect 6289 19066 6345 19068
rect 6369 19066 6425 19068
rect 6449 19066 6505 19068
rect 6529 19066 6585 19068
rect 6289 19014 6315 19066
rect 6315 19014 6345 19066
rect 6369 19014 6379 19066
rect 6379 19014 6425 19066
rect 6449 19014 6495 19066
rect 6495 19014 6505 19066
rect 6529 19014 6559 19066
rect 6559 19014 6585 19066
rect 6289 19012 6345 19014
rect 6369 19012 6425 19014
rect 6449 19012 6505 19014
rect 6529 19012 6585 19014
rect 6289 17978 6345 17980
rect 6369 17978 6425 17980
rect 6449 17978 6505 17980
rect 6529 17978 6585 17980
rect 6289 17926 6315 17978
rect 6315 17926 6345 17978
rect 6369 17926 6379 17978
rect 6379 17926 6425 17978
rect 6449 17926 6495 17978
rect 6495 17926 6505 17978
rect 6529 17926 6559 17978
rect 6559 17926 6585 17978
rect 6289 17924 6345 17926
rect 6369 17924 6425 17926
rect 6449 17924 6505 17926
rect 6529 17924 6585 17926
rect 6289 16890 6345 16892
rect 6369 16890 6425 16892
rect 6449 16890 6505 16892
rect 6529 16890 6585 16892
rect 6289 16838 6315 16890
rect 6315 16838 6345 16890
rect 6369 16838 6379 16890
rect 6379 16838 6425 16890
rect 6449 16838 6495 16890
rect 6495 16838 6505 16890
rect 6529 16838 6559 16890
rect 6559 16838 6585 16890
rect 6289 16836 6345 16838
rect 6369 16836 6425 16838
rect 6449 16836 6505 16838
rect 6529 16836 6585 16838
rect 6289 15802 6345 15804
rect 6369 15802 6425 15804
rect 6449 15802 6505 15804
rect 6529 15802 6585 15804
rect 6289 15750 6315 15802
rect 6315 15750 6345 15802
rect 6369 15750 6379 15802
rect 6379 15750 6425 15802
rect 6449 15750 6495 15802
rect 6495 15750 6505 15802
rect 6529 15750 6559 15802
rect 6559 15750 6585 15802
rect 6289 15748 6345 15750
rect 6369 15748 6425 15750
rect 6449 15748 6505 15750
rect 6529 15748 6585 15750
rect 6289 14714 6345 14716
rect 6369 14714 6425 14716
rect 6449 14714 6505 14716
rect 6529 14714 6585 14716
rect 6289 14662 6315 14714
rect 6315 14662 6345 14714
rect 6369 14662 6379 14714
rect 6379 14662 6425 14714
rect 6449 14662 6495 14714
rect 6495 14662 6505 14714
rect 6529 14662 6559 14714
rect 6559 14662 6585 14714
rect 6289 14660 6345 14662
rect 6369 14660 6425 14662
rect 6449 14660 6505 14662
rect 6529 14660 6585 14662
rect 6289 13626 6345 13628
rect 6369 13626 6425 13628
rect 6449 13626 6505 13628
rect 6529 13626 6585 13628
rect 6289 13574 6315 13626
rect 6315 13574 6345 13626
rect 6369 13574 6379 13626
rect 6379 13574 6425 13626
rect 6449 13574 6495 13626
rect 6495 13574 6505 13626
rect 6529 13574 6559 13626
rect 6559 13574 6585 13626
rect 6289 13572 6345 13574
rect 6369 13572 6425 13574
rect 6449 13572 6505 13574
rect 6529 13572 6585 13574
rect 6289 12538 6345 12540
rect 6369 12538 6425 12540
rect 6449 12538 6505 12540
rect 6529 12538 6585 12540
rect 6289 12486 6315 12538
rect 6315 12486 6345 12538
rect 6369 12486 6379 12538
rect 6379 12486 6425 12538
rect 6449 12486 6495 12538
rect 6495 12486 6505 12538
rect 6529 12486 6559 12538
rect 6559 12486 6585 12538
rect 6289 12484 6345 12486
rect 6369 12484 6425 12486
rect 6449 12484 6505 12486
rect 6529 12484 6585 12486
rect 6289 11450 6345 11452
rect 6369 11450 6425 11452
rect 6449 11450 6505 11452
rect 6529 11450 6585 11452
rect 6289 11398 6315 11450
rect 6315 11398 6345 11450
rect 6369 11398 6379 11450
rect 6379 11398 6425 11450
rect 6449 11398 6495 11450
rect 6495 11398 6505 11450
rect 6529 11398 6559 11450
rect 6559 11398 6585 11450
rect 6289 11396 6345 11398
rect 6369 11396 6425 11398
rect 6449 11396 6505 11398
rect 6529 11396 6585 11398
rect 6289 10362 6345 10364
rect 6369 10362 6425 10364
rect 6449 10362 6505 10364
rect 6529 10362 6585 10364
rect 6289 10310 6315 10362
rect 6315 10310 6345 10362
rect 6369 10310 6379 10362
rect 6379 10310 6425 10362
rect 6449 10310 6495 10362
rect 6495 10310 6505 10362
rect 6529 10310 6559 10362
rect 6559 10310 6585 10362
rect 6289 10308 6345 10310
rect 6369 10308 6425 10310
rect 6449 10308 6505 10310
rect 6529 10308 6585 10310
rect 6289 9274 6345 9276
rect 6369 9274 6425 9276
rect 6449 9274 6505 9276
rect 6529 9274 6585 9276
rect 6289 9222 6315 9274
rect 6315 9222 6345 9274
rect 6369 9222 6379 9274
rect 6379 9222 6425 9274
rect 6449 9222 6495 9274
rect 6495 9222 6505 9274
rect 6529 9222 6559 9274
rect 6559 9222 6585 9274
rect 6289 9220 6345 9222
rect 6369 9220 6425 9222
rect 6449 9220 6505 9222
rect 6529 9220 6585 9222
rect 6289 8186 6345 8188
rect 6369 8186 6425 8188
rect 6449 8186 6505 8188
rect 6529 8186 6585 8188
rect 6289 8134 6315 8186
rect 6315 8134 6345 8186
rect 6369 8134 6379 8186
rect 6379 8134 6425 8186
rect 6449 8134 6495 8186
rect 6495 8134 6505 8186
rect 6529 8134 6559 8186
rect 6559 8134 6585 8186
rect 6289 8132 6345 8134
rect 6369 8132 6425 8134
rect 6449 8132 6505 8134
rect 6529 8132 6585 8134
rect 6826 33088 6882 33144
rect 6826 23468 6828 23488
rect 6828 23468 6880 23488
rect 6880 23468 6882 23488
rect 6826 23432 6882 23468
rect 7654 28600 7710 28656
rect 8022 24656 8078 24712
rect 7470 22480 7526 22536
rect 7378 20204 7380 20224
rect 7380 20204 7432 20224
rect 7432 20204 7434 20224
rect 7378 20168 7434 20204
rect 7194 16088 7250 16144
rect 6918 15544 6974 15600
rect 7194 15272 7250 15328
rect 6289 7098 6345 7100
rect 6369 7098 6425 7100
rect 6449 7098 6505 7100
rect 6529 7098 6585 7100
rect 6289 7046 6315 7098
rect 6315 7046 6345 7098
rect 6369 7046 6379 7098
rect 6379 7046 6425 7098
rect 6449 7046 6495 7098
rect 6495 7046 6505 7098
rect 6529 7046 6559 7098
rect 6559 7046 6585 7098
rect 6289 7044 6345 7046
rect 6369 7044 6425 7046
rect 6449 7044 6505 7046
rect 6529 7044 6585 7046
rect 6182 6840 6238 6896
rect 6090 3984 6146 4040
rect 6090 3032 6146 3088
rect 5814 2760 5870 2816
rect 6289 6010 6345 6012
rect 6369 6010 6425 6012
rect 6449 6010 6505 6012
rect 6529 6010 6585 6012
rect 6289 5958 6315 6010
rect 6315 5958 6345 6010
rect 6369 5958 6379 6010
rect 6379 5958 6425 6010
rect 6449 5958 6495 6010
rect 6495 5958 6505 6010
rect 6529 5958 6559 6010
rect 6559 5958 6585 6010
rect 6289 5956 6345 5958
rect 6369 5956 6425 5958
rect 6449 5956 6505 5958
rect 6529 5956 6585 5958
rect 6289 4922 6345 4924
rect 6369 4922 6425 4924
rect 6449 4922 6505 4924
rect 6529 4922 6585 4924
rect 6289 4870 6315 4922
rect 6315 4870 6345 4922
rect 6369 4870 6379 4922
rect 6379 4870 6425 4922
rect 6449 4870 6495 4922
rect 6495 4870 6505 4922
rect 6529 4870 6559 4922
rect 6559 4870 6585 4922
rect 6289 4868 6345 4870
rect 6369 4868 6425 4870
rect 6449 4868 6505 4870
rect 6529 4868 6585 4870
rect 6289 3834 6345 3836
rect 6369 3834 6425 3836
rect 6449 3834 6505 3836
rect 6529 3834 6585 3836
rect 6289 3782 6315 3834
rect 6315 3782 6345 3834
rect 6369 3782 6379 3834
rect 6379 3782 6425 3834
rect 6449 3782 6495 3834
rect 6495 3782 6505 3834
rect 6529 3782 6559 3834
rect 6559 3782 6585 3834
rect 6289 3780 6345 3782
rect 6369 3780 6425 3782
rect 6449 3780 6505 3782
rect 6529 3780 6585 3782
rect 6289 2746 6345 2748
rect 6369 2746 6425 2748
rect 6449 2746 6505 2748
rect 6529 2746 6585 2748
rect 6289 2694 6315 2746
rect 6315 2694 6345 2746
rect 6369 2694 6379 2746
rect 6379 2694 6425 2746
rect 6449 2694 6495 2746
rect 6495 2694 6505 2746
rect 6529 2694 6559 2746
rect 6559 2694 6585 2746
rect 6289 2692 6345 2694
rect 6369 2692 6425 2694
rect 6449 2692 6505 2694
rect 6529 2692 6585 2694
rect 7654 20460 7710 20496
rect 7654 20440 7656 20460
rect 7656 20440 7708 20460
rect 7708 20440 7710 20460
rect 7562 14864 7618 14920
rect 8022 14612 8078 14648
rect 8022 14592 8024 14612
rect 8024 14592 8076 14612
rect 8076 14592 8078 14612
rect 7930 12688 7986 12744
rect 8390 15000 8446 15056
rect 8298 14592 8354 14648
rect 7838 9560 7894 9616
rect 7010 7248 7066 7304
rect 6826 6704 6882 6760
rect 6918 3712 6974 3768
rect 6734 2624 6790 2680
rect 7746 3576 7802 3632
rect 7378 2760 7434 2816
rect 7102 2488 7158 2544
rect 7562 1944 7618 2000
rect 8114 2352 8170 2408
rect 8956 37018 9012 37020
rect 9036 37018 9092 37020
rect 9116 37018 9172 37020
rect 9196 37018 9252 37020
rect 8956 36966 8982 37018
rect 8982 36966 9012 37018
rect 9036 36966 9046 37018
rect 9046 36966 9092 37018
rect 9116 36966 9162 37018
rect 9162 36966 9172 37018
rect 9196 36966 9226 37018
rect 9226 36966 9252 37018
rect 8956 36964 9012 36966
rect 9036 36964 9092 36966
rect 9116 36964 9172 36966
rect 9196 36964 9252 36966
rect 8956 35930 9012 35932
rect 9036 35930 9092 35932
rect 9116 35930 9172 35932
rect 9196 35930 9252 35932
rect 8956 35878 8982 35930
rect 8982 35878 9012 35930
rect 9036 35878 9046 35930
rect 9046 35878 9092 35930
rect 9116 35878 9162 35930
rect 9162 35878 9172 35930
rect 9196 35878 9226 35930
rect 9226 35878 9252 35930
rect 8956 35876 9012 35878
rect 9036 35876 9092 35878
rect 9116 35876 9172 35878
rect 9196 35876 9252 35878
rect 9402 35672 9458 35728
rect 8666 35536 8722 35592
rect 8574 16632 8630 16688
rect 8574 3304 8630 3360
rect 8956 34842 9012 34844
rect 9036 34842 9092 34844
rect 9116 34842 9172 34844
rect 9196 34842 9252 34844
rect 8956 34790 8982 34842
rect 8982 34790 9012 34842
rect 9036 34790 9046 34842
rect 9046 34790 9092 34842
rect 9116 34790 9162 34842
rect 9162 34790 9172 34842
rect 9196 34790 9226 34842
rect 9226 34790 9252 34842
rect 8956 34788 9012 34790
rect 9036 34788 9092 34790
rect 9116 34788 9172 34790
rect 9196 34788 9252 34790
rect 8956 33754 9012 33756
rect 9036 33754 9092 33756
rect 9116 33754 9172 33756
rect 9196 33754 9252 33756
rect 8956 33702 8982 33754
rect 8982 33702 9012 33754
rect 9036 33702 9046 33754
rect 9046 33702 9092 33754
rect 9116 33702 9162 33754
rect 9162 33702 9172 33754
rect 9196 33702 9226 33754
rect 9226 33702 9252 33754
rect 8956 33700 9012 33702
rect 9036 33700 9092 33702
rect 9116 33700 9172 33702
rect 9196 33700 9252 33702
rect 8758 33088 8814 33144
rect 8956 32666 9012 32668
rect 9036 32666 9092 32668
rect 9116 32666 9172 32668
rect 9196 32666 9252 32668
rect 8956 32614 8982 32666
rect 8982 32614 9012 32666
rect 9036 32614 9046 32666
rect 9046 32614 9092 32666
rect 9116 32614 9162 32666
rect 9162 32614 9172 32666
rect 9196 32614 9226 32666
rect 9226 32614 9252 32666
rect 8956 32612 9012 32614
rect 9036 32612 9092 32614
rect 9116 32612 9172 32614
rect 9196 32612 9252 32614
rect 8956 31578 9012 31580
rect 9036 31578 9092 31580
rect 9116 31578 9172 31580
rect 9196 31578 9252 31580
rect 8956 31526 8982 31578
rect 8982 31526 9012 31578
rect 9036 31526 9046 31578
rect 9046 31526 9092 31578
rect 9116 31526 9162 31578
rect 9162 31526 9172 31578
rect 9196 31526 9226 31578
rect 9226 31526 9252 31578
rect 8956 31524 9012 31526
rect 9036 31524 9092 31526
rect 9116 31524 9172 31526
rect 9196 31524 9252 31526
rect 8956 30490 9012 30492
rect 9036 30490 9092 30492
rect 9116 30490 9172 30492
rect 9196 30490 9252 30492
rect 8956 30438 8982 30490
rect 8982 30438 9012 30490
rect 9036 30438 9046 30490
rect 9046 30438 9092 30490
rect 9116 30438 9162 30490
rect 9162 30438 9172 30490
rect 9196 30438 9226 30490
rect 9226 30438 9252 30490
rect 8956 30436 9012 30438
rect 9036 30436 9092 30438
rect 9116 30436 9172 30438
rect 9196 30436 9252 30438
rect 8956 29402 9012 29404
rect 9036 29402 9092 29404
rect 9116 29402 9172 29404
rect 9196 29402 9252 29404
rect 8956 29350 8982 29402
rect 8982 29350 9012 29402
rect 9036 29350 9046 29402
rect 9046 29350 9092 29402
rect 9116 29350 9162 29402
rect 9162 29350 9172 29402
rect 9196 29350 9226 29402
rect 9226 29350 9252 29402
rect 8956 29348 9012 29350
rect 9036 29348 9092 29350
rect 9116 29348 9172 29350
rect 9196 29348 9252 29350
rect 8956 28314 9012 28316
rect 9036 28314 9092 28316
rect 9116 28314 9172 28316
rect 9196 28314 9252 28316
rect 8956 28262 8982 28314
rect 8982 28262 9012 28314
rect 9036 28262 9046 28314
rect 9046 28262 9092 28314
rect 9116 28262 9162 28314
rect 9162 28262 9172 28314
rect 9196 28262 9226 28314
rect 9226 28262 9252 28314
rect 8956 28260 9012 28262
rect 9036 28260 9092 28262
rect 9116 28260 9172 28262
rect 9196 28260 9252 28262
rect 8956 27226 9012 27228
rect 9036 27226 9092 27228
rect 9116 27226 9172 27228
rect 9196 27226 9252 27228
rect 8956 27174 8982 27226
rect 8982 27174 9012 27226
rect 9036 27174 9046 27226
rect 9046 27174 9092 27226
rect 9116 27174 9162 27226
rect 9162 27174 9172 27226
rect 9196 27174 9226 27226
rect 9226 27174 9252 27226
rect 8956 27172 9012 27174
rect 9036 27172 9092 27174
rect 9116 27172 9172 27174
rect 9196 27172 9252 27174
rect 8956 26138 9012 26140
rect 9036 26138 9092 26140
rect 9116 26138 9172 26140
rect 9196 26138 9252 26140
rect 8956 26086 8982 26138
rect 8982 26086 9012 26138
rect 9036 26086 9046 26138
rect 9046 26086 9092 26138
rect 9116 26086 9162 26138
rect 9162 26086 9172 26138
rect 9196 26086 9226 26138
rect 9226 26086 9252 26138
rect 8956 26084 9012 26086
rect 9036 26084 9092 26086
rect 9116 26084 9172 26086
rect 9196 26084 9252 26086
rect 8956 25050 9012 25052
rect 9036 25050 9092 25052
rect 9116 25050 9172 25052
rect 9196 25050 9252 25052
rect 8956 24998 8982 25050
rect 8982 24998 9012 25050
rect 9036 24998 9046 25050
rect 9046 24998 9092 25050
rect 9116 24998 9162 25050
rect 9162 24998 9172 25050
rect 9196 24998 9226 25050
rect 9226 24998 9252 25050
rect 8956 24996 9012 24998
rect 9036 24996 9092 24998
rect 9116 24996 9172 24998
rect 9196 24996 9252 24998
rect 8956 23962 9012 23964
rect 9036 23962 9092 23964
rect 9116 23962 9172 23964
rect 9196 23962 9252 23964
rect 8956 23910 8982 23962
rect 8982 23910 9012 23962
rect 9036 23910 9046 23962
rect 9046 23910 9092 23962
rect 9116 23910 9162 23962
rect 9162 23910 9172 23962
rect 9196 23910 9226 23962
rect 9226 23910 9252 23962
rect 8956 23908 9012 23910
rect 9036 23908 9092 23910
rect 9116 23908 9172 23910
rect 9196 23908 9252 23910
rect 8758 23432 8814 23488
rect 8956 22874 9012 22876
rect 9036 22874 9092 22876
rect 9116 22874 9172 22876
rect 9196 22874 9252 22876
rect 8956 22822 8982 22874
rect 8982 22822 9012 22874
rect 9036 22822 9046 22874
rect 9046 22822 9092 22874
rect 9116 22822 9162 22874
rect 9162 22822 9172 22874
rect 9196 22822 9226 22874
rect 9226 22822 9252 22874
rect 8956 22820 9012 22822
rect 9036 22820 9092 22822
rect 9116 22820 9172 22822
rect 9196 22820 9252 22822
rect 8956 21786 9012 21788
rect 9036 21786 9092 21788
rect 9116 21786 9172 21788
rect 9196 21786 9252 21788
rect 8956 21734 8982 21786
rect 8982 21734 9012 21786
rect 9036 21734 9046 21786
rect 9046 21734 9092 21786
rect 9116 21734 9162 21786
rect 9162 21734 9172 21786
rect 9196 21734 9226 21786
rect 9226 21734 9252 21786
rect 8956 21732 9012 21734
rect 9036 21732 9092 21734
rect 9116 21732 9172 21734
rect 9196 21732 9252 21734
rect 8956 20698 9012 20700
rect 9036 20698 9092 20700
rect 9116 20698 9172 20700
rect 9196 20698 9252 20700
rect 8956 20646 8982 20698
rect 8982 20646 9012 20698
rect 9036 20646 9046 20698
rect 9046 20646 9092 20698
rect 9116 20646 9162 20698
rect 9162 20646 9172 20698
rect 9196 20646 9226 20698
rect 9226 20646 9252 20698
rect 8956 20644 9012 20646
rect 9036 20644 9092 20646
rect 9116 20644 9172 20646
rect 9196 20644 9252 20646
rect 8956 19610 9012 19612
rect 9036 19610 9092 19612
rect 9116 19610 9172 19612
rect 9196 19610 9252 19612
rect 8956 19558 8982 19610
rect 8982 19558 9012 19610
rect 9036 19558 9046 19610
rect 9046 19558 9092 19610
rect 9116 19558 9162 19610
rect 9162 19558 9172 19610
rect 9196 19558 9226 19610
rect 9226 19558 9252 19610
rect 8956 19556 9012 19558
rect 9036 19556 9092 19558
rect 9116 19556 9172 19558
rect 9196 19556 9252 19558
rect 8956 18522 9012 18524
rect 9036 18522 9092 18524
rect 9116 18522 9172 18524
rect 9196 18522 9252 18524
rect 8956 18470 8982 18522
rect 8982 18470 9012 18522
rect 9036 18470 9046 18522
rect 9046 18470 9092 18522
rect 9116 18470 9162 18522
rect 9162 18470 9172 18522
rect 9196 18470 9226 18522
rect 9226 18470 9252 18522
rect 8956 18468 9012 18470
rect 9036 18468 9092 18470
rect 9116 18468 9172 18470
rect 9196 18468 9252 18470
rect 8956 17434 9012 17436
rect 9036 17434 9092 17436
rect 9116 17434 9172 17436
rect 9196 17434 9252 17436
rect 8956 17382 8982 17434
rect 8982 17382 9012 17434
rect 9036 17382 9046 17434
rect 9046 17382 9092 17434
rect 9116 17382 9162 17434
rect 9162 17382 9172 17434
rect 9196 17382 9226 17434
rect 9226 17382 9252 17434
rect 8956 17380 9012 17382
rect 9036 17380 9092 17382
rect 9116 17380 9172 17382
rect 9196 17380 9252 17382
rect 8956 16346 9012 16348
rect 9036 16346 9092 16348
rect 9116 16346 9172 16348
rect 9196 16346 9252 16348
rect 8956 16294 8982 16346
rect 8982 16294 9012 16346
rect 9036 16294 9046 16346
rect 9046 16294 9092 16346
rect 9116 16294 9162 16346
rect 9162 16294 9172 16346
rect 9196 16294 9226 16346
rect 9226 16294 9252 16346
rect 8956 16292 9012 16294
rect 9036 16292 9092 16294
rect 9116 16292 9172 16294
rect 9196 16292 9252 16294
rect 8956 15258 9012 15260
rect 9036 15258 9092 15260
rect 9116 15258 9172 15260
rect 9196 15258 9252 15260
rect 8956 15206 8982 15258
rect 8982 15206 9012 15258
rect 9036 15206 9046 15258
rect 9046 15206 9092 15258
rect 9116 15206 9162 15258
rect 9162 15206 9172 15258
rect 9196 15206 9226 15258
rect 9226 15206 9252 15258
rect 8956 15204 9012 15206
rect 9036 15204 9092 15206
rect 9116 15204 9172 15206
rect 9196 15204 9252 15206
rect 9770 30232 9826 30288
rect 9862 25336 9918 25392
rect 9402 21800 9458 21856
rect 10966 35128 11022 35184
rect 11334 34992 11390 35048
rect 11622 37562 11678 37564
rect 11702 37562 11758 37564
rect 11782 37562 11838 37564
rect 11862 37562 11918 37564
rect 11622 37510 11648 37562
rect 11648 37510 11678 37562
rect 11702 37510 11712 37562
rect 11712 37510 11758 37562
rect 11782 37510 11828 37562
rect 11828 37510 11838 37562
rect 11862 37510 11892 37562
rect 11892 37510 11918 37562
rect 11622 37508 11678 37510
rect 11702 37508 11758 37510
rect 11782 37508 11838 37510
rect 11862 37508 11918 37510
rect 11622 36474 11678 36476
rect 11702 36474 11758 36476
rect 11782 36474 11838 36476
rect 11862 36474 11918 36476
rect 11622 36422 11648 36474
rect 11648 36422 11678 36474
rect 11702 36422 11712 36474
rect 11712 36422 11758 36474
rect 11782 36422 11828 36474
rect 11828 36422 11838 36474
rect 11862 36422 11892 36474
rect 11892 36422 11918 36474
rect 11622 36420 11678 36422
rect 11702 36420 11758 36422
rect 11782 36420 11838 36422
rect 11862 36420 11918 36422
rect 11622 35386 11678 35388
rect 11702 35386 11758 35388
rect 11782 35386 11838 35388
rect 11862 35386 11918 35388
rect 11622 35334 11648 35386
rect 11648 35334 11678 35386
rect 11702 35334 11712 35386
rect 11712 35334 11758 35386
rect 11782 35334 11828 35386
rect 11828 35334 11838 35386
rect 11862 35334 11892 35386
rect 11892 35334 11918 35386
rect 11622 35332 11678 35334
rect 11702 35332 11758 35334
rect 11782 35332 11838 35334
rect 11862 35332 11918 35334
rect 11518 34584 11574 34640
rect 11622 34298 11678 34300
rect 11702 34298 11758 34300
rect 11782 34298 11838 34300
rect 11862 34298 11918 34300
rect 11622 34246 11648 34298
rect 11648 34246 11678 34298
rect 11702 34246 11712 34298
rect 11712 34246 11758 34298
rect 11782 34246 11828 34298
rect 11828 34246 11838 34298
rect 11862 34246 11892 34298
rect 11892 34246 11918 34298
rect 11622 34244 11678 34246
rect 11702 34244 11758 34246
rect 11782 34244 11838 34246
rect 11862 34244 11918 34246
rect 11622 33210 11678 33212
rect 11702 33210 11758 33212
rect 11782 33210 11838 33212
rect 11862 33210 11918 33212
rect 11622 33158 11648 33210
rect 11648 33158 11678 33210
rect 11702 33158 11712 33210
rect 11712 33158 11758 33210
rect 11782 33158 11828 33210
rect 11828 33158 11838 33210
rect 11862 33158 11892 33210
rect 11892 33158 11918 33210
rect 11622 33156 11678 33158
rect 11702 33156 11758 33158
rect 11782 33156 11838 33158
rect 11862 33156 11918 33158
rect 11622 32122 11678 32124
rect 11702 32122 11758 32124
rect 11782 32122 11838 32124
rect 11862 32122 11918 32124
rect 11622 32070 11648 32122
rect 11648 32070 11678 32122
rect 11702 32070 11712 32122
rect 11712 32070 11758 32122
rect 11782 32070 11828 32122
rect 11828 32070 11838 32122
rect 11862 32070 11892 32122
rect 11892 32070 11918 32122
rect 11622 32068 11678 32070
rect 11702 32068 11758 32070
rect 11782 32068 11838 32070
rect 11862 32068 11918 32070
rect 11622 31034 11678 31036
rect 11702 31034 11758 31036
rect 11782 31034 11838 31036
rect 11862 31034 11918 31036
rect 11622 30982 11648 31034
rect 11648 30982 11678 31034
rect 11702 30982 11712 31034
rect 11712 30982 11758 31034
rect 11782 30982 11828 31034
rect 11828 30982 11838 31034
rect 11862 30982 11892 31034
rect 11892 30982 11918 31034
rect 11622 30980 11678 30982
rect 11702 30980 11758 30982
rect 11782 30980 11838 30982
rect 11862 30980 11918 30982
rect 11622 29946 11678 29948
rect 11702 29946 11758 29948
rect 11782 29946 11838 29948
rect 11862 29946 11918 29948
rect 11622 29894 11648 29946
rect 11648 29894 11678 29946
rect 11702 29894 11712 29946
rect 11712 29894 11758 29946
rect 11782 29894 11828 29946
rect 11828 29894 11838 29946
rect 11862 29894 11892 29946
rect 11892 29894 11918 29946
rect 11622 29892 11678 29894
rect 11702 29892 11758 29894
rect 11782 29892 11838 29894
rect 11862 29892 11918 29894
rect 9954 23024 10010 23080
rect 9862 22480 9918 22536
rect 9770 21800 9826 21856
rect 9770 20984 9826 21040
rect 9310 14456 9366 14512
rect 8956 14170 9012 14172
rect 9036 14170 9092 14172
rect 9116 14170 9172 14172
rect 9196 14170 9252 14172
rect 8956 14118 8982 14170
rect 8982 14118 9012 14170
rect 9036 14118 9046 14170
rect 9046 14118 9092 14170
rect 9116 14118 9162 14170
rect 9162 14118 9172 14170
rect 9196 14118 9226 14170
rect 9226 14118 9252 14170
rect 8956 14116 9012 14118
rect 9036 14116 9092 14118
rect 9116 14116 9172 14118
rect 9196 14116 9252 14118
rect 8956 13082 9012 13084
rect 9036 13082 9092 13084
rect 9116 13082 9172 13084
rect 9196 13082 9252 13084
rect 8956 13030 8982 13082
rect 8982 13030 9012 13082
rect 9036 13030 9046 13082
rect 9046 13030 9092 13082
rect 9116 13030 9162 13082
rect 9162 13030 9172 13082
rect 9196 13030 9226 13082
rect 9226 13030 9252 13082
rect 8956 13028 9012 13030
rect 9036 13028 9092 13030
rect 9116 13028 9172 13030
rect 9196 13028 9252 13030
rect 8956 11994 9012 11996
rect 9036 11994 9092 11996
rect 9116 11994 9172 11996
rect 9196 11994 9252 11996
rect 8956 11942 8982 11994
rect 8982 11942 9012 11994
rect 9036 11942 9046 11994
rect 9046 11942 9092 11994
rect 9116 11942 9162 11994
rect 9162 11942 9172 11994
rect 9196 11942 9226 11994
rect 9226 11942 9252 11994
rect 8956 11940 9012 11942
rect 9036 11940 9092 11942
rect 9116 11940 9172 11942
rect 9196 11940 9252 11942
rect 8956 10906 9012 10908
rect 9036 10906 9092 10908
rect 9116 10906 9172 10908
rect 9196 10906 9252 10908
rect 8956 10854 8982 10906
rect 8982 10854 9012 10906
rect 9036 10854 9046 10906
rect 9046 10854 9092 10906
rect 9116 10854 9162 10906
rect 9162 10854 9172 10906
rect 9196 10854 9226 10906
rect 9226 10854 9252 10906
rect 8956 10852 9012 10854
rect 9036 10852 9092 10854
rect 9116 10852 9172 10854
rect 9196 10852 9252 10854
rect 8956 9818 9012 9820
rect 9036 9818 9092 9820
rect 9116 9818 9172 9820
rect 9196 9818 9252 9820
rect 8956 9766 8982 9818
rect 8982 9766 9012 9818
rect 9036 9766 9046 9818
rect 9046 9766 9092 9818
rect 9116 9766 9162 9818
rect 9162 9766 9172 9818
rect 9196 9766 9226 9818
rect 9226 9766 9252 9818
rect 8956 9764 9012 9766
rect 9036 9764 9092 9766
rect 9116 9764 9172 9766
rect 9196 9764 9252 9766
rect 8956 8730 9012 8732
rect 9036 8730 9092 8732
rect 9116 8730 9172 8732
rect 9196 8730 9252 8732
rect 8956 8678 8982 8730
rect 8982 8678 9012 8730
rect 9036 8678 9046 8730
rect 9046 8678 9092 8730
rect 9116 8678 9162 8730
rect 9162 8678 9172 8730
rect 9196 8678 9226 8730
rect 9226 8678 9252 8730
rect 8956 8676 9012 8678
rect 9036 8676 9092 8678
rect 9116 8676 9172 8678
rect 9196 8676 9252 8678
rect 8956 7642 9012 7644
rect 9036 7642 9092 7644
rect 9116 7642 9172 7644
rect 9196 7642 9252 7644
rect 8956 7590 8982 7642
rect 8982 7590 9012 7642
rect 9036 7590 9046 7642
rect 9046 7590 9092 7642
rect 9116 7590 9162 7642
rect 9162 7590 9172 7642
rect 9196 7590 9226 7642
rect 9226 7590 9252 7642
rect 8956 7588 9012 7590
rect 9036 7588 9092 7590
rect 9116 7588 9172 7590
rect 9196 7588 9252 7590
rect 8850 6840 8906 6896
rect 8956 6554 9012 6556
rect 9036 6554 9092 6556
rect 9116 6554 9172 6556
rect 9196 6554 9252 6556
rect 8956 6502 8982 6554
rect 8982 6502 9012 6554
rect 9036 6502 9046 6554
rect 9046 6502 9092 6554
rect 9116 6502 9162 6554
rect 9162 6502 9172 6554
rect 9196 6502 9226 6554
rect 9226 6502 9252 6554
rect 8956 6500 9012 6502
rect 9036 6500 9092 6502
rect 9116 6500 9172 6502
rect 9196 6500 9252 6502
rect 8850 6332 8852 6352
rect 8852 6332 8904 6352
rect 8904 6332 8906 6352
rect 8850 6296 8906 6332
rect 8956 5466 9012 5468
rect 9036 5466 9092 5468
rect 9116 5466 9172 5468
rect 9196 5466 9252 5468
rect 8956 5414 8982 5466
rect 8982 5414 9012 5466
rect 9036 5414 9046 5466
rect 9046 5414 9092 5466
rect 9116 5414 9162 5466
rect 9162 5414 9172 5466
rect 9196 5414 9226 5466
rect 9226 5414 9252 5466
rect 8956 5412 9012 5414
rect 9036 5412 9092 5414
rect 9116 5412 9172 5414
rect 9196 5412 9252 5414
rect 8956 4378 9012 4380
rect 9036 4378 9092 4380
rect 9116 4378 9172 4380
rect 9196 4378 9252 4380
rect 8956 4326 8982 4378
rect 8982 4326 9012 4378
rect 9036 4326 9046 4378
rect 9046 4326 9092 4378
rect 9116 4326 9162 4378
rect 9162 4326 9172 4378
rect 9196 4326 9226 4378
rect 9226 4326 9252 4378
rect 8956 4324 9012 4326
rect 9036 4324 9092 4326
rect 9116 4324 9172 4326
rect 9196 4324 9252 4326
rect 8956 3290 9012 3292
rect 9036 3290 9092 3292
rect 9116 3290 9172 3292
rect 9196 3290 9252 3292
rect 8956 3238 8982 3290
rect 8982 3238 9012 3290
rect 9036 3238 9046 3290
rect 9046 3238 9092 3290
rect 9116 3238 9162 3290
rect 9162 3238 9172 3290
rect 9196 3238 9226 3290
rect 9226 3238 9252 3290
rect 8956 3236 9012 3238
rect 9036 3236 9092 3238
rect 9116 3236 9172 3238
rect 9196 3236 9252 3238
rect 8850 2896 8906 2952
rect 8758 2252 8760 2272
rect 8760 2252 8812 2272
rect 8812 2252 8814 2272
rect 8758 2216 8814 2252
rect 8956 2202 9012 2204
rect 9036 2202 9092 2204
rect 9116 2202 9172 2204
rect 9196 2202 9252 2204
rect 8956 2150 8982 2202
rect 8982 2150 9012 2202
rect 9036 2150 9046 2202
rect 9046 2150 9092 2202
rect 9116 2150 9162 2202
rect 9162 2150 9172 2202
rect 9196 2150 9226 2202
rect 9226 2150 9252 2202
rect 8956 2148 9012 2150
rect 9036 2148 9092 2150
rect 9116 2148 9172 2150
rect 9196 2148 9252 2150
rect 9678 14592 9734 14648
rect 9402 3304 9458 3360
rect 9402 2252 9404 2272
rect 9404 2252 9456 2272
rect 9456 2252 9458 2272
rect 9402 2216 9458 2252
rect 9402 1808 9458 1864
rect 10046 20440 10102 20496
rect 11622 28858 11678 28860
rect 11702 28858 11758 28860
rect 11782 28858 11838 28860
rect 11862 28858 11918 28860
rect 11622 28806 11648 28858
rect 11648 28806 11678 28858
rect 11702 28806 11712 28858
rect 11712 28806 11758 28858
rect 11782 28806 11828 28858
rect 11828 28806 11838 28858
rect 11862 28806 11892 28858
rect 11892 28806 11918 28858
rect 11622 28804 11678 28806
rect 11702 28804 11758 28806
rect 11782 28804 11838 28806
rect 11862 28804 11918 28806
rect 11622 27770 11678 27772
rect 11702 27770 11758 27772
rect 11782 27770 11838 27772
rect 11862 27770 11918 27772
rect 11622 27718 11648 27770
rect 11648 27718 11678 27770
rect 11702 27718 11712 27770
rect 11712 27718 11758 27770
rect 11782 27718 11828 27770
rect 11828 27718 11838 27770
rect 11862 27718 11892 27770
rect 11892 27718 11918 27770
rect 11622 27716 11678 27718
rect 11702 27716 11758 27718
rect 11782 27716 11838 27718
rect 11862 27716 11918 27718
rect 11622 26682 11678 26684
rect 11702 26682 11758 26684
rect 11782 26682 11838 26684
rect 11862 26682 11918 26684
rect 11622 26630 11648 26682
rect 11648 26630 11678 26682
rect 11702 26630 11712 26682
rect 11712 26630 11758 26682
rect 11782 26630 11828 26682
rect 11828 26630 11838 26682
rect 11862 26630 11892 26682
rect 11892 26630 11918 26682
rect 11622 26628 11678 26630
rect 11702 26628 11758 26630
rect 11782 26628 11838 26630
rect 11862 26628 11918 26630
rect 11622 25594 11678 25596
rect 11702 25594 11758 25596
rect 11782 25594 11838 25596
rect 11862 25594 11918 25596
rect 11622 25542 11648 25594
rect 11648 25542 11678 25594
rect 11702 25542 11712 25594
rect 11712 25542 11758 25594
rect 11782 25542 11828 25594
rect 11828 25542 11838 25594
rect 11862 25542 11892 25594
rect 11892 25542 11918 25594
rect 11622 25540 11678 25542
rect 11702 25540 11758 25542
rect 11782 25540 11838 25542
rect 11862 25540 11918 25542
rect 11622 24506 11678 24508
rect 11702 24506 11758 24508
rect 11782 24506 11838 24508
rect 11862 24506 11918 24508
rect 11622 24454 11648 24506
rect 11648 24454 11678 24506
rect 11702 24454 11712 24506
rect 11712 24454 11758 24506
rect 11782 24454 11828 24506
rect 11828 24454 11838 24506
rect 11862 24454 11892 24506
rect 11892 24454 11918 24506
rect 11622 24452 11678 24454
rect 11702 24452 11758 24454
rect 11782 24452 11838 24454
rect 11862 24452 11918 24454
rect 11622 23418 11678 23420
rect 11702 23418 11758 23420
rect 11782 23418 11838 23420
rect 11862 23418 11918 23420
rect 11622 23366 11648 23418
rect 11648 23366 11678 23418
rect 11702 23366 11712 23418
rect 11712 23366 11758 23418
rect 11782 23366 11828 23418
rect 11828 23366 11838 23418
rect 11862 23366 11892 23418
rect 11892 23366 11918 23418
rect 11622 23364 11678 23366
rect 11702 23364 11758 23366
rect 11782 23364 11838 23366
rect 11862 23364 11918 23366
rect 12346 34584 12402 34640
rect 12254 25200 12310 25256
rect 12070 24656 12126 24712
rect 12070 23468 12072 23488
rect 12072 23468 12124 23488
rect 12124 23468 12126 23488
rect 12070 23432 12126 23468
rect 11058 23160 11114 23216
rect 11622 22330 11678 22332
rect 11702 22330 11758 22332
rect 11782 22330 11838 22332
rect 11862 22330 11918 22332
rect 11622 22278 11648 22330
rect 11648 22278 11678 22330
rect 11702 22278 11712 22330
rect 11712 22278 11758 22330
rect 11782 22278 11828 22330
rect 11828 22278 11838 22330
rect 11862 22278 11892 22330
rect 11892 22278 11918 22330
rect 11622 22276 11678 22278
rect 11702 22276 11758 22278
rect 11782 22276 11838 22278
rect 11862 22276 11918 22278
rect 11058 22072 11114 22128
rect 11622 21242 11678 21244
rect 11702 21242 11758 21244
rect 11782 21242 11838 21244
rect 11862 21242 11918 21244
rect 11622 21190 11648 21242
rect 11648 21190 11678 21242
rect 11702 21190 11712 21242
rect 11712 21190 11758 21242
rect 11782 21190 11828 21242
rect 11828 21190 11838 21242
rect 11862 21190 11892 21242
rect 11892 21190 11918 21242
rect 11622 21188 11678 21190
rect 11702 21188 11758 21190
rect 11782 21188 11838 21190
rect 11862 21188 11918 21190
rect 11150 20168 11206 20224
rect 10138 9016 10194 9072
rect 9954 3440 10010 3496
rect 9954 1400 10010 1456
rect 11622 20154 11678 20156
rect 11702 20154 11758 20156
rect 11782 20154 11838 20156
rect 11862 20154 11918 20156
rect 11622 20102 11648 20154
rect 11648 20102 11678 20154
rect 11702 20102 11712 20154
rect 11712 20102 11758 20154
rect 11782 20102 11828 20154
rect 11828 20102 11838 20154
rect 11862 20102 11892 20154
rect 11892 20102 11918 20154
rect 11622 20100 11678 20102
rect 11702 20100 11758 20102
rect 11782 20100 11838 20102
rect 11862 20100 11918 20102
rect 11622 19066 11678 19068
rect 11702 19066 11758 19068
rect 11782 19066 11838 19068
rect 11862 19066 11918 19068
rect 11622 19014 11648 19066
rect 11648 19014 11678 19066
rect 11702 19014 11712 19066
rect 11712 19014 11758 19066
rect 11782 19014 11828 19066
rect 11828 19014 11838 19066
rect 11862 19014 11892 19066
rect 11892 19014 11918 19066
rect 11622 19012 11678 19014
rect 11702 19012 11758 19014
rect 11782 19012 11838 19014
rect 11862 19012 11918 19014
rect 11622 17978 11678 17980
rect 11702 17978 11758 17980
rect 11782 17978 11838 17980
rect 11862 17978 11918 17980
rect 11622 17926 11648 17978
rect 11648 17926 11678 17978
rect 11702 17926 11712 17978
rect 11712 17926 11758 17978
rect 11782 17926 11828 17978
rect 11828 17926 11838 17978
rect 11862 17926 11892 17978
rect 11892 17926 11918 17978
rect 11622 17924 11678 17926
rect 11702 17924 11758 17926
rect 11782 17924 11838 17926
rect 11862 17924 11918 17926
rect 13358 35536 13414 35592
rect 12438 22072 12494 22128
rect 12254 17176 12310 17232
rect 11622 16890 11678 16892
rect 11702 16890 11758 16892
rect 11782 16890 11838 16892
rect 11862 16890 11918 16892
rect 11622 16838 11648 16890
rect 11648 16838 11678 16890
rect 11702 16838 11712 16890
rect 11712 16838 11758 16890
rect 11782 16838 11828 16890
rect 11828 16838 11838 16890
rect 11862 16838 11892 16890
rect 11892 16838 11918 16890
rect 11622 16836 11678 16838
rect 11702 16836 11758 16838
rect 11782 16836 11838 16838
rect 11862 16836 11918 16838
rect 11518 16652 11574 16688
rect 11518 16632 11520 16652
rect 11520 16632 11572 16652
rect 11572 16632 11574 16652
rect 11622 15802 11678 15804
rect 11702 15802 11758 15804
rect 11782 15802 11838 15804
rect 11862 15802 11918 15804
rect 11622 15750 11648 15802
rect 11648 15750 11678 15802
rect 11702 15750 11712 15802
rect 11712 15750 11758 15802
rect 11782 15750 11828 15802
rect 11828 15750 11838 15802
rect 11862 15750 11892 15802
rect 11892 15750 11918 15802
rect 11622 15748 11678 15750
rect 11702 15748 11758 15750
rect 11782 15748 11838 15750
rect 11862 15748 11918 15750
rect 10598 9424 10654 9480
rect 10414 6704 10470 6760
rect 10322 6160 10378 6216
rect 10598 4664 10654 4720
rect 10506 4120 10562 4176
rect 10598 3984 10654 4040
rect 10414 3188 10470 3224
rect 10414 3168 10416 3188
rect 10416 3168 10468 3188
rect 10468 3168 10470 3188
rect 10414 2508 10470 2544
rect 10414 2488 10416 2508
rect 10416 2488 10468 2508
rect 10468 2488 10470 2508
rect 10966 3440 11022 3496
rect 10966 3304 11022 3360
rect 11622 14714 11678 14716
rect 11702 14714 11758 14716
rect 11782 14714 11838 14716
rect 11862 14714 11918 14716
rect 11622 14662 11648 14714
rect 11648 14662 11678 14714
rect 11702 14662 11712 14714
rect 11712 14662 11758 14714
rect 11782 14662 11828 14714
rect 11828 14662 11838 14714
rect 11862 14662 11892 14714
rect 11892 14662 11918 14714
rect 11622 14660 11678 14662
rect 11702 14660 11758 14662
rect 11782 14660 11838 14662
rect 11862 14660 11918 14662
rect 11622 13626 11678 13628
rect 11702 13626 11758 13628
rect 11782 13626 11838 13628
rect 11862 13626 11918 13628
rect 11622 13574 11648 13626
rect 11648 13574 11678 13626
rect 11702 13574 11712 13626
rect 11712 13574 11758 13626
rect 11782 13574 11828 13626
rect 11828 13574 11838 13626
rect 11862 13574 11892 13626
rect 11892 13574 11918 13626
rect 11622 13572 11678 13574
rect 11702 13572 11758 13574
rect 11782 13572 11838 13574
rect 11862 13572 11918 13574
rect 11622 12538 11678 12540
rect 11702 12538 11758 12540
rect 11782 12538 11838 12540
rect 11862 12538 11918 12540
rect 11622 12486 11648 12538
rect 11648 12486 11678 12538
rect 11702 12486 11712 12538
rect 11712 12486 11758 12538
rect 11782 12486 11828 12538
rect 11828 12486 11838 12538
rect 11862 12486 11892 12538
rect 11892 12486 11918 12538
rect 11622 12484 11678 12486
rect 11702 12484 11758 12486
rect 11782 12484 11838 12486
rect 11862 12484 11918 12486
rect 11622 11450 11678 11452
rect 11702 11450 11758 11452
rect 11782 11450 11838 11452
rect 11862 11450 11918 11452
rect 11622 11398 11648 11450
rect 11648 11398 11678 11450
rect 11702 11398 11712 11450
rect 11712 11398 11758 11450
rect 11782 11398 11828 11450
rect 11828 11398 11838 11450
rect 11862 11398 11892 11450
rect 11892 11398 11918 11450
rect 11622 11396 11678 11398
rect 11702 11396 11758 11398
rect 11782 11396 11838 11398
rect 11862 11396 11918 11398
rect 11622 10362 11678 10364
rect 11702 10362 11758 10364
rect 11782 10362 11838 10364
rect 11862 10362 11918 10364
rect 11622 10310 11648 10362
rect 11648 10310 11678 10362
rect 11702 10310 11712 10362
rect 11712 10310 11758 10362
rect 11782 10310 11828 10362
rect 11828 10310 11838 10362
rect 11862 10310 11892 10362
rect 11892 10310 11918 10362
rect 11622 10308 11678 10310
rect 11702 10308 11758 10310
rect 11782 10308 11838 10310
rect 11862 10308 11918 10310
rect 11622 9274 11678 9276
rect 11702 9274 11758 9276
rect 11782 9274 11838 9276
rect 11862 9274 11918 9276
rect 11622 9222 11648 9274
rect 11648 9222 11678 9274
rect 11702 9222 11712 9274
rect 11712 9222 11758 9274
rect 11782 9222 11828 9274
rect 11828 9222 11838 9274
rect 11862 9222 11892 9274
rect 11892 9222 11918 9274
rect 11622 9220 11678 9222
rect 11702 9220 11758 9222
rect 11782 9220 11838 9222
rect 11862 9220 11918 9222
rect 11622 8186 11678 8188
rect 11702 8186 11758 8188
rect 11782 8186 11838 8188
rect 11862 8186 11918 8188
rect 11622 8134 11648 8186
rect 11648 8134 11678 8186
rect 11702 8134 11712 8186
rect 11712 8134 11758 8186
rect 11782 8134 11828 8186
rect 11828 8134 11838 8186
rect 11862 8134 11892 8186
rect 11892 8134 11918 8186
rect 11622 8132 11678 8134
rect 11702 8132 11758 8134
rect 11782 8132 11838 8134
rect 11862 8132 11918 8134
rect 11622 7098 11678 7100
rect 11702 7098 11758 7100
rect 11782 7098 11838 7100
rect 11862 7098 11918 7100
rect 11622 7046 11648 7098
rect 11648 7046 11678 7098
rect 11702 7046 11712 7098
rect 11712 7046 11758 7098
rect 11782 7046 11828 7098
rect 11828 7046 11838 7098
rect 11862 7046 11892 7098
rect 11892 7046 11918 7098
rect 11622 7044 11678 7046
rect 11702 7044 11758 7046
rect 11782 7044 11838 7046
rect 11862 7044 11918 7046
rect 11622 6010 11678 6012
rect 11702 6010 11758 6012
rect 11782 6010 11838 6012
rect 11862 6010 11918 6012
rect 11622 5958 11648 6010
rect 11648 5958 11678 6010
rect 11702 5958 11712 6010
rect 11712 5958 11758 6010
rect 11782 5958 11828 6010
rect 11828 5958 11838 6010
rect 11862 5958 11892 6010
rect 11892 5958 11918 6010
rect 11622 5956 11678 5958
rect 11702 5956 11758 5958
rect 11782 5956 11838 5958
rect 11862 5956 11918 5958
rect 11334 5752 11390 5808
rect 11150 3712 11206 3768
rect 11150 3304 11206 3360
rect 12346 4936 12402 4992
rect 11622 4922 11678 4924
rect 11702 4922 11758 4924
rect 11782 4922 11838 4924
rect 11862 4922 11918 4924
rect 11622 4870 11648 4922
rect 11648 4870 11678 4922
rect 11702 4870 11712 4922
rect 11712 4870 11758 4922
rect 11782 4870 11828 4922
rect 11828 4870 11838 4922
rect 11862 4870 11892 4922
rect 11892 4870 11918 4922
rect 11622 4868 11678 4870
rect 11702 4868 11758 4870
rect 11782 4868 11838 4870
rect 11862 4868 11918 4870
rect 11426 3848 11482 3904
rect 11426 3068 11428 3088
rect 11428 3068 11480 3088
rect 11480 3068 11482 3088
rect 11426 3032 11482 3068
rect 11426 2644 11482 2680
rect 11426 2624 11428 2644
rect 11428 2624 11480 2644
rect 11480 2624 11482 2644
rect 11622 3834 11678 3836
rect 11702 3834 11758 3836
rect 11782 3834 11838 3836
rect 11862 3834 11918 3836
rect 11622 3782 11648 3834
rect 11648 3782 11678 3834
rect 11702 3782 11712 3834
rect 11712 3782 11758 3834
rect 11782 3782 11828 3834
rect 11828 3782 11838 3834
rect 11862 3782 11892 3834
rect 11892 3782 11918 3834
rect 11622 3780 11678 3782
rect 11702 3780 11758 3782
rect 11782 3780 11838 3782
rect 11862 3780 11918 3782
rect 11610 3576 11666 3632
rect 12530 9560 12586 9616
rect 12622 3304 12678 3360
rect 11610 3032 11666 3088
rect 12438 3032 12494 3088
rect 12622 2896 12678 2952
rect 11622 2746 11678 2748
rect 11702 2746 11758 2748
rect 11782 2746 11838 2748
rect 11862 2746 11918 2748
rect 11622 2694 11648 2746
rect 11648 2694 11678 2746
rect 11702 2694 11712 2746
rect 11712 2694 11758 2746
rect 11782 2694 11828 2746
rect 11828 2694 11838 2746
rect 11862 2694 11892 2746
rect 11892 2694 11918 2746
rect 11622 2692 11678 2694
rect 11702 2692 11758 2694
rect 11782 2692 11838 2694
rect 11862 2692 11918 2694
rect 13082 8356 13138 8392
rect 13082 8336 13084 8356
rect 13084 8336 13136 8356
rect 13136 8336 13138 8356
rect 14289 37018 14345 37020
rect 14369 37018 14425 37020
rect 14449 37018 14505 37020
rect 14529 37018 14585 37020
rect 14289 36966 14315 37018
rect 14315 36966 14345 37018
rect 14369 36966 14379 37018
rect 14379 36966 14425 37018
rect 14449 36966 14495 37018
rect 14495 36966 14505 37018
rect 14529 36966 14559 37018
rect 14559 36966 14585 37018
rect 14289 36964 14345 36966
rect 14369 36964 14425 36966
rect 14449 36964 14505 36966
rect 14529 36964 14585 36966
rect 14289 35930 14345 35932
rect 14369 35930 14425 35932
rect 14449 35930 14505 35932
rect 14529 35930 14585 35932
rect 14289 35878 14315 35930
rect 14315 35878 14345 35930
rect 14369 35878 14379 35930
rect 14379 35878 14425 35930
rect 14449 35878 14495 35930
rect 14495 35878 14505 35930
rect 14529 35878 14559 35930
rect 14559 35878 14585 35930
rect 14289 35876 14345 35878
rect 14369 35876 14425 35878
rect 14449 35876 14505 35878
rect 14529 35876 14585 35878
rect 14289 34842 14345 34844
rect 14369 34842 14425 34844
rect 14449 34842 14505 34844
rect 14529 34842 14585 34844
rect 14289 34790 14315 34842
rect 14315 34790 14345 34842
rect 14369 34790 14379 34842
rect 14379 34790 14425 34842
rect 14449 34790 14495 34842
rect 14495 34790 14505 34842
rect 14529 34790 14559 34842
rect 14559 34790 14585 34842
rect 14289 34788 14345 34790
rect 14369 34788 14425 34790
rect 14449 34788 14505 34790
rect 14529 34788 14585 34790
rect 14289 33754 14345 33756
rect 14369 33754 14425 33756
rect 14449 33754 14505 33756
rect 14529 33754 14585 33756
rect 14289 33702 14315 33754
rect 14315 33702 14345 33754
rect 14369 33702 14379 33754
rect 14379 33702 14425 33754
rect 14449 33702 14495 33754
rect 14495 33702 14505 33754
rect 14529 33702 14559 33754
rect 14559 33702 14585 33754
rect 14289 33700 14345 33702
rect 14369 33700 14425 33702
rect 14449 33700 14505 33702
rect 14529 33700 14585 33702
rect 14289 32666 14345 32668
rect 14369 32666 14425 32668
rect 14449 32666 14505 32668
rect 14529 32666 14585 32668
rect 14289 32614 14315 32666
rect 14315 32614 14345 32666
rect 14369 32614 14379 32666
rect 14379 32614 14425 32666
rect 14449 32614 14495 32666
rect 14495 32614 14505 32666
rect 14529 32614 14559 32666
rect 14559 32614 14585 32666
rect 14289 32612 14345 32614
rect 14369 32612 14425 32614
rect 14449 32612 14505 32614
rect 14529 32612 14585 32614
rect 14289 31578 14345 31580
rect 14369 31578 14425 31580
rect 14449 31578 14505 31580
rect 14529 31578 14585 31580
rect 14289 31526 14315 31578
rect 14315 31526 14345 31578
rect 14369 31526 14379 31578
rect 14379 31526 14425 31578
rect 14449 31526 14495 31578
rect 14495 31526 14505 31578
rect 14529 31526 14559 31578
rect 14559 31526 14585 31578
rect 14289 31524 14345 31526
rect 14369 31524 14425 31526
rect 14449 31524 14505 31526
rect 14529 31524 14585 31526
rect 14289 30490 14345 30492
rect 14369 30490 14425 30492
rect 14449 30490 14505 30492
rect 14529 30490 14585 30492
rect 14289 30438 14315 30490
rect 14315 30438 14345 30490
rect 14369 30438 14379 30490
rect 14379 30438 14425 30490
rect 14449 30438 14495 30490
rect 14495 30438 14505 30490
rect 14529 30438 14559 30490
rect 14559 30438 14585 30490
rect 14289 30436 14345 30438
rect 14369 30436 14425 30438
rect 14449 30436 14505 30438
rect 14529 30436 14585 30438
rect 14646 30232 14702 30288
rect 14289 29402 14345 29404
rect 14369 29402 14425 29404
rect 14449 29402 14505 29404
rect 14529 29402 14585 29404
rect 14289 29350 14315 29402
rect 14315 29350 14345 29402
rect 14369 29350 14379 29402
rect 14379 29350 14425 29402
rect 14449 29350 14495 29402
rect 14495 29350 14505 29402
rect 14529 29350 14559 29402
rect 14559 29350 14585 29402
rect 14289 29348 14345 29350
rect 14369 29348 14425 29350
rect 14449 29348 14505 29350
rect 14529 29348 14585 29350
rect 14289 28314 14345 28316
rect 14369 28314 14425 28316
rect 14449 28314 14505 28316
rect 14529 28314 14585 28316
rect 14289 28262 14315 28314
rect 14315 28262 14345 28314
rect 14369 28262 14379 28314
rect 14379 28262 14425 28314
rect 14449 28262 14495 28314
rect 14495 28262 14505 28314
rect 14529 28262 14559 28314
rect 14559 28262 14585 28314
rect 14289 28260 14345 28262
rect 14369 28260 14425 28262
rect 14449 28260 14505 28262
rect 14529 28260 14585 28262
rect 14289 27226 14345 27228
rect 14369 27226 14425 27228
rect 14449 27226 14505 27228
rect 14529 27226 14585 27228
rect 14289 27174 14315 27226
rect 14315 27174 14345 27226
rect 14369 27174 14379 27226
rect 14379 27174 14425 27226
rect 14449 27174 14495 27226
rect 14495 27174 14505 27226
rect 14529 27174 14559 27226
rect 14559 27174 14585 27226
rect 14289 27172 14345 27174
rect 14369 27172 14425 27174
rect 14449 27172 14505 27174
rect 14529 27172 14585 27174
rect 13818 21800 13874 21856
rect 13358 4120 13414 4176
rect 13174 3168 13230 3224
rect 13266 2760 13322 2816
rect 12898 2488 12954 2544
rect 12806 2372 12862 2408
rect 12806 2352 12808 2372
rect 12808 2352 12860 2372
rect 12860 2352 12862 2372
rect 12530 2216 12586 2272
rect 12990 1944 13046 2000
rect 13726 3440 13782 3496
rect 14289 26138 14345 26140
rect 14369 26138 14425 26140
rect 14449 26138 14505 26140
rect 14529 26138 14585 26140
rect 14289 26086 14315 26138
rect 14315 26086 14345 26138
rect 14369 26086 14379 26138
rect 14379 26086 14425 26138
rect 14449 26086 14495 26138
rect 14495 26086 14505 26138
rect 14529 26086 14559 26138
rect 14559 26086 14585 26138
rect 14289 26084 14345 26086
rect 14369 26084 14425 26086
rect 14449 26084 14505 26086
rect 14529 26084 14585 26086
rect 14289 25050 14345 25052
rect 14369 25050 14425 25052
rect 14449 25050 14505 25052
rect 14529 25050 14585 25052
rect 14289 24998 14315 25050
rect 14315 24998 14345 25050
rect 14369 24998 14379 25050
rect 14379 24998 14425 25050
rect 14449 24998 14495 25050
rect 14495 24998 14505 25050
rect 14529 24998 14559 25050
rect 14559 24998 14585 25050
rect 14289 24996 14345 24998
rect 14369 24996 14425 24998
rect 14449 24996 14505 24998
rect 14529 24996 14585 24998
rect 14289 23962 14345 23964
rect 14369 23962 14425 23964
rect 14449 23962 14505 23964
rect 14529 23962 14585 23964
rect 14289 23910 14315 23962
rect 14315 23910 14345 23962
rect 14369 23910 14379 23962
rect 14379 23910 14425 23962
rect 14449 23910 14495 23962
rect 14495 23910 14505 23962
rect 14529 23910 14559 23962
rect 14559 23910 14585 23962
rect 14289 23908 14345 23910
rect 14369 23908 14425 23910
rect 14449 23908 14505 23910
rect 14529 23908 14585 23910
rect 14186 23432 14242 23488
rect 14289 22874 14345 22876
rect 14369 22874 14425 22876
rect 14449 22874 14505 22876
rect 14529 22874 14585 22876
rect 14289 22822 14315 22874
rect 14315 22822 14345 22874
rect 14369 22822 14379 22874
rect 14379 22822 14425 22874
rect 14449 22822 14495 22874
rect 14495 22822 14505 22874
rect 14529 22822 14559 22874
rect 14559 22822 14585 22874
rect 14289 22820 14345 22822
rect 14369 22820 14425 22822
rect 14449 22820 14505 22822
rect 14529 22820 14585 22822
rect 14289 21786 14345 21788
rect 14369 21786 14425 21788
rect 14449 21786 14505 21788
rect 14529 21786 14585 21788
rect 14289 21734 14315 21786
rect 14315 21734 14345 21786
rect 14369 21734 14379 21786
rect 14379 21734 14425 21786
rect 14449 21734 14495 21786
rect 14495 21734 14505 21786
rect 14529 21734 14559 21786
rect 14559 21734 14585 21786
rect 14289 21732 14345 21734
rect 14369 21732 14425 21734
rect 14449 21732 14505 21734
rect 14529 21732 14585 21734
rect 14289 20698 14345 20700
rect 14369 20698 14425 20700
rect 14449 20698 14505 20700
rect 14529 20698 14585 20700
rect 14289 20646 14315 20698
rect 14315 20646 14345 20698
rect 14369 20646 14379 20698
rect 14379 20646 14425 20698
rect 14449 20646 14495 20698
rect 14495 20646 14505 20698
rect 14529 20646 14559 20698
rect 14559 20646 14585 20698
rect 14289 20644 14345 20646
rect 14369 20644 14425 20646
rect 14449 20644 14505 20646
rect 14529 20644 14585 20646
rect 14289 19610 14345 19612
rect 14369 19610 14425 19612
rect 14449 19610 14505 19612
rect 14529 19610 14585 19612
rect 14289 19558 14315 19610
rect 14315 19558 14345 19610
rect 14369 19558 14379 19610
rect 14379 19558 14425 19610
rect 14449 19558 14495 19610
rect 14495 19558 14505 19610
rect 14529 19558 14559 19610
rect 14559 19558 14585 19610
rect 14289 19556 14345 19558
rect 14369 19556 14425 19558
rect 14449 19556 14505 19558
rect 14529 19556 14585 19558
rect 14289 18522 14345 18524
rect 14369 18522 14425 18524
rect 14449 18522 14505 18524
rect 14529 18522 14585 18524
rect 14289 18470 14315 18522
rect 14315 18470 14345 18522
rect 14369 18470 14379 18522
rect 14379 18470 14425 18522
rect 14449 18470 14495 18522
rect 14495 18470 14505 18522
rect 14529 18470 14559 18522
rect 14559 18470 14585 18522
rect 14289 18468 14345 18470
rect 14369 18468 14425 18470
rect 14449 18468 14505 18470
rect 14529 18468 14585 18470
rect 14289 17434 14345 17436
rect 14369 17434 14425 17436
rect 14449 17434 14505 17436
rect 14529 17434 14585 17436
rect 14289 17382 14315 17434
rect 14315 17382 14345 17434
rect 14369 17382 14379 17434
rect 14379 17382 14425 17434
rect 14449 17382 14495 17434
rect 14495 17382 14505 17434
rect 14529 17382 14559 17434
rect 14559 17382 14585 17434
rect 14289 17380 14345 17382
rect 14369 17380 14425 17382
rect 14449 17380 14505 17382
rect 14529 17380 14585 17382
rect 14289 16346 14345 16348
rect 14369 16346 14425 16348
rect 14449 16346 14505 16348
rect 14529 16346 14585 16348
rect 14289 16294 14315 16346
rect 14315 16294 14345 16346
rect 14369 16294 14379 16346
rect 14379 16294 14425 16346
rect 14449 16294 14495 16346
rect 14495 16294 14505 16346
rect 14529 16294 14559 16346
rect 14559 16294 14585 16346
rect 14289 16292 14345 16294
rect 14369 16292 14425 16294
rect 14449 16292 14505 16294
rect 14529 16292 14585 16294
rect 14289 15258 14345 15260
rect 14369 15258 14425 15260
rect 14449 15258 14505 15260
rect 14529 15258 14585 15260
rect 14289 15206 14315 15258
rect 14315 15206 14345 15258
rect 14369 15206 14379 15258
rect 14379 15206 14425 15258
rect 14449 15206 14495 15258
rect 14495 15206 14505 15258
rect 14529 15206 14559 15258
rect 14559 15206 14585 15258
rect 14289 15204 14345 15206
rect 14369 15204 14425 15206
rect 14449 15204 14505 15206
rect 14529 15204 14585 15206
rect 14289 14170 14345 14172
rect 14369 14170 14425 14172
rect 14449 14170 14505 14172
rect 14529 14170 14585 14172
rect 14289 14118 14315 14170
rect 14315 14118 14345 14170
rect 14369 14118 14379 14170
rect 14379 14118 14425 14170
rect 14449 14118 14495 14170
rect 14495 14118 14505 14170
rect 14529 14118 14559 14170
rect 14559 14118 14585 14170
rect 14289 14116 14345 14118
rect 14369 14116 14425 14118
rect 14449 14116 14505 14118
rect 14529 14116 14585 14118
rect 14289 13082 14345 13084
rect 14369 13082 14425 13084
rect 14449 13082 14505 13084
rect 14529 13082 14585 13084
rect 14289 13030 14315 13082
rect 14315 13030 14345 13082
rect 14369 13030 14379 13082
rect 14379 13030 14425 13082
rect 14449 13030 14495 13082
rect 14495 13030 14505 13082
rect 14529 13030 14559 13082
rect 14559 13030 14585 13082
rect 14289 13028 14345 13030
rect 14369 13028 14425 13030
rect 14449 13028 14505 13030
rect 14529 13028 14585 13030
rect 14289 11994 14345 11996
rect 14369 11994 14425 11996
rect 14449 11994 14505 11996
rect 14529 11994 14585 11996
rect 14289 11942 14315 11994
rect 14315 11942 14345 11994
rect 14369 11942 14379 11994
rect 14379 11942 14425 11994
rect 14449 11942 14495 11994
rect 14495 11942 14505 11994
rect 14529 11942 14559 11994
rect 14559 11942 14585 11994
rect 14289 11940 14345 11942
rect 14369 11940 14425 11942
rect 14449 11940 14505 11942
rect 14529 11940 14585 11942
rect 14289 10906 14345 10908
rect 14369 10906 14425 10908
rect 14449 10906 14505 10908
rect 14529 10906 14585 10908
rect 14289 10854 14315 10906
rect 14315 10854 14345 10906
rect 14369 10854 14379 10906
rect 14379 10854 14425 10906
rect 14449 10854 14495 10906
rect 14495 10854 14505 10906
rect 14529 10854 14559 10906
rect 14559 10854 14585 10906
rect 14289 10852 14345 10854
rect 14369 10852 14425 10854
rect 14449 10852 14505 10854
rect 14529 10852 14585 10854
rect 14289 9818 14345 9820
rect 14369 9818 14425 9820
rect 14449 9818 14505 9820
rect 14529 9818 14585 9820
rect 14289 9766 14315 9818
rect 14315 9766 14345 9818
rect 14369 9766 14379 9818
rect 14379 9766 14425 9818
rect 14449 9766 14495 9818
rect 14495 9766 14505 9818
rect 14529 9766 14559 9818
rect 14559 9766 14585 9818
rect 14289 9764 14345 9766
rect 14369 9764 14425 9766
rect 14449 9764 14505 9766
rect 14529 9764 14585 9766
rect 14289 8730 14345 8732
rect 14369 8730 14425 8732
rect 14449 8730 14505 8732
rect 14529 8730 14585 8732
rect 14289 8678 14315 8730
rect 14315 8678 14345 8730
rect 14369 8678 14379 8730
rect 14379 8678 14425 8730
rect 14449 8678 14495 8730
rect 14495 8678 14505 8730
rect 14529 8678 14559 8730
rect 14559 8678 14585 8730
rect 14289 8676 14345 8678
rect 14369 8676 14425 8678
rect 14449 8676 14505 8678
rect 14529 8676 14585 8678
rect 14289 7642 14345 7644
rect 14369 7642 14425 7644
rect 14449 7642 14505 7644
rect 14529 7642 14585 7644
rect 14289 7590 14315 7642
rect 14315 7590 14345 7642
rect 14369 7590 14379 7642
rect 14379 7590 14425 7642
rect 14449 7590 14495 7642
rect 14495 7590 14505 7642
rect 14529 7590 14559 7642
rect 14559 7590 14585 7642
rect 14289 7588 14345 7590
rect 14369 7588 14425 7590
rect 14449 7588 14505 7590
rect 14529 7588 14585 7590
rect 14289 6554 14345 6556
rect 14369 6554 14425 6556
rect 14449 6554 14505 6556
rect 14529 6554 14585 6556
rect 14289 6502 14315 6554
rect 14315 6502 14345 6554
rect 14369 6502 14379 6554
rect 14379 6502 14425 6554
rect 14449 6502 14495 6554
rect 14495 6502 14505 6554
rect 14529 6502 14559 6554
rect 14559 6502 14585 6554
rect 14289 6500 14345 6502
rect 14369 6500 14425 6502
rect 14449 6500 14505 6502
rect 14529 6500 14585 6502
rect 14289 5466 14345 5468
rect 14369 5466 14425 5468
rect 14449 5466 14505 5468
rect 14529 5466 14585 5468
rect 14289 5414 14315 5466
rect 14315 5414 14345 5466
rect 14369 5414 14379 5466
rect 14379 5414 14425 5466
rect 14449 5414 14495 5466
rect 14495 5414 14505 5466
rect 14529 5414 14559 5466
rect 14559 5414 14585 5466
rect 14289 5412 14345 5414
rect 14369 5412 14425 5414
rect 14449 5412 14505 5414
rect 14529 5412 14585 5414
rect 14289 4378 14345 4380
rect 14369 4378 14425 4380
rect 14449 4378 14505 4380
rect 14529 4378 14585 4380
rect 14289 4326 14315 4378
rect 14315 4326 14345 4378
rect 14369 4326 14379 4378
rect 14379 4326 14425 4378
rect 14449 4326 14495 4378
rect 14495 4326 14505 4378
rect 14529 4326 14559 4378
rect 14559 4326 14585 4378
rect 14289 4324 14345 4326
rect 14369 4324 14425 4326
rect 14449 4324 14505 4326
rect 14529 4324 14585 4326
rect 14289 3290 14345 3292
rect 14369 3290 14425 3292
rect 14449 3290 14505 3292
rect 14529 3290 14585 3292
rect 14289 3238 14315 3290
rect 14315 3238 14345 3290
rect 14369 3238 14379 3290
rect 14379 3238 14425 3290
rect 14449 3238 14495 3290
rect 14495 3238 14505 3290
rect 14529 3238 14559 3290
rect 14559 3238 14585 3290
rect 14289 3236 14345 3238
rect 14369 3236 14425 3238
rect 14449 3236 14505 3238
rect 14529 3236 14585 3238
rect 15750 8336 15806 8392
rect 15382 2760 15438 2816
rect 14289 2202 14345 2204
rect 14369 2202 14425 2204
rect 14449 2202 14505 2204
rect 14529 2202 14585 2204
rect 14289 2150 14315 2202
rect 14315 2150 14345 2202
rect 14369 2150 14379 2202
rect 14379 2150 14425 2202
rect 14449 2150 14495 2202
rect 14495 2150 14505 2202
rect 14529 2150 14559 2202
rect 14559 2150 14585 2202
rect 14289 2148 14345 2150
rect 14369 2148 14425 2150
rect 14449 2148 14505 2150
rect 14529 2148 14585 2150
<< metal3 >>
rect 6277 37568 6597 37569
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 37503 6597 37504
rect 11610 37568 11930 37569
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 37503 11930 37504
rect 3610 37024 3930 37025
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3930 37024
rect 3610 36959 3930 36960
rect 8944 37024 9264 37025
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 36959 9264 36960
rect 14277 37024 14597 37025
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 36959 14597 36960
rect 0 36682 480 36712
rect 1945 36682 2011 36685
rect 0 36680 2011 36682
rect 0 36624 1950 36680
rect 2006 36624 2011 36680
rect 0 36622 2011 36624
rect 0 36592 480 36622
rect 1945 36619 2011 36622
rect 6277 36480 6597 36481
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 36415 6597 36416
rect 11610 36480 11930 36481
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 36415 11930 36416
rect 3610 35936 3930 35937
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3930 35936
rect 3610 35871 3930 35872
rect 8944 35936 9264 35937
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 35871 9264 35872
rect 14277 35936 14597 35937
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 35871 14597 35872
rect 9397 35730 9463 35733
rect 6134 35728 9463 35730
rect 6134 35672 9402 35728
rect 9458 35672 9463 35728
rect 6134 35670 9463 35672
rect 2313 35594 2379 35597
rect 6134 35594 6194 35670
rect 9397 35667 9463 35670
rect 2313 35592 6194 35594
rect 2313 35536 2318 35592
rect 2374 35536 6194 35592
rect 2313 35534 6194 35536
rect 8661 35594 8727 35597
rect 13353 35594 13419 35597
rect 8661 35592 13419 35594
rect 8661 35536 8666 35592
rect 8722 35536 13358 35592
rect 13414 35536 13419 35592
rect 8661 35534 13419 35536
rect 2313 35531 2379 35534
rect 8661 35531 8727 35534
rect 13353 35531 13419 35534
rect 6277 35392 6597 35393
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 35327 6597 35328
rect 11610 35392 11930 35393
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 35327 11930 35328
rect 5993 35186 6059 35189
rect 10961 35186 11027 35189
rect 5993 35184 11027 35186
rect 5993 35128 5998 35184
rect 6054 35128 10966 35184
rect 11022 35128 11027 35184
rect 5993 35126 11027 35128
rect 5993 35123 6059 35126
rect 10961 35123 11027 35126
rect 5809 35050 5875 35053
rect 11329 35050 11395 35053
rect 5809 35048 11395 35050
rect 5809 34992 5814 35048
rect 5870 34992 11334 35048
rect 11390 34992 11395 35048
rect 5809 34990 11395 34992
rect 5809 34987 5875 34990
rect 11329 34987 11395 34990
rect 15520 34914 16000 34944
rect 14782 34854 16000 34914
rect 3610 34848 3930 34849
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3930 34848
rect 3610 34783 3930 34784
rect 8944 34848 9264 34849
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 34783 9264 34784
rect 14277 34848 14597 34849
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 34783 14597 34784
rect 4429 34642 4495 34645
rect 11513 34642 11579 34645
rect 4429 34640 11579 34642
rect 4429 34584 4434 34640
rect 4490 34584 11518 34640
rect 11574 34584 11579 34640
rect 4429 34582 11579 34584
rect 4429 34579 4495 34582
rect 11513 34579 11579 34582
rect 12341 34642 12407 34645
rect 14782 34642 14842 34854
rect 15520 34824 16000 34854
rect 12341 34640 14842 34642
rect 12341 34584 12346 34640
rect 12402 34584 14842 34640
rect 12341 34582 14842 34584
rect 12341 34579 12407 34582
rect 6277 34304 6597 34305
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 34239 6597 34240
rect 11610 34304 11930 34305
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 34239 11930 34240
rect 3610 33760 3930 33761
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3930 33760
rect 3610 33695 3930 33696
rect 8944 33760 9264 33761
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 33695 9264 33696
rect 14277 33760 14597 33761
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 33695 14597 33696
rect 6277 33216 6597 33217
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 33151 6597 33152
rect 11610 33216 11930 33217
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 33151 11930 33152
rect 6821 33146 6887 33149
rect 8753 33146 8819 33149
rect 6821 33144 8819 33146
rect 6821 33088 6826 33144
rect 6882 33088 8758 33144
rect 8814 33088 8819 33144
rect 6821 33086 8819 33088
rect 6821 33083 6887 33086
rect 8753 33083 8819 33086
rect 3610 32672 3930 32673
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3930 32672
rect 3610 32607 3930 32608
rect 8944 32672 9264 32673
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 32607 9264 32608
rect 14277 32672 14597 32673
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 32607 14597 32608
rect 6277 32128 6597 32129
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 32063 6597 32064
rect 11610 32128 11930 32129
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 32063 11930 32064
rect 3610 31584 3930 31585
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3930 31584
rect 3610 31519 3930 31520
rect 8944 31584 9264 31585
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 31519 9264 31520
rect 14277 31584 14597 31585
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 31519 14597 31520
rect 6277 31040 6597 31041
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 30975 6597 30976
rect 11610 31040 11930 31041
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 30975 11930 30976
rect 3610 30496 3930 30497
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3930 30496
rect 3610 30431 3930 30432
rect 8944 30496 9264 30497
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 30431 9264 30432
rect 14277 30496 14597 30497
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 30431 14597 30432
rect 9765 30290 9831 30293
rect 14641 30290 14707 30293
rect 9765 30288 14707 30290
rect 9765 30232 9770 30288
rect 9826 30232 14646 30288
rect 14702 30232 14707 30288
rect 9765 30230 14707 30232
rect 9765 30227 9831 30230
rect 14641 30227 14707 30230
rect 0 30018 480 30048
rect 1577 30018 1643 30021
rect 0 30016 1643 30018
rect 0 29960 1582 30016
rect 1638 29960 1643 30016
rect 0 29958 1643 29960
rect 0 29928 480 29958
rect 1577 29955 1643 29958
rect 6277 29952 6597 29953
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 29887 6597 29888
rect 11610 29952 11930 29953
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 29887 11930 29888
rect 3610 29408 3930 29409
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3930 29408
rect 3610 29343 3930 29344
rect 8944 29408 9264 29409
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 29343 9264 29344
rect 14277 29408 14597 29409
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 29343 14597 29344
rect 4429 29066 4495 29069
rect 4429 29064 4538 29066
rect 4429 29008 4434 29064
rect 4490 29032 4538 29064
rect 4613 29032 4679 29035
rect 4490 29030 4679 29032
rect 4490 29008 4618 29030
rect 4429 29003 4618 29008
rect 4478 28974 4618 29003
rect 4674 28974 4679 29030
rect 4478 28972 4679 28974
rect 4613 28969 4679 28972
rect 6277 28864 6597 28865
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 28799 6597 28800
rect 11610 28864 11930 28865
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 28799 11930 28800
rect 5349 28658 5415 28661
rect 7649 28658 7715 28661
rect 5349 28656 7715 28658
rect 5349 28600 5354 28656
rect 5410 28600 7654 28656
rect 7710 28600 7715 28656
rect 5349 28598 7715 28600
rect 5349 28595 5415 28598
rect 7649 28595 7715 28598
rect 2405 28522 2471 28525
rect 4521 28522 4587 28525
rect 2405 28520 4587 28522
rect 2405 28464 2410 28520
rect 2466 28464 4526 28520
rect 4582 28464 4587 28520
rect 2405 28462 4587 28464
rect 2405 28459 2471 28462
rect 4521 28459 4587 28462
rect 3610 28320 3930 28321
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3930 28320
rect 3610 28255 3930 28256
rect 8944 28320 9264 28321
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 28255 9264 28256
rect 14277 28320 14597 28321
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 28255 14597 28256
rect 6277 27776 6597 27777
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 27711 6597 27712
rect 11610 27776 11930 27777
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 27711 11930 27712
rect 3610 27232 3930 27233
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3930 27232
rect 3610 27167 3930 27168
rect 8944 27232 9264 27233
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 27167 9264 27168
rect 14277 27232 14597 27233
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 27167 14597 27168
rect 6277 26688 6597 26689
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 26623 6597 26624
rect 11610 26688 11930 26689
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 26623 11930 26624
rect 3610 26144 3930 26145
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3930 26144
rect 3610 26079 3930 26080
rect 8944 26144 9264 26145
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 26079 9264 26080
rect 14277 26144 14597 26145
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 26079 14597 26080
rect 6277 25600 6597 25601
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 25535 6597 25536
rect 11610 25600 11930 25601
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 25535 11930 25536
rect 4061 25394 4127 25397
rect 9857 25394 9923 25397
rect 4061 25392 9923 25394
rect 4061 25336 4066 25392
rect 4122 25336 9862 25392
rect 9918 25336 9923 25392
rect 4061 25334 9923 25336
rect 4061 25331 4127 25334
rect 9857 25331 9923 25334
rect 2129 25258 2195 25261
rect 4245 25258 4311 25261
rect 2129 25256 4311 25258
rect 2129 25200 2134 25256
rect 2190 25200 4250 25256
rect 4306 25200 4311 25256
rect 2129 25198 4311 25200
rect 2129 25195 2195 25198
rect 4245 25195 4311 25198
rect 12249 25258 12315 25261
rect 12249 25256 14842 25258
rect 12249 25200 12254 25256
rect 12310 25200 14842 25256
rect 12249 25198 14842 25200
rect 12249 25195 12315 25198
rect 3610 25056 3930 25057
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3930 25056
rect 3610 24991 3930 24992
rect 8944 25056 9264 25057
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 24991 9264 24992
rect 14277 25056 14597 25057
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 24991 14597 24992
rect 14782 24986 14842 25198
rect 15520 24986 16000 25016
rect 14782 24926 16000 24986
rect 15520 24896 16000 24926
rect 8017 24714 8083 24717
rect 12065 24714 12131 24717
rect 8017 24712 12131 24714
rect 8017 24656 8022 24712
rect 8078 24656 12070 24712
rect 12126 24656 12131 24712
rect 8017 24654 12131 24656
rect 8017 24651 8083 24654
rect 12065 24651 12131 24654
rect 6277 24512 6597 24513
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 24447 6597 24448
rect 11610 24512 11930 24513
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 24447 11930 24448
rect 3610 23968 3930 23969
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3930 23968
rect 3610 23903 3930 23904
rect 8944 23968 9264 23969
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 23903 9264 23904
rect 14277 23968 14597 23969
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 23903 14597 23904
rect 6821 23490 6887 23493
rect 8753 23490 8819 23493
rect 6821 23488 8819 23490
rect 6821 23432 6826 23488
rect 6882 23432 8758 23488
rect 8814 23432 8819 23488
rect 6821 23430 8819 23432
rect 6821 23427 6887 23430
rect 8753 23427 8819 23430
rect 12065 23490 12131 23493
rect 14181 23490 14247 23493
rect 12065 23488 14247 23490
rect 12065 23432 12070 23488
rect 12126 23432 14186 23488
rect 14242 23432 14247 23488
rect 12065 23430 14247 23432
rect 12065 23427 12131 23430
rect 14181 23427 14247 23430
rect 6277 23424 6597 23425
rect 0 23354 480 23384
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 23359 6597 23360
rect 11610 23424 11930 23425
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 23359 11930 23360
rect 0 23294 6194 23354
rect 0 23264 480 23294
rect 6134 23218 6194 23294
rect 11053 23218 11119 23221
rect 6134 23216 11119 23218
rect 6134 23160 11058 23216
rect 11114 23160 11119 23216
rect 6134 23158 11119 23160
rect 11053 23155 11119 23158
rect 5993 23082 6059 23085
rect 9949 23082 10015 23085
rect 5993 23080 10015 23082
rect 5993 23024 5998 23080
rect 6054 23024 9954 23080
rect 10010 23024 10015 23080
rect 5993 23022 10015 23024
rect 5993 23019 6059 23022
rect 9949 23019 10015 23022
rect 3610 22880 3930 22881
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3930 22880
rect 3610 22815 3930 22816
rect 8944 22880 9264 22881
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 22815 9264 22816
rect 14277 22880 14597 22881
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 22815 14597 22816
rect 7465 22538 7531 22541
rect 9857 22538 9923 22541
rect 7465 22536 9923 22538
rect 7465 22480 7470 22536
rect 7526 22480 9862 22536
rect 9918 22480 9923 22536
rect 7465 22478 9923 22480
rect 7465 22475 7531 22478
rect 9857 22475 9923 22478
rect 6277 22336 6597 22337
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 22271 6597 22272
rect 11610 22336 11930 22337
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 22271 11930 22272
rect 1853 22130 1919 22133
rect 5993 22130 6059 22133
rect 1853 22128 6059 22130
rect 1853 22072 1858 22128
rect 1914 22072 5998 22128
rect 6054 22072 6059 22128
rect 1853 22070 6059 22072
rect 1853 22067 1919 22070
rect 5993 22067 6059 22070
rect 11053 22130 11119 22133
rect 12433 22130 12499 22133
rect 11053 22128 12499 22130
rect 11053 22072 11058 22128
rect 11114 22072 12438 22128
rect 12494 22072 12499 22128
rect 11053 22070 12499 22072
rect 11053 22067 11119 22070
rect 12433 22067 12499 22070
rect 4429 21994 4495 21997
rect 6269 21994 6335 21997
rect 4429 21992 6335 21994
rect 4429 21936 4434 21992
rect 4490 21936 6274 21992
rect 6330 21936 6335 21992
rect 4429 21934 6335 21936
rect 4429 21931 4495 21934
rect 6269 21931 6335 21934
rect 4153 21858 4219 21861
rect 6085 21858 6151 21861
rect 4153 21856 6151 21858
rect 4153 21800 4158 21856
rect 4214 21800 6090 21856
rect 6146 21800 6151 21856
rect 4153 21798 6151 21800
rect 4153 21795 4219 21798
rect 6085 21795 6151 21798
rect 9397 21858 9463 21861
rect 9765 21858 9831 21861
rect 13813 21858 13879 21861
rect 9397 21856 13879 21858
rect 9397 21800 9402 21856
rect 9458 21800 9770 21856
rect 9826 21800 13818 21856
rect 13874 21800 13879 21856
rect 9397 21798 13879 21800
rect 9397 21795 9463 21798
rect 9765 21795 9831 21798
rect 13813 21795 13879 21798
rect 3610 21792 3930 21793
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3930 21792
rect 3610 21727 3930 21728
rect 8944 21792 9264 21793
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 21727 9264 21728
rect 14277 21792 14597 21793
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 21727 14597 21728
rect 6277 21248 6597 21249
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 21183 6597 21184
rect 11610 21248 11930 21249
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 21183 11930 21184
rect 5993 21042 6059 21045
rect 9765 21042 9831 21045
rect 5993 21040 9831 21042
rect 5993 20984 5998 21040
rect 6054 20984 9770 21040
rect 9826 20984 9831 21040
rect 5993 20982 9831 20984
rect 5993 20979 6059 20982
rect 9765 20979 9831 20982
rect 3610 20704 3930 20705
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3930 20704
rect 3610 20639 3930 20640
rect 8944 20704 9264 20705
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 20639 9264 20640
rect 14277 20704 14597 20705
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 20639 14597 20640
rect 5717 20498 5783 20501
rect 7649 20498 7715 20501
rect 10041 20498 10107 20501
rect 5717 20496 10107 20498
rect 5717 20440 5722 20496
rect 5778 20440 7654 20496
rect 7710 20440 10046 20496
rect 10102 20440 10107 20496
rect 5717 20438 10107 20440
rect 5717 20435 5783 20438
rect 7649 20435 7715 20438
rect 10041 20435 10107 20438
rect 7373 20226 7439 20229
rect 11145 20226 11211 20229
rect 7373 20224 11211 20226
rect 7373 20168 7378 20224
rect 7434 20168 11150 20224
rect 11206 20168 11211 20224
rect 7373 20166 11211 20168
rect 7373 20163 7439 20166
rect 11145 20163 11211 20166
rect 6277 20160 6597 20161
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 20095 6597 20096
rect 11610 20160 11930 20161
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 20095 11930 20096
rect 3610 19616 3930 19617
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3930 19616
rect 3610 19551 3930 19552
rect 8944 19616 9264 19617
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 19551 9264 19552
rect 14277 19616 14597 19617
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 19551 14597 19552
rect 6277 19072 6597 19073
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 19007 6597 19008
rect 11610 19072 11930 19073
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 19007 11930 19008
rect 3610 18528 3930 18529
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3930 18528
rect 3610 18463 3930 18464
rect 8944 18528 9264 18529
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 18463 9264 18464
rect 14277 18528 14597 18529
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 18463 14597 18464
rect 6277 17984 6597 17985
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 17919 6597 17920
rect 11610 17984 11930 17985
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 17919 11930 17920
rect 3610 17440 3930 17441
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3930 17440
rect 3610 17375 3930 17376
rect 8944 17440 9264 17441
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 17375 9264 17376
rect 14277 17440 14597 17441
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 17375 14597 17376
rect 2037 17234 2103 17237
rect 12249 17234 12315 17237
rect 2037 17232 12315 17234
rect 2037 17176 2042 17232
rect 2098 17176 12254 17232
rect 12310 17176 12315 17232
rect 2037 17174 12315 17176
rect 2037 17171 2103 17174
rect 12249 17171 12315 17174
rect 6277 16896 6597 16897
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 16831 6597 16832
rect 11610 16896 11930 16897
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 16831 11930 16832
rect 0 16690 480 16720
rect 1577 16690 1643 16693
rect 0 16688 1643 16690
rect 0 16632 1582 16688
rect 1638 16632 1643 16688
rect 0 16630 1643 16632
rect 0 16600 480 16630
rect 1577 16627 1643 16630
rect 8569 16690 8635 16693
rect 11513 16690 11579 16693
rect 8569 16688 11579 16690
rect 8569 16632 8574 16688
rect 8630 16632 11518 16688
rect 11574 16632 11579 16688
rect 8569 16630 11579 16632
rect 8569 16627 8635 16630
rect 11513 16627 11579 16630
rect 3610 16352 3930 16353
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3930 16352
rect 3610 16287 3930 16288
rect 8944 16352 9264 16353
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 16287 9264 16288
rect 14277 16352 14597 16353
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 16287 14597 16288
rect 2313 16146 2379 16149
rect 4797 16146 4863 16149
rect 7189 16146 7255 16149
rect 2313 16144 7255 16146
rect 2313 16088 2318 16144
rect 2374 16088 4802 16144
rect 4858 16088 7194 16144
rect 7250 16088 7255 16144
rect 2313 16086 7255 16088
rect 2313 16083 2379 16086
rect 4797 16083 4863 16086
rect 7189 16083 7255 16086
rect 1945 16010 2011 16013
rect 4337 16010 4403 16013
rect 1945 16008 4403 16010
rect 1945 15952 1950 16008
rect 2006 15952 4342 16008
rect 4398 15952 4403 16008
rect 1945 15950 4403 15952
rect 1945 15947 2011 15950
rect 4337 15947 4403 15950
rect 6277 15808 6597 15809
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 15743 6597 15744
rect 11610 15808 11930 15809
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 15743 11930 15744
rect 4889 15602 4955 15605
rect 6913 15602 6979 15605
rect 4889 15600 6979 15602
rect 4889 15544 4894 15600
rect 4950 15544 6918 15600
rect 6974 15544 6979 15600
rect 4889 15542 6979 15544
rect 4889 15539 4955 15542
rect 6913 15539 6979 15542
rect 5165 15330 5231 15333
rect 7189 15330 7255 15333
rect 5165 15328 7255 15330
rect 5165 15272 5170 15328
rect 5226 15272 7194 15328
rect 7250 15272 7255 15328
rect 5165 15270 7255 15272
rect 5165 15267 5231 15270
rect 7189 15267 7255 15270
rect 3610 15264 3930 15265
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3930 15264
rect 3610 15199 3930 15200
rect 8944 15264 9264 15265
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 15199 9264 15200
rect 14277 15264 14597 15265
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 15199 14597 15200
rect 1669 15058 1735 15061
rect 4337 15058 4403 15061
rect 1669 15056 4403 15058
rect 1669 15000 1674 15056
rect 1730 15000 4342 15056
rect 4398 15000 4403 15056
rect 1669 14998 4403 15000
rect 1669 14995 1735 14998
rect 4337 14995 4403 14998
rect 4797 15058 4863 15061
rect 8385 15058 8451 15061
rect 4797 15056 8451 15058
rect 4797 15000 4802 15056
rect 4858 15000 8390 15056
rect 8446 15000 8451 15056
rect 4797 14998 8451 15000
rect 4797 14995 4863 14998
rect 8385 14995 8451 14998
rect 7557 14922 7623 14925
rect 15520 14922 16000 14952
rect 7557 14920 16000 14922
rect 7557 14864 7562 14920
rect 7618 14864 16000 14920
rect 7557 14862 16000 14864
rect 7557 14859 7623 14862
rect 15520 14832 16000 14862
rect 6277 14720 6597 14721
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 14655 6597 14656
rect 11610 14720 11930 14721
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 14655 11930 14656
rect 8017 14650 8083 14653
rect 8293 14650 8359 14653
rect 9673 14650 9739 14653
rect 8017 14648 9739 14650
rect 8017 14592 8022 14648
rect 8078 14592 8298 14648
rect 8354 14592 9678 14648
rect 9734 14592 9739 14648
rect 8017 14590 9739 14592
rect 8017 14587 8083 14590
rect 8293 14587 8359 14590
rect 9673 14587 9739 14590
rect 4889 14514 4955 14517
rect 9305 14514 9371 14517
rect 4889 14512 9371 14514
rect 4889 14456 4894 14512
rect 4950 14456 9310 14512
rect 9366 14456 9371 14512
rect 4889 14454 9371 14456
rect 4889 14451 4955 14454
rect 9305 14451 9371 14454
rect 3610 14176 3930 14177
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3930 14176
rect 3610 14111 3930 14112
rect 8944 14176 9264 14177
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 14111 9264 14112
rect 14277 14176 14597 14177
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 14111 14597 14112
rect 2037 13970 2103 13973
rect 4797 13970 4863 13973
rect 2037 13968 4863 13970
rect 2037 13912 2042 13968
rect 2098 13912 4802 13968
rect 4858 13912 4863 13968
rect 2037 13910 4863 13912
rect 2037 13907 2103 13910
rect 4797 13907 4863 13910
rect 6277 13632 6597 13633
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 13567 6597 13568
rect 11610 13632 11930 13633
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 13567 11930 13568
rect 3610 13088 3930 13089
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3930 13088
rect 3610 13023 3930 13024
rect 8944 13088 9264 13089
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 13023 9264 13024
rect 14277 13088 14597 13089
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 13023 14597 13024
rect 1393 12746 1459 12749
rect 7925 12746 7991 12749
rect 1393 12744 7991 12746
rect 1393 12688 1398 12744
rect 1454 12688 7930 12744
rect 7986 12688 7991 12744
rect 1393 12686 7991 12688
rect 1393 12683 1459 12686
rect 7925 12683 7991 12686
rect 6277 12544 6597 12545
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 12479 6597 12480
rect 11610 12544 11930 12545
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 12479 11930 12480
rect 3610 12000 3930 12001
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3930 12000
rect 3610 11935 3930 11936
rect 8944 12000 9264 12001
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 11935 9264 11936
rect 14277 12000 14597 12001
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 11935 14597 11936
rect 6277 11456 6597 11457
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 11391 6597 11392
rect 11610 11456 11930 11457
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 11391 11930 11392
rect 3610 10912 3930 10913
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3930 10912
rect 3610 10847 3930 10848
rect 8944 10912 9264 10913
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 10847 9264 10848
rect 14277 10912 14597 10913
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 10847 14597 10848
rect 6277 10368 6597 10369
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 10303 6597 10304
rect 11610 10368 11930 10369
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 10303 11930 10304
rect 0 10026 480 10056
rect 1577 10026 1643 10029
rect 0 10024 1643 10026
rect 0 9968 1582 10024
rect 1638 9968 1643 10024
rect 0 9966 1643 9968
rect 0 9936 480 9966
rect 1577 9963 1643 9966
rect 3610 9824 3930 9825
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3930 9824
rect 3610 9759 3930 9760
rect 8944 9824 9264 9825
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 9759 9264 9760
rect 14277 9824 14597 9825
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 9759 14597 9760
rect 7833 9618 7899 9621
rect 12525 9618 12591 9621
rect 7833 9616 12591 9618
rect 7833 9560 7838 9616
rect 7894 9560 12530 9616
rect 12586 9560 12591 9616
rect 7833 9558 12591 9560
rect 7833 9555 7899 9558
rect 12525 9555 12591 9558
rect 5073 9482 5139 9485
rect 10593 9482 10659 9485
rect 5073 9480 10659 9482
rect 5073 9424 5078 9480
rect 5134 9424 10598 9480
rect 10654 9424 10659 9480
rect 5073 9422 10659 9424
rect 5073 9419 5139 9422
rect 10593 9419 10659 9422
rect 6277 9280 6597 9281
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 9215 6597 9216
rect 11610 9280 11930 9281
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 9215 11930 9216
rect 3509 9074 3575 9077
rect 10133 9074 10199 9077
rect 3509 9072 10199 9074
rect 3509 9016 3514 9072
rect 3570 9016 10138 9072
rect 10194 9016 10199 9072
rect 3509 9014 10199 9016
rect 3509 9011 3575 9014
rect 10133 9011 10199 9014
rect 3610 8736 3930 8737
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3930 8736
rect 3610 8671 3930 8672
rect 8944 8736 9264 8737
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 8671 9264 8672
rect 14277 8736 14597 8737
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 8671 14597 8672
rect 13077 8394 13143 8397
rect 15745 8394 15811 8397
rect 13077 8392 15811 8394
rect 13077 8336 13082 8392
rect 13138 8336 15750 8392
rect 15806 8336 15811 8392
rect 13077 8334 15811 8336
rect 13077 8331 13143 8334
rect 15745 8331 15811 8334
rect 6277 8192 6597 8193
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 8127 6597 8128
rect 11610 8192 11930 8193
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 8127 11930 8128
rect 3610 7648 3930 7649
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3930 7648
rect 3610 7583 3930 7584
rect 8944 7648 9264 7649
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 7583 9264 7584
rect 14277 7648 14597 7649
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 7583 14597 7584
rect 4245 7306 4311 7309
rect 7005 7306 7071 7309
rect 4245 7304 7071 7306
rect 4245 7248 4250 7304
rect 4306 7248 7010 7304
rect 7066 7248 7071 7304
rect 4245 7246 7071 7248
rect 4245 7243 4311 7246
rect 7005 7243 7071 7246
rect 6277 7104 6597 7105
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 7039 6597 7040
rect 11610 7104 11930 7105
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 7039 11930 7040
rect 2681 6898 2747 6901
rect 6177 6898 6243 6901
rect 8845 6898 8911 6901
rect 2681 6896 6243 6898
rect 2681 6840 2686 6896
rect 2742 6840 6182 6896
rect 6238 6840 6243 6896
rect 2681 6838 6243 6840
rect 2681 6835 2747 6838
rect 6177 6835 6243 6838
rect 6318 6896 8911 6898
rect 6318 6840 8850 6896
rect 8906 6840 8911 6896
rect 6318 6838 8911 6840
rect 1577 6762 1643 6765
rect 6318 6762 6378 6838
rect 8845 6835 8911 6838
rect 1577 6760 6378 6762
rect 1577 6704 1582 6760
rect 1638 6704 6378 6760
rect 1577 6702 6378 6704
rect 6821 6762 6887 6765
rect 10409 6762 10475 6765
rect 6821 6760 10475 6762
rect 6821 6704 6826 6760
rect 6882 6704 10414 6760
rect 10470 6704 10475 6760
rect 6821 6702 10475 6704
rect 1577 6699 1643 6702
rect 6821 6699 6887 6702
rect 10409 6699 10475 6702
rect 3610 6560 3930 6561
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3930 6560
rect 3610 6495 3930 6496
rect 8944 6560 9264 6561
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 6495 9264 6496
rect 14277 6560 14597 6561
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 6495 14597 6496
rect 3325 6354 3391 6357
rect 8845 6354 8911 6357
rect 3325 6352 8911 6354
rect 3325 6296 3330 6352
rect 3386 6296 8850 6352
rect 8906 6296 8911 6352
rect 3325 6294 8911 6296
rect 3325 6291 3391 6294
rect 8845 6291 8911 6294
rect 4797 6218 4863 6221
rect 10317 6218 10383 6221
rect 4797 6216 10383 6218
rect 4797 6160 4802 6216
rect 4858 6160 10322 6216
rect 10378 6160 10383 6216
rect 4797 6158 10383 6160
rect 4797 6155 4863 6158
rect 10317 6155 10383 6158
rect 6277 6016 6597 6017
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 5951 6597 5952
rect 11610 6016 11930 6017
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 5951 11930 5952
rect 4889 5810 4955 5813
rect 11329 5810 11395 5813
rect 4889 5808 11395 5810
rect 4889 5752 4894 5808
rect 4950 5752 11334 5808
rect 11390 5752 11395 5808
rect 4889 5750 11395 5752
rect 4889 5747 4955 5750
rect 11329 5747 11395 5750
rect 2589 5674 2655 5677
rect 4337 5674 4403 5677
rect 2589 5672 4403 5674
rect 2589 5616 2594 5672
rect 2650 5616 4342 5672
rect 4398 5616 4403 5672
rect 2589 5614 4403 5616
rect 2589 5611 2655 5614
rect 4337 5611 4403 5614
rect 3610 5472 3930 5473
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3930 5472
rect 3610 5407 3930 5408
rect 8944 5472 9264 5473
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 5407 9264 5408
rect 14277 5472 14597 5473
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 5407 14597 5408
rect 12341 4994 12407 4997
rect 15520 4994 16000 5024
rect 12341 4992 16000 4994
rect 12341 4936 12346 4992
rect 12402 4936 16000 4992
rect 12341 4934 16000 4936
rect 12341 4931 12407 4934
rect 6277 4928 6597 4929
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 4863 6597 4864
rect 11610 4928 11930 4929
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 15520 4904 16000 4934
rect 11610 4863 11930 4864
rect 5717 4722 5783 4725
rect 10593 4722 10659 4725
rect 5717 4720 10659 4722
rect 5717 4664 5722 4720
rect 5778 4664 10598 4720
rect 10654 4664 10659 4720
rect 5717 4662 10659 4664
rect 5717 4659 5783 4662
rect 10593 4659 10659 4662
rect 3610 4384 3930 4385
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3930 4384
rect 3610 4319 3930 4320
rect 8944 4384 9264 4385
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 4319 9264 4320
rect 14277 4384 14597 4385
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 4319 14597 4320
rect 10501 4178 10567 4181
rect 13353 4178 13419 4181
rect 10501 4176 13419 4178
rect 10501 4120 10506 4176
rect 10562 4120 13358 4176
rect 13414 4120 13419 4176
rect 10501 4118 13419 4120
rect 10501 4115 10567 4118
rect 13353 4115 13419 4118
rect 6085 4042 6151 4045
rect 10593 4042 10659 4045
rect 6085 4040 10659 4042
rect 6085 3984 6090 4040
rect 6146 3984 10598 4040
rect 10654 3984 10659 4040
rect 6085 3982 10659 3984
rect 6085 3979 6151 3982
rect 10593 3979 10659 3982
rect 11421 3906 11487 3909
rect 6686 3904 11487 3906
rect 6686 3848 11426 3904
rect 11482 3848 11487 3904
rect 6686 3846 11487 3848
rect 6277 3840 6597 3841
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 3775 6597 3776
rect 4705 3634 4771 3637
rect 6686 3634 6746 3846
rect 11421 3843 11487 3846
rect 11610 3840 11930 3841
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 3775 11930 3776
rect 6913 3770 6979 3773
rect 11145 3770 11211 3773
rect 6913 3768 11211 3770
rect 6913 3712 6918 3768
rect 6974 3712 11150 3768
rect 11206 3712 11211 3768
rect 6913 3710 11211 3712
rect 6913 3707 6979 3710
rect 11145 3707 11211 3710
rect 4705 3632 6746 3634
rect 4705 3576 4710 3632
rect 4766 3576 6746 3632
rect 4705 3574 6746 3576
rect 7741 3634 7807 3637
rect 11605 3634 11671 3637
rect 7741 3632 11671 3634
rect 7741 3576 7746 3632
rect 7802 3576 11610 3632
rect 11666 3576 11671 3632
rect 7741 3574 11671 3576
rect 4705 3571 4771 3574
rect 7741 3571 7807 3574
rect 11605 3571 11671 3574
rect 1669 3498 1735 3501
rect 4429 3498 4495 3501
rect 9949 3498 10015 3501
rect 1669 3496 4354 3498
rect 1669 3440 1674 3496
rect 1730 3440 4354 3496
rect 1669 3438 4354 3440
rect 1669 3435 1735 3438
rect 0 3362 480 3392
rect 1761 3362 1827 3365
rect 0 3360 1827 3362
rect 0 3304 1766 3360
rect 1822 3304 1827 3360
rect 0 3302 1827 3304
rect 4294 3362 4354 3438
rect 4429 3496 10015 3498
rect 4429 3440 4434 3496
rect 4490 3440 9954 3496
rect 10010 3440 10015 3496
rect 4429 3438 10015 3440
rect 4429 3435 4495 3438
rect 9949 3435 10015 3438
rect 10961 3498 11027 3501
rect 13721 3498 13787 3501
rect 10961 3496 13787 3498
rect 10961 3440 10966 3496
rect 11022 3440 13726 3496
rect 13782 3440 13787 3496
rect 10961 3438 13787 3440
rect 10961 3435 11027 3438
rect 13721 3435 13787 3438
rect 8569 3362 8635 3365
rect 4294 3360 8635 3362
rect 4294 3304 8574 3360
rect 8630 3304 8635 3360
rect 4294 3302 8635 3304
rect 0 3272 480 3302
rect 1761 3299 1827 3302
rect 8569 3299 8635 3302
rect 9397 3362 9463 3365
rect 10961 3362 11027 3365
rect 9397 3360 11027 3362
rect 9397 3304 9402 3360
rect 9458 3304 10966 3360
rect 11022 3304 11027 3360
rect 9397 3302 11027 3304
rect 9397 3299 9463 3302
rect 10961 3299 11027 3302
rect 11145 3362 11211 3365
rect 12617 3362 12683 3365
rect 11145 3360 12683 3362
rect 11145 3304 11150 3360
rect 11206 3304 12622 3360
rect 12678 3304 12683 3360
rect 11145 3302 12683 3304
rect 11145 3299 11211 3302
rect 12617 3299 12683 3302
rect 3610 3296 3930 3297
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3930 3296
rect 3610 3231 3930 3232
rect 8944 3296 9264 3297
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 3231 9264 3232
rect 14277 3296 14597 3297
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 3231 14597 3232
rect 10409 3226 10475 3229
rect 13169 3226 13235 3229
rect 10409 3224 13235 3226
rect 10409 3168 10414 3224
rect 10470 3168 13174 3224
rect 13230 3168 13235 3224
rect 10409 3166 13235 3168
rect 10409 3163 10475 3166
rect 13169 3163 13235 3166
rect 6085 3090 6151 3093
rect 11421 3090 11487 3093
rect 6085 3088 11487 3090
rect 6085 3032 6090 3088
rect 6146 3032 11426 3088
rect 11482 3032 11487 3088
rect 6085 3030 11487 3032
rect 6085 3027 6151 3030
rect 11421 3027 11487 3030
rect 11605 3090 11671 3093
rect 12433 3090 12499 3093
rect 11605 3088 12499 3090
rect 11605 3032 11610 3088
rect 11666 3032 12438 3088
rect 12494 3032 12499 3088
rect 11605 3030 12499 3032
rect 11605 3027 11671 3030
rect 12433 3027 12499 3030
rect 5349 2954 5415 2957
rect 8845 2954 8911 2957
rect 12617 2954 12683 2957
rect 5349 2952 8911 2954
rect 5349 2896 5354 2952
rect 5410 2896 8850 2952
rect 8906 2896 8911 2952
rect 5349 2894 8911 2896
rect 5349 2891 5415 2894
rect 8845 2891 8911 2894
rect 9078 2952 12683 2954
rect 9078 2896 12622 2952
rect 12678 2896 12683 2952
rect 9078 2894 12683 2896
rect 2957 2818 3023 2821
rect 5809 2818 5875 2821
rect 2957 2816 5875 2818
rect 2957 2760 2962 2816
rect 3018 2760 5814 2816
rect 5870 2760 5875 2816
rect 2957 2758 5875 2760
rect 2957 2755 3023 2758
rect 5809 2755 5875 2758
rect 7373 2818 7439 2821
rect 9078 2818 9138 2894
rect 12617 2891 12683 2894
rect 7373 2816 9138 2818
rect 7373 2760 7378 2816
rect 7434 2760 9138 2816
rect 7373 2758 9138 2760
rect 13261 2818 13327 2821
rect 15377 2818 15443 2821
rect 13261 2816 15443 2818
rect 13261 2760 13266 2816
rect 13322 2760 15382 2816
rect 15438 2760 15443 2816
rect 13261 2758 15443 2760
rect 7373 2755 7439 2758
rect 13261 2755 13327 2758
rect 15377 2755 15443 2758
rect 6277 2752 6597 2753
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2687 6597 2688
rect 11610 2752 11930 2753
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2687 11930 2688
rect 6729 2682 6795 2685
rect 11421 2682 11487 2685
rect 6729 2680 11487 2682
rect 6729 2624 6734 2680
rect 6790 2624 11426 2680
rect 11482 2624 11487 2680
rect 6729 2622 11487 2624
rect 6729 2619 6795 2622
rect 11421 2619 11487 2622
rect 5257 2546 5323 2549
rect 7097 2546 7163 2549
rect 5257 2544 7163 2546
rect 5257 2488 5262 2544
rect 5318 2488 7102 2544
rect 7158 2488 7163 2544
rect 5257 2486 7163 2488
rect 5257 2483 5323 2486
rect 7097 2483 7163 2486
rect 10409 2546 10475 2549
rect 12893 2546 12959 2549
rect 10409 2544 12959 2546
rect 10409 2488 10414 2544
rect 10470 2488 12898 2544
rect 12954 2488 12959 2544
rect 10409 2486 12959 2488
rect 10409 2483 10475 2486
rect 12893 2483 12959 2486
rect 8109 2410 8175 2413
rect 12801 2410 12867 2413
rect 8109 2408 12867 2410
rect 8109 2352 8114 2408
rect 8170 2352 12806 2408
rect 12862 2352 12867 2408
rect 8109 2350 12867 2352
rect 8109 2347 8175 2350
rect 12801 2347 12867 2350
rect 5441 2274 5507 2277
rect 8753 2274 8819 2277
rect 5441 2272 8819 2274
rect 5441 2216 5446 2272
rect 5502 2216 8758 2272
rect 8814 2216 8819 2272
rect 5441 2214 8819 2216
rect 5441 2211 5507 2214
rect 8753 2211 8819 2214
rect 9397 2274 9463 2277
rect 12525 2274 12591 2277
rect 9397 2272 12591 2274
rect 9397 2216 9402 2272
rect 9458 2216 12530 2272
rect 12586 2216 12591 2272
rect 9397 2214 12591 2216
rect 9397 2211 9463 2214
rect 12525 2211 12591 2214
rect 3610 2208 3930 2209
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3930 2208
rect 3610 2143 3930 2144
rect 8944 2208 9264 2209
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2143 9264 2144
rect 14277 2208 14597 2209
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2143 14597 2144
rect 7557 2002 7623 2005
rect 12985 2002 13051 2005
rect 7557 2000 13051 2002
rect 7557 1944 7562 2000
rect 7618 1944 12990 2000
rect 13046 1944 13051 2000
rect 7557 1942 13051 1944
rect 7557 1939 7623 1942
rect 12985 1939 13051 1942
rect 3509 1866 3575 1869
rect 9397 1866 9463 1869
rect 3509 1864 9463 1866
rect 3509 1808 3514 1864
rect 3570 1808 9402 1864
rect 9458 1808 9463 1864
rect 3509 1806 9463 1808
rect 3509 1803 3575 1806
rect 9397 1803 9463 1806
rect 4981 1458 5047 1461
rect 9949 1458 10015 1461
rect 4981 1456 10015 1458
rect 4981 1400 4986 1456
rect 5042 1400 9954 1456
rect 10010 1400 10015 1456
rect 4981 1398 10015 1400
rect 4981 1395 5047 1398
rect 9949 1395 10015 1398
<< via3 >>
rect 6285 37564 6349 37568
rect 6285 37508 6289 37564
rect 6289 37508 6345 37564
rect 6345 37508 6349 37564
rect 6285 37504 6349 37508
rect 6365 37564 6429 37568
rect 6365 37508 6369 37564
rect 6369 37508 6425 37564
rect 6425 37508 6429 37564
rect 6365 37504 6429 37508
rect 6445 37564 6509 37568
rect 6445 37508 6449 37564
rect 6449 37508 6505 37564
rect 6505 37508 6509 37564
rect 6445 37504 6509 37508
rect 6525 37564 6589 37568
rect 6525 37508 6529 37564
rect 6529 37508 6585 37564
rect 6585 37508 6589 37564
rect 6525 37504 6589 37508
rect 11618 37564 11682 37568
rect 11618 37508 11622 37564
rect 11622 37508 11678 37564
rect 11678 37508 11682 37564
rect 11618 37504 11682 37508
rect 11698 37564 11762 37568
rect 11698 37508 11702 37564
rect 11702 37508 11758 37564
rect 11758 37508 11762 37564
rect 11698 37504 11762 37508
rect 11778 37564 11842 37568
rect 11778 37508 11782 37564
rect 11782 37508 11838 37564
rect 11838 37508 11842 37564
rect 11778 37504 11842 37508
rect 11858 37564 11922 37568
rect 11858 37508 11862 37564
rect 11862 37508 11918 37564
rect 11918 37508 11922 37564
rect 11858 37504 11922 37508
rect 3618 37020 3682 37024
rect 3618 36964 3622 37020
rect 3622 36964 3678 37020
rect 3678 36964 3682 37020
rect 3618 36960 3682 36964
rect 3698 37020 3762 37024
rect 3698 36964 3702 37020
rect 3702 36964 3758 37020
rect 3758 36964 3762 37020
rect 3698 36960 3762 36964
rect 3778 37020 3842 37024
rect 3778 36964 3782 37020
rect 3782 36964 3838 37020
rect 3838 36964 3842 37020
rect 3778 36960 3842 36964
rect 3858 37020 3922 37024
rect 3858 36964 3862 37020
rect 3862 36964 3918 37020
rect 3918 36964 3922 37020
rect 3858 36960 3922 36964
rect 8952 37020 9016 37024
rect 8952 36964 8956 37020
rect 8956 36964 9012 37020
rect 9012 36964 9016 37020
rect 8952 36960 9016 36964
rect 9032 37020 9096 37024
rect 9032 36964 9036 37020
rect 9036 36964 9092 37020
rect 9092 36964 9096 37020
rect 9032 36960 9096 36964
rect 9112 37020 9176 37024
rect 9112 36964 9116 37020
rect 9116 36964 9172 37020
rect 9172 36964 9176 37020
rect 9112 36960 9176 36964
rect 9192 37020 9256 37024
rect 9192 36964 9196 37020
rect 9196 36964 9252 37020
rect 9252 36964 9256 37020
rect 9192 36960 9256 36964
rect 14285 37020 14349 37024
rect 14285 36964 14289 37020
rect 14289 36964 14345 37020
rect 14345 36964 14349 37020
rect 14285 36960 14349 36964
rect 14365 37020 14429 37024
rect 14365 36964 14369 37020
rect 14369 36964 14425 37020
rect 14425 36964 14429 37020
rect 14365 36960 14429 36964
rect 14445 37020 14509 37024
rect 14445 36964 14449 37020
rect 14449 36964 14505 37020
rect 14505 36964 14509 37020
rect 14445 36960 14509 36964
rect 14525 37020 14589 37024
rect 14525 36964 14529 37020
rect 14529 36964 14585 37020
rect 14585 36964 14589 37020
rect 14525 36960 14589 36964
rect 6285 36476 6349 36480
rect 6285 36420 6289 36476
rect 6289 36420 6345 36476
rect 6345 36420 6349 36476
rect 6285 36416 6349 36420
rect 6365 36476 6429 36480
rect 6365 36420 6369 36476
rect 6369 36420 6425 36476
rect 6425 36420 6429 36476
rect 6365 36416 6429 36420
rect 6445 36476 6509 36480
rect 6445 36420 6449 36476
rect 6449 36420 6505 36476
rect 6505 36420 6509 36476
rect 6445 36416 6509 36420
rect 6525 36476 6589 36480
rect 6525 36420 6529 36476
rect 6529 36420 6585 36476
rect 6585 36420 6589 36476
rect 6525 36416 6589 36420
rect 11618 36476 11682 36480
rect 11618 36420 11622 36476
rect 11622 36420 11678 36476
rect 11678 36420 11682 36476
rect 11618 36416 11682 36420
rect 11698 36476 11762 36480
rect 11698 36420 11702 36476
rect 11702 36420 11758 36476
rect 11758 36420 11762 36476
rect 11698 36416 11762 36420
rect 11778 36476 11842 36480
rect 11778 36420 11782 36476
rect 11782 36420 11838 36476
rect 11838 36420 11842 36476
rect 11778 36416 11842 36420
rect 11858 36476 11922 36480
rect 11858 36420 11862 36476
rect 11862 36420 11918 36476
rect 11918 36420 11922 36476
rect 11858 36416 11922 36420
rect 3618 35932 3682 35936
rect 3618 35876 3622 35932
rect 3622 35876 3678 35932
rect 3678 35876 3682 35932
rect 3618 35872 3682 35876
rect 3698 35932 3762 35936
rect 3698 35876 3702 35932
rect 3702 35876 3758 35932
rect 3758 35876 3762 35932
rect 3698 35872 3762 35876
rect 3778 35932 3842 35936
rect 3778 35876 3782 35932
rect 3782 35876 3838 35932
rect 3838 35876 3842 35932
rect 3778 35872 3842 35876
rect 3858 35932 3922 35936
rect 3858 35876 3862 35932
rect 3862 35876 3918 35932
rect 3918 35876 3922 35932
rect 3858 35872 3922 35876
rect 8952 35932 9016 35936
rect 8952 35876 8956 35932
rect 8956 35876 9012 35932
rect 9012 35876 9016 35932
rect 8952 35872 9016 35876
rect 9032 35932 9096 35936
rect 9032 35876 9036 35932
rect 9036 35876 9092 35932
rect 9092 35876 9096 35932
rect 9032 35872 9096 35876
rect 9112 35932 9176 35936
rect 9112 35876 9116 35932
rect 9116 35876 9172 35932
rect 9172 35876 9176 35932
rect 9112 35872 9176 35876
rect 9192 35932 9256 35936
rect 9192 35876 9196 35932
rect 9196 35876 9252 35932
rect 9252 35876 9256 35932
rect 9192 35872 9256 35876
rect 14285 35932 14349 35936
rect 14285 35876 14289 35932
rect 14289 35876 14345 35932
rect 14345 35876 14349 35932
rect 14285 35872 14349 35876
rect 14365 35932 14429 35936
rect 14365 35876 14369 35932
rect 14369 35876 14425 35932
rect 14425 35876 14429 35932
rect 14365 35872 14429 35876
rect 14445 35932 14509 35936
rect 14445 35876 14449 35932
rect 14449 35876 14505 35932
rect 14505 35876 14509 35932
rect 14445 35872 14509 35876
rect 14525 35932 14589 35936
rect 14525 35876 14529 35932
rect 14529 35876 14585 35932
rect 14585 35876 14589 35932
rect 14525 35872 14589 35876
rect 6285 35388 6349 35392
rect 6285 35332 6289 35388
rect 6289 35332 6345 35388
rect 6345 35332 6349 35388
rect 6285 35328 6349 35332
rect 6365 35388 6429 35392
rect 6365 35332 6369 35388
rect 6369 35332 6425 35388
rect 6425 35332 6429 35388
rect 6365 35328 6429 35332
rect 6445 35388 6509 35392
rect 6445 35332 6449 35388
rect 6449 35332 6505 35388
rect 6505 35332 6509 35388
rect 6445 35328 6509 35332
rect 6525 35388 6589 35392
rect 6525 35332 6529 35388
rect 6529 35332 6585 35388
rect 6585 35332 6589 35388
rect 6525 35328 6589 35332
rect 11618 35388 11682 35392
rect 11618 35332 11622 35388
rect 11622 35332 11678 35388
rect 11678 35332 11682 35388
rect 11618 35328 11682 35332
rect 11698 35388 11762 35392
rect 11698 35332 11702 35388
rect 11702 35332 11758 35388
rect 11758 35332 11762 35388
rect 11698 35328 11762 35332
rect 11778 35388 11842 35392
rect 11778 35332 11782 35388
rect 11782 35332 11838 35388
rect 11838 35332 11842 35388
rect 11778 35328 11842 35332
rect 11858 35388 11922 35392
rect 11858 35332 11862 35388
rect 11862 35332 11918 35388
rect 11918 35332 11922 35388
rect 11858 35328 11922 35332
rect 3618 34844 3682 34848
rect 3618 34788 3622 34844
rect 3622 34788 3678 34844
rect 3678 34788 3682 34844
rect 3618 34784 3682 34788
rect 3698 34844 3762 34848
rect 3698 34788 3702 34844
rect 3702 34788 3758 34844
rect 3758 34788 3762 34844
rect 3698 34784 3762 34788
rect 3778 34844 3842 34848
rect 3778 34788 3782 34844
rect 3782 34788 3838 34844
rect 3838 34788 3842 34844
rect 3778 34784 3842 34788
rect 3858 34844 3922 34848
rect 3858 34788 3862 34844
rect 3862 34788 3918 34844
rect 3918 34788 3922 34844
rect 3858 34784 3922 34788
rect 8952 34844 9016 34848
rect 8952 34788 8956 34844
rect 8956 34788 9012 34844
rect 9012 34788 9016 34844
rect 8952 34784 9016 34788
rect 9032 34844 9096 34848
rect 9032 34788 9036 34844
rect 9036 34788 9092 34844
rect 9092 34788 9096 34844
rect 9032 34784 9096 34788
rect 9112 34844 9176 34848
rect 9112 34788 9116 34844
rect 9116 34788 9172 34844
rect 9172 34788 9176 34844
rect 9112 34784 9176 34788
rect 9192 34844 9256 34848
rect 9192 34788 9196 34844
rect 9196 34788 9252 34844
rect 9252 34788 9256 34844
rect 9192 34784 9256 34788
rect 14285 34844 14349 34848
rect 14285 34788 14289 34844
rect 14289 34788 14345 34844
rect 14345 34788 14349 34844
rect 14285 34784 14349 34788
rect 14365 34844 14429 34848
rect 14365 34788 14369 34844
rect 14369 34788 14425 34844
rect 14425 34788 14429 34844
rect 14365 34784 14429 34788
rect 14445 34844 14509 34848
rect 14445 34788 14449 34844
rect 14449 34788 14505 34844
rect 14505 34788 14509 34844
rect 14445 34784 14509 34788
rect 14525 34844 14589 34848
rect 14525 34788 14529 34844
rect 14529 34788 14585 34844
rect 14585 34788 14589 34844
rect 14525 34784 14589 34788
rect 6285 34300 6349 34304
rect 6285 34244 6289 34300
rect 6289 34244 6345 34300
rect 6345 34244 6349 34300
rect 6285 34240 6349 34244
rect 6365 34300 6429 34304
rect 6365 34244 6369 34300
rect 6369 34244 6425 34300
rect 6425 34244 6429 34300
rect 6365 34240 6429 34244
rect 6445 34300 6509 34304
rect 6445 34244 6449 34300
rect 6449 34244 6505 34300
rect 6505 34244 6509 34300
rect 6445 34240 6509 34244
rect 6525 34300 6589 34304
rect 6525 34244 6529 34300
rect 6529 34244 6585 34300
rect 6585 34244 6589 34300
rect 6525 34240 6589 34244
rect 11618 34300 11682 34304
rect 11618 34244 11622 34300
rect 11622 34244 11678 34300
rect 11678 34244 11682 34300
rect 11618 34240 11682 34244
rect 11698 34300 11762 34304
rect 11698 34244 11702 34300
rect 11702 34244 11758 34300
rect 11758 34244 11762 34300
rect 11698 34240 11762 34244
rect 11778 34300 11842 34304
rect 11778 34244 11782 34300
rect 11782 34244 11838 34300
rect 11838 34244 11842 34300
rect 11778 34240 11842 34244
rect 11858 34300 11922 34304
rect 11858 34244 11862 34300
rect 11862 34244 11918 34300
rect 11918 34244 11922 34300
rect 11858 34240 11922 34244
rect 3618 33756 3682 33760
rect 3618 33700 3622 33756
rect 3622 33700 3678 33756
rect 3678 33700 3682 33756
rect 3618 33696 3682 33700
rect 3698 33756 3762 33760
rect 3698 33700 3702 33756
rect 3702 33700 3758 33756
rect 3758 33700 3762 33756
rect 3698 33696 3762 33700
rect 3778 33756 3842 33760
rect 3778 33700 3782 33756
rect 3782 33700 3838 33756
rect 3838 33700 3842 33756
rect 3778 33696 3842 33700
rect 3858 33756 3922 33760
rect 3858 33700 3862 33756
rect 3862 33700 3918 33756
rect 3918 33700 3922 33756
rect 3858 33696 3922 33700
rect 8952 33756 9016 33760
rect 8952 33700 8956 33756
rect 8956 33700 9012 33756
rect 9012 33700 9016 33756
rect 8952 33696 9016 33700
rect 9032 33756 9096 33760
rect 9032 33700 9036 33756
rect 9036 33700 9092 33756
rect 9092 33700 9096 33756
rect 9032 33696 9096 33700
rect 9112 33756 9176 33760
rect 9112 33700 9116 33756
rect 9116 33700 9172 33756
rect 9172 33700 9176 33756
rect 9112 33696 9176 33700
rect 9192 33756 9256 33760
rect 9192 33700 9196 33756
rect 9196 33700 9252 33756
rect 9252 33700 9256 33756
rect 9192 33696 9256 33700
rect 14285 33756 14349 33760
rect 14285 33700 14289 33756
rect 14289 33700 14345 33756
rect 14345 33700 14349 33756
rect 14285 33696 14349 33700
rect 14365 33756 14429 33760
rect 14365 33700 14369 33756
rect 14369 33700 14425 33756
rect 14425 33700 14429 33756
rect 14365 33696 14429 33700
rect 14445 33756 14509 33760
rect 14445 33700 14449 33756
rect 14449 33700 14505 33756
rect 14505 33700 14509 33756
rect 14445 33696 14509 33700
rect 14525 33756 14589 33760
rect 14525 33700 14529 33756
rect 14529 33700 14585 33756
rect 14585 33700 14589 33756
rect 14525 33696 14589 33700
rect 6285 33212 6349 33216
rect 6285 33156 6289 33212
rect 6289 33156 6345 33212
rect 6345 33156 6349 33212
rect 6285 33152 6349 33156
rect 6365 33212 6429 33216
rect 6365 33156 6369 33212
rect 6369 33156 6425 33212
rect 6425 33156 6429 33212
rect 6365 33152 6429 33156
rect 6445 33212 6509 33216
rect 6445 33156 6449 33212
rect 6449 33156 6505 33212
rect 6505 33156 6509 33212
rect 6445 33152 6509 33156
rect 6525 33212 6589 33216
rect 6525 33156 6529 33212
rect 6529 33156 6585 33212
rect 6585 33156 6589 33212
rect 6525 33152 6589 33156
rect 11618 33212 11682 33216
rect 11618 33156 11622 33212
rect 11622 33156 11678 33212
rect 11678 33156 11682 33212
rect 11618 33152 11682 33156
rect 11698 33212 11762 33216
rect 11698 33156 11702 33212
rect 11702 33156 11758 33212
rect 11758 33156 11762 33212
rect 11698 33152 11762 33156
rect 11778 33212 11842 33216
rect 11778 33156 11782 33212
rect 11782 33156 11838 33212
rect 11838 33156 11842 33212
rect 11778 33152 11842 33156
rect 11858 33212 11922 33216
rect 11858 33156 11862 33212
rect 11862 33156 11918 33212
rect 11918 33156 11922 33212
rect 11858 33152 11922 33156
rect 3618 32668 3682 32672
rect 3618 32612 3622 32668
rect 3622 32612 3678 32668
rect 3678 32612 3682 32668
rect 3618 32608 3682 32612
rect 3698 32668 3762 32672
rect 3698 32612 3702 32668
rect 3702 32612 3758 32668
rect 3758 32612 3762 32668
rect 3698 32608 3762 32612
rect 3778 32668 3842 32672
rect 3778 32612 3782 32668
rect 3782 32612 3838 32668
rect 3838 32612 3842 32668
rect 3778 32608 3842 32612
rect 3858 32668 3922 32672
rect 3858 32612 3862 32668
rect 3862 32612 3918 32668
rect 3918 32612 3922 32668
rect 3858 32608 3922 32612
rect 8952 32668 9016 32672
rect 8952 32612 8956 32668
rect 8956 32612 9012 32668
rect 9012 32612 9016 32668
rect 8952 32608 9016 32612
rect 9032 32668 9096 32672
rect 9032 32612 9036 32668
rect 9036 32612 9092 32668
rect 9092 32612 9096 32668
rect 9032 32608 9096 32612
rect 9112 32668 9176 32672
rect 9112 32612 9116 32668
rect 9116 32612 9172 32668
rect 9172 32612 9176 32668
rect 9112 32608 9176 32612
rect 9192 32668 9256 32672
rect 9192 32612 9196 32668
rect 9196 32612 9252 32668
rect 9252 32612 9256 32668
rect 9192 32608 9256 32612
rect 14285 32668 14349 32672
rect 14285 32612 14289 32668
rect 14289 32612 14345 32668
rect 14345 32612 14349 32668
rect 14285 32608 14349 32612
rect 14365 32668 14429 32672
rect 14365 32612 14369 32668
rect 14369 32612 14425 32668
rect 14425 32612 14429 32668
rect 14365 32608 14429 32612
rect 14445 32668 14509 32672
rect 14445 32612 14449 32668
rect 14449 32612 14505 32668
rect 14505 32612 14509 32668
rect 14445 32608 14509 32612
rect 14525 32668 14589 32672
rect 14525 32612 14529 32668
rect 14529 32612 14585 32668
rect 14585 32612 14589 32668
rect 14525 32608 14589 32612
rect 6285 32124 6349 32128
rect 6285 32068 6289 32124
rect 6289 32068 6345 32124
rect 6345 32068 6349 32124
rect 6285 32064 6349 32068
rect 6365 32124 6429 32128
rect 6365 32068 6369 32124
rect 6369 32068 6425 32124
rect 6425 32068 6429 32124
rect 6365 32064 6429 32068
rect 6445 32124 6509 32128
rect 6445 32068 6449 32124
rect 6449 32068 6505 32124
rect 6505 32068 6509 32124
rect 6445 32064 6509 32068
rect 6525 32124 6589 32128
rect 6525 32068 6529 32124
rect 6529 32068 6585 32124
rect 6585 32068 6589 32124
rect 6525 32064 6589 32068
rect 11618 32124 11682 32128
rect 11618 32068 11622 32124
rect 11622 32068 11678 32124
rect 11678 32068 11682 32124
rect 11618 32064 11682 32068
rect 11698 32124 11762 32128
rect 11698 32068 11702 32124
rect 11702 32068 11758 32124
rect 11758 32068 11762 32124
rect 11698 32064 11762 32068
rect 11778 32124 11842 32128
rect 11778 32068 11782 32124
rect 11782 32068 11838 32124
rect 11838 32068 11842 32124
rect 11778 32064 11842 32068
rect 11858 32124 11922 32128
rect 11858 32068 11862 32124
rect 11862 32068 11918 32124
rect 11918 32068 11922 32124
rect 11858 32064 11922 32068
rect 3618 31580 3682 31584
rect 3618 31524 3622 31580
rect 3622 31524 3678 31580
rect 3678 31524 3682 31580
rect 3618 31520 3682 31524
rect 3698 31580 3762 31584
rect 3698 31524 3702 31580
rect 3702 31524 3758 31580
rect 3758 31524 3762 31580
rect 3698 31520 3762 31524
rect 3778 31580 3842 31584
rect 3778 31524 3782 31580
rect 3782 31524 3838 31580
rect 3838 31524 3842 31580
rect 3778 31520 3842 31524
rect 3858 31580 3922 31584
rect 3858 31524 3862 31580
rect 3862 31524 3918 31580
rect 3918 31524 3922 31580
rect 3858 31520 3922 31524
rect 8952 31580 9016 31584
rect 8952 31524 8956 31580
rect 8956 31524 9012 31580
rect 9012 31524 9016 31580
rect 8952 31520 9016 31524
rect 9032 31580 9096 31584
rect 9032 31524 9036 31580
rect 9036 31524 9092 31580
rect 9092 31524 9096 31580
rect 9032 31520 9096 31524
rect 9112 31580 9176 31584
rect 9112 31524 9116 31580
rect 9116 31524 9172 31580
rect 9172 31524 9176 31580
rect 9112 31520 9176 31524
rect 9192 31580 9256 31584
rect 9192 31524 9196 31580
rect 9196 31524 9252 31580
rect 9252 31524 9256 31580
rect 9192 31520 9256 31524
rect 14285 31580 14349 31584
rect 14285 31524 14289 31580
rect 14289 31524 14345 31580
rect 14345 31524 14349 31580
rect 14285 31520 14349 31524
rect 14365 31580 14429 31584
rect 14365 31524 14369 31580
rect 14369 31524 14425 31580
rect 14425 31524 14429 31580
rect 14365 31520 14429 31524
rect 14445 31580 14509 31584
rect 14445 31524 14449 31580
rect 14449 31524 14505 31580
rect 14505 31524 14509 31580
rect 14445 31520 14509 31524
rect 14525 31580 14589 31584
rect 14525 31524 14529 31580
rect 14529 31524 14585 31580
rect 14585 31524 14589 31580
rect 14525 31520 14589 31524
rect 6285 31036 6349 31040
rect 6285 30980 6289 31036
rect 6289 30980 6345 31036
rect 6345 30980 6349 31036
rect 6285 30976 6349 30980
rect 6365 31036 6429 31040
rect 6365 30980 6369 31036
rect 6369 30980 6425 31036
rect 6425 30980 6429 31036
rect 6365 30976 6429 30980
rect 6445 31036 6509 31040
rect 6445 30980 6449 31036
rect 6449 30980 6505 31036
rect 6505 30980 6509 31036
rect 6445 30976 6509 30980
rect 6525 31036 6589 31040
rect 6525 30980 6529 31036
rect 6529 30980 6585 31036
rect 6585 30980 6589 31036
rect 6525 30976 6589 30980
rect 11618 31036 11682 31040
rect 11618 30980 11622 31036
rect 11622 30980 11678 31036
rect 11678 30980 11682 31036
rect 11618 30976 11682 30980
rect 11698 31036 11762 31040
rect 11698 30980 11702 31036
rect 11702 30980 11758 31036
rect 11758 30980 11762 31036
rect 11698 30976 11762 30980
rect 11778 31036 11842 31040
rect 11778 30980 11782 31036
rect 11782 30980 11838 31036
rect 11838 30980 11842 31036
rect 11778 30976 11842 30980
rect 11858 31036 11922 31040
rect 11858 30980 11862 31036
rect 11862 30980 11918 31036
rect 11918 30980 11922 31036
rect 11858 30976 11922 30980
rect 3618 30492 3682 30496
rect 3618 30436 3622 30492
rect 3622 30436 3678 30492
rect 3678 30436 3682 30492
rect 3618 30432 3682 30436
rect 3698 30492 3762 30496
rect 3698 30436 3702 30492
rect 3702 30436 3758 30492
rect 3758 30436 3762 30492
rect 3698 30432 3762 30436
rect 3778 30492 3842 30496
rect 3778 30436 3782 30492
rect 3782 30436 3838 30492
rect 3838 30436 3842 30492
rect 3778 30432 3842 30436
rect 3858 30492 3922 30496
rect 3858 30436 3862 30492
rect 3862 30436 3918 30492
rect 3918 30436 3922 30492
rect 3858 30432 3922 30436
rect 8952 30492 9016 30496
rect 8952 30436 8956 30492
rect 8956 30436 9012 30492
rect 9012 30436 9016 30492
rect 8952 30432 9016 30436
rect 9032 30492 9096 30496
rect 9032 30436 9036 30492
rect 9036 30436 9092 30492
rect 9092 30436 9096 30492
rect 9032 30432 9096 30436
rect 9112 30492 9176 30496
rect 9112 30436 9116 30492
rect 9116 30436 9172 30492
rect 9172 30436 9176 30492
rect 9112 30432 9176 30436
rect 9192 30492 9256 30496
rect 9192 30436 9196 30492
rect 9196 30436 9252 30492
rect 9252 30436 9256 30492
rect 9192 30432 9256 30436
rect 14285 30492 14349 30496
rect 14285 30436 14289 30492
rect 14289 30436 14345 30492
rect 14345 30436 14349 30492
rect 14285 30432 14349 30436
rect 14365 30492 14429 30496
rect 14365 30436 14369 30492
rect 14369 30436 14425 30492
rect 14425 30436 14429 30492
rect 14365 30432 14429 30436
rect 14445 30492 14509 30496
rect 14445 30436 14449 30492
rect 14449 30436 14505 30492
rect 14505 30436 14509 30492
rect 14445 30432 14509 30436
rect 14525 30492 14589 30496
rect 14525 30436 14529 30492
rect 14529 30436 14585 30492
rect 14585 30436 14589 30492
rect 14525 30432 14589 30436
rect 6285 29948 6349 29952
rect 6285 29892 6289 29948
rect 6289 29892 6345 29948
rect 6345 29892 6349 29948
rect 6285 29888 6349 29892
rect 6365 29948 6429 29952
rect 6365 29892 6369 29948
rect 6369 29892 6425 29948
rect 6425 29892 6429 29948
rect 6365 29888 6429 29892
rect 6445 29948 6509 29952
rect 6445 29892 6449 29948
rect 6449 29892 6505 29948
rect 6505 29892 6509 29948
rect 6445 29888 6509 29892
rect 6525 29948 6589 29952
rect 6525 29892 6529 29948
rect 6529 29892 6585 29948
rect 6585 29892 6589 29948
rect 6525 29888 6589 29892
rect 11618 29948 11682 29952
rect 11618 29892 11622 29948
rect 11622 29892 11678 29948
rect 11678 29892 11682 29948
rect 11618 29888 11682 29892
rect 11698 29948 11762 29952
rect 11698 29892 11702 29948
rect 11702 29892 11758 29948
rect 11758 29892 11762 29948
rect 11698 29888 11762 29892
rect 11778 29948 11842 29952
rect 11778 29892 11782 29948
rect 11782 29892 11838 29948
rect 11838 29892 11842 29948
rect 11778 29888 11842 29892
rect 11858 29948 11922 29952
rect 11858 29892 11862 29948
rect 11862 29892 11918 29948
rect 11918 29892 11922 29948
rect 11858 29888 11922 29892
rect 3618 29404 3682 29408
rect 3618 29348 3622 29404
rect 3622 29348 3678 29404
rect 3678 29348 3682 29404
rect 3618 29344 3682 29348
rect 3698 29404 3762 29408
rect 3698 29348 3702 29404
rect 3702 29348 3758 29404
rect 3758 29348 3762 29404
rect 3698 29344 3762 29348
rect 3778 29404 3842 29408
rect 3778 29348 3782 29404
rect 3782 29348 3838 29404
rect 3838 29348 3842 29404
rect 3778 29344 3842 29348
rect 3858 29404 3922 29408
rect 3858 29348 3862 29404
rect 3862 29348 3918 29404
rect 3918 29348 3922 29404
rect 3858 29344 3922 29348
rect 8952 29404 9016 29408
rect 8952 29348 8956 29404
rect 8956 29348 9012 29404
rect 9012 29348 9016 29404
rect 8952 29344 9016 29348
rect 9032 29404 9096 29408
rect 9032 29348 9036 29404
rect 9036 29348 9092 29404
rect 9092 29348 9096 29404
rect 9032 29344 9096 29348
rect 9112 29404 9176 29408
rect 9112 29348 9116 29404
rect 9116 29348 9172 29404
rect 9172 29348 9176 29404
rect 9112 29344 9176 29348
rect 9192 29404 9256 29408
rect 9192 29348 9196 29404
rect 9196 29348 9252 29404
rect 9252 29348 9256 29404
rect 9192 29344 9256 29348
rect 14285 29404 14349 29408
rect 14285 29348 14289 29404
rect 14289 29348 14345 29404
rect 14345 29348 14349 29404
rect 14285 29344 14349 29348
rect 14365 29404 14429 29408
rect 14365 29348 14369 29404
rect 14369 29348 14425 29404
rect 14425 29348 14429 29404
rect 14365 29344 14429 29348
rect 14445 29404 14509 29408
rect 14445 29348 14449 29404
rect 14449 29348 14505 29404
rect 14505 29348 14509 29404
rect 14445 29344 14509 29348
rect 14525 29404 14589 29408
rect 14525 29348 14529 29404
rect 14529 29348 14585 29404
rect 14585 29348 14589 29404
rect 14525 29344 14589 29348
rect 6285 28860 6349 28864
rect 6285 28804 6289 28860
rect 6289 28804 6345 28860
rect 6345 28804 6349 28860
rect 6285 28800 6349 28804
rect 6365 28860 6429 28864
rect 6365 28804 6369 28860
rect 6369 28804 6425 28860
rect 6425 28804 6429 28860
rect 6365 28800 6429 28804
rect 6445 28860 6509 28864
rect 6445 28804 6449 28860
rect 6449 28804 6505 28860
rect 6505 28804 6509 28860
rect 6445 28800 6509 28804
rect 6525 28860 6589 28864
rect 6525 28804 6529 28860
rect 6529 28804 6585 28860
rect 6585 28804 6589 28860
rect 6525 28800 6589 28804
rect 11618 28860 11682 28864
rect 11618 28804 11622 28860
rect 11622 28804 11678 28860
rect 11678 28804 11682 28860
rect 11618 28800 11682 28804
rect 11698 28860 11762 28864
rect 11698 28804 11702 28860
rect 11702 28804 11758 28860
rect 11758 28804 11762 28860
rect 11698 28800 11762 28804
rect 11778 28860 11842 28864
rect 11778 28804 11782 28860
rect 11782 28804 11838 28860
rect 11838 28804 11842 28860
rect 11778 28800 11842 28804
rect 11858 28860 11922 28864
rect 11858 28804 11862 28860
rect 11862 28804 11918 28860
rect 11918 28804 11922 28860
rect 11858 28800 11922 28804
rect 3618 28316 3682 28320
rect 3618 28260 3622 28316
rect 3622 28260 3678 28316
rect 3678 28260 3682 28316
rect 3618 28256 3682 28260
rect 3698 28316 3762 28320
rect 3698 28260 3702 28316
rect 3702 28260 3758 28316
rect 3758 28260 3762 28316
rect 3698 28256 3762 28260
rect 3778 28316 3842 28320
rect 3778 28260 3782 28316
rect 3782 28260 3838 28316
rect 3838 28260 3842 28316
rect 3778 28256 3842 28260
rect 3858 28316 3922 28320
rect 3858 28260 3862 28316
rect 3862 28260 3918 28316
rect 3918 28260 3922 28316
rect 3858 28256 3922 28260
rect 8952 28316 9016 28320
rect 8952 28260 8956 28316
rect 8956 28260 9012 28316
rect 9012 28260 9016 28316
rect 8952 28256 9016 28260
rect 9032 28316 9096 28320
rect 9032 28260 9036 28316
rect 9036 28260 9092 28316
rect 9092 28260 9096 28316
rect 9032 28256 9096 28260
rect 9112 28316 9176 28320
rect 9112 28260 9116 28316
rect 9116 28260 9172 28316
rect 9172 28260 9176 28316
rect 9112 28256 9176 28260
rect 9192 28316 9256 28320
rect 9192 28260 9196 28316
rect 9196 28260 9252 28316
rect 9252 28260 9256 28316
rect 9192 28256 9256 28260
rect 14285 28316 14349 28320
rect 14285 28260 14289 28316
rect 14289 28260 14345 28316
rect 14345 28260 14349 28316
rect 14285 28256 14349 28260
rect 14365 28316 14429 28320
rect 14365 28260 14369 28316
rect 14369 28260 14425 28316
rect 14425 28260 14429 28316
rect 14365 28256 14429 28260
rect 14445 28316 14509 28320
rect 14445 28260 14449 28316
rect 14449 28260 14505 28316
rect 14505 28260 14509 28316
rect 14445 28256 14509 28260
rect 14525 28316 14589 28320
rect 14525 28260 14529 28316
rect 14529 28260 14585 28316
rect 14585 28260 14589 28316
rect 14525 28256 14589 28260
rect 6285 27772 6349 27776
rect 6285 27716 6289 27772
rect 6289 27716 6345 27772
rect 6345 27716 6349 27772
rect 6285 27712 6349 27716
rect 6365 27772 6429 27776
rect 6365 27716 6369 27772
rect 6369 27716 6425 27772
rect 6425 27716 6429 27772
rect 6365 27712 6429 27716
rect 6445 27772 6509 27776
rect 6445 27716 6449 27772
rect 6449 27716 6505 27772
rect 6505 27716 6509 27772
rect 6445 27712 6509 27716
rect 6525 27772 6589 27776
rect 6525 27716 6529 27772
rect 6529 27716 6585 27772
rect 6585 27716 6589 27772
rect 6525 27712 6589 27716
rect 11618 27772 11682 27776
rect 11618 27716 11622 27772
rect 11622 27716 11678 27772
rect 11678 27716 11682 27772
rect 11618 27712 11682 27716
rect 11698 27772 11762 27776
rect 11698 27716 11702 27772
rect 11702 27716 11758 27772
rect 11758 27716 11762 27772
rect 11698 27712 11762 27716
rect 11778 27772 11842 27776
rect 11778 27716 11782 27772
rect 11782 27716 11838 27772
rect 11838 27716 11842 27772
rect 11778 27712 11842 27716
rect 11858 27772 11922 27776
rect 11858 27716 11862 27772
rect 11862 27716 11918 27772
rect 11918 27716 11922 27772
rect 11858 27712 11922 27716
rect 3618 27228 3682 27232
rect 3618 27172 3622 27228
rect 3622 27172 3678 27228
rect 3678 27172 3682 27228
rect 3618 27168 3682 27172
rect 3698 27228 3762 27232
rect 3698 27172 3702 27228
rect 3702 27172 3758 27228
rect 3758 27172 3762 27228
rect 3698 27168 3762 27172
rect 3778 27228 3842 27232
rect 3778 27172 3782 27228
rect 3782 27172 3838 27228
rect 3838 27172 3842 27228
rect 3778 27168 3842 27172
rect 3858 27228 3922 27232
rect 3858 27172 3862 27228
rect 3862 27172 3918 27228
rect 3918 27172 3922 27228
rect 3858 27168 3922 27172
rect 8952 27228 9016 27232
rect 8952 27172 8956 27228
rect 8956 27172 9012 27228
rect 9012 27172 9016 27228
rect 8952 27168 9016 27172
rect 9032 27228 9096 27232
rect 9032 27172 9036 27228
rect 9036 27172 9092 27228
rect 9092 27172 9096 27228
rect 9032 27168 9096 27172
rect 9112 27228 9176 27232
rect 9112 27172 9116 27228
rect 9116 27172 9172 27228
rect 9172 27172 9176 27228
rect 9112 27168 9176 27172
rect 9192 27228 9256 27232
rect 9192 27172 9196 27228
rect 9196 27172 9252 27228
rect 9252 27172 9256 27228
rect 9192 27168 9256 27172
rect 14285 27228 14349 27232
rect 14285 27172 14289 27228
rect 14289 27172 14345 27228
rect 14345 27172 14349 27228
rect 14285 27168 14349 27172
rect 14365 27228 14429 27232
rect 14365 27172 14369 27228
rect 14369 27172 14425 27228
rect 14425 27172 14429 27228
rect 14365 27168 14429 27172
rect 14445 27228 14509 27232
rect 14445 27172 14449 27228
rect 14449 27172 14505 27228
rect 14505 27172 14509 27228
rect 14445 27168 14509 27172
rect 14525 27228 14589 27232
rect 14525 27172 14529 27228
rect 14529 27172 14585 27228
rect 14585 27172 14589 27228
rect 14525 27168 14589 27172
rect 6285 26684 6349 26688
rect 6285 26628 6289 26684
rect 6289 26628 6345 26684
rect 6345 26628 6349 26684
rect 6285 26624 6349 26628
rect 6365 26684 6429 26688
rect 6365 26628 6369 26684
rect 6369 26628 6425 26684
rect 6425 26628 6429 26684
rect 6365 26624 6429 26628
rect 6445 26684 6509 26688
rect 6445 26628 6449 26684
rect 6449 26628 6505 26684
rect 6505 26628 6509 26684
rect 6445 26624 6509 26628
rect 6525 26684 6589 26688
rect 6525 26628 6529 26684
rect 6529 26628 6585 26684
rect 6585 26628 6589 26684
rect 6525 26624 6589 26628
rect 11618 26684 11682 26688
rect 11618 26628 11622 26684
rect 11622 26628 11678 26684
rect 11678 26628 11682 26684
rect 11618 26624 11682 26628
rect 11698 26684 11762 26688
rect 11698 26628 11702 26684
rect 11702 26628 11758 26684
rect 11758 26628 11762 26684
rect 11698 26624 11762 26628
rect 11778 26684 11842 26688
rect 11778 26628 11782 26684
rect 11782 26628 11838 26684
rect 11838 26628 11842 26684
rect 11778 26624 11842 26628
rect 11858 26684 11922 26688
rect 11858 26628 11862 26684
rect 11862 26628 11918 26684
rect 11918 26628 11922 26684
rect 11858 26624 11922 26628
rect 3618 26140 3682 26144
rect 3618 26084 3622 26140
rect 3622 26084 3678 26140
rect 3678 26084 3682 26140
rect 3618 26080 3682 26084
rect 3698 26140 3762 26144
rect 3698 26084 3702 26140
rect 3702 26084 3758 26140
rect 3758 26084 3762 26140
rect 3698 26080 3762 26084
rect 3778 26140 3842 26144
rect 3778 26084 3782 26140
rect 3782 26084 3838 26140
rect 3838 26084 3842 26140
rect 3778 26080 3842 26084
rect 3858 26140 3922 26144
rect 3858 26084 3862 26140
rect 3862 26084 3918 26140
rect 3918 26084 3922 26140
rect 3858 26080 3922 26084
rect 8952 26140 9016 26144
rect 8952 26084 8956 26140
rect 8956 26084 9012 26140
rect 9012 26084 9016 26140
rect 8952 26080 9016 26084
rect 9032 26140 9096 26144
rect 9032 26084 9036 26140
rect 9036 26084 9092 26140
rect 9092 26084 9096 26140
rect 9032 26080 9096 26084
rect 9112 26140 9176 26144
rect 9112 26084 9116 26140
rect 9116 26084 9172 26140
rect 9172 26084 9176 26140
rect 9112 26080 9176 26084
rect 9192 26140 9256 26144
rect 9192 26084 9196 26140
rect 9196 26084 9252 26140
rect 9252 26084 9256 26140
rect 9192 26080 9256 26084
rect 14285 26140 14349 26144
rect 14285 26084 14289 26140
rect 14289 26084 14345 26140
rect 14345 26084 14349 26140
rect 14285 26080 14349 26084
rect 14365 26140 14429 26144
rect 14365 26084 14369 26140
rect 14369 26084 14425 26140
rect 14425 26084 14429 26140
rect 14365 26080 14429 26084
rect 14445 26140 14509 26144
rect 14445 26084 14449 26140
rect 14449 26084 14505 26140
rect 14505 26084 14509 26140
rect 14445 26080 14509 26084
rect 14525 26140 14589 26144
rect 14525 26084 14529 26140
rect 14529 26084 14585 26140
rect 14585 26084 14589 26140
rect 14525 26080 14589 26084
rect 6285 25596 6349 25600
rect 6285 25540 6289 25596
rect 6289 25540 6345 25596
rect 6345 25540 6349 25596
rect 6285 25536 6349 25540
rect 6365 25596 6429 25600
rect 6365 25540 6369 25596
rect 6369 25540 6425 25596
rect 6425 25540 6429 25596
rect 6365 25536 6429 25540
rect 6445 25596 6509 25600
rect 6445 25540 6449 25596
rect 6449 25540 6505 25596
rect 6505 25540 6509 25596
rect 6445 25536 6509 25540
rect 6525 25596 6589 25600
rect 6525 25540 6529 25596
rect 6529 25540 6585 25596
rect 6585 25540 6589 25596
rect 6525 25536 6589 25540
rect 11618 25596 11682 25600
rect 11618 25540 11622 25596
rect 11622 25540 11678 25596
rect 11678 25540 11682 25596
rect 11618 25536 11682 25540
rect 11698 25596 11762 25600
rect 11698 25540 11702 25596
rect 11702 25540 11758 25596
rect 11758 25540 11762 25596
rect 11698 25536 11762 25540
rect 11778 25596 11842 25600
rect 11778 25540 11782 25596
rect 11782 25540 11838 25596
rect 11838 25540 11842 25596
rect 11778 25536 11842 25540
rect 11858 25596 11922 25600
rect 11858 25540 11862 25596
rect 11862 25540 11918 25596
rect 11918 25540 11922 25596
rect 11858 25536 11922 25540
rect 3618 25052 3682 25056
rect 3618 24996 3622 25052
rect 3622 24996 3678 25052
rect 3678 24996 3682 25052
rect 3618 24992 3682 24996
rect 3698 25052 3762 25056
rect 3698 24996 3702 25052
rect 3702 24996 3758 25052
rect 3758 24996 3762 25052
rect 3698 24992 3762 24996
rect 3778 25052 3842 25056
rect 3778 24996 3782 25052
rect 3782 24996 3838 25052
rect 3838 24996 3842 25052
rect 3778 24992 3842 24996
rect 3858 25052 3922 25056
rect 3858 24996 3862 25052
rect 3862 24996 3918 25052
rect 3918 24996 3922 25052
rect 3858 24992 3922 24996
rect 8952 25052 9016 25056
rect 8952 24996 8956 25052
rect 8956 24996 9012 25052
rect 9012 24996 9016 25052
rect 8952 24992 9016 24996
rect 9032 25052 9096 25056
rect 9032 24996 9036 25052
rect 9036 24996 9092 25052
rect 9092 24996 9096 25052
rect 9032 24992 9096 24996
rect 9112 25052 9176 25056
rect 9112 24996 9116 25052
rect 9116 24996 9172 25052
rect 9172 24996 9176 25052
rect 9112 24992 9176 24996
rect 9192 25052 9256 25056
rect 9192 24996 9196 25052
rect 9196 24996 9252 25052
rect 9252 24996 9256 25052
rect 9192 24992 9256 24996
rect 14285 25052 14349 25056
rect 14285 24996 14289 25052
rect 14289 24996 14345 25052
rect 14345 24996 14349 25052
rect 14285 24992 14349 24996
rect 14365 25052 14429 25056
rect 14365 24996 14369 25052
rect 14369 24996 14425 25052
rect 14425 24996 14429 25052
rect 14365 24992 14429 24996
rect 14445 25052 14509 25056
rect 14445 24996 14449 25052
rect 14449 24996 14505 25052
rect 14505 24996 14509 25052
rect 14445 24992 14509 24996
rect 14525 25052 14589 25056
rect 14525 24996 14529 25052
rect 14529 24996 14585 25052
rect 14585 24996 14589 25052
rect 14525 24992 14589 24996
rect 6285 24508 6349 24512
rect 6285 24452 6289 24508
rect 6289 24452 6345 24508
rect 6345 24452 6349 24508
rect 6285 24448 6349 24452
rect 6365 24508 6429 24512
rect 6365 24452 6369 24508
rect 6369 24452 6425 24508
rect 6425 24452 6429 24508
rect 6365 24448 6429 24452
rect 6445 24508 6509 24512
rect 6445 24452 6449 24508
rect 6449 24452 6505 24508
rect 6505 24452 6509 24508
rect 6445 24448 6509 24452
rect 6525 24508 6589 24512
rect 6525 24452 6529 24508
rect 6529 24452 6585 24508
rect 6585 24452 6589 24508
rect 6525 24448 6589 24452
rect 11618 24508 11682 24512
rect 11618 24452 11622 24508
rect 11622 24452 11678 24508
rect 11678 24452 11682 24508
rect 11618 24448 11682 24452
rect 11698 24508 11762 24512
rect 11698 24452 11702 24508
rect 11702 24452 11758 24508
rect 11758 24452 11762 24508
rect 11698 24448 11762 24452
rect 11778 24508 11842 24512
rect 11778 24452 11782 24508
rect 11782 24452 11838 24508
rect 11838 24452 11842 24508
rect 11778 24448 11842 24452
rect 11858 24508 11922 24512
rect 11858 24452 11862 24508
rect 11862 24452 11918 24508
rect 11918 24452 11922 24508
rect 11858 24448 11922 24452
rect 3618 23964 3682 23968
rect 3618 23908 3622 23964
rect 3622 23908 3678 23964
rect 3678 23908 3682 23964
rect 3618 23904 3682 23908
rect 3698 23964 3762 23968
rect 3698 23908 3702 23964
rect 3702 23908 3758 23964
rect 3758 23908 3762 23964
rect 3698 23904 3762 23908
rect 3778 23964 3842 23968
rect 3778 23908 3782 23964
rect 3782 23908 3838 23964
rect 3838 23908 3842 23964
rect 3778 23904 3842 23908
rect 3858 23964 3922 23968
rect 3858 23908 3862 23964
rect 3862 23908 3918 23964
rect 3918 23908 3922 23964
rect 3858 23904 3922 23908
rect 8952 23964 9016 23968
rect 8952 23908 8956 23964
rect 8956 23908 9012 23964
rect 9012 23908 9016 23964
rect 8952 23904 9016 23908
rect 9032 23964 9096 23968
rect 9032 23908 9036 23964
rect 9036 23908 9092 23964
rect 9092 23908 9096 23964
rect 9032 23904 9096 23908
rect 9112 23964 9176 23968
rect 9112 23908 9116 23964
rect 9116 23908 9172 23964
rect 9172 23908 9176 23964
rect 9112 23904 9176 23908
rect 9192 23964 9256 23968
rect 9192 23908 9196 23964
rect 9196 23908 9252 23964
rect 9252 23908 9256 23964
rect 9192 23904 9256 23908
rect 14285 23964 14349 23968
rect 14285 23908 14289 23964
rect 14289 23908 14345 23964
rect 14345 23908 14349 23964
rect 14285 23904 14349 23908
rect 14365 23964 14429 23968
rect 14365 23908 14369 23964
rect 14369 23908 14425 23964
rect 14425 23908 14429 23964
rect 14365 23904 14429 23908
rect 14445 23964 14509 23968
rect 14445 23908 14449 23964
rect 14449 23908 14505 23964
rect 14505 23908 14509 23964
rect 14445 23904 14509 23908
rect 14525 23964 14589 23968
rect 14525 23908 14529 23964
rect 14529 23908 14585 23964
rect 14585 23908 14589 23964
rect 14525 23904 14589 23908
rect 6285 23420 6349 23424
rect 6285 23364 6289 23420
rect 6289 23364 6345 23420
rect 6345 23364 6349 23420
rect 6285 23360 6349 23364
rect 6365 23420 6429 23424
rect 6365 23364 6369 23420
rect 6369 23364 6425 23420
rect 6425 23364 6429 23420
rect 6365 23360 6429 23364
rect 6445 23420 6509 23424
rect 6445 23364 6449 23420
rect 6449 23364 6505 23420
rect 6505 23364 6509 23420
rect 6445 23360 6509 23364
rect 6525 23420 6589 23424
rect 6525 23364 6529 23420
rect 6529 23364 6585 23420
rect 6585 23364 6589 23420
rect 6525 23360 6589 23364
rect 11618 23420 11682 23424
rect 11618 23364 11622 23420
rect 11622 23364 11678 23420
rect 11678 23364 11682 23420
rect 11618 23360 11682 23364
rect 11698 23420 11762 23424
rect 11698 23364 11702 23420
rect 11702 23364 11758 23420
rect 11758 23364 11762 23420
rect 11698 23360 11762 23364
rect 11778 23420 11842 23424
rect 11778 23364 11782 23420
rect 11782 23364 11838 23420
rect 11838 23364 11842 23420
rect 11778 23360 11842 23364
rect 11858 23420 11922 23424
rect 11858 23364 11862 23420
rect 11862 23364 11918 23420
rect 11918 23364 11922 23420
rect 11858 23360 11922 23364
rect 3618 22876 3682 22880
rect 3618 22820 3622 22876
rect 3622 22820 3678 22876
rect 3678 22820 3682 22876
rect 3618 22816 3682 22820
rect 3698 22876 3762 22880
rect 3698 22820 3702 22876
rect 3702 22820 3758 22876
rect 3758 22820 3762 22876
rect 3698 22816 3762 22820
rect 3778 22876 3842 22880
rect 3778 22820 3782 22876
rect 3782 22820 3838 22876
rect 3838 22820 3842 22876
rect 3778 22816 3842 22820
rect 3858 22876 3922 22880
rect 3858 22820 3862 22876
rect 3862 22820 3918 22876
rect 3918 22820 3922 22876
rect 3858 22816 3922 22820
rect 8952 22876 9016 22880
rect 8952 22820 8956 22876
rect 8956 22820 9012 22876
rect 9012 22820 9016 22876
rect 8952 22816 9016 22820
rect 9032 22876 9096 22880
rect 9032 22820 9036 22876
rect 9036 22820 9092 22876
rect 9092 22820 9096 22876
rect 9032 22816 9096 22820
rect 9112 22876 9176 22880
rect 9112 22820 9116 22876
rect 9116 22820 9172 22876
rect 9172 22820 9176 22876
rect 9112 22816 9176 22820
rect 9192 22876 9256 22880
rect 9192 22820 9196 22876
rect 9196 22820 9252 22876
rect 9252 22820 9256 22876
rect 9192 22816 9256 22820
rect 14285 22876 14349 22880
rect 14285 22820 14289 22876
rect 14289 22820 14345 22876
rect 14345 22820 14349 22876
rect 14285 22816 14349 22820
rect 14365 22876 14429 22880
rect 14365 22820 14369 22876
rect 14369 22820 14425 22876
rect 14425 22820 14429 22876
rect 14365 22816 14429 22820
rect 14445 22876 14509 22880
rect 14445 22820 14449 22876
rect 14449 22820 14505 22876
rect 14505 22820 14509 22876
rect 14445 22816 14509 22820
rect 14525 22876 14589 22880
rect 14525 22820 14529 22876
rect 14529 22820 14585 22876
rect 14585 22820 14589 22876
rect 14525 22816 14589 22820
rect 6285 22332 6349 22336
rect 6285 22276 6289 22332
rect 6289 22276 6345 22332
rect 6345 22276 6349 22332
rect 6285 22272 6349 22276
rect 6365 22332 6429 22336
rect 6365 22276 6369 22332
rect 6369 22276 6425 22332
rect 6425 22276 6429 22332
rect 6365 22272 6429 22276
rect 6445 22332 6509 22336
rect 6445 22276 6449 22332
rect 6449 22276 6505 22332
rect 6505 22276 6509 22332
rect 6445 22272 6509 22276
rect 6525 22332 6589 22336
rect 6525 22276 6529 22332
rect 6529 22276 6585 22332
rect 6585 22276 6589 22332
rect 6525 22272 6589 22276
rect 11618 22332 11682 22336
rect 11618 22276 11622 22332
rect 11622 22276 11678 22332
rect 11678 22276 11682 22332
rect 11618 22272 11682 22276
rect 11698 22332 11762 22336
rect 11698 22276 11702 22332
rect 11702 22276 11758 22332
rect 11758 22276 11762 22332
rect 11698 22272 11762 22276
rect 11778 22332 11842 22336
rect 11778 22276 11782 22332
rect 11782 22276 11838 22332
rect 11838 22276 11842 22332
rect 11778 22272 11842 22276
rect 11858 22332 11922 22336
rect 11858 22276 11862 22332
rect 11862 22276 11918 22332
rect 11918 22276 11922 22332
rect 11858 22272 11922 22276
rect 3618 21788 3682 21792
rect 3618 21732 3622 21788
rect 3622 21732 3678 21788
rect 3678 21732 3682 21788
rect 3618 21728 3682 21732
rect 3698 21788 3762 21792
rect 3698 21732 3702 21788
rect 3702 21732 3758 21788
rect 3758 21732 3762 21788
rect 3698 21728 3762 21732
rect 3778 21788 3842 21792
rect 3778 21732 3782 21788
rect 3782 21732 3838 21788
rect 3838 21732 3842 21788
rect 3778 21728 3842 21732
rect 3858 21788 3922 21792
rect 3858 21732 3862 21788
rect 3862 21732 3918 21788
rect 3918 21732 3922 21788
rect 3858 21728 3922 21732
rect 8952 21788 9016 21792
rect 8952 21732 8956 21788
rect 8956 21732 9012 21788
rect 9012 21732 9016 21788
rect 8952 21728 9016 21732
rect 9032 21788 9096 21792
rect 9032 21732 9036 21788
rect 9036 21732 9092 21788
rect 9092 21732 9096 21788
rect 9032 21728 9096 21732
rect 9112 21788 9176 21792
rect 9112 21732 9116 21788
rect 9116 21732 9172 21788
rect 9172 21732 9176 21788
rect 9112 21728 9176 21732
rect 9192 21788 9256 21792
rect 9192 21732 9196 21788
rect 9196 21732 9252 21788
rect 9252 21732 9256 21788
rect 9192 21728 9256 21732
rect 14285 21788 14349 21792
rect 14285 21732 14289 21788
rect 14289 21732 14345 21788
rect 14345 21732 14349 21788
rect 14285 21728 14349 21732
rect 14365 21788 14429 21792
rect 14365 21732 14369 21788
rect 14369 21732 14425 21788
rect 14425 21732 14429 21788
rect 14365 21728 14429 21732
rect 14445 21788 14509 21792
rect 14445 21732 14449 21788
rect 14449 21732 14505 21788
rect 14505 21732 14509 21788
rect 14445 21728 14509 21732
rect 14525 21788 14589 21792
rect 14525 21732 14529 21788
rect 14529 21732 14585 21788
rect 14585 21732 14589 21788
rect 14525 21728 14589 21732
rect 6285 21244 6349 21248
rect 6285 21188 6289 21244
rect 6289 21188 6345 21244
rect 6345 21188 6349 21244
rect 6285 21184 6349 21188
rect 6365 21244 6429 21248
rect 6365 21188 6369 21244
rect 6369 21188 6425 21244
rect 6425 21188 6429 21244
rect 6365 21184 6429 21188
rect 6445 21244 6509 21248
rect 6445 21188 6449 21244
rect 6449 21188 6505 21244
rect 6505 21188 6509 21244
rect 6445 21184 6509 21188
rect 6525 21244 6589 21248
rect 6525 21188 6529 21244
rect 6529 21188 6585 21244
rect 6585 21188 6589 21244
rect 6525 21184 6589 21188
rect 11618 21244 11682 21248
rect 11618 21188 11622 21244
rect 11622 21188 11678 21244
rect 11678 21188 11682 21244
rect 11618 21184 11682 21188
rect 11698 21244 11762 21248
rect 11698 21188 11702 21244
rect 11702 21188 11758 21244
rect 11758 21188 11762 21244
rect 11698 21184 11762 21188
rect 11778 21244 11842 21248
rect 11778 21188 11782 21244
rect 11782 21188 11838 21244
rect 11838 21188 11842 21244
rect 11778 21184 11842 21188
rect 11858 21244 11922 21248
rect 11858 21188 11862 21244
rect 11862 21188 11918 21244
rect 11918 21188 11922 21244
rect 11858 21184 11922 21188
rect 3618 20700 3682 20704
rect 3618 20644 3622 20700
rect 3622 20644 3678 20700
rect 3678 20644 3682 20700
rect 3618 20640 3682 20644
rect 3698 20700 3762 20704
rect 3698 20644 3702 20700
rect 3702 20644 3758 20700
rect 3758 20644 3762 20700
rect 3698 20640 3762 20644
rect 3778 20700 3842 20704
rect 3778 20644 3782 20700
rect 3782 20644 3838 20700
rect 3838 20644 3842 20700
rect 3778 20640 3842 20644
rect 3858 20700 3922 20704
rect 3858 20644 3862 20700
rect 3862 20644 3918 20700
rect 3918 20644 3922 20700
rect 3858 20640 3922 20644
rect 8952 20700 9016 20704
rect 8952 20644 8956 20700
rect 8956 20644 9012 20700
rect 9012 20644 9016 20700
rect 8952 20640 9016 20644
rect 9032 20700 9096 20704
rect 9032 20644 9036 20700
rect 9036 20644 9092 20700
rect 9092 20644 9096 20700
rect 9032 20640 9096 20644
rect 9112 20700 9176 20704
rect 9112 20644 9116 20700
rect 9116 20644 9172 20700
rect 9172 20644 9176 20700
rect 9112 20640 9176 20644
rect 9192 20700 9256 20704
rect 9192 20644 9196 20700
rect 9196 20644 9252 20700
rect 9252 20644 9256 20700
rect 9192 20640 9256 20644
rect 14285 20700 14349 20704
rect 14285 20644 14289 20700
rect 14289 20644 14345 20700
rect 14345 20644 14349 20700
rect 14285 20640 14349 20644
rect 14365 20700 14429 20704
rect 14365 20644 14369 20700
rect 14369 20644 14425 20700
rect 14425 20644 14429 20700
rect 14365 20640 14429 20644
rect 14445 20700 14509 20704
rect 14445 20644 14449 20700
rect 14449 20644 14505 20700
rect 14505 20644 14509 20700
rect 14445 20640 14509 20644
rect 14525 20700 14589 20704
rect 14525 20644 14529 20700
rect 14529 20644 14585 20700
rect 14585 20644 14589 20700
rect 14525 20640 14589 20644
rect 6285 20156 6349 20160
rect 6285 20100 6289 20156
rect 6289 20100 6345 20156
rect 6345 20100 6349 20156
rect 6285 20096 6349 20100
rect 6365 20156 6429 20160
rect 6365 20100 6369 20156
rect 6369 20100 6425 20156
rect 6425 20100 6429 20156
rect 6365 20096 6429 20100
rect 6445 20156 6509 20160
rect 6445 20100 6449 20156
rect 6449 20100 6505 20156
rect 6505 20100 6509 20156
rect 6445 20096 6509 20100
rect 6525 20156 6589 20160
rect 6525 20100 6529 20156
rect 6529 20100 6585 20156
rect 6585 20100 6589 20156
rect 6525 20096 6589 20100
rect 11618 20156 11682 20160
rect 11618 20100 11622 20156
rect 11622 20100 11678 20156
rect 11678 20100 11682 20156
rect 11618 20096 11682 20100
rect 11698 20156 11762 20160
rect 11698 20100 11702 20156
rect 11702 20100 11758 20156
rect 11758 20100 11762 20156
rect 11698 20096 11762 20100
rect 11778 20156 11842 20160
rect 11778 20100 11782 20156
rect 11782 20100 11838 20156
rect 11838 20100 11842 20156
rect 11778 20096 11842 20100
rect 11858 20156 11922 20160
rect 11858 20100 11862 20156
rect 11862 20100 11918 20156
rect 11918 20100 11922 20156
rect 11858 20096 11922 20100
rect 3618 19612 3682 19616
rect 3618 19556 3622 19612
rect 3622 19556 3678 19612
rect 3678 19556 3682 19612
rect 3618 19552 3682 19556
rect 3698 19612 3762 19616
rect 3698 19556 3702 19612
rect 3702 19556 3758 19612
rect 3758 19556 3762 19612
rect 3698 19552 3762 19556
rect 3778 19612 3842 19616
rect 3778 19556 3782 19612
rect 3782 19556 3838 19612
rect 3838 19556 3842 19612
rect 3778 19552 3842 19556
rect 3858 19612 3922 19616
rect 3858 19556 3862 19612
rect 3862 19556 3918 19612
rect 3918 19556 3922 19612
rect 3858 19552 3922 19556
rect 8952 19612 9016 19616
rect 8952 19556 8956 19612
rect 8956 19556 9012 19612
rect 9012 19556 9016 19612
rect 8952 19552 9016 19556
rect 9032 19612 9096 19616
rect 9032 19556 9036 19612
rect 9036 19556 9092 19612
rect 9092 19556 9096 19612
rect 9032 19552 9096 19556
rect 9112 19612 9176 19616
rect 9112 19556 9116 19612
rect 9116 19556 9172 19612
rect 9172 19556 9176 19612
rect 9112 19552 9176 19556
rect 9192 19612 9256 19616
rect 9192 19556 9196 19612
rect 9196 19556 9252 19612
rect 9252 19556 9256 19612
rect 9192 19552 9256 19556
rect 14285 19612 14349 19616
rect 14285 19556 14289 19612
rect 14289 19556 14345 19612
rect 14345 19556 14349 19612
rect 14285 19552 14349 19556
rect 14365 19612 14429 19616
rect 14365 19556 14369 19612
rect 14369 19556 14425 19612
rect 14425 19556 14429 19612
rect 14365 19552 14429 19556
rect 14445 19612 14509 19616
rect 14445 19556 14449 19612
rect 14449 19556 14505 19612
rect 14505 19556 14509 19612
rect 14445 19552 14509 19556
rect 14525 19612 14589 19616
rect 14525 19556 14529 19612
rect 14529 19556 14585 19612
rect 14585 19556 14589 19612
rect 14525 19552 14589 19556
rect 6285 19068 6349 19072
rect 6285 19012 6289 19068
rect 6289 19012 6345 19068
rect 6345 19012 6349 19068
rect 6285 19008 6349 19012
rect 6365 19068 6429 19072
rect 6365 19012 6369 19068
rect 6369 19012 6425 19068
rect 6425 19012 6429 19068
rect 6365 19008 6429 19012
rect 6445 19068 6509 19072
rect 6445 19012 6449 19068
rect 6449 19012 6505 19068
rect 6505 19012 6509 19068
rect 6445 19008 6509 19012
rect 6525 19068 6589 19072
rect 6525 19012 6529 19068
rect 6529 19012 6585 19068
rect 6585 19012 6589 19068
rect 6525 19008 6589 19012
rect 11618 19068 11682 19072
rect 11618 19012 11622 19068
rect 11622 19012 11678 19068
rect 11678 19012 11682 19068
rect 11618 19008 11682 19012
rect 11698 19068 11762 19072
rect 11698 19012 11702 19068
rect 11702 19012 11758 19068
rect 11758 19012 11762 19068
rect 11698 19008 11762 19012
rect 11778 19068 11842 19072
rect 11778 19012 11782 19068
rect 11782 19012 11838 19068
rect 11838 19012 11842 19068
rect 11778 19008 11842 19012
rect 11858 19068 11922 19072
rect 11858 19012 11862 19068
rect 11862 19012 11918 19068
rect 11918 19012 11922 19068
rect 11858 19008 11922 19012
rect 3618 18524 3682 18528
rect 3618 18468 3622 18524
rect 3622 18468 3678 18524
rect 3678 18468 3682 18524
rect 3618 18464 3682 18468
rect 3698 18524 3762 18528
rect 3698 18468 3702 18524
rect 3702 18468 3758 18524
rect 3758 18468 3762 18524
rect 3698 18464 3762 18468
rect 3778 18524 3842 18528
rect 3778 18468 3782 18524
rect 3782 18468 3838 18524
rect 3838 18468 3842 18524
rect 3778 18464 3842 18468
rect 3858 18524 3922 18528
rect 3858 18468 3862 18524
rect 3862 18468 3918 18524
rect 3918 18468 3922 18524
rect 3858 18464 3922 18468
rect 8952 18524 9016 18528
rect 8952 18468 8956 18524
rect 8956 18468 9012 18524
rect 9012 18468 9016 18524
rect 8952 18464 9016 18468
rect 9032 18524 9096 18528
rect 9032 18468 9036 18524
rect 9036 18468 9092 18524
rect 9092 18468 9096 18524
rect 9032 18464 9096 18468
rect 9112 18524 9176 18528
rect 9112 18468 9116 18524
rect 9116 18468 9172 18524
rect 9172 18468 9176 18524
rect 9112 18464 9176 18468
rect 9192 18524 9256 18528
rect 9192 18468 9196 18524
rect 9196 18468 9252 18524
rect 9252 18468 9256 18524
rect 9192 18464 9256 18468
rect 14285 18524 14349 18528
rect 14285 18468 14289 18524
rect 14289 18468 14345 18524
rect 14345 18468 14349 18524
rect 14285 18464 14349 18468
rect 14365 18524 14429 18528
rect 14365 18468 14369 18524
rect 14369 18468 14425 18524
rect 14425 18468 14429 18524
rect 14365 18464 14429 18468
rect 14445 18524 14509 18528
rect 14445 18468 14449 18524
rect 14449 18468 14505 18524
rect 14505 18468 14509 18524
rect 14445 18464 14509 18468
rect 14525 18524 14589 18528
rect 14525 18468 14529 18524
rect 14529 18468 14585 18524
rect 14585 18468 14589 18524
rect 14525 18464 14589 18468
rect 6285 17980 6349 17984
rect 6285 17924 6289 17980
rect 6289 17924 6345 17980
rect 6345 17924 6349 17980
rect 6285 17920 6349 17924
rect 6365 17980 6429 17984
rect 6365 17924 6369 17980
rect 6369 17924 6425 17980
rect 6425 17924 6429 17980
rect 6365 17920 6429 17924
rect 6445 17980 6509 17984
rect 6445 17924 6449 17980
rect 6449 17924 6505 17980
rect 6505 17924 6509 17980
rect 6445 17920 6509 17924
rect 6525 17980 6589 17984
rect 6525 17924 6529 17980
rect 6529 17924 6585 17980
rect 6585 17924 6589 17980
rect 6525 17920 6589 17924
rect 11618 17980 11682 17984
rect 11618 17924 11622 17980
rect 11622 17924 11678 17980
rect 11678 17924 11682 17980
rect 11618 17920 11682 17924
rect 11698 17980 11762 17984
rect 11698 17924 11702 17980
rect 11702 17924 11758 17980
rect 11758 17924 11762 17980
rect 11698 17920 11762 17924
rect 11778 17980 11842 17984
rect 11778 17924 11782 17980
rect 11782 17924 11838 17980
rect 11838 17924 11842 17980
rect 11778 17920 11842 17924
rect 11858 17980 11922 17984
rect 11858 17924 11862 17980
rect 11862 17924 11918 17980
rect 11918 17924 11922 17980
rect 11858 17920 11922 17924
rect 3618 17436 3682 17440
rect 3618 17380 3622 17436
rect 3622 17380 3678 17436
rect 3678 17380 3682 17436
rect 3618 17376 3682 17380
rect 3698 17436 3762 17440
rect 3698 17380 3702 17436
rect 3702 17380 3758 17436
rect 3758 17380 3762 17436
rect 3698 17376 3762 17380
rect 3778 17436 3842 17440
rect 3778 17380 3782 17436
rect 3782 17380 3838 17436
rect 3838 17380 3842 17436
rect 3778 17376 3842 17380
rect 3858 17436 3922 17440
rect 3858 17380 3862 17436
rect 3862 17380 3918 17436
rect 3918 17380 3922 17436
rect 3858 17376 3922 17380
rect 8952 17436 9016 17440
rect 8952 17380 8956 17436
rect 8956 17380 9012 17436
rect 9012 17380 9016 17436
rect 8952 17376 9016 17380
rect 9032 17436 9096 17440
rect 9032 17380 9036 17436
rect 9036 17380 9092 17436
rect 9092 17380 9096 17436
rect 9032 17376 9096 17380
rect 9112 17436 9176 17440
rect 9112 17380 9116 17436
rect 9116 17380 9172 17436
rect 9172 17380 9176 17436
rect 9112 17376 9176 17380
rect 9192 17436 9256 17440
rect 9192 17380 9196 17436
rect 9196 17380 9252 17436
rect 9252 17380 9256 17436
rect 9192 17376 9256 17380
rect 14285 17436 14349 17440
rect 14285 17380 14289 17436
rect 14289 17380 14345 17436
rect 14345 17380 14349 17436
rect 14285 17376 14349 17380
rect 14365 17436 14429 17440
rect 14365 17380 14369 17436
rect 14369 17380 14425 17436
rect 14425 17380 14429 17436
rect 14365 17376 14429 17380
rect 14445 17436 14509 17440
rect 14445 17380 14449 17436
rect 14449 17380 14505 17436
rect 14505 17380 14509 17436
rect 14445 17376 14509 17380
rect 14525 17436 14589 17440
rect 14525 17380 14529 17436
rect 14529 17380 14585 17436
rect 14585 17380 14589 17436
rect 14525 17376 14589 17380
rect 6285 16892 6349 16896
rect 6285 16836 6289 16892
rect 6289 16836 6345 16892
rect 6345 16836 6349 16892
rect 6285 16832 6349 16836
rect 6365 16892 6429 16896
rect 6365 16836 6369 16892
rect 6369 16836 6425 16892
rect 6425 16836 6429 16892
rect 6365 16832 6429 16836
rect 6445 16892 6509 16896
rect 6445 16836 6449 16892
rect 6449 16836 6505 16892
rect 6505 16836 6509 16892
rect 6445 16832 6509 16836
rect 6525 16892 6589 16896
rect 6525 16836 6529 16892
rect 6529 16836 6585 16892
rect 6585 16836 6589 16892
rect 6525 16832 6589 16836
rect 11618 16892 11682 16896
rect 11618 16836 11622 16892
rect 11622 16836 11678 16892
rect 11678 16836 11682 16892
rect 11618 16832 11682 16836
rect 11698 16892 11762 16896
rect 11698 16836 11702 16892
rect 11702 16836 11758 16892
rect 11758 16836 11762 16892
rect 11698 16832 11762 16836
rect 11778 16892 11842 16896
rect 11778 16836 11782 16892
rect 11782 16836 11838 16892
rect 11838 16836 11842 16892
rect 11778 16832 11842 16836
rect 11858 16892 11922 16896
rect 11858 16836 11862 16892
rect 11862 16836 11918 16892
rect 11918 16836 11922 16892
rect 11858 16832 11922 16836
rect 3618 16348 3682 16352
rect 3618 16292 3622 16348
rect 3622 16292 3678 16348
rect 3678 16292 3682 16348
rect 3618 16288 3682 16292
rect 3698 16348 3762 16352
rect 3698 16292 3702 16348
rect 3702 16292 3758 16348
rect 3758 16292 3762 16348
rect 3698 16288 3762 16292
rect 3778 16348 3842 16352
rect 3778 16292 3782 16348
rect 3782 16292 3838 16348
rect 3838 16292 3842 16348
rect 3778 16288 3842 16292
rect 3858 16348 3922 16352
rect 3858 16292 3862 16348
rect 3862 16292 3918 16348
rect 3918 16292 3922 16348
rect 3858 16288 3922 16292
rect 8952 16348 9016 16352
rect 8952 16292 8956 16348
rect 8956 16292 9012 16348
rect 9012 16292 9016 16348
rect 8952 16288 9016 16292
rect 9032 16348 9096 16352
rect 9032 16292 9036 16348
rect 9036 16292 9092 16348
rect 9092 16292 9096 16348
rect 9032 16288 9096 16292
rect 9112 16348 9176 16352
rect 9112 16292 9116 16348
rect 9116 16292 9172 16348
rect 9172 16292 9176 16348
rect 9112 16288 9176 16292
rect 9192 16348 9256 16352
rect 9192 16292 9196 16348
rect 9196 16292 9252 16348
rect 9252 16292 9256 16348
rect 9192 16288 9256 16292
rect 14285 16348 14349 16352
rect 14285 16292 14289 16348
rect 14289 16292 14345 16348
rect 14345 16292 14349 16348
rect 14285 16288 14349 16292
rect 14365 16348 14429 16352
rect 14365 16292 14369 16348
rect 14369 16292 14425 16348
rect 14425 16292 14429 16348
rect 14365 16288 14429 16292
rect 14445 16348 14509 16352
rect 14445 16292 14449 16348
rect 14449 16292 14505 16348
rect 14505 16292 14509 16348
rect 14445 16288 14509 16292
rect 14525 16348 14589 16352
rect 14525 16292 14529 16348
rect 14529 16292 14585 16348
rect 14585 16292 14589 16348
rect 14525 16288 14589 16292
rect 6285 15804 6349 15808
rect 6285 15748 6289 15804
rect 6289 15748 6345 15804
rect 6345 15748 6349 15804
rect 6285 15744 6349 15748
rect 6365 15804 6429 15808
rect 6365 15748 6369 15804
rect 6369 15748 6425 15804
rect 6425 15748 6429 15804
rect 6365 15744 6429 15748
rect 6445 15804 6509 15808
rect 6445 15748 6449 15804
rect 6449 15748 6505 15804
rect 6505 15748 6509 15804
rect 6445 15744 6509 15748
rect 6525 15804 6589 15808
rect 6525 15748 6529 15804
rect 6529 15748 6585 15804
rect 6585 15748 6589 15804
rect 6525 15744 6589 15748
rect 11618 15804 11682 15808
rect 11618 15748 11622 15804
rect 11622 15748 11678 15804
rect 11678 15748 11682 15804
rect 11618 15744 11682 15748
rect 11698 15804 11762 15808
rect 11698 15748 11702 15804
rect 11702 15748 11758 15804
rect 11758 15748 11762 15804
rect 11698 15744 11762 15748
rect 11778 15804 11842 15808
rect 11778 15748 11782 15804
rect 11782 15748 11838 15804
rect 11838 15748 11842 15804
rect 11778 15744 11842 15748
rect 11858 15804 11922 15808
rect 11858 15748 11862 15804
rect 11862 15748 11918 15804
rect 11918 15748 11922 15804
rect 11858 15744 11922 15748
rect 3618 15260 3682 15264
rect 3618 15204 3622 15260
rect 3622 15204 3678 15260
rect 3678 15204 3682 15260
rect 3618 15200 3682 15204
rect 3698 15260 3762 15264
rect 3698 15204 3702 15260
rect 3702 15204 3758 15260
rect 3758 15204 3762 15260
rect 3698 15200 3762 15204
rect 3778 15260 3842 15264
rect 3778 15204 3782 15260
rect 3782 15204 3838 15260
rect 3838 15204 3842 15260
rect 3778 15200 3842 15204
rect 3858 15260 3922 15264
rect 3858 15204 3862 15260
rect 3862 15204 3918 15260
rect 3918 15204 3922 15260
rect 3858 15200 3922 15204
rect 8952 15260 9016 15264
rect 8952 15204 8956 15260
rect 8956 15204 9012 15260
rect 9012 15204 9016 15260
rect 8952 15200 9016 15204
rect 9032 15260 9096 15264
rect 9032 15204 9036 15260
rect 9036 15204 9092 15260
rect 9092 15204 9096 15260
rect 9032 15200 9096 15204
rect 9112 15260 9176 15264
rect 9112 15204 9116 15260
rect 9116 15204 9172 15260
rect 9172 15204 9176 15260
rect 9112 15200 9176 15204
rect 9192 15260 9256 15264
rect 9192 15204 9196 15260
rect 9196 15204 9252 15260
rect 9252 15204 9256 15260
rect 9192 15200 9256 15204
rect 14285 15260 14349 15264
rect 14285 15204 14289 15260
rect 14289 15204 14345 15260
rect 14345 15204 14349 15260
rect 14285 15200 14349 15204
rect 14365 15260 14429 15264
rect 14365 15204 14369 15260
rect 14369 15204 14425 15260
rect 14425 15204 14429 15260
rect 14365 15200 14429 15204
rect 14445 15260 14509 15264
rect 14445 15204 14449 15260
rect 14449 15204 14505 15260
rect 14505 15204 14509 15260
rect 14445 15200 14509 15204
rect 14525 15260 14589 15264
rect 14525 15204 14529 15260
rect 14529 15204 14585 15260
rect 14585 15204 14589 15260
rect 14525 15200 14589 15204
rect 6285 14716 6349 14720
rect 6285 14660 6289 14716
rect 6289 14660 6345 14716
rect 6345 14660 6349 14716
rect 6285 14656 6349 14660
rect 6365 14716 6429 14720
rect 6365 14660 6369 14716
rect 6369 14660 6425 14716
rect 6425 14660 6429 14716
rect 6365 14656 6429 14660
rect 6445 14716 6509 14720
rect 6445 14660 6449 14716
rect 6449 14660 6505 14716
rect 6505 14660 6509 14716
rect 6445 14656 6509 14660
rect 6525 14716 6589 14720
rect 6525 14660 6529 14716
rect 6529 14660 6585 14716
rect 6585 14660 6589 14716
rect 6525 14656 6589 14660
rect 11618 14716 11682 14720
rect 11618 14660 11622 14716
rect 11622 14660 11678 14716
rect 11678 14660 11682 14716
rect 11618 14656 11682 14660
rect 11698 14716 11762 14720
rect 11698 14660 11702 14716
rect 11702 14660 11758 14716
rect 11758 14660 11762 14716
rect 11698 14656 11762 14660
rect 11778 14716 11842 14720
rect 11778 14660 11782 14716
rect 11782 14660 11838 14716
rect 11838 14660 11842 14716
rect 11778 14656 11842 14660
rect 11858 14716 11922 14720
rect 11858 14660 11862 14716
rect 11862 14660 11918 14716
rect 11918 14660 11922 14716
rect 11858 14656 11922 14660
rect 3618 14172 3682 14176
rect 3618 14116 3622 14172
rect 3622 14116 3678 14172
rect 3678 14116 3682 14172
rect 3618 14112 3682 14116
rect 3698 14172 3762 14176
rect 3698 14116 3702 14172
rect 3702 14116 3758 14172
rect 3758 14116 3762 14172
rect 3698 14112 3762 14116
rect 3778 14172 3842 14176
rect 3778 14116 3782 14172
rect 3782 14116 3838 14172
rect 3838 14116 3842 14172
rect 3778 14112 3842 14116
rect 3858 14172 3922 14176
rect 3858 14116 3862 14172
rect 3862 14116 3918 14172
rect 3918 14116 3922 14172
rect 3858 14112 3922 14116
rect 8952 14172 9016 14176
rect 8952 14116 8956 14172
rect 8956 14116 9012 14172
rect 9012 14116 9016 14172
rect 8952 14112 9016 14116
rect 9032 14172 9096 14176
rect 9032 14116 9036 14172
rect 9036 14116 9092 14172
rect 9092 14116 9096 14172
rect 9032 14112 9096 14116
rect 9112 14172 9176 14176
rect 9112 14116 9116 14172
rect 9116 14116 9172 14172
rect 9172 14116 9176 14172
rect 9112 14112 9176 14116
rect 9192 14172 9256 14176
rect 9192 14116 9196 14172
rect 9196 14116 9252 14172
rect 9252 14116 9256 14172
rect 9192 14112 9256 14116
rect 14285 14172 14349 14176
rect 14285 14116 14289 14172
rect 14289 14116 14345 14172
rect 14345 14116 14349 14172
rect 14285 14112 14349 14116
rect 14365 14172 14429 14176
rect 14365 14116 14369 14172
rect 14369 14116 14425 14172
rect 14425 14116 14429 14172
rect 14365 14112 14429 14116
rect 14445 14172 14509 14176
rect 14445 14116 14449 14172
rect 14449 14116 14505 14172
rect 14505 14116 14509 14172
rect 14445 14112 14509 14116
rect 14525 14172 14589 14176
rect 14525 14116 14529 14172
rect 14529 14116 14585 14172
rect 14585 14116 14589 14172
rect 14525 14112 14589 14116
rect 6285 13628 6349 13632
rect 6285 13572 6289 13628
rect 6289 13572 6345 13628
rect 6345 13572 6349 13628
rect 6285 13568 6349 13572
rect 6365 13628 6429 13632
rect 6365 13572 6369 13628
rect 6369 13572 6425 13628
rect 6425 13572 6429 13628
rect 6365 13568 6429 13572
rect 6445 13628 6509 13632
rect 6445 13572 6449 13628
rect 6449 13572 6505 13628
rect 6505 13572 6509 13628
rect 6445 13568 6509 13572
rect 6525 13628 6589 13632
rect 6525 13572 6529 13628
rect 6529 13572 6585 13628
rect 6585 13572 6589 13628
rect 6525 13568 6589 13572
rect 11618 13628 11682 13632
rect 11618 13572 11622 13628
rect 11622 13572 11678 13628
rect 11678 13572 11682 13628
rect 11618 13568 11682 13572
rect 11698 13628 11762 13632
rect 11698 13572 11702 13628
rect 11702 13572 11758 13628
rect 11758 13572 11762 13628
rect 11698 13568 11762 13572
rect 11778 13628 11842 13632
rect 11778 13572 11782 13628
rect 11782 13572 11838 13628
rect 11838 13572 11842 13628
rect 11778 13568 11842 13572
rect 11858 13628 11922 13632
rect 11858 13572 11862 13628
rect 11862 13572 11918 13628
rect 11918 13572 11922 13628
rect 11858 13568 11922 13572
rect 3618 13084 3682 13088
rect 3618 13028 3622 13084
rect 3622 13028 3678 13084
rect 3678 13028 3682 13084
rect 3618 13024 3682 13028
rect 3698 13084 3762 13088
rect 3698 13028 3702 13084
rect 3702 13028 3758 13084
rect 3758 13028 3762 13084
rect 3698 13024 3762 13028
rect 3778 13084 3842 13088
rect 3778 13028 3782 13084
rect 3782 13028 3838 13084
rect 3838 13028 3842 13084
rect 3778 13024 3842 13028
rect 3858 13084 3922 13088
rect 3858 13028 3862 13084
rect 3862 13028 3918 13084
rect 3918 13028 3922 13084
rect 3858 13024 3922 13028
rect 8952 13084 9016 13088
rect 8952 13028 8956 13084
rect 8956 13028 9012 13084
rect 9012 13028 9016 13084
rect 8952 13024 9016 13028
rect 9032 13084 9096 13088
rect 9032 13028 9036 13084
rect 9036 13028 9092 13084
rect 9092 13028 9096 13084
rect 9032 13024 9096 13028
rect 9112 13084 9176 13088
rect 9112 13028 9116 13084
rect 9116 13028 9172 13084
rect 9172 13028 9176 13084
rect 9112 13024 9176 13028
rect 9192 13084 9256 13088
rect 9192 13028 9196 13084
rect 9196 13028 9252 13084
rect 9252 13028 9256 13084
rect 9192 13024 9256 13028
rect 14285 13084 14349 13088
rect 14285 13028 14289 13084
rect 14289 13028 14345 13084
rect 14345 13028 14349 13084
rect 14285 13024 14349 13028
rect 14365 13084 14429 13088
rect 14365 13028 14369 13084
rect 14369 13028 14425 13084
rect 14425 13028 14429 13084
rect 14365 13024 14429 13028
rect 14445 13084 14509 13088
rect 14445 13028 14449 13084
rect 14449 13028 14505 13084
rect 14505 13028 14509 13084
rect 14445 13024 14509 13028
rect 14525 13084 14589 13088
rect 14525 13028 14529 13084
rect 14529 13028 14585 13084
rect 14585 13028 14589 13084
rect 14525 13024 14589 13028
rect 6285 12540 6349 12544
rect 6285 12484 6289 12540
rect 6289 12484 6345 12540
rect 6345 12484 6349 12540
rect 6285 12480 6349 12484
rect 6365 12540 6429 12544
rect 6365 12484 6369 12540
rect 6369 12484 6425 12540
rect 6425 12484 6429 12540
rect 6365 12480 6429 12484
rect 6445 12540 6509 12544
rect 6445 12484 6449 12540
rect 6449 12484 6505 12540
rect 6505 12484 6509 12540
rect 6445 12480 6509 12484
rect 6525 12540 6589 12544
rect 6525 12484 6529 12540
rect 6529 12484 6585 12540
rect 6585 12484 6589 12540
rect 6525 12480 6589 12484
rect 11618 12540 11682 12544
rect 11618 12484 11622 12540
rect 11622 12484 11678 12540
rect 11678 12484 11682 12540
rect 11618 12480 11682 12484
rect 11698 12540 11762 12544
rect 11698 12484 11702 12540
rect 11702 12484 11758 12540
rect 11758 12484 11762 12540
rect 11698 12480 11762 12484
rect 11778 12540 11842 12544
rect 11778 12484 11782 12540
rect 11782 12484 11838 12540
rect 11838 12484 11842 12540
rect 11778 12480 11842 12484
rect 11858 12540 11922 12544
rect 11858 12484 11862 12540
rect 11862 12484 11918 12540
rect 11918 12484 11922 12540
rect 11858 12480 11922 12484
rect 3618 11996 3682 12000
rect 3618 11940 3622 11996
rect 3622 11940 3678 11996
rect 3678 11940 3682 11996
rect 3618 11936 3682 11940
rect 3698 11996 3762 12000
rect 3698 11940 3702 11996
rect 3702 11940 3758 11996
rect 3758 11940 3762 11996
rect 3698 11936 3762 11940
rect 3778 11996 3842 12000
rect 3778 11940 3782 11996
rect 3782 11940 3838 11996
rect 3838 11940 3842 11996
rect 3778 11936 3842 11940
rect 3858 11996 3922 12000
rect 3858 11940 3862 11996
rect 3862 11940 3918 11996
rect 3918 11940 3922 11996
rect 3858 11936 3922 11940
rect 8952 11996 9016 12000
rect 8952 11940 8956 11996
rect 8956 11940 9012 11996
rect 9012 11940 9016 11996
rect 8952 11936 9016 11940
rect 9032 11996 9096 12000
rect 9032 11940 9036 11996
rect 9036 11940 9092 11996
rect 9092 11940 9096 11996
rect 9032 11936 9096 11940
rect 9112 11996 9176 12000
rect 9112 11940 9116 11996
rect 9116 11940 9172 11996
rect 9172 11940 9176 11996
rect 9112 11936 9176 11940
rect 9192 11996 9256 12000
rect 9192 11940 9196 11996
rect 9196 11940 9252 11996
rect 9252 11940 9256 11996
rect 9192 11936 9256 11940
rect 14285 11996 14349 12000
rect 14285 11940 14289 11996
rect 14289 11940 14345 11996
rect 14345 11940 14349 11996
rect 14285 11936 14349 11940
rect 14365 11996 14429 12000
rect 14365 11940 14369 11996
rect 14369 11940 14425 11996
rect 14425 11940 14429 11996
rect 14365 11936 14429 11940
rect 14445 11996 14509 12000
rect 14445 11940 14449 11996
rect 14449 11940 14505 11996
rect 14505 11940 14509 11996
rect 14445 11936 14509 11940
rect 14525 11996 14589 12000
rect 14525 11940 14529 11996
rect 14529 11940 14585 11996
rect 14585 11940 14589 11996
rect 14525 11936 14589 11940
rect 6285 11452 6349 11456
rect 6285 11396 6289 11452
rect 6289 11396 6345 11452
rect 6345 11396 6349 11452
rect 6285 11392 6349 11396
rect 6365 11452 6429 11456
rect 6365 11396 6369 11452
rect 6369 11396 6425 11452
rect 6425 11396 6429 11452
rect 6365 11392 6429 11396
rect 6445 11452 6509 11456
rect 6445 11396 6449 11452
rect 6449 11396 6505 11452
rect 6505 11396 6509 11452
rect 6445 11392 6509 11396
rect 6525 11452 6589 11456
rect 6525 11396 6529 11452
rect 6529 11396 6585 11452
rect 6585 11396 6589 11452
rect 6525 11392 6589 11396
rect 11618 11452 11682 11456
rect 11618 11396 11622 11452
rect 11622 11396 11678 11452
rect 11678 11396 11682 11452
rect 11618 11392 11682 11396
rect 11698 11452 11762 11456
rect 11698 11396 11702 11452
rect 11702 11396 11758 11452
rect 11758 11396 11762 11452
rect 11698 11392 11762 11396
rect 11778 11452 11842 11456
rect 11778 11396 11782 11452
rect 11782 11396 11838 11452
rect 11838 11396 11842 11452
rect 11778 11392 11842 11396
rect 11858 11452 11922 11456
rect 11858 11396 11862 11452
rect 11862 11396 11918 11452
rect 11918 11396 11922 11452
rect 11858 11392 11922 11396
rect 3618 10908 3682 10912
rect 3618 10852 3622 10908
rect 3622 10852 3678 10908
rect 3678 10852 3682 10908
rect 3618 10848 3682 10852
rect 3698 10908 3762 10912
rect 3698 10852 3702 10908
rect 3702 10852 3758 10908
rect 3758 10852 3762 10908
rect 3698 10848 3762 10852
rect 3778 10908 3842 10912
rect 3778 10852 3782 10908
rect 3782 10852 3838 10908
rect 3838 10852 3842 10908
rect 3778 10848 3842 10852
rect 3858 10908 3922 10912
rect 3858 10852 3862 10908
rect 3862 10852 3918 10908
rect 3918 10852 3922 10908
rect 3858 10848 3922 10852
rect 8952 10908 9016 10912
rect 8952 10852 8956 10908
rect 8956 10852 9012 10908
rect 9012 10852 9016 10908
rect 8952 10848 9016 10852
rect 9032 10908 9096 10912
rect 9032 10852 9036 10908
rect 9036 10852 9092 10908
rect 9092 10852 9096 10908
rect 9032 10848 9096 10852
rect 9112 10908 9176 10912
rect 9112 10852 9116 10908
rect 9116 10852 9172 10908
rect 9172 10852 9176 10908
rect 9112 10848 9176 10852
rect 9192 10908 9256 10912
rect 9192 10852 9196 10908
rect 9196 10852 9252 10908
rect 9252 10852 9256 10908
rect 9192 10848 9256 10852
rect 14285 10908 14349 10912
rect 14285 10852 14289 10908
rect 14289 10852 14345 10908
rect 14345 10852 14349 10908
rect 14285 10848 14349 10852
rect 14365 10908 14429 10912
rect 14365 10852 14369 10908
rect 14369 10852 14425 10908
rect 14425 10852 14429 10908
rect 14365 10848 14429 10852
rect 14445 10908 14509 10912
rect 14445 10852 14449 10908
rect 14449 10852 14505 10908
rect 14505 10852 14509 10908
rect 14445 10848 14509 10852
rect 14525 10908 14589 10912
rect 14525 10852 14529 10908
rect 14529 10852 14585 10908
rect 14585 10852 14589 10908
rect 14525 10848 14589 10852
rect 6285 10364 6349 10368
rect 6285 10308 6289 10364
rect 6289 10308 6345 10364
rect 6345 10308 6349 10364
rect 6285 10304 6349 10308
rect 6365 10364 6429 10368
rect 6365 10308 6369 10364
rect 6369 10308 6425 10364
rect 6425 10308 6429 10364
rect 6365 10304 6429 10308
rect 6445 10364 6509 10368
rect 6445 10308 6449 10364
rect 6449 10308 6505 10364
rect 6505 10308 6509 10364
rect 6445 10304 6509 10308
rect 6525 10364 6589 10368
rect 6525 10308 6529 10364
rect 6529 10308 6585 10364
rect 6585 10308 6589 10364
rect 6525 10304 6589 10308
rect 11618 10364 11682 10368
rect 11618 10308 11622 10364
rect 11622 10308 11678 10364
rect 11678 10308 11682 10364
rect 11618 10304 11682 10308
rect 11698 10364 11762 10368
rect 11698 10308 11702 10364
rect 11702 10308 11758 10364
rect 11758 10308 11762 10364
rect 11698 10304 11762 10308
rect 11778 10364 11842 10368
rect 11778 10308 11782 10364
rect 11782 10308 11838 10364
rect 11838 10308 11842 10364
rect 11778 10304 11842 10308
rect 11858 10364 11922 10368
rect 11858 10308 11862 10364
rect 11862 10308 11918 10364
rect 11918 10308 11922 10364
rect 11858 10304 11922 10308
rect 3618 9820 3682 9824
rect 3618 9764 3622 9820
rect 3622 9764 3678 9820
rect 3678 9764 3682 9820
rect 3618 9760 3682 9764
rect 3698 9820 3762 9824
rect 3698 9764 3702 9820
rect 3702 9764 3758 9820
rect 3758 9764 3762 9820
rect 3698 9760 3762 9764
rect 3778 9820 3842 9824
rect 3778 9764 3782 9820
rect 3782 9764 3838 9820
rect 3838 9764 3842 9820
rect 3778 9760 3842 9764
rect 3858 9820 3922 9824
rect 3858 9764 3862 9820
rect 3862 9764 3918 9820
rect 3918 9764 3922 9820
rect 3858 9760 3922 9764
rect 8952 9820 9016 9824
rect 8952 9764 8956 9820
rect 8956 9764 9012 9820
rect 9012 9764 9016 9820
rect 8952 9760 9016 9764
rect 9032 9820 9096 9824
rect 9032 9764 9036 9820
rect 9036 9764 9092 9820
rect 9092 9764 9096 9820
rect 9032 9760 9096 9764
rect 9112 9820 9176 9824
rect 9112 9764 9116 9820
rect 9116 9764 9172 9820
rect 9172 9764 9176 9820
rect 9112 9760 9176 9764
rect 9192 9820 9256 9824
rect 9192 9764 9196 9820
rect 9196 9764 9252 9820
rect 9252 9764 9256 9820
rect 9192 9760 9256 9764
rect 14285 9820 14349 9824
rect 14285 9764 14289 9820
rect 14289 9764 14345 9820
rect 14345 9764 14349 9820
rect 14285 9760 14349 9764
rect 14365 9820 14429 9824
rect 14365 9764 14369 9820
rect 14369 9764 14425 9820
rect 14425 9764 14429 9820
rect 14365 9760 14429 9764
rect 14445 9820 14509 9824
rect 14445 9764 14449 9820
rect 14449 9764 14505 9820
rect 14505 9764 14509 9820
rect 14445 9760 14509 9764
rect 14525 9820 14589 9824
rect 14525 9764 14529 9820
rect 14529 9764 14585 9820
rect 14585 9764 14589 9820
rect 14525 9760 14589 9764
rect 6285 9276 6349 9280
rect 6285 9220 6289 9276
rect 6289 9220 6345 9276
rect 6345 9220 6349 9276
rect 6285 9216 6349 9220
rect 6365 9276 6429 9280
rect 6365 9220 6369 9276
rect 6369 9220 6425 9276
rect 6425 9220 6429 9276
rect 6365 9216 6429 9220
rect 6445 9276 6509 9280
rect 6445 9220 6449 9276
rect 6449 9220 6505 9276
rect 6505 9220 6509 9276
rect 6445 9216 6509 9220
rect 6525 9276 6589 9280
rect 6525 9220 6529 9276
rect 6529 9220 6585 9276
rect 6585 9220 6589 9276
rect 6525 9216 6589 9220
rect 11618 9276 11682 9280
rect 11618 9220 11622 9276
rect 11622 9220 11678 9276
rect 11678 9220 11682 9276
rect 11618 9216 11682 9220
rect 11698 9276 11762 9280
rect 11698 9220 11702 9276
rect 11702 9220 11758 9276
rect 11758 9220 11762 9276
rect 11698 9216 11762 9220
rect 11778 9276 11842 9280
rect 11778 9220 11782 9276
rect 11782 9220 11838 9276
rect 11838 9220 11842 9276
rect 11778 9216 11842 9220
rect 11858 9276 11922 9280
rect 11858 9220 11862 9276
rect 11862 9220 11918 9276
rect 11918 9220 11922 9276
rect 11858 9216 11922 9220
rect 3618 8732 3682 8736
rect 3618 8676 3622 8732
rect 3622 8676 3678 8732
rect 3678 8676 3682 8732
rect 3618 8672 3682 8676
rect 3698 8732 3762 8736
rect 3698 8676 3702 8732
rect 3702 8676 3758 8732
rect 3758 8676 3762 8732
rect 3698 8672 3762 8676
rect 3778 8732 3842 8736
rect 3778 8676 3782 8732
rect 3782 8676 3838 8732
rect 3838 8676 3842 8732
rect 3778 8672 3842 8676
rect 3858 8732 3922 8736
rect 3858 8676 3862 8732
rect 3862 8676 3918 8732
rect 3918 8676 3922 8732
rect 3858 8672 3922 8676
rect 8952 8732 9016 8736
rect 8952 8676 8956 8732
rect 8956 8676 9012 8732
rect 9012 8676 9016 8732
rect 8952 8672 9016 8676
rect 9032 8732 9096 8736
rect 9032 8676 9036 8732
rect 9036 8676 9092 8732
rect 9092 8676 9096 8732
rect 9032 8672 9096 8676
rect 9112 8732 9176 8736
rect 9112 8676 9116 8732
rect 9116 8676 9172 8732
rect 9172 8676 9176 8732
rect 9112 8672 9176 8676
rect 9192 8732 9256 8736
rect 9192 8676 9196 8732
rect 9196 8676 9252 8732
rect 9252 8676 9256 8732
rect 9192 8672 9256 8676
rect 14285 8732 14349 8736
rect 14285 8676 14289 8732
rect 14289 8676 14345 8732
rect 14345 8676 14349 8732
rect 14285 8672 14349 8676
rect 14365 8732 14429 8736
rect 14365 8676 14369 8732
rect 14369 8676 14425 8732
rect 14425 8676 14429 8732
rect 14365 8672 14429 8676
rect 14445 8732 14509 8736
rect 14445 8676 14449 8732
rect 14449 8676 14505 8732
rect 14505 8676 14509 8732
rect 14445 8672 14509 8676
rect 14525 8732 14589 8736
rect 14525 8676 14529 8732
rect 14529 8676 14585 8732
rect 14585 8676 14589 8732
rect 14525 8672 14589 8676
rect 6285 8188 6349 8192
rect 6285 8132 6289 8188
rect 6289 8132 6345 8188
rect 6345 8132 6349 8188
rect 6285 8128 6349 8132
rect 6365 8188 6429 8192
rect 6365 8132 6369 8188
rect 6369 8132 6425 8188
rect 6425 8132 6429 8188
rect 6365 8128 6429 8132
rect 6445 8188 6509 8192
rect 6445 8132 6449 8188
rect 6449 8132 6505 8188
rect 6505 8132 6509 8188
rect 6445 8128 6509 8132
rect 6525 8188 6589 8192
rect 6525 8132 6529 8188
rect 6529 8132 6585 8188
rect 6585 8132 6589 8188
rect 6525 8128 6589 8132
rect 11618 8188 11682 8192
rect 11618 8132 11622 8188
rect 11622 8132 11678 8188
rect 11678 8132 11682 8188
rect 11618 8128 11682 8132
rect 11698 8188 11762 8192
rect 11698 8132 11702 8188
rect 11702 8132 11758 8188
rect 11758 8132 11762 8188
rect 11698 8128 11762 8132
rect 11778 8188 11842 8192
rect 11778 8132 11782 8188
rect 11782 8132 11838 8188
rect 11838 8132 11842 8188
rect 11778 8128 11842 8132
rect 11858 8188 11922 8192
rect 11858 8132 11862 8188
rect 11862 8132 11918 8188
rect 11918 8132 11922 8188
rect 11858 8128 11922 8132
rect 3618 7644 3682 7648
rect 3618 7588 3622 7644
rect 3622 7588 3678 7644
rect 3678 7588 3682 7644
rect 3618 7584 3682 7588
rect 3698 7644 3762 7648
rect 3698 7588 3702 7644
rect 3702 7588 3758 7644
rect 3758 7588 3762 7644
rect 3698 7584 3762 7588
rect 3778 7644 3842 7648
rect 3778 7588 3782 7644
rect 3782 7588 3838 7644
rect 3838 7588 3842 7644
rect 3778 7584 3842 7588
rect 3858 7644 3922 7648
rect 3858 7588 3862 7644
rect 3862 7588 3918 7644
rect 3918 7588 3922 7644
rect 3858 7584 3922 7588
rect 8952 7644 9016 7648
rect 8952 7588 8956 7644
rect 8956 7588 9012 7644
rect 9012 7588 9016 7644
rect 8952 7584 9016 7588
rect 9032 7644 9096 7648
rect 9032 7588 9036 7644
rect 9036 7588 9092 7644
rect 9092 7588 9096 7644
rect 9032 7584 9096 7588
rect 9112 7644 9176 7648
rect 9112 7588 9116 7644
rect 9116 7588 9172 7644
rect 9172 7588 9176 7644
rect 9112 7584 9176 7588
rect 9192 7644 9256 7648
rect 9192 7588 9196 7644
rect 9196 7588 9252 7644
rect 9252 7588 9256 7644
rect 9192 7584 9256 7588
rect 14285 7644 14349 7648
rect 14285 7588 14289 7644
rect 14289 7588 14345 7644
rect 14345 7588 14349 7644
rect 14285 7584 14349 7588
rect 14365 7644 14429 7648
rect 14365 7588 14369 7644
rect 14369 7588 14425 7644
rect 14425 7588 14429 7644
rect 14365 7584 14429 7588
rect 14445 7644 14509 7648
rect 14445 7588 14449 7644
rect 14449 7588 14505 7644
rect 14505 7588 14509 7644
rect 14445 7584 14509 7588
rect 14525 7644 14589 7648
rect 14525 7588 14529 7644
rect 14529 7588 14585 7644
rect 14585 7588 14589 7644
rect 14525 7584 14589 7588
rect 6285 7100 6349 7104
rect 6285 7044 6289 7100
rect 6289 7044 6345 7100
rect 6345 7044 6349 7100
rect 6285 7040 6349 7044
rect 6365 7100 6429 7104
rect 6365 7044 6369 7100
rect 6369 7044 6425 7100
rect 6425 7044 6429 7100
rect 6365 7040 6429 7044
rect 6445 7100 6509 7104
rect 6445 7044 6449 7100
rect 6449 7044 6505 7100
rect 6505 7044 6509 7100
rect 6445 7040 6509 7044
rect 6525 7100 6589 7104
rect 6525 7044 6529 7100
rect 6529 7044 6585 7100
rect 6585 7044 6589 7100
rect 6525 7040 6589 7044
rect 11618 7100 11682 7104
rect 11618 7044 11622 7100
rect 11622 7044 11678 7100
rect 11678 7044 11682 7100
rect 11618 7040 11682 7044
rect 11698 7100 11762 7104
rect 11698 7044 11702 7100
rect 11702 7044 11758 7100
rect 11758 7044 11762 7100
rect 11698 7040 11762 7044
rect 11778 7100 11842 7104
rect 11778 7044 11782 7100
rect 11782 7044 11838 7100
rect 11838 7044 11842 7100
rect 11778 7040 11842 7044
rect 11858 7100 11922 7104
rect 11858 7044 11862 7100
rect 11862 7044 11918 7100
rect 11918 7044 11922 7100
rect 11858 7040 11922 7044
rect 3618 6556 3682 6560
rect 3618 6500 3622 6556
rect 3622 6500 3678 6556
rect 3678 6500 3682 6556
rect 3618 6496 3682 6500
rect 3698 6556 3762 6560
rect 3698 6500 3702 6556
rect 3702 6500 3758 6556
rect 3758 6500 3762 6556
rect 3698 6496 3762 6500
rect 3778 6556 3842 6560
rect 3778 6500 3782 6556
rect 3782 6500 3838 6556
rect 3838 6500 3842 6556
rect 3778 6496 3842 6500
rect 3858 6556 3922 6560
rect 3858 6500 3862 6556
rect 3862 6500 3918 6556
rect 3918 6500 3922 6556
rect 3858 6496 3922 6500
rect 8952 6556 9016 6560
rect 8952 6500 8956 6556
rect 8956 6500 9012 6556
rect 9012 6500 9016 6556
rect 8952 6496 9016 6500
rect 9032 6556 9096 6560
rect 9032 6500 9036 6556
rect 9036 6500 9092 6556
rect 9092 6500 9096 6556
rect 9032 6496 9096 6500
rect 9112 6556 9176 6560
rect 9112 6500 9116 6556
rect 9116 6500 9172 6556
rect 9172 6500 9176 6556
rect 9112 6496 9176 6500
rect 9192 6556 9256 6560
rect 9192 6500 9196 6556
rect 9196 6500 9252 6556
rect 9252 6500 9256 6556
rect 9192 6496 9256 6500
rect 14285 6556 14349 6560
rect 14285 6500 14289 6556
rect 14289 6500 14345 6556
rect 14345 6500 14349 6556
rect 14285 6496 14349 6500
rect 14365 6556 14429 6560
rect 14365 6500 14369 6556
rect 14369 6500 14425 6556
rect 14425 6500 14429 6556
rect 14365 6496 14429 6500
rect 14445 6556 14509 6560
rect 14445 6500 14449 6556
rect 14449 6500 14505 6556
rect 14505 6500 14509 6556
rect 14445 6496 14509 6500
rect 14525 6556 14589 6560
rect 14525 6500 14529 6556
rect 14529 6500 14585 6556
rect 14585 6500 14589 6556
rect 14525 6496 14589 6500
rect 6285 6012 6349 6016
rect 6285 5956 6289 6012
rect 6289 5956 6345 6012
rect 6345 5956 6349 6012
rect 6285 5952 6349 5956
rect 6365 6012 6429 6016
rect 6365 5956 6369 6012
rect 6369 5956 6425 6012
rect 6425 5956 6429 6012
rect 6365 5952 6429 5956
rect 6445 6012 6509 6016
rect 6445 5956 6449 6012
rect 6449 5956 6505 6012
rect 6505 5956 6509 6012
rect 6445 5952 6509 5956
rect 6525 6012 6589 6016
rect 6525 5956 6529 6012
rect 6529 5956 6585 6012
rect 6585 5956 6589 6012
rect 6525 5952 6589 5956
rect 11618 6012 11682 6016
rect 11618 5956 11622 6012
rect 11622 5956 11678 6012
rect 11678 5956 11682 6012
rect 11618 5952 11682 5956
rect 11698 6012 11762 6016
rect 11698 5956 11702 6012
rect 11702 5956 11758 6012
rect 11758 5956 11762 6012
rect 11698 5952 11762 5956
rect 11778 6012 11842 6016
rect 11778 5956 11782 6012
rect 11782 5956 11838 6012
rect 11838 5956 11842 6012
rect 11778 5952 11842 5956
rect 11858 6012 11922 6016
rect 11858 5956 11862 6012
rect 11862 5956 11918 6012
rect 11918 5956 11922 6012
rect 11858 5952 11922 5956
rect 3618 5468 3682 5472
rect 3618 5412 3622 5468
rect 3622 5412 3678 5468
rect 3678 5412 3682 5468
rect 3618 5408 3682 5412
rect 3698 5468 3762 5472
rect 3698 5412 3702 5468
rect 3702 5412 3758 5468
rect 3758 5412 3762 5468
rect 3698 5408 3762 5412
rect 3778 5468 3842 5472
rect 3778 5412 3782 5468
rect 3782 5412 3838 5468
rect 3838 5412 3842 5468
rect 3778 5408 3842 5412
rect 3858 5468 3922 5472
rect 3858 5412 3862 5468
rect 3862 5412 3918 5468
rect 3918 5412 3922 5468
rect 3858 5408 3922 5412
rect 8952 5468 9016 5472
rect 8952 5412 8956 5468
rect 8956 5412 9012 5468
rect 9012 5412 9016 5468
rect 8952 5408 9016 5412
rect 9032 5468 9096 5472
rect 9032 5412 9036 5468
rect 9036 5412 9092 5468
rect 9092 5412 9096 5468
rect 9032 5408 9096 5412
rect 9112 5468 9176 5472
rect 9112 5412 9116 5468
rect 9116 5412 9172 5468
rect 9172 5412 9176 5468
rect 9112 5408 9176 5412
rect 9192 5468 9256 5472
rect 9192 5412 9196 5468
rect 9196 5412 9252 5468
rect 9252 5412 9256 5468
rect 9192 5408 9256 5412
rect 14285 5468 14349 5472
rect 14285 5412 14289 5468
rect 14289 5412 14345 5468
rect 14345 5412 14349 5468
rect 14285 5408 14349 5412
rect 14365 5468 14429 5472
rect 14365 5412 14369 5468
rect 14369 5412 14425 5468
rect 14425 5412 14429 5468
rect 14365 5408 14429 5412
rect 14445 5468 14509 5472
rect 14445 5412 14449 5468
rect 14449 5412 14505 5468
rect 14505 5412 14509 5468
rect 14445 5408 14509 5412
rect 14525 5468 14589 5472
rect 14525 5412 14529 5468
rect 14529 5412 14585 5468
rect 14585 5412 14589 5468
rect 14525 5408 14589 5412
rect 6285 4924 6349 4928
rect 6285 4868 6289 4924
rect 6289 4868 6345 4924
rect 6345 4868 6349 4924
rect 6285 4864 6349 4868
rect 6365 4924 6429 4928
rect 6365 4868 6369 4924
rect 6369 4868 6425 4924
rect 6425 4868 6429 4924
rect 6365 4864 6429 4868
rect 6445 4924 6509 4928
rect 6445 4868 6449 4924
rect 6449 4868 6505 4924
rect 6505 4868 6509 4924
rect 6445 4864 6509 4868
rect 6525 4924 6589 4928
rect 6525 4868 6529 4924
rect 6529 4868 6585 4924
rect 6585 4868 6589 4924
rect 6525 4864 6589 4868
rect 11618 4924 11682 4928
rect 11618 4868 11622 4924
rect 11622 4868 11678 4924
rect 11678 4868 11682 4924
rect 11618 4864 11682 4868
rect 11698 4924 11762 4928
rect 11698 4868 11702 4924
rect 11702 4868 11758 4924
rect 11758 4868 11762 4924
rect 11698 4864 11762 4868
rect 11778 4924 11842 4928
rect 11778 4868 11782 4924
rect 11782 4868 11838 4924
rect 11838 4868 11842 4924
rect 11778 4864 11842 4868
rect 11858 4924 11922 4928
rect 11858 4868 11862 4924
rect 11862 4868 11918 4924
rect 11918 4868 11922 4924
rect 11858 4864 11922 4868
rect 3618 4380 3682 4384
rect 3618 4324 3622 4380
rect 3622 4324 3678 4380
rect 3678 4324 3682 4380
rect 3618 4320 3682 4324
rect 3698 4380 3762 4384
rect 3698 4324 3702 4380
rect 3702 4324 3758 4380
rect 3758 4324 3762 4380
rect 3698 4320 3762 4324
rect 3778 4380 3842 4384
rect 3778 4324 3782 4380
rect 3782 4324 3838 4380
rect 3838 4324 3842 4380
rect 3778 4320 3842 4324
rect 3858 4380 3922 4384
rect 3858 4324 3862 4380
rect 3862 4324 3918 4380
rect 3918 4324 3922 4380
rect 3858 4320 3922 4324
rect 8952 4380 9016 4384
rect 8952 4324 8956 4380
rect 8956 4324 9012 4380
rect 9012 4324 9016 4380
rect 8952 4320 9016 4324
rect 9032 4380 9096 4384
rect 9032 4324 9036 4380
rect 9036 4324 9092 4380
rect 9092 4324 9096 4380
rect 9032 4320 9096 4324
rect 9112 4380 9176 4384
rect 9112 4324 9116 4380
rect 9116 4324 9172 4380
rect 9172 4324 9176 4380
rect 9112 4320 9176 4324
rect 9192 4380 9256 4384
rect 9192 4324 9196 4380
rect 9196 4324 9252 4380
rect 9252 4324 9256 4380
rect 9192 4320 9256 4324
rect 14285 4380 14349 4384
rect 14285 4324 14289 4380
rect 14289 4324 14345 4380
rect 14345 4324 14349 4380
rect 14285 4320 14349 4324
rect 14365 4380 14429 4384
rect 14365 4324 14369 4380
rect 14369 4324 14425 4380
rect 14425 4324 14429 4380
rect 14365 4320 14429 4324
rect 14445 4380 14509 4384
rect 14445 4324 14449 4380
rect 14449 4324 14505 4380
rect 14505 4324 14509 4380
rect 14445 4320 14509 4324
rect 14525 4380 14589 4384
rect 14525 4324 14529 4380
rect 14529 4324 14585 4380
rect 14585 4324 14589 4380
rect 14525 4320 14589 4324
rect 6285 3836 6349 3840
rect 6285 3780 6289 3836
rect 6289 3780 6345 3836
rect 6345 3780 6349 3836
rect 6285 3776 6349 3780
rect 6365 3836 6429 3840
rect 6365 3780 6369 3836
rect 6369 3780 6425 3836
rect 6425 3780 6429 3836
rect 6365 3776 6429 3780
rect 6445 3836 6509 3840
rect 6445 3780 6449 3836
rect 6449 3780 6505 3836
rect 6505 3780 6509 3836
rect 6445 3776 6509 3780
rect 6525 3836 6589 3840
rect 6525 3780 6529 3836
rect 6529 3780 6585 3836
rect 6585 3780 6589 3836
rect 6525 3776 6589 3780
rect 11618 3836 11682 3840
rect 11618 3780 11622 3836
rect 11622 3780 11678 3836
rect 11678 3780 11682 3836
rect 11618 3776 11682 3780
rect 11698 3836 11762 3840
rect 11698 3780 11702 3836
rect 11702 3780 11758 3836
rect 11758 3780 11762 3836
rect 11698 3776 11762 3780
rect 11778 3836 11842 3840
rect 11778 3780 11782 3836
rect 11782 3780 11838 3836
rect 11838 3780 11842 3836
rect 11778 3776 11842 3780
rect 11858 3836 11922 3840
rect 11858 3780 11862 3836
rect 11862 3780 11918 3836
rect 11918 3780 11922 3836
rect 11858 3776 11922 3780
rect 3618 3292 3682 3296
rect 3618 3236 3622 3292
rect 3622 3236 3678 3292
rect 3678 3236 3682 3292
rect 3618 3232 3682 3236
rect 3698 3292 3762 3296
rect 3698 3236 3702 3292
rect 3702 3236 3758 3292
rect 3758 3236 3762 3292
rect 3698 3232 3762 3236
rect 3778 3292 3842 3296
rect 3778 3236 3782 3292
rect 3782 3236 3838 3292
rect 3838 3236 3842 3292
rect 3778 3232 3842 3236
rect 3858 3292 3922 3296
rect 3858 3236 3862 3292
rect 3862 3236 3918 3292
rect 3918 3236 3922 3292
rect 3858 3232 3922 3236
rect 8952 3292 9016 3296
rect 8952 3236 8956 3292
rect 8956 3236 9012 3292
rect 9012 3236 9016 3292
rect 8952 3232 9016 3236
rect 9032 3292 9096 3296
rect 9032 3236 9036 3292
rect 9036 3236 9092 3292
rect 9092 3236 9096 3292
rect 9032 3232 9096 3236
rect 9112 3292 9176 3296
rect 9112 3236 9116 3292
rect 9116 3236 9172 3292
rect 9172 3236 9176 3292
rect 9112 3232 9176 3236
rect 9192 3292 9256 3296
rect 9192 3236 9196 3292
rect 9196 3236 9252 3292
rect 9252 3236 9256 3292
rect 9192 3232 9256 3236
rect 14285 3292 14349 3296
rect 14285 3236 14289 3292
rect 14289 3236 14345 3292
rect 14345 3236 14349 3292
rect 14285 3232 14349 3236
rect 14365 3292 14429 3296
rect 14365 3236 14369 3292
rect 14369 3236 14425 3292
rect 14425 3236 14429 3292
rect 14365 3232 14429 3236
rect 14445 3292 14509 3296
rect 14445 3236 14449 3292
rect 14449 3236 14505 3292
rect 14505 3236 14509 3292
rect 14445 3232 14509 3236
rect 14525 3292 14589 3296
rect 14525 3236 14529 3292
rect 14529 3236 14585 3292
rect 14585 3236 14589 3292
rect 14525 3232 14589 3236
rect 6285 2748 6349 2752
rect 6285 2692 6289 2748
rect 6289 2692 6345 2748
rect 6345 2692 6349 2748
rect 6285 2688 6349 2692
rect 6365 2748 6429 2752
rect 6365 2692 6369 2748
rect 6369 2692 6425 2748
rect 6425 2692 6429 2748
rect 6365 2688 6429 2692
rect 6445 2748 6509 2752
rect 6445 2692 6449 2748
rect 6449 2692 6505 2748
rect 6505 2692 6509 2748
rect 6445 2688 6509 2692
rect 6525 2748 6589 2752
rect 6525 2692 6529 2748
rect 6529 2692 6585 2748
rect 6585 2692 6589 2748
rect 6525 2688 6589 2692
rect 11618 2748 11682 2752
rect 11618 2692 11622 2748
rect 11622 2692 11678 2748
rect 11678 2692 11682 2748
rect 11618 2688 11682 2692
rect 11698 2748 11762 2752
rect 11698 2692 11702 2748
rect 11702 2692 11758 2748
rect 11758 2692 11762 2748
rect 11698 2688 11762 2692
rect 11778 2748 11842 2752
rect 11778 2692 11782 2748
rect 11782 2692 11838 2748
rect 11838 2692 11842 2748
rect 11778 2688 11842 2692
rect 11858 2748 11922 2752
rect 11858 2692 11862 2748
rect 11862 2692 11918 2748
rect 11918 2692 11922 2748
rect 11858 2688 11922 2692
rect 3618 2204 3682 2208
rect 3618 2148 3622 2204
rect 3622 2148 3678 2204
rect 3678 2148 3682 2204
rect 3618 2144 3682 2148
rect 3698 2204 3762 2208
rect 3698 2148 3702 2204
rect 3702 2148 3758 2204
rect 3758 2148 3762 2204
rect 3698 2144 3762 2148
rect 3778 2204 3842 2208
rect 3778 2148 3782 2204
rect 3782 2148 3838 2204
rect 3838 2148 3842 2204
rect 3778 2144 3842 2148
rect 3858 2204 3922 2208
rect 3858 2148 3862 2204
rect 3862 2148 3918 2204
rect 3918 2148 3922 2204
rect 3858 2144 3922 2148
rect 8952 2204 9016 2208
rect 8952 2148 8956 2204
rect 8956 2148 9012 2204
rect 9012 2148 9016 2204
rect 8952 2144 9016 2148
rect 9032 2204 9096 2208
rect 9032 2148 9036 2204
rect 9036 2148 9092 2204
rect 9092 2148 9096 2204
rect 9032 2144 9096 2148
rect 9112 2204 9176 2208
rect 9112 2148 9116 2204
rect 9116 2148 9172 2204
rect 9172 2148 9176 2204
rect 9112 2144 9176 2148
rect 9192 2204 9256 2208
rect 9192 2148 9196 2204
rect 9196 2148 9252 2204
rect 9252 2148 9256 2204
rect 9192 2144 9256 2148
rect 14285 2204 14349 2208
rect 14285 2148 14289 2204
rect 14289 2148 14345 2204
rect 14345 2148 14349 2204
rect 14285 2144 14349 2148
rect 14365 2204 14429 2208
rect 14365 2148 14369 2204
rect 14369 2148 14425 2204
rect 14425 2148 14429 2204
rect 14365 2144 14429 2148
rect 14445 2204 14509 2208
rect 14445 2148 14449 2204
rect 14449 2148 14505 2204
rect 14505 2148 14509 2204
rect 14445 2144 14509 2148
rect 14525 2204 14589 2208
rect 14525 2148 14529 2204
rect 14529 2148 14585 2204
rect 14585 2148 14589 2204
rect 14525 2144 14589 2148
<< metal4 >>
rect 3610 37024 3931 37584
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3931 37024
rect 3610 35936 3931 36960
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3931 35936
rect 3610 34848 3931 35872
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3931 34848
rect 3610 33760 3931 34784
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3931 33760
rect 3610 32672 3931 33696
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3931 32672
rect 3610 31584 3931 32608
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3931 31584
rect 3610 30496 3931 31520
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3931 30496
rect 3610 29408 3931 30432
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3931 29408
rect 3610 28320 3931 29344
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3931 28320
rect 3610 27232 3931 28256
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3931 27232
rect 3610 26144 3931 27168
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3931 26144
rect 3610 25056 3931 26080
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3931 25056
rect 3610 23968 3931 24992
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3931 23968
rect 3610 22880 3931 23904
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3931 22880
rect 3610 21792 3931 22816
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3931 21792
rect 3610 20704 3931 21728
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3931 20704
rect 3610 19616 3931 20640
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3931 19616
rect 3610 18528 3931 19552
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3931 18528
rect 3610 17440 3931 18464
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3931 17440
rect 3610 16352 3931 17376
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3931 16352
rect 3610 15264 3931 16288
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3931 15264
rect 3610 14176 3931 15200
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3931 14176
rect 3610 13088 3931 14112
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3931 13088
rect 3610 12000 3931 13024
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3931 12000
rect 3610 10912 3931 11936
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3931 10912
rect 3610 9824 3931 10848
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3931 9824
rect 3610 8736 3931 9760
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3931 8736
rect 3610 7648 3931 8672
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3931 7648
rect 3610 6560 3931 7584
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3931 6560
rect 3610 5472 3931 6496
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3931 5472
rect 3610 4384 3931 5408
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3931 4384
rect 3610 3296 3931 4320
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3931 3296
rect 3610 2208 3931 3232
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3931 2208
rect 3610 2128 3931 2144
rect 6277 37568 6597 37584
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 36480 6597 37504
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 35392 6597 36416
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 34304 6597 35328
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 33216 6597 34240
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 32128 6597 33152
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 31040 6597 32064
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 29952 6597 30976
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 28864 6597 29888
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 27776 6597 28800
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 26688 6597 27712
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 25600 6597 26624
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 24512 6597 25536
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 23424 6597 24448
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 22336 6597 23360
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 21248 6597 22272
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 20160 6597 21184
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 19072 6597 20096
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 17984 6597 19008
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 16896 6597 17920
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 15808 6597 16832
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 14720 6597 15744
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 13632 6597 14656
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 12544 6597 13568
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 11456 6597 12480
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 10368 6597 11392
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 9280 6597 10304
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 8192 6597 9216
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 7104 6597 8128
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 6016 6597 7040
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 4928 6597 5952
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 3840 6597 4864
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 2752 6597 3776
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2128 6597 2688
rect 8944 37024 9264 37584
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 35936 9264 36960
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 34848 9264 35872
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 33760 9264 34784
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 32672 9264 33696
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 31584 9264 32608
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 30496 9264 31520
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 29408 9264 30432
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 28320 9264 29344
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 27232 9264 28256
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 26144 9264 27168
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 25056 9264 26080
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 23968 9264 24992
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 22880 9264 23904
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 21792 9264 22816
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 20704 9264 21728
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 19616 9264 20640
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 18528 9264 19552
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 17440 9264 18464
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 16352 9264 17376
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 15264 9264 16288
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 14176 9264 15200
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 13088 9264 14112
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 12000 9264 13024
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 10912 9264 11936
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 9824 9264 10848
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 8736 9264 9760
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 7648 9264 8672
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 6560 9264 7584
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 5472 9264 6496
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 4384 9264 5408
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 3296 9264 4320
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 2208 9264 3232
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2128 9264 2144
rect 11610 37568 11930 37584
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 36480 11930 37504
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 35392 11930 36416
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 34304 11930 35328
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 33216 11930 34240
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 32128 11930 33152
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 31040 11930 32064
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 29952 11930 30976
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 28864 11930 29888
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 27776 11930 28800
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 26688 11930 27712
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 25600 11930 26624
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 24512 11930 25536
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 23424 11930 24448
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 22336 11930 23360
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 21248 11930 22272
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 20160 11930 21184
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 19072 11930 20096
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 17984 11930 19008
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 16896 11930 17920
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 15808 11930 16832
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 14720 11930 15744
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 13632 11930 14656
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 12544 11930 13568
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 11456 11930 12480
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 10368 11930 11392
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 9280 11930 10304
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 8192 11930 9216
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 7104 11930 8128
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 6016 11930 7040
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 4928 11930 5952
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 3840 11930 4864
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 2752 11930 3776
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2128 11930 2688
rect 14277 37024 14597 37584
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 35936 14597 36960
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 34848 14597 35872
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 33760 14597 34784
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 32672 14597 33696
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 31584 14597 32608
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 30496 14597 31520
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 29408 14597 30432
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 28320 14597 29344
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 27232 14597 28256
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 26144 14597 27168
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 25056 14597 26080
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 23968 14597 24992
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 22880 14597 23904
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 21792 14597 22816
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 20704 14597 21728
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 19616 14597 20640
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 18528 14597 19552
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 17440 14597 18464
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 16352 14597 17376
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 15264 14597 16288
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 14176 14597 15200
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 13088 14597 14112
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 12000 14597 13024
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 10912 14597 11936
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 9824 14597 10848
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 8736 14597 9760
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 7648 14597 8672
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 6560 14597 7584
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 5472 14597 6496
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 4384 14597 5408
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 3296 14597 4320
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 2208 14597 3232
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2128 14597 2144
use sky130_fd_sc_hd__fill_1  FILLER_1_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1748 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__15__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1564 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _38_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1604681595
transform 1 0 1840 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_12
timestamp 1604681595
transform 1 0 2208 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15
timestamp 1604681595
transform 1 0 2484 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11
timestamp 1604681595
transform 1 0 2116 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1604681595
transform 1 0 2392 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1604681595
transform 1 0 2300 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _13_
timestamp 1604681595
transform 1 0 2852 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_16 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2576 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_28 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3680 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1604681595
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__13__A
timestamp 1604681595
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_36
timestamp 1604681595
transform 1 0 4416 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36
timestamp 1604681595
transform 1 0 4416 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__07__A
timestamp 1604681595
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _31_
timestamp 1604681595
transform 1 0 4508 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_39
timestamp 1604681595
transform 1 0 4692 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41
timestamp 1604681595
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_50
timestamp 1604681595
transform 1 0 5704 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_46
timestamp 1604681595
transform 1 0 5336 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45
timestamp 1604681595
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__31__A
timestamp 1604681595
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1604681595
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1604681595
transform 1 0 5612 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1604681595
transform 1 0 4968 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_58
timestamp 1604681595
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1604681595
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1604681595
transform 1 0 6348 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53
timestamp 1604681595
transform 1 0 5980 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1604681595
transform 1 0 6164 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _04_
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _05_
timestamp 1604681595
transform 1 0 8556 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _27_
timestamp 1604681595
transform 1 0 8648 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__04__A
timestamp 1604681595
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67
timestamp 1604681595
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71
timestamp 1604681595
transform 1 0 7636 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_79
timestamp 1604681595
transform 1 0 8372 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_74
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_90
timestamp 1604681595
transform 1 0 9384 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_86
timestamp 1604681595
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89
timestamp 1604681595
transform 1 0 9292 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__27__A
timestamp 1604681595
transform 1 0 9200 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__05__A
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_98
timestamp 1604681595
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_98
timestamp 1604681595
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__28__A
timestamp 1604681595
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__29__A
timestamp 1604681595
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _29_
timestamp 1604681595
transform 1 0 9752 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _28_
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_102
timestamp 1604681595
transform 1 0 10488 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_102
timestamp 1604681595
transform 1 0 10488 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1604681595
transform 1 0 11224 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1604681595
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _25_
timestamp 1604681595
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_118
timestamp 1604681595
transform 1 0 11960 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604681595
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__25__A
timestamp 1604681595
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _22_
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1604681595
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__22__A
timestamp 1604681595
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_129
timestamp 1604681595
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_133
timestamp 1604681595
transform 1 0 13340 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145
timestamp 1604681595
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_127
timestamp 1604681595
transform 1 0 12788 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_131
timestamp 1604681595
transform 1 0 13156 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_143
timestamp 1604681595
transform 1 0 14260 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _15_
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_7
timestamp 1604681595
transform 1 0 1748 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_19
timestamp 1604681595
transform 1 0 2852 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _07_
timestamp 1604681595
transform 1 0 4508 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_36
timestamp 1604681595
transform 1 0 4416 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1604681595
transform 1 0 4876 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1604681595
transform 1 0 5980 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1604681595
transform 1 0 7084 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_77
timestamp 1604681595
transform 1 0 8188 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_89
timestamp 1604681595
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1604681595
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1604681595
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1604681595
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1604681595
transform 1 0 14076 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_145
timestamp 1604681595
transform 1 0 14444 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 14812 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604681595
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1604681595
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1604681595
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_135
timestamp 1604681595
transform 1 0 13524 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_143
timestamp 1604681595
transform 1 0 14260 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604681595
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1604681595
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1604681595
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1604681595
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1604681595
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1604681595
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1604681595
transform 1 0 14076 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_145
timestamp 1604681595
transform 1 0 14444 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 14812 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1604681595
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1604681595
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1604681595
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1604681595
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1604681595
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1604681595
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1604681595
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_135
timestamp 1604681595
transform 1 0 13524 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_143
timestamp 1604681595
transform 1 0 14260 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1604681595
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1604681595
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_7
timestamp 1604681595
transform 1 0 1748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_19
timestamp 1604681595
transform 1 0 2852 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1604681595
transform 1 0 4140 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1604681595
transform 1 0 4692 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_31
timestamp 1604681595
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_37
timestamp 1604681595
transform 1 0 4508 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_41
timestamp 1604681595
transform 1 0 4876 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__10__A
timestamp 1604681595
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604681595
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_55 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6164 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _09_
timestamp 1604681595
transform 1 0 8648 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _24_
timestamp 1604681595
transform 1 0 7544 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__24__A
timestamp 1604681595
transform 1 0 8096 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1604681595
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_74
timestamp 1604681595
transform 1 0 7912 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_78
timestamp 1604681595
transform 1 0 8280 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _02_
timestamp 1604681595
transform 1 0 10304 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__09__A
timestamp 1604681595
transform 1 0 9200 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_86
timestamp 1604681595
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_90
timestamp 1604681595
transform 1 0 9384 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_98
timestamp 1604681595
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_104
timestamp 1604681595
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__02__A
timestamp 1604681595
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__26__A
timestamp 1604681595
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1604681595
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1604681595
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_108
timestamp 1604681595
transform 1 0 11040 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_112
timestamp 1604681595
transform 1 0 11408 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1604681595
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1604681595
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp 1604681595
transform 1 0 14076 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_145
timestamp 1604681595
transform 1 0 14444 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_135
timestamp 1604681595
transform 1 0 13524 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_143
timestamp 1604681595
transform 1 0 14260 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 14812 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1604681595
transform 1 0 1564 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_9
timestamp 1604681595
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_21
timestamp 1604681595
transform 1 0 3036 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1604681595
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _10_
timestamp 1604681595
transform 1 0 5980 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_44
timestamp 1604681595
transform 1 0 5152 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_52
timestamp 1604681595
transform 1 0 5888 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_57
timestamp 1604681595
transform 1 0 6348 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_69
timestamp 1604681595
transform 1 0 7452 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_81
timestamp 1604681595
transform 1 0 8556 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _26_
timestamp 1604681595
transform 1 0 10396 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_89
timestamp 1604681595
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1604681595
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1604681595
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1604681595
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1604681595
transform 1 0 14076 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_145
timestamp 1604681595
transform 1 0 14444 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 14812 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1604681595
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__08__A
timestamp 1604681595
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_41
timestamp 1604681595
transform 1 0 4876 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _30_
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_53
timestamp 1604681595
transform 1 0 5980 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__30__A
timestamp 1604681595
transform 1 0 7360 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_66
timestamp 1604681595
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_70
timestamp 1604681595
transform 1 0 7544 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_82
timestamp 1604681595
transform 1 0 8648 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_94
timestamp 1604681595
transform 1 0 9752 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_106
timestamp 1604681595
transform 1 0 10856 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1604681595
transform 1 0 11960 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_135
timestamp 1604681595
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_143
timestamp 1604681595
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 14812 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1604681595
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _08_
timestamp 1604681595
transform 1 0 4692 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_38
timestamp 1604681595
transform 1 0 4600 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_43
timestamp 1604681595
transform 1 0 5060 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_55
timestamp 1604681595
transform 1 0 6164 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_67
timestamp 1604681595
transform 1 0 7268 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_79
timestamp 1604681595
transform 1 0 8372 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1604681595
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1604681595
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1604681595
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1604681595
transform 1 0 14076 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_145
timestamp 1604681595
transform 1 0 14444 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1604681595
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1604681595
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1604681595
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1604681595
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__03__A
timestamp 1604681595
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_86
timestamp 1604681595
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_98
timestamp 1604681595
transform 1 0 10120 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_103
timestamp 1604681595
transform 1 0 10580 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _23_
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__23__A
timestamp 1604681595
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_115
timestamp 1604681595
transform 1 0 11684 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_119
timestamp 1604681595
transform 1 0 12052 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1604681595
transform 1 0 12972 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_127
timestamp 1604681595
transform 1 0 12788 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_131
timestamp 1604681595
transform 1 0 13156 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_143
timestamp 1604681595
transform 1 0 14260 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 14812 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1604681595
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1604681595
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1604681595
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1604681595
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1604681595
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _03_
timestamp 1604681595
transform 1 0 10396 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604681595
transform 1 0 12328 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1604681595
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_117
timestamp 1604681595
transform 1 0 11868 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_121
timestamp 1604681595
transform 1 0 12236 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_126
timestamp 1604681595
transform 1 0 12696 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_138
timestamp 1604681595
transform 1 0 13800 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 14812 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _11_
timestamp 1604681595
transform 1 0 2668 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_15
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1604681595
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__11__A
timestamp 1604681595
transform 1 0 3220 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_21
timestamp 1604681595
transform 1 0 3036 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_25
timestamp 1604681595
transform 1 0 3404 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_37
timestamp 1604681595
transform 1 0 4508 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604681595
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_49
timestamp 1604681595
transform 1 0 5612 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1604681595
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1604681595
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1604681595
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1604681595
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1604681595
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_86
timestamp 1604681595
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_98
timestamp 1604681595
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_110
timestamp 1604681595
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1604681595
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_117
timestamp 1604681595
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_135
timestamp 1604681595
transform 1 0 13524 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_143
timestamp 1604681595
transform 1 0 14260 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_129
timestamp 1604681595
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1604681595
transform 1 0 14076 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_145
timestamp 1604681595
transform 1 0 14444 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 14812 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 14812 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1604681595
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_11
timestamp 1604681595
transform 1 0 2116 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_23
timestamp 1604681595
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_35
timestamp 1604681595
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_47
timestamp 1604681595
transform 1 0 5428 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1604681595
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_98
timestamp 1604681595
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _21_
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_110
timestamp 1604681595
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__21__A
timestamp 1604681595
transform 1 0 12972 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_127
timestamp 1604681595
transform 1 0 12788 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_131
timestamp 1604681595
transform 1 0 13156 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_143
timestamp 1604681595
transform 1 0 14260 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 14812 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1604681595
transform 1 0 1932 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_3
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_13
timestamp 1604681595
transform 1 0 2300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_25
timestamp 1604681595
transform 1 0 3404 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1604681595
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1604681595
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1604681595
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1604681595
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_117
timestamp 1604681595
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_129
timestamp 1604681595
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1604681595
transform 1 0 14076 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_145
timestamp 1604681595
transform 1 0 14444 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 14812 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_7
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_19
timestamp 1604681595
transform 1 0 2852 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_31
timestamp 1604681595
transform 1 0 3956 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_43
timestamp 1604681595
transform 1 0 5060 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_55
timestamp 1604681595
transform 1 0 6164 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1604681595
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1604681595
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_98
timestamp 1604681595
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_110
timestamp 1604681595
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_135
timestamp 1604681595
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_143
timestamp 1604681595
transform 1 0 14260 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 14812 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_9
timestamp 1604681595
transform 1 0 1932 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_21
timestamp 1604681595
transform 1 0 3036 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1604681595
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1604681595
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1604681595
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1604681595
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1604681595
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1604681595
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1604681595
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1604681595
transform 1 0 14076 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_145
timestamp 1604681595
transform 1 0 14444 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 14812 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1604681595
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1604681595
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1604681595
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1604681595
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1604681595
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1604681595
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1604681595
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 7912 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1604681595
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_68
timestamp 1604681595
transform 1 0 7360 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_76
timestamp 1604681595
transform 1 0 8096 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1604681595
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1604681595
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_88
timestamp 1604681595
transform 1 0 9200 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1604681595
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1604681595
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1604681595
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_135
timestamp 1604681595
transform 1 0 13524 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_143
timestamp 1604681595
transform 1 0 14260 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1604681595
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1604681595
transform 1 0 14076 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_145
timestamp 1604681595
transform 1 0 14444 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 14812 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 14812 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1604681595
transform 1 0 2024 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1604681595
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_9
timestamp 1604681595
transform 1 0 1932 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_14
timestamp 1604681595
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_18
timestamp 1604681595
transform 1 0 2760 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_30
timestamp 1604681595
transform 1 0 3864 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_42
timestamp 1604681595
transform 1 0 4968 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_54
timestamp 1604681595
transform 1 0 6072 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp 1604681595
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7912 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 7728 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_70
timestamp 1604681595
transform 1 0 7544 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_83
timestamp 1604681595
transform 1 0 8740 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_95
timestamp 1604681595
transform 1 0 9844 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_107
timestamp 1604681595
transform 1 0 10948 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_119
timestamp 1604681595
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_135
timestamp 1604681595
transform 1 0 13524 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_143
timestamp 1604681595
transform 1 0 14260 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 14812 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604681595
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 4416 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1604681595
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_38
timestamp 1604681595
transform 1 0 4600 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_46
timestamp 1604681595
transform 1 0 5336 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_58
timestamp 1604681595
transform 1 0 6440 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 7912 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_66
timestamp 1604681595
transform 1 0 7176 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_69
timestamp 1604681595
transform 1 0 7452 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_73
timestamp 1604681595
transform 1 0 7820 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_76
timestamp 1604681595
transform 1 0 8096 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_88
timestamp 1604681595
transform 1 0 9200 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1604681595
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1604681595
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1604681595
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1604681595
transform 1 0 14076 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_145
timestamp 1604681595
transform 1 0 14444 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 14812 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _17_
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__17__A
timestamp 1604681595
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_7
timestamp 1604681595
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_11
timestamp 1604681595
transform 1 0 2116 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 4416 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_23
timestamp 1604681595
transform 1 0 3220 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_29
timestamp 1604681595
transform 1 0 3772 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_32
timestamp 1604681595
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 5428 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_45
timestamp 1604681595
transform 1 0 5244 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_49
timestamp 1604681595
transform 1 0 5612 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_53
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7268 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7084 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_76
timestamp 1604681595
transform 1 0 8096 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9476 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 9292 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_84
timestamp 1604681595
transform 1 0 8832 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_87
timestamp 1604681595
transform 1 0 9108 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_107
timestamp 1604681595
transform 1 0 10948 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_119
timestamp 1604681595
transform 1 0 12052 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_135
timestamp 1604681595
transform 1 0 13524 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_143
timestamp 1604681595
transform 1 0 14260 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 14812 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604681595
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_38
timestamp 1604681595
transform 1 0 4600 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5152 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1604681595
transform 1 0 5980 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7268 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_65
timestamp 1604681595
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_69
timestamp 1604681595
transform 1 0 7452 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_81
timestamp 1604681595
transform 1 0 8556 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_89
timestamp 1604681595
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1604681595
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1604681595
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1604681595
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1604681595
transform 1 0 14076 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1604681595
transform 1 0 14444 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 14812 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1604681595
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4416 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_27
timestamp 1604681595
transform 1 0 3588 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_33
timestamp 1604681595
transform 1 0 4140 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_45
timestamp 1604681595
transform 1 0 5244 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1604681595
transform 1 0 6348 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1604681595
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1604681595
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1604681595
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11500 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 11868 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_110
timestamp 1604681595
transform 1 0 11224 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_115
timestamp 1604681595
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_119
timestamp 1604681595
transform 1 0 12052 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_135
timestamp 1604681595
transform 1 0 13524 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_143
timestamp 1604681595
transform 1 0 14260 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 14812 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1604681595
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1604681595
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4416 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_38
timestamp 1604681595
transform 1 0 4600 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1604681595
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1604681595
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_50
timestamp 1604681595
transform 1 0 5704 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_62
timestamp 1604681595
transform 1 0 6808 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1604681595
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1604681595
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_74
timestamp 1604681595
transform 1 0 7912 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1604681595
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_86
timestamp 1604681595
transform 1 0 9016 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1604681595
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1604681595
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11500 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_105
timestamp 1604681595
transform 1 0 10764 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1604681595
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1604681595
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_141
timestamp 1604681595
transform 1 0 14076 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_145
timestamp 1604681595
transform 1 0 14444 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_135
timestamp 1604681595
transform 1 0 13524 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_143
timestamp 1604681595
transform 1 0 14260 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 14812 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 14812 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1604681595
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1604681595
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1604681595
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1604681595
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1604681595
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1604681595
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1604681595
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1604681595
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_141
timestamp 1604681595
transform 1 0 14076 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_145
timestamp 1604681595
transform 1 0 14444 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 14812 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1604681595
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1604681595
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1604681595
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1604681595
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1604681595
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1604681595
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1604681595
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_110
timestamp 1604681595
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_135
timestamp 1604681595
transform 1 0 13524 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_143
timestamp 1604681595
transform 1 0 14260 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 14812 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604681595
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1604681595
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1604681595
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1604681595
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1604681595
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1604681595
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1604681595
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1604681595
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1604681595
transform 1 0 14076 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_145
timestamp 1604681595
transform 1 0 14444 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 14812 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1604681595
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1604681595
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1604681595
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1604681595
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1604681595
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__19__A
timestamp 1604681595
transform 1 0 12604 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1604681595
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_127
timestamp 1604681595
transform 1 0 12788 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_139
timestamp 1604681595
transform 1 0 13892 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_145
timestamp 1604681595
transform 1 0 14444 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 14812 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_56
timestamp 1604681595
transform 1 0 6256 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 6992 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_66
timestamp 1604681595
transform 1 0 7176 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_78
timestamp 1604681595
transform 1 0 8280 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_90
timestamp 1604681595
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _19_
timestamp 1604681595
transform 1 0 12328 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1604681595
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_117
timestamp 1604681595
transform 1 0 11868 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_121
timestamp 1604681595
transform 1 0 12236 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_126
timestamp 1604681595
transform 1 0 12696 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_138
timestamp 1604681595
transform 1 0 13800 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 14812 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1604681595
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604681595
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_56
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 6992 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8556 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6992 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_73
timestamp 1604681595
transform 1 0 7820 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_66
timestamp 1604681595
transform 1 0 7176 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_78
timestamp 1604681595
transform 1 0 8280 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 9016 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_84
timestamp 1604681595
transform 1 0 8832 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_88
timestamp 1604681595
transform 1 0 9200 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_100
timestamp 1604681595
transform 1 0 10304 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_90
timestamp 1604681595
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_112
timestamp 1604681595
transform 1 0 11408 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_120
timestamp 1604681595
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604681595
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1604681595
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_135
timestamp 1604681595
transform 1 0 13524 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_143
timestamp 1604681595
transform 1 0 14260 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1604681595
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1604681595
transform 1 0 14076 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1604681595
transform 1 0 14444 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 14812 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 14812 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_39
timestamp 1604681595
transform 1 0 4692 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 5612 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 5980 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 6348 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_47
timestamp 1604681595
transform 1 0 5428 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_51
timestamp 1604681595
transform 1 0 5796 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_55
timestamp 1604681595
transform 1 0 6164 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1604681595
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_74
timestamp 1604681595
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_86
timestamp 1604681595
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_98
timestamp 1604681595
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_110
timestamp 1604681595
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_123
timestamp 1604681595
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_135
timestamp 1604681595
transform 1 0 13524 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_143
timestamp 1604681595
transform 1 0 14260 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 14812 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604681595
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1604681595
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1604681595
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1604681595
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1604681595
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 5612 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_36_44
timestamp 1604681595
transform 1 0 5152 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_48
timestamp 1604681595
transform 1 0 5520 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_58
timestamp 1604681595
transform 1 0 6440 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_70
timestamp 1604681595
transform 1 0 7544 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_82
timestamp 1604681595
transform 1 0 8648 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 9844 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 10212 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_93
timestamp 1604681595
transform 1 0 9660 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_97
timestamp 1604681595
transform 1 0 10028 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_101
timestamp 1604681595
transform 1 0 10396 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_113
timestamp 1604681595
transform 1 0 11500 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_125
timestamp 1604681595
transform 1 0 12604 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_137
timestamp 1604681595
transform 1 0 13708 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_145
timestamp 1604681595
transform 1 0 14444 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604681595
transform -1 0 14812 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604681595
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1604681595
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1604681595
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1604681595
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1604681595
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_51
timestamp 1604681595
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1604681595
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_62
timestamp 1604681595
transform 1 0 6808 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7544 0 1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 7360 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 9384 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 10396 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_99
timestamp 1604681595
transform 1 0 10212 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_103
timestamp 1604681595
transform 1 0 10580 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 10764 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_107
timestamp 1604681595
transform 1 0 10948 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_119
timestamp 1604681595
transform 1 0 12052 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_123
timestamp 1604681595
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_135
timestamp 1604681595
transform 1 0 13524 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_143
timestamp 1604681595
transform 1 0 14260 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604681595
transform -1 0 14812 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604681595
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1604681595
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1604681595
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1604681595
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1604681595
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1604681595
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1604681595
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1604681595
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_80
timestamp 1604681595
transform 1 0 8464 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_88
timestamp 1604681595
transform 1 0 9200 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_102
timestamp 1604681595
transform 1 0 10488 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_114
timestamp 1604681595
transform 1 0 11592 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_126
timestamp 1604681595
transform 1 0 12696 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_138
timestamp 1604681595
transform 1 0 13800 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604681595
transform -1 0 14812 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604681595
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604681595
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1604681595
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1604681595
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1604681595
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1604681595
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1604681595
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1604681595
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1604681595
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1604681595
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1604681595
transform 1 0 6256 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 6256 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1604681595
transform 1 0 5796 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1604681595
transform 1 0 6164 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_58
timestamp 1604681595
transform 1 0 6440 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1604681595
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1604681595
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_59
timestamp 1604681595
transform 1 0 6532 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_74
timestamp 1604681595
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_71
timestamp 1604681595
transform 1 0 7636 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_83
timestamp 1604681595
transform 1 0 8740 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_86
timestamp 1604681595
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_98
timestamp 1604681595
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_91
timestamp 1604681595
transform 1 0 9476 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_93
timestamp 1604681595
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1604681595
transform 1 0 11868 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1604681595
transform 1 0 11868 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_110
timestamp 1604681595
transform 1 0 11224 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_116
timestamp 1604681595
transform 1 0 11776 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_119
timestamp 1604681595
transform 1 0 12052 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1604681595
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_105
timestamp 1604681595
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1604681595
transform 1 0 12236 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_135
timestamp 1604681595
transform 1 0 13524 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_143
timestamp 1604681595
transform 1 0 14260 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_133
timestamp 1604681595
transform 1 0 13340 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_145
timestamp 1604681595
transform 1 0 14444 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604681595
transform -1 0 14812 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604681595
transform -1 0 14812 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604681595
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1604681595
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1604681595
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1604681595
transform 1 0 4048 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_27
timestamp 1604681595
transform 1 0 3588 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_31
timestamp 1604681595
transform 1 0 3956 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_34
timestamp 1604681595
transform 1 0 4232 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_46
timestamp 1604681595
transform 1 0 5336 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_58
timestamp 1604681595
transform 1 0 6440 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1604681595
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_74
timestamp 1604681595
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_86
timestamp 1604681595
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_98
timestamp 1604681595
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_110
timestamp 1604681595
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1604681595
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_135
timestamp 1604681595
transform 1 0 13524 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_143
timestamp 1604681595
transform 1 0 14260 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604681595
transform -1 0 14812 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604681595
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1604681595
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1604681595
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1604681595
transform 1 0 4048 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1604681595
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_36
timestamp 1604681595
transform 1 0 4416 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_48
timestamp 1604681595
transform 1 0 5520 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_60
timestamp 1604681595
transform 1 0 6624 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_72
timestamp 1604681595
transform 1 0 7728 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_84
timestamp 1604681595
transform 1 0 8832 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_93
timestamp 1604681595
transform 1 0 9660 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_105
timestamp 1604681595
transform 1 0 10764 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_117
timestamp 1604681595
transform 1 0 11868 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_129
timestamp 1604681595
transform 1 0 12972 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_141
timestamp 1604681595
transform 1 0 14076 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_145
timestamp 1604681595
transform 1 0 14444 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604681595
transform -1 0 14812 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _18_
timestamp 1604681595
transform 1 0 1380 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1604681595
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__18__A
timestamp 1604681595
transform 1 0 1932 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_7
timestamp 1604681595
transform 1 0 1748 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_11
timestamp 1604681595
transform 1 0 2116 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_23
timestamp 1604681595
transform 1 0 3220 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_35
timestamp 1604681595
transform 1 0 4324 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_47
timestamp 1604681595
transform 1 0 5428 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_59
timestamp 1604681595
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_62
timestamp 1604681595
transform 1 0 6808 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_74
timestamp 1604681595
transform 1 0 7912 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_86
timestamp 1604681595
transform 1 0 9016 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_98
timestamp 1604681595
transform 1 0 10120 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_110
timestamp 1604681595
transform 1 0 11224 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_123
timestamp 1604681595
transform 1 0 12420 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_135
timestamp 1604681595
transform 1 0 13524 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_143
timestamp 1604681595
transform 1 0 14260 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1604681595
transform -1 0 14812 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1604681595
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1604681595
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1604681595
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_27
timestamp 1604681595
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_32
timestamp 1604681595
transform 1 0 4048 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_44
timestamp 1604681595
transform 1 0 5152 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_56
timestamp 1604681595
transform 1 0 6256 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_68
timestamp 1604681595
transform 1 0 7360 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_80
timestamp 1604681595
transform 1 0 8464 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_93
timestamp 1604681595
transform 1 0 9660 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_105
timestamp 1604681595
transform 1 0 10764 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_117
timestamp 1604681595
transform 1 0 11868 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_129
timestamp 1604681595
transform 1 0 12972 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_141
timestamp 1604681595
transform 1 0 14076 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_145
timestamp 1604681595
transform 1 0 14444 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1604681595
transform -1 0 14812 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1604681595
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1604681595
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1604681595
transform 1 0 2484 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1604681595
transform 1 0 3588 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1604681595
transform 1 0 4692 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_51
timestamp 1604681595
transform 1 0 5796 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_59
timestamp 1604681595
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_62
timestamp 1604681595
transform 1 0 6808 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_74
timestamp 1604681595
transform 1 0 7912 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_86
timestamp 1604681595
transform 1 0 9016 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_98
timestamp 1604681595
transform 1 0 10120 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_110
timestamp 1604681595
transform 1 0 11224 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_123
timestamp 1604681595
transform 1 0 12420 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_135
timestamp 1604681595
transform 1 0 13524 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_143
timestamp 1604681595
transform 1 0 14260 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1604681595
transform -1 0 14812 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1604681595
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1604681595
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1604681595
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1604681595
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1604681595
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1604681595
transform 1 0 2484 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 4508 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 4324 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 4508 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_27
timestamp 1604681595
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_32
timestamp 1604681595
transform 1 0 4048 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_36
timestamp 1604681595
transform 1 0 4416 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_39
timestamp 1604681595
transform 1 0 4692 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_27
timestamp 1604681595
transform 1 0 3588 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_51
timestamp 1604681595
transform 1 0 5796 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_53
timestamp 1604681595
transform 1 0 5980 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_62
timestamp 1604681595
transform 1 0 6808 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_63
timestamp 1604681595
transform 1 0 6900 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_75
timestamp 1604681595
transform 1 0 8004 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_74
timestamp 1604681595
transform 1 0 7912 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_87
timestamp 1604681595
transform 1 0 9108 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_91
timestamp 1604681595
transform 1 0 9476 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_93
timestamp 1604681595
transform 1 0 9660 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_86
timestamp 1604681595
transform 1 0 9016 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_98
timestamp 1604681595
transform 1 0 10120 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_105
timestamp 1604681595
transform 1 0 10764 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_117
timestamp 1604681595
transform 1 0 11868 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_110
timestamp 1604681595
transform 1 0 11224 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_123
timestamp 1604681595
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_129
timestamp 1604681595
transform 1 0 12972 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_141
timestamp 1604681595
transform 1 0 14076 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_145
timestamp 1604681595
transform 1 0 14444 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_135
timestamp 1604681595
transform 1 0 13524 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_143
timestamp 1604681595
transform 1 0 14260 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1604681595
transform -1 0 14812 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1604681595
transform -1 0 14812 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1604681595
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 2392 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_3
timestamp 1604681595
transform 1 0 1380 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_11
timestamp 1604681595
transform 1 0 2116 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_16
timestamp 1604681595
transform 1 0 2576 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_28
timestamp 1604681595
transform 1 0 3680 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_32
timestamp 1604681595
transform 1 0 4048 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_44
timestamp 1604681595
transform 1 0 5152 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_56
timestamp 1604681595
transform 1 0 6256 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_68
timestamp 1604681595
transform 1 0 7360 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_80
timestamp 1604681595
transform 1 0 8464 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_93
timestamp 1604681595
transform 1 0 9660 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_105
timestamp 1604681595
transform 1 0 10764 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_117
timestamp 1604681595
transform 1 0 11868 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_129
timestamp 1604681595
transform 1 0 12972 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_141
timestamp 1604681595
transform 1 0 14076 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_145
timestamp 1604681595
transform 1 0 14444 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1604681595
transform -1 0 14812 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 2392 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1604681595
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 2208 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_3
timestamp 1604681595
transform 1 0 1380 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_11
timestamp 1604681595
transform 1 0 2116 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_30
timestamp 1604681595
transform 1 0 3864 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_42
timestamp 1604681595
transform 1 0 4968 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_54
timestamp 1604681595
transform 1 0 6072 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_60
timestamp 1604681595
transform 1 0 6624 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_62
timestamp 1604681595
transform 1 0 6808 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 7268 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 7636 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_66
timestamp 1604681595
transform 1 0 7176 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_69
timestamp 1604681595
transform 1 0 7452 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_73
timestamp 1604681595
transform 1 0 7820 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_85
timestamp 1604681595
transform 1 0 8924 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_97
timestamp 1604681595
transform 1 0 10028 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_109
timestamp 1604681595
transform 1 0 11132 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_121
timestamp 1604681595
transform 1 0 12236 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_123
timestamp 1604681595
transform 1 0 12420 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_135
timestamp 1604681595
transform 1 0 13524 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_143
timestamp 1604681595
transform 1 0 14260 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1604681595
transform -1 0 14812 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1604681595
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1604681595
transform 1 0 1380 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1604681595
transform 1 0 2484 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_27
timestamp 1604681595
transform 1 0 3588 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_32
timestamp 1604681595
transform 1 0 4048 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_44
timestamp 1604681595
transform 1 0 5152 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_56
timestamp 1604681595
transform 1 0 6256 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 7268 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_50_64
timestamp 1604681595
transform 1 0 6992 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_50_83
timestamp 1604681595
transform 1 0 8740 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 9292 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_91
timestamp 1604681595
transform 1 0 9476 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_93
timestamp 1604681595
transform 1 0 9660 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_105
timestamp 1604681595
transform 1 0 10764 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_117
timestamp 1604681595
transform 1 0 11868 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_129
timestamp 1604681595
transform 1 0 12972 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_141
timestamp 1604681595
transform 1 0 14076 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_145
timestamp 1604681595
transform 1 0 14444 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1604681595
transform -1 0 14812 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1604681595
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1604681595
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1604681595
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1604681595
transform 1 0 3588 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1604681595
transform 1 0 4692 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_51
timestamp 1604681595
transform 1 0 5796 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_59
timestamp 1604681595
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_62
timestamp 1604681595
transform 1 0 6808 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_74
timestamp 1604681595
transform 1 0 7912 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 9292 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 9108 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_86
timestamp 1604681595
transform 1 0 9016 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_98
timestamp 1604681595
transform 1 0 10120 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_110
timestamp 1604681595
transform 1 0 11224 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_123
timestamp 1604681595
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_135
timestamp 1604681595
transform 1 0 13524 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_143
timestamp 1604681595
transform 1 0 14260 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1604681595
transform -1 0 14812 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_7
timestamp 1604681595
transform 1 0 1748 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1604681595
transform 1 0 1380 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__14__A
timestamp 1604681595
transform 1 0 1564 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__16__A
timestamp 1604681595
transform 1 0 1932 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1604681595
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1604681595
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _14_
timestamp 1604681595
transform 1 0 1380 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_11
timestamp 1604681595
transform 1 0 2116 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_19
timestamp 1604681595
transform 1 0 2852 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_7
timestamp 1604681595
transform 1 0 1748 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__12__A
timestamp 1604681595
transform 1 0 4048 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_32
timestamp 1604681595
transform 1 0 4048 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_23
timestamp 1604681595
transform 1 0 3220 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_31
timestamp 1604681595
transform 1 0 3956 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_34
timestamp 1604681595
transform 1 0 4232 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__06__A
timestamp 1604681595
transform 1 0 5152 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_44
timestamp 1604681595
transform 1 0 5152 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_56
timestamp 1604681595
transform 1 0 6256 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_42
timestamp 1604681595
transform 1 0 4968 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_46
timestamp 1604681595
transform 1 0 5336 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_58
timestamp 1604681595
transform 1 0 6440 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_62
timestamp 1604681595
transform 1 0 6808 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1604681595
transform 1 0 8556 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_68
timestamp 1604681595
transform 1 0 7360 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_80
timestamp 1604681595
transform 1 0 8464 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_53_74
timestamp 1604681595
transform 1 0 7912 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_80
timestamp 1604681595
transform 1 0 8464 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_85
timestamp 1604681595
transform 1 0 8924 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_91
timestamp 1604681595
transform 1 0 9476 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_88
timestamp 1604681595
transform 1 0 9200 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 9292 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1604681595
transform 1 0 9108 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _01_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9660 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_101
timestamp 1604681595
transform 1 0 10396 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_89
timestamp 1604681595
transform 1 0 9292 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_96
timestamp 1604681595
transform 1 0 9936 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _20_
timestamp 1604681595
transform 1 0 12420 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_108
timestamp 1604681595
transform 1 0 11040 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_120
timestamp 1604681595
transform 1 0 12144 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_113
timestamp 1604681595
transform 1 0 11500 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_121
timestamp 1604681595
transform 1 0 12236 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__20__A
timestamp 1604681595
transform 1 0 12972 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_132
timestamp 1604681595
transform 1 0 13248 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_144
timestamp 1604681595
transform 1 0 14352 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_127
timestamp 1604681595
transform 1 0 12788 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_131
timestamp 1604681595
transform 1 0 13156 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_143
timestamp 1604681595
transform 1 0 14260 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1604681595
transform -1 0 14812 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1604681595
transform -1 0 14812 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _16_
timestamp 1604681595
transform 1 0 1380 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1604681595
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_7
timestamp 1604681595
transform 1 0 1748 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_19
timestamp 1604681595
transform 1 0 2852 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _12_
timestamp 1604681595
transform 1 0 4048 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_36
timestamp 1604681595
transform 1 0 4416 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _06_
timestamp 1604681595
transform 1 0 5152 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_48
timestamp 1604681595
transform 1 0 5520 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_60
timestamp 1604681595
transform 1 0 6624 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_72
timestamp 1604681595
transform 1 0 7728 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_84
timestamp 1604681595
transform 1 0 8832 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_93
timestamp 1604681595
transform 1 0 9660 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_105
timestamp 1604681595
transform 1 0 10764 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_117
timestamp 1604681595
transform 1 0 11868 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_129
timestamp 1604681595
transform 1 0 12972 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_141
timestamp 1604681595
transform 1 0 14076 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_145
timestamp 1604681595
transform 1 0 14444 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1604681595
transform -1 0 14812 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1604681595
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1604681595
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1604681595
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1604681595
transform 1 0 3588 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1604681595
transform 1 0 4692 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_51
timestamp 1604681595
transform 1 0 5796 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_59
timestamp 1604681595
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_62
timestamp 1604681595
transform 1 0 6808 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_74
timestamp 1604681595
transform 1 0 7912 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_86
timestamp 1604681595
transform 1 0 9016 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_98
timestamp 1604681595
transform 1 0 10120 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604681595
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_110
timestamp 1604681595
transform 1 0 11224 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_123
timestamp 1604681595
transform 1 0 12420 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_135
timestamp 1604681595
transform 1 0 13524 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_143
timestamp 1604681595
transform 1 0 14260 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1604681595
transform -1 0 14812 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1604681595
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1604681595
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1604681595
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604681595
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_27
timestamp 1604681595
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_32
timestamp 1604681595
transform 1 0 4048 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_44
timestamp 1604681595
transform 1 0 5152 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_56
timestamp 1604681595
transform 1 0 6256 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_68
timestamp 1604681595
transform 1 0 7360 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_80
timestamp 1604681595
transform 1 0 8464 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604681595
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_93
timestamp 1604681595
transform 1 0 9660 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_105
timestamp 1604681595
transform 1 0 10764 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_117
timestamp 1604681595
transform 1 0 11868 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_129
timestamp 1604681595
transform 1 0 12972 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_141
timestamp 1604681595
transform 1 0 14076 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_145
timestamp 1604681595
transform 1 0 14444 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1604681595
transform -1 0 14812 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1604681595
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1604681595
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1604681595
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1604681595
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1604681595
transform 1 0 4692 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604681595
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_51
timestamp 1604681595
transform 1 0 5796 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_59
timestamp 1604681595
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_62
timestamp 1604681595
transform 1 0 6808 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_74
timestamp 1604681595
transform 1 0 7912 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_86
timestamp 1604681595
transform 1 0 9016 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_98
timestamp 1604681595
transform 1 0 10120 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604681595
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_110
timestamp 1604681595
transform 1 0 11224 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_123
timestamp 1604681595
transform 1 0 12420 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_135
timestamp 1604681595
transform 1 0 13524 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_143
timestamp 1604681595
transform 1 0 14260 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1604681595
transform -1 0 14812 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1604681595
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1604681595
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1604681595
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604681595
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_27
timestamp 1604681595
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_32
timestamp 1604681595
transform 1 0 4048 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_44
timestamp 1604681595
transform 1 0 5152 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_56
timestamp 1604681595
transform 1 0 6256 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_68
timestamp 1604681595
transform 1 0 7360 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_80
timestamp 1604681595
transform 1 0 8464 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604681595
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_93
timestamp 1604681595
transform 1 0 9660 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_105
timestamp 1604681595
transform 1 0 10764 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_117
timestamp 1604681595
transform 1 0 11868 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_129
timestamp 1604681595
transform 1 0 12972 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_141
timestamp 1604681595
transform 1 0 14076 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_145
timestamp 1604681595
transform 1 0 14444 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1604681595
transform -1 0 14812 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1604681595
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1604681595
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1604681595
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1604681595
transform 1 0 2484 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1604681595
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1604681595
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604681595
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1604681595
transform 1 0 3588 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1604681595
transform 1 0 4692 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_27
timestamp 1604681595
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_32
timestamp 1604681595
transform 1 0 4048 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604681595
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_51
timestamp 1604681595
transform 1 0 5796 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_59
timestamp 1604681595
transform 1 0 6532 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_62
timestamp 1604681595
transform 1 0 6808 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_44
timestamp 1604681595
transform 1 0 5152 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_56
timestamp 1604681595
transform 1 0 6256 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_74
timestamp 1604681595
transform 1 0 7912 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_68
timestamp 1604681595
transform 1 0 7360 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_80
timestamp 1604681595
transform 1 0 8464 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604681595
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_86
timestamp 1604681595
transform 1 0 9016 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_98
timestamp 1604681595
transform 1 0 10120 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_93
timestamp 1604681595
transform 1 0 9660 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604681595
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_110
timestamp 1604681595
transform 1 0 11224 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_123
timestamp 1604681595
transform 1 0 12420 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_105
timestamp 1604681595
transform 1 0 10764 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_117
timestamp 1604681595
transform 1 0 11868 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_135
timestamp 1604681595
transform 1 0 13524 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_143
timestamp 1604681595
transform 1 0 14260 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_129
timestamp 1604681595
transform 1 0 12972 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_141
timestamp 1604681595
transform 1 0 14076 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_145
timestamp 1604681595
transform 1 0 14444 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1604681595
transform -1 0 14812 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1604681595
transform -1 0 14812 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1604681595
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1604681595
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1604681595
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1604681595
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1604681595
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604681595
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_51
timestamp 1604681595
transform 1 0 5796 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_59
timestamp 1604681595
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_62
timestamp 1604681595
transform 1 0 6808 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_74
timestamp 1604681595
transform 1 0 7912 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_86
timestamp 1604681595
transform 1 0 9016 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_98
timestamp 1604681595
transform 1 0 10120 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604681595
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_110
timestamp 1604681595
transform 1 0 11224 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_123
timestamp 1604681595
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_135
timestamp 1604681595
transform 1 0 13524 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_143
timestamp 1604681595
transform 1 0 14260 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1604681595
transform -1 0 14812 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1604681595
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1604681595
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1604681595
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604681595
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_27
timestamp 1604681595
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_32
timestamp 1604681595
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_44
timestamp 1604681595
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_56
timestamp 1604681595
transform 1 0 6256 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_68
timestamp 1604681595
transform 1 0 7360 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_80
timestamp 1604681595
transform 1 0 8464 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604681595
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_93
timestamp 1604681595
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_105
timestamp 1604681595
transform 1 0 10764 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_117
timestamp 1604681595
transform 1 0 11868 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_129
timestamp 1604681595
transform 1 0 12972 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_141
timestamp 1604681595
transform 1 0 14076 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_145
timestamp 1604681595
transform 1 0 14444 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1604681595
transform -1 0 14812 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1604681595
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1604681595
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1604681595
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1604681595
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1604681595
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604681595
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_51
timestamp 1604681595
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_59
timestamp 1604681595
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_62
timestamp 1604681595
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_74
timestamp 1604681595
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_86
timestamp 1604681595
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_98
timestamp 1604681595
transform 1 0 10120 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604681595
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_110
timestamp 1604681595
transform 1 0 11224 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_123
timestamp 1604681595
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_135
timestamp 1604681595
transform 1 0 13524 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_143
timestamp 1604681595
transform 1 0 14260 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1604681595
transform -1 0 14812 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1604681595
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1604681595
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1604681595
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604681595
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_27
timestamp 1604681595
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_32
timestamp 1604681595
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604681595
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_44
timestamp 1604681595
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_56
timestamp 1604681595
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_63
timestamp 1604681595
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_75
timestamp 1604681595
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604681595
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_87
timestamp 1604681595
transform 1 0 9108 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_94
timestamp 1604681595
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604681595
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_106
timestamp 1604681595
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_118
timestamp 1604681595
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_125
timestamp 1604681595
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_137
timestamp 1604681595
transform 1 0 13708 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_145
timestamp 1604681595
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1604681595
transform -1 0 14812 0 -1 37536
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 36592 480 36712 6 ccff_head
port 0 nsew default input
rlabel metal3 s 15520 24896 16000 25016 6 ccff_tail
port 1 nsew default tristate
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[0]
port 2 nsew default input
rlabel metal2 s 12162 0 12218 480 6 chany_bottom_in[10]
port 3 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[11]
port 4 nsew default input
rlabel metal2 s 12990 0 13046 480 6 chany_bottom_in[12]
port 5 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[13]
port 6 nsew default input
rlabel metal2 s 13726 0 13782 480 6 chany_bottom_in[14]
port 7 nsew default input
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_in[15]
port 8 nsew default input
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_in[16]
port 9 nsew default input
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_in[17]
port 10 nsew default input
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_in[18]
port 11 nsew default input
rlabel metal2 s 15750 0 15806 480 6 chany_bottom_in[19]
port 12 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[1]
port 13 nsew default input
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_in[2]
port 14 nsew default input
rlabel metal2 s 9402 0 9458 480 6 chany_bottom_in[3]
port 15 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[4]
port 16 nsew default input
rlabel metal2 s 10138 0 10194 480 6 chany_bottom_in[5]
port 17 nsew default input
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_in[6]
port 18 nsew default input
rlabel metal2 s 10966 0 11022 480 6 chany_bottom_in[7]
port 19 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[8]
port 20 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_in[9]
port 21 nsew default input
rlabel metal2 s 202 0 258 480 6 chany_bottom_out[0]
port 22 nsew default tristate
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_out[10]
port 23 nsew default tristate
rlabel metal2 s 4526 0 4582 480 6 chany_bottom_out[11]
port 24 nsew default tristate
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_out[12]
port 25 nsew default tristate
rlabel metal2 s 5354 0 5410 480 6 chany_bottom_out[13]
port 26 nsew default tristate
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_out[14]
port 27 nsew default tristate
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_out[15]
port 28 nsew default tristate
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_out[16]
port 29 nsew default tristate
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_out[17]
port 30 nsew default tristate
rlabel metal2 s 7378 0 7434 480 6 chany_bottom_out[18]
port 31 nsew default tristate
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_out[19]
port 32 nsew default tristate
rlabel metal2 s 570 0 626 480 6 chany_bottom_out[1]
port 33 nsew default tristate
rlabel metal2 s 938 0 994 480 6 chany_bottom_out[2]
port 34 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_out[3]
port 35 nsew default tristate
rlabel metal2 s 1766 0 1822 480 6 chany_bottom_out[4]
port 36 nsew default tristate
rlabel metal2 s 2134 0 2190 480 6 chany_bottom_out[5]
port 37 nsew default tristate
rlabel metal2 s 2594 0 2650 480 6 chany_bottom_out[6]
port 38 nsew default tristate
rlabel metal2 s 2962 0 3018 480 6 chany_bottom_out[7]
port 39 nsew default tristate
rlabel metal2 s 3330 0 3386 480 6 chany_bottom_out[8]
port 40 nsew default tristate
rlabel metal2 s 3790 0 3846 480 6 chany_bottom_out[9]
port 41 nsew default tristate
rlabel metal2 s 8206 39520 8262 40000 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 12162 39520 12218 40000 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 12530 39520 12586 40000 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 12990 39520 13046 40000 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 13358 39520 13414 40000 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 13726 39520 13782 40000 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 14186 39520 14242 40000 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 14554 39520 14610 40000 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 14922 39520 14978 40000 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 15382 39520 15438 40000 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 15750 39520 15806 40000 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 8574 39520 8630 40000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 8942 39520 8998 40000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 9402 39520 9458 40000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 9770 39520 9826 40000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 10138 39520 10194 40000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 10598 39520 10654 40000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 10966 39520 11022 40000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 11334 39520 11390 40000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 11794 39520 11850 40000 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 202 39520 258 40000 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 4158 39520 4214 40000 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 4526 39520 4582 40000 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 4986 39520 5042 40000 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 5354 39520 5410 40000 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 5722 39520 5778 40000 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 6182 39520 6238 40000 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 6550 39520 6606 40000 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 6918 39520 6974 40000 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 7378 39520 7434 40000 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 7746 39520 7802 40000 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 570 39520 626 40000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 938 39520 994 40000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 1398 39520 1454 40000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 1766 39520 1822 40000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 2134 39520 2190 40000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 2594 39520 2650 40000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 2962 39520 3018 40000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 3330 39520 3386 40000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 3790 39520 3846 40000 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 gfpga_pad_EMBEDDED_IO_SOC_DIR
port 82 nsew default tristate
rlabel metal3 s 0 23264 480 23384 6 gfpga_pad_EMBEDDED_IO_SOC_IN
port 83 nsew default input
rlabel metal3 s 0 29928 480 30048 6 gfpga_pad_EMBEDDED_IO_SOC_OUT
port 84 nsew default tristate
rlabel metal3 s 0 9936 480 10056 6 left_grid_pin_0_
port 85 nsew default tristate
rlabel metal3 s 15520 14832 16000 14952 6 prog_clk
port 86 nsew default input
rlabel metal3 s 0 3272 480 3392 6 right_width_0_height_0__pin_0_
port 87 nsew default input
rlabel metal3 s 15520 4904 16000 5024 6 right_width_0_height_0__pin_1_lower
port 88 nsew default tristate
rlabel metal3 s 15520 34824 16000 34944 6 right_width_0_height_0__pin_1_upper
port 89 nsew default tristate
rlabel metal4 s 3611 2128 3931 37584 6 VPWR
port 90 nsew default input
rlabel metal4 s 6277 2128 6597 37584 6 VGND
port 91 nsew default input
<< properties >>
string FIXED_BBOX 0 0 16000 40000
<< end >>
