magic
tech sky130A
magscale 1 2
timestamp 1605173470
<< locali >>
rect 12725 19839 12759 20009
rect 22293 11543 22327 11713
rect 10977 8279 11011 8585
rect 15853 6103 15887 6205
<< viali >>
rect 10057 20961 10091 20995
rect 22549 20961 22583 20995
rect 10149 20893 10183 20927
rect 10241 20893 10275 20927
rect 19809 20893 19843 20927
rect 22293 20893 22327 20927
rect 8769 20757 8803 20791
rect 9689 20757 9723 20791
rect 23673 20757 23707 20791
rect 7113 20553 7147 20587
rect 10793 20553 10827 20587
rect 22385 20553 22419 20587
rect 27169 20553 27203 20587
rect 12173 20485 12207 20519
rect 22661 20485 22695 20519
rect 8769 20417 8803 20451
rect 12449 20417 12483 20451
rect 16129 20417 16163 20451
rect 19717 20417 19751 20451
rect 10977 20349 11011 20383
rect 15853 20349 15887 20383
rect 16589 20349 16623 20383
rect 25881 20349 25915 20383
rect 26985 20349 27019 20383
rect 8677 20281 8711 20315
rect 9036 20281 9070 20315
rect 11437 20281 11471 20315
rect 12716 20281 12750 20315
rect 19625 20281 19659 20315
rect 19962 20281 19996 20315
rect 10149 20213 10183 20247
rect 10425 20213 10459 20247
rect 13829 20213 13863 20247
rect 21097 20213 21131 20247
rect 26065 20213 26099 20247
rect 26525 20213 26559 20247
rect 27537 20213 27571 20247
rect 8033 20009 8067 20043
rect 8401 20009 8435 20043
rect 10517 20009 10551 20043
rect 12449 20009 12483 20043
rect 12725 20009 12759 20043
rect 21097 20009 21131 20043
rect 5897 19873 5931 19907
rect 8493 19873 8527 19907
rect 10885 19873 10919 19907
rect 13073 19873 13107 19907
rect 20913 19873 20947 19907
rect 22845 19873 22879 19907
rect 23112 19873 23146 19907
rect 5641 19805 5675 19839
rect 8585 19805 8619 19839
rect 10977 19805 11011 19839
rect 11069 19805 11103 19839
rect 12725 19805 12759 19839
rect 12817 19805 12851 19839
rect 14197 19737 14231 19771
rect 7021 19669 7055 19703
rect 10241 19669 10275 19703
rect 16221 19669 16255 19703
rect 19625 19669 19659 19703
rect 22109 19669 22143 19703
rect 24225 19669 24259 19703
rect 25513 19669 25547 19703
rect 27077 19669 27111 19703
rect 5733 19465 5767 19499
rect 10149 19465 10183 19499
rect 21281 19465 21315 19499
rect 23397 19465 23431 19499
rect 11161 19397 11195 19431
rect 25513 19397 25547 19431
rect 9321 19329 9355 19363
rect 9689 19329 9723 19363
rect 10793 19329 10827 19363
rect 16681 19329 16715 19363
rect 19625 19329 19659 19363
rect 22661 19329 22695 19363
rect 24501 19329 24535 19363
rect 26065 19329 26099 19363
rect 27629 19329 27663 19363
rect 6653 19261 6687 19295
rect 6837 19261 6871 19295
rect 9965 19261 9999 19295
rect 10517 19261 10551 19295
rect 16497 19261 16531 19295
rect 21833 19261 21867 19295
rect 22385 19261 22419 19295
rect 24317 19261 24351 19295
rect 27537 19261 27571 19295
rect 7104 19193 7138 19227
rect 13185 19193 13219 19227
rect 19533 19193 19567 19227
rect 19870 19193 19904 19227
rect 24409 19193 24443 19227
rect 25973 19193 26007 19227
rect 26985 19193 27019 19227
rect 6101 19125 6135 19159
rect 8217 19125 8251 19159
rect 8493 19125 8527 19159
rect 8861 19125 8895 19159
rect 10609 19125 10643 19159
rect 12817 19125 12851 19159
rect 15577 19125 15611 19159
rect 15945 19125 15979 19159
rect 16129 19125 16163 19159
rect 16589 19125 16623 19159
rect 21005 19125 21039 19159
rect 22017 19125 22051 19159
rect 22477 19125 22511 19159
rect 23121 19125 23155 19159
rect 23949 19125 23983 19159
rect 25329 19125 25363 19159
rect 25881 19125 25915 19159
rect 27077 19125 27111 19159
rect 27445 19125 27479 19159
rect 8493 18921 8527 18955
rect 10793 18921 10827 18955
rect 22109 18921 22143 18955
rect 23029 18921 23063 18955
rect 24133 18921 24167 18955
rect 24501 18921 24535 18955
rect 26525 18921 26559 18955
rect 27169 18921 27203 18955
rect 22845 18853 22879 18887
rect 4445 18785 4479 18819
rect 10057 18785 10091 18819
rect 15557 18785 15591 18819
rect 23397 18785 23431 18819
rect 23489 18785 23523 18819
rect 4537 18717 4571 18751
rect 4721 18717 4755 18751
rect 10149 18717 10183 18751
rect 10333 18717 10367 18751
rect 15301 18717 15335 18751
rect 19441 18717 19475 18751
rect 23581 18717 23615 18751
rect 8217 18649 8251 18683
rect 9689 18649 9723 18683
rect 4077 18581 4111 18615
rect 5089 18581 5123 18615
rect 6929 18581 6963 18615
rect 12817 18581 12851 18615
rect 16681 18581 16715 18615
rect 25605 18581 25639 18615
rect 5365 18377 5399 18411
rect 8125 18377 8159 18411
rect 9229 18377 9263 18411
rect 10793 18377 10827 18411
rect 18889 18377 18923 18411
rect 20453 18377 20487 18411
rect 23121 18377 23155 18411
rect 9689 18309 9723 18343
rect 21005 18309 21039 18343
rect 4997 18241 5031 18275
rect 5733 18241 5767 18275
rect 8585 18241 8619 18275
rect 8769 18241 8803 18275
rect 10241 18241 10275 18275
rect 14565 18241 14599 18275
rect 15853 18241 15887 18275
rect 16037 18241 16071 18275
rect 19901 18241 19935 18275
rect 19993 18241 20027 18275
rect 21557 18241 21591 18275
rect 2145 18173 2179 18207
rect 4721 18173 4755 18207
rect 8493 18173 8527 18207
rect 10149 18173 10183 18207
rect 11069 18173 11103 18207
rect 12817 18173 12851 18207
rect 13084 18173 13118 18207
rect 14933 18173 14967 18207
rect 19349 18173 19383 18207
rect 19809 18173 19843 18207
rect 21373 18173 21407 18207
rect 2053 18105 2087 18139
rect 2390 18105 2424 18139
rect 4169 18105 4203 18139
rect 8033 18105 8067 18139
rect 10057 18105 10091 18139
rect 11437 18105 11471 18139
rect 12725 18105 12759 18139
rect 15761 18105 15795 18139
rect 18613 18105 18647 18139
rect 23857 18105 23891 18139
rect 3525 18037 3559 18071
rect 4353 18037 4387 18071
rect 4813 18037 4847 18071
rect 9597 18037 9631 18071
rect 14197 18037 14231 18071
rect 15209 18037 15243 18071
rect 15393 18037 15427 18071
rect 16405 18037 16439 18071
rect 16957 18037 16991 18071
rect 19441 18037 19475 18071
rect 20913 18037 20947 18071
rect 21465 18037 21499 18071
rect 23489 18037 23523 18071
rect 2973 17833 3007 17867
rect 4537 17833 4571 17867
rect 8217 17833 8251 17867
rect 10241 17833 10275 17867
rect 13277 17833 13311 17867
rect 16221 17833 16255 17867
rect 19717 17833 19751 17867
rect 21097 17833 21131 17867
rect 23029 17833 23063 17867
rect 24869 17833 24903 17867
rect 3893 17765 3927 17799
rect 16681 17765 16715 17799
rect 25329 17765 25363 17799
rect 1409 17697 1443 17731
rect 4445 17697 4479 17731
rect 6368 17697 6402 17731
rect 9505 17697 9539 17731
rect 10609 17697 10643 17731
rect 10701 17697 10735 17731
rect 16589 17697 16623 17731
rect 19625 17697 19659 17731
rect 23397 17697 23431 17731
rect 24777 17697 24811 17731
rect 25237 17697 25271 17731
rect 4721 17629 4755 17663
rect 5181 17629 5215 17663
rect 6101 17629 6135 17663
rect 10885 17629 10919 17663
rect 13369 17629 13403 17663
rect 13553 17629 13587 17663
rect 16773 17629 16807 17663
rect 19901 17629 19935 17663
rect 22937 17629 22971 17663
rect 23489 17629 23523 17663
rect 23581 17629 23615 17663
rect 25421 17629 25455 17663
rect 15669 17561 15703 17595
rect 1593 17493 1627 17527
rect 2237 17493 2271 17527
rect 4077 17493 4111 17527
rect 7481 17493 7515 17527
rect 10149 17493 10183 17527
rect 12909 17493 12943 17527
rect 13921 17493 13955 17527
rect 16037 17493 16071 17527
rect 19165 17493 19199 17527
rect 19257 17493 19291 17527
rect 25881 17493 25915 17527
rect 2053 17289 2087 17323
rect 4353 17289 4387 17323
rect 4997 17289 5031 17323
rect 6193 17289 6227 17323
rect 10057 17289 10091 17323
rect 13369 17289 13403 17323
rect 14473 17289 14507 17323
rect 16681 17289 16715 17323
rect 16957 17289 16991 17323
rect 20177 17289 20211 17323
rect 22753 17289 22787 17323
rect 23673 17289 23707 17323
rect 27077 17289 27111 17323
rect 1593 17221 1627 17255
rect 4629 17221 4663 17255
rect 9597 17221 9631 17255
rect 11529 17221 11563 17255
rect 13001 17221 13035 17255
rect 17325 17221 17359 17255
rect 19165 17221 19199 17255
rect 20637 17221 20671 17255
rect 21281 17221 21315 17255
rect 24869 17221 24903 17255
rect 3157 17153 3191 17187
rect 3893 17153 3927 17187
rect 9229 17153 9263 17187
rect 10701 17153 10735 17187
rect 12265 17153 12299 17187
rect 14013 17153 14047 17187
rect 16221 17153 16255 17187
rect 19073 17153 19107 17187
rect 19809 17153 19843 17187
rect 24225 17153 24259 17187
rect 25513 17153 25547 17187
rect 1409 17085 1443 17119
rect 7205 17085 7239 17119
rect 19533 17085 19567 17119
rect 21373 17085 21407 17119
rect 21629 17085 21663 17119
rect 25697 17085 25731 17119
rect 25953 17085 25987 17119
rect 2789 17017 2823 17051
rect 3617 17017 3651 17051
rect 7450 17017 7484 17051
rect 10517 17017 10551 17051
rect 13737 17017 13771 17051
rect 14749 17017 14783 17051
rect 16037 17017 16071 17051
rect 18705 17017 18739 17051
rect 23489 17017 23523 17051
rect 24133 17017 24167 17051
rect 3249 16949 3283 16983
rect 3709 16949 3743 16983
rect 6469 16949 6503 16983
rect 7021 16949 7055 16983
rect 8585 16949 8619 16983
rect 9873 16949 9907 16983
rect 10425 16949 10459 16983
rect 11069 16949 11103 16983
rect 13829 16949 13863 16983
rect 15393 16949 15427 16983
rect 15577 16949 15611 16983
rect 15945 16949 15979 16983
rect 18337 16949 18371 16983
rect 19625 16949 19659 16983
rect 23121 16949 23155 16983
rect 24041 16949 24075 16983
rect 1593 16745 1627 16779
rect 3341 16745 3375 16779
rect 4077 16745 4111 16779
rect 4445 16745 4479 16779
rect 6837 16745 6871 16779
rect 7389 16745 7423 16779
rect 10149 16745 10183 16779
rect 13461 16745 13495 16779
rect 17509 16745 17543 16779
rect 19165 16745 19199 16779
rect 21373 16745 21407 16779
rect 23121 16745 23155 16779
rect 24133 16745 24167 16779
rect 24869 16745 24903 16779
rect 26709 16745 26743 16779
rect 6745 16677 6779 16711
rect 13001 16677 13035 16711
rect 13829 16677 13863 16711
rect 19073 16677 19107 16711
rect 25329 16677 25363 16711
rect 4537 16609 4571 16643
rect 10517 16609 10551 16643
rect 16129 16609 16163 16643
rect 16396 16609 16430 16643
rect 19533 16609 19567 16643
rect 19625 16609 19659 16643
rect 23673 16609 23707 16643
rect 25237 16609 25271 16643
rect 26525 16609 26559 16643
rect 4629 16541 4663 16575
rect 6929 16541 6963 16575
rect 10609 16541 10643 16575
rect 10793 16541 10827 16575
rect 13921 16541 13955 16575
rect 14013 16541 14047 16575
rect 19809 16541 19843 16575
rect 25513 16541 25547 16575
rect 25881 16473 25915 16507
rect 2053 16405 2087 16439
rect 3709 16405 3743 16439
rect 6377 16405 6411 16439
rect 15117 16405 15151 16439
rect 15669 16405 15703 16439
rect 24685 16405 24719 16439
rect 3617 16201 3651 16235
rect 4721 16201 4755 16235
rect 5089 16201 5123 16235
rect 6009 16201 6043 16235
rect 6469 16201 6503 16235
rect 7021 16201 7055 16235
rect 10517 16201 10551 16235
rect 10885 16201 10919 16235
rect 13277 16201 13311 16235
rect 15025 16201 15059 16235
rect 18613 16201 18647 16235
rect 20453 16201 20487 16235
rect 21005 16201 21039 16235
rect 23029 16201 23063 16235
rect 25053 16201 25087 16235
rect 25697 16201 25731 16235
rect 26893 16201 26927 16235
rect 2789 16133 2823 16167
rect 5365 16133 5399 16167
rect 10241 16133 10275 16167
rect 16129 16133 16163 16167
rect 19349 16133 19383 16167
rect 25881 16133 25915 16167
rect 4077 16065 4111 16099
rect 4261 16065 4295 16099
rect 13921 16065 13955 16099
rect 14381 16065 14415 16099
rect 15485 16065 15519 16099
rect 15577 16065 15611 16099
rect 20085 16065 20119 16099
rect 21557 16065 21591 16099
rect 23673 16065 23707 16099
rect 26341 16065 26375 16099
rect 26433 16065 26467 16099
rect 1409 15997 1443 16031
rect 9321 15997 9355 16031
rect 9597 15997 9631 16031
rect 14841 15997 14875 16031
rect 15393 15997 15427 16031
rect 19809 15997 19843 16031
rect 25329 15997 25363 16031
rect 1676 15929 1710 15963
rect 13829 15929 13863 15963
rect 19901 15929 19935 15963
rect 23918 15929 23952 15963
rect 3525 15861 3559 15895
rect 3985 15861 4019 15895
rect 9413 15861 9447 15895
rect 12817 15861 12851 15895
rect 13369 15861 13403 15895
rect 13737 15861 13771 15895
rect 16589 15861 16623 15895
rect 18889 15861 18923 15895
rect 19441 15861 19475 15895
rect 20821 15861 20855 15895
rect 21373 15861 21407 15895
rect 21465 15861 21499 15895
rect 23489 15861 23523 15895
rect 26249 15861 26283 15895
rect 4077 15657 4111 15691
rect 4445 15657 4479 15691
rect 4537 15657 4571 15691
rect 13277 15657 13311 15691
rect 14289 15657 14323 15691
rect 15577 15657 15611 15691
rect 15945 15657 15979 15691
rect 16037 15657 16071 15691
rect 18797 15657 18831 15691
rect 19717 15657 19751 15691
rect 21649 15657 21683 15691
rect 25329 15657 25363 15691
rect 3709 15589 3743 15623
rect 12142 15589 12176 15623
rect 14013 15589 14047 15623
rect 15117 15589 15151 15623
rect 19165 15589 19199 15623
rect 22906 15589 22940 15623
rect 5917 15521 5951 15555
rect 6276 15521 6310 15555
rect 9689 15521 9723 15555
rect 9956 15521 9990 15555
rect 13645 15521 13679 15555
rect 18061 15521 18095 15555
rect 19625 15521 19659 15555
rect 21833 15521 21867 15555
rect 22661 15521 22695 15555
rect 26525 15521 26559 15555
rect 1869 15453 1903 15487
rect 4721 15453 4755 15487
rect 6009 15453 6043 15487
rect 11897 15453 11931 15487
rect 16129 15453 16163 15487
rect 19809 15453 19843 15487
rect 1685 15385 1719 15419
rect 19257 15385 19291 15419
rect 21097 15385 21131 15419
rect 24869 15385 24903 15419
rect 2421 15317 2455 15351
rect 5733 15317 5767 15351
rect 7389 15317 7423 15351
rect 8401 15317 8435 15351
rect 11069 15317 11103 15351
rect 17877 15317 17911 15351
rect 24041 15317 24075 15351
rect 25973 15317 26007 15351
rect 26709 15317 26743 15351
rect 4445 15113 4479 15147
rect 4905 15113 4939 15147
rect 5733 15113 5767 15147
rect 6469 15113 6503 15147
rect 8309 15113 8343 15147
rect 10425 15113 10459 15147
rect 12633 15113 12667 15147
rect 13461 15113 13495 15147
rect 15945 15113 15979 15147
rect 16313 15113 16347 15147
rect 17877 15113 17911 15147
rect 18889 15113 18923 15147
rect 19165 15113 19199 15147
rect 20729 15113 20763 15147
rect 21741 15113 21775 15147
rect 22753 15113 22787 15147
rect 27353 15113 27387 15147
rect 15669 15045 15703 15079
rect 21005 15045 21039 15079
rect 23029 15045 23063 15079
rect 25145 15045 25179 15079
rect 2329 14977 2363 15011
rect 4169 14977 4203 15011
rect 8401 14977 8435 15011
rect 19349 14977 19383 15011
rect 25697 14977 25731 15011
rect 13553 14909 13587 14943
rect 13820 14909 13854 14943
rect 2237 14841 2271 14875
rect 2574 14841 2608 14875
rect 6101 14841 6135 14875
rect 8646 14841 8680 14875
rect 18521 14841 18555 14875
rect 19594 14841 19628 14875
rect 25605 14841 25639 14875
rect 25942 14841 25976 14875
rect 1685 14773 1719 14807
rect 3709 14773 3743 14807
rect 9781 14773 9815 14807
rect 10057 14773 10091 14807
rect 11897 14773 11931 14807
rect 14933 14773 14967 14807
rect 27077 14773 27111 14807
rect 1685 14569 1719 14603
rect 2237 14569 2271 14603
rect 8125 14569 8159 14603
rect 19809 14569 19843 14603
rect 20085 14569 20119 14603
rect 25513 14569 25547 14603
rect 2329 14501 2363 14535
rect 5816 14501 5850 14535
rect 10854 14501 10888 14535
rect 15761 14501 15795 14535
rect 5549 14433 5583 14467
rect 8309 14433 8343 14467
rect 10609 14433 10643 14467
rect 15669 14433 15703 14467
rect 18685 14433 18719 14467
rect 22293 14433 22327 14467
rect 22560 14433 22594 14467
rect 2513 14365 2547 14399
rect 15853 14365 15887 14399
rect 18429 14365 18463 14399
rect 1869 14229 1903 14263
rect 5089 14229 5123 14263
rect 6929 14229 6963 14263
rect 8677 14229 8711 14263
rect 11989 14229 12023 14263
rect 13645 14229 13679 14263
rect 15301 14229 15335 14263
rect 23673 14229 23707 14263
rect 2605 14025 2639 14059
rect 2973 14025 3007 14059
rect 6009 14025 6043 14059
rect 10977 14025 11011 14059
rect 14841 14025 14875 14059
rect 18889 14025 18923 14059
rect 19533 14025 19567 14059
rect 22385 14025 22419 14059
rect 22661 14025 22695 14059
rect 25329 14025 25363 14059
rect 4997 13957 5031 13991
rect 6377 13957 6411 13991
rect 16681 13957 16715 13991
rect 2053 13889 2087 13923
rect 2145 13889 2179 13923
rect 5457 13889 5491 13923
rect 5641 13889 5675 13923
rect 7757 13889 7791 13923
rect 9229 13889 9263 13923
rect 3433 13821 3467 13855
rect 4905 13821 4939 13855
rect 8125 13821 8159 13855
rect 9045 13821 9079 13855
rect 10701 13821 10735 13855
rect 15209 13821 15243 13855
rect 15301 13821 15335 13855
rect 16957 13821 16991 13855
rect 19717 13821 19751 13855
rect 19993 13821 20027 13855
rect 25513 13821 25547 13855
rect 25769 13821 25803 13855
rect 4537 13753 4571 13787
rect 5365 13753 5399 13787
rect 8401 13753 8435 13787
rect 8953 13753 8987 13787
rect 15546 13753 15580 13787
rect 1593 13685 1627 13719
rect 1961 13685 1995 13719
rect 8585 13685 8619 13719
rect 14381 13685 14415 13719
rect 18429 13685 18463 13719
rect 26893 13685 26927 13719
rect 1869 13481 1903 13515
rect 2881 13481 2915 13515
rect 3525 13481 3559 13515
rect 4445 13481 4479 13515
rect 4997 13481 5031 13515
rect 6101 13481 6135 13515
rect 6469 13481 6503 13515
rect 8033 13481 8067 13515
rect 15025 13481 15059 13515
rect 19165 13481 19199 13515
rect 4905 13413 4939 13447
rect 5641 13413 5675 13447
rect 11253 13413 11287 13447
rect 15761 13413 15795 13447
rect 23673 13413 23707 13447
rect 2237 13345 2271 13379
rect 2329 13345 2363 13379
rect 8401 13345 8435 13379
rect 14013 13345 14047 13379
rect 14105 13345 14139 13379
rect 15669 13345 15703 13379
rect 17785 13345 17819 13379
rect 18052 13345 18086 13379
rect 21281 13345 21315 13379
rect 23581 13345 23615 13379
rect 25237 13345 25271 13379
rect 2513 13277 2547 13311
rect 5089 13277 5123 13311
rect 6561 13277 6595 13311
rect 6653 13277 6687 13311
rect 8493 13277 8527 13311
rect 8677 13277 8711 13311
rect 11345 13277 11379 13311
rect 11437 13277 11471 13311
rect 12449 13277 12483 13311
rect 14197 13277 14231 13311
rect 15853 13277 15887 13311
rect 21373 13277 21407 13311
rect 21465 13277 21499 13311
rect 23765 13277 23799 13311
rect 24777 13277 24811 13311
rect 25329 13277 25363 13311
rect 25513 13277 25547 13311
rect 27077 13277 27111 13311
rect 1777 13209 1811 13243
rect 4537 13141 4571 13175
rect 9137 13141 9171 13175
rect 10149 13141 10183 13175
rect 10885 13141 10919 13175
rect 13645 13141 13679 13175
rect 15301 13141 15335 13175
rect 20913 13141 20947 13175
rect 23213 13141 23247 13175
rect 24317 13141 24351 13175
rect 24869 13141 24903 13175
rect 4629 12937 4663 12971
rect 5181 12937 5215 12971
rect 6285 12937 6319 12971
rect 7021 12937 7055 12971
rect 8585 12937 8619 12971
rect 11529 12937 11563 12971
rect 14841 12937 14875 12971
rect 15669 12937 15703 12971
rect 16313 12937 16347 12971
rect 22385 12937 22419 12971
rect 22937 12937 22971 12971
rect 23949 12937 23983 12971
rect 25513 12937 25547 12971
rect 26525 12937 26559 12971
rect 3433 12869 3467 12903
rect 4997 12869 5031 12903
rect 7757 12869 7791 12903
rect 10149 12869 10183 12903
rect 13001 12869 13035 12903
rect 16037 12869 16071 12903
rect 22017 12869 22051 12903
rect 23305 12869 23339 12903
rect 27077 12869 27111 12903
rect 2237 12801 2271 12835
rect 2421 12801 2455 12835
rect 3157 12801 3191 12835
rect 3985 12801 4019 12835
rect 5641 12801 5675 12835
rect 5825 12801 5859 12835
rect 9045 12801 9079 12835
rect 9137 12801 9171 12835
rect 10609 12801 10643 12835
rect 10701 12801 10735 12835
rect 17509 12801 17543 12835
rect 17877 12801 17911 12835
rect 18797 12801 18831 12835
rect 20361 12801 20395 12835
rect 24593 12801 24627 12835
rect 26065 12801 26099 12835
rect 27629 12801 27663 12835
rect 2145 12733 2179 12767
rect 3801 12733 3835 12767
rect 9689 12733 9723 12767
rect 10517 12733 10551 12767
rect 11161 12733 11195 12767
rect 13553 12733 13587 12767
rect 24317 12733 24351 12767
rect 25881 12733 25915 12767
rect 27537 12733 27571 12767
rect 1685 12665 1719 12699
rect 8953 12665 8987 12699
rect 10057 12665 10091 12699
rect 18521 12665 18555 12699
rect 19533 12665 19567 12699
rect 20269 12665 20303 12699
rect 20628 12665 20662 12699
rect 1777 12597 1811 12631
rect 2881 12597 2915 12631
rect 3893 12597 3927 12631
rect 5549 12597 5583 12631
rect 6653 12597 6687 12631
rect 8033 12597 8067 12631
rect 8493 12597 8527 12631
rect 13461 12597 13495 12631
rect 18153 12597 18187 12631
rect 18613 12597 18647 12631
rect 19165 12597 19199 12631
rect 21741 12597 21775 12631
rect 24409 12597 24443 12631
rect 24961 12597 24995 12631
rect 25421 12597 25455 12631
rect 25973 12597 26007 12631
rect 26893 12597 26927 12631
rect 27445 12597 27479 12631
rect 3893 12393 3927 12427
rect 4629 12393 4663 12427
rect 5641 12393 5675 12427
rect 8677 12393 8711 12427
rect 8953 12393 8987 12427
rect 9689 12393 9723 12427
rect 10793 12393 10827 12427
rect 11161 12393 11195 12427
rect 11437 12393 11471 12427
rect 11805 12393 11839 12427
rect 12449 12393 12483 12427
rect 14105 12393 14139 12427
rect 17417 12393 17451 12427
rect 17969 12393 18003 12427
rect 18521 12393 18555 12427
rect 20361 12393 20395 12427
rect 21097 12393 21131 12427
rect 21465 12393 21499 12427
rect 21925 12393 21959 12427
rect 23581 12393 23615 12427
rect 24501 12393 24535 12427
rect 24961 12393 24995 12427
rect 25881 12393 25915 12427
rect 27169 12393 27203 12427
rect 1838 12325 1872 12359
rect 3525 12325 3559 12359
rect 6101 12325 6135 12359
rect 15669 12325 15703 12359
rect 18889 12325 18923 12359
rect 24041 12325 24075 12359
rect 24869 12325 24903 12359
rect 1593 12257 1627 12291
rect 6009 12257 6043 12291
rect 10057 12257 10091 12291
rect 12817 12257 12851 12291
rect 13645 12257 13679 12291
rect 14657 12257 14691 12291
rect 15761 12257 15795 12291
rect 16681 12257 16715 12291
rect 17325 12257 17359 12291
rect 21833 12257 21867 12291
rect 26525 12257 26559 12291
rect 6193 12189 6227 12223
rect 10149 12189 10183 12223
rect 10241 12189 10275 12223
rect 11897 12189 11931 12223
rect 11989 12189 12023 12223
rect 12909 12189 12943 12223
rect 13001 12189 13035 12223
rect 14749 12189 14783 12223
rect 14933 12189 14967 12223
rect 15853 12189 15887 12223
rect 17601 12189 17635 12223
rect 18429 12189 18463 12223
rect 18981 12189 19015 12223
rect 19165 12189 19199 12223
rect 22109 12189 22143 12223
rect 23029 12189 23063 12223
rect 25053 12189 25087 12223
rect 2973 12053 3007 12087
rect 5273 12053 5307 12087
rect 14289 12053 14323 12087
rect 15301 12053 15335 12087
rect 16405 12053 16439 12087
rect 16957 12053 16991 12087
rect 24317 12053 24351 12087
rect 25513 12053 25547 12087
rect 26709 12053 26743 12087
rect 2421 11849 2455 11883
rect 2789 11849 2823 11883
rect 5641 11849 5675 11883
rect 6377 11849 6411 11883
rect 9781 11849 9815 11883
rect 11897 11849 11931 11883
rect 13001 11849 13035 11883
rect 15393 11849 15427 11883
rect 17049 11849 17083 11883
rect 17417 11849 17451 11883
rect 18521 11849 18555 11883
rect 20913 11849 20947 11883
rect 21465 11849 21499 11883
rect 24133 11849 24167 11883
rect 25329 11849 25363 11883
rect 26617 11849 26651 11883
rect 2053 11781 2087 11815
rect 6101 11781 6135 11815
rect 12725 11781 12759 11815
rect 16681 11781 16715 11815
rect 19625 11781 19659 11815
rect 24869 11781 24903 11815
rect 9045 11713 9079 11747
rect 10701 11713 10735 11747
rect 14565 11713 14599 11747
rect 16129 11713 16163 11747
rect 17785 11713 17819 11747
rect 19165 11713 19199 11747
rect 21925 11713 21959 11747
rect 22109 11713 22143 11747
rect 22293 11713 22327 11747
rect 25145 11713 25179 11747
rect 25789 11713 25823 11747
rect 25881 11713 25915 11747
rect 27445 11713 27479 11747
rect 1409 11645 1443 11679
rect 10517 11645 10551 11679
rect 14473 11645 14507 11679
rect 15945 11645 15979 11679
rect 9413 11577 9447 11611
rect 14381 11577 14415 11611
rect 16037 11577 16071 11611
rect 18981 11577 19015 11611
rect 19901 11577 19935 11611
rect 20637 11577 20671 11611
rect 21833 11577 21867 11611
rect 25697 11645 25731 11679
rect 27353 11645 27387 11679
rect 24501 11577 24535 11611
rect 27905 11577 27939 11611
rect 1593 11509 1627 11543
rect 10149 11509 10183 11543
rect 10609 11509 10643 11543
rect 11437 11509 11471 11543
rect 12265 11509 12299 11543
rect 13553 11509 13587 11543
rect 13829 11509 13863 11543
rect 14013 11509 14047 11543
rect 15577 11509 15611 11543
rect 18429 11509 18463 11543
rect 18889 11509 18923 11543
rect 21281 11509 21315 11543
rect 22293 11509 22327 11543
rect 22569 11509 22603 11543
rect 22937 11509 22971 11543
rect 26893 11509 26927 11543
rect 27261 11509 27295 11543
rect 2053 11305 2087 11339
rect 2329 11305 2363 11339
rect 2697 11305 2731 11339
rect 6561 11305 6595 11339
rect 9505 11305 9539 11339
rect 12449 11305 12483 11339
rect 14565 11305 14599 11339
rect 17049 11305 17083 11339
rect 18981 11305 19015 11339
rect 21557 11305 21591 11339
rect 23305 11305 23339 11339
rect 24593 11305 24627 11339
rect 24961 11305 24995 11339
rect 25421 11305 25455 11339
rect 27445 11305 27479 11339
rect 7634 11237 7668 11271
rect 9873 11237 9907 11271
rect 15853 11237 15887 11271
rect 22170 11237 22204 11271
rect 27077 11237 27111 11271
rect 1409 11169 1443 11203
rect 2513 11169 2547 11203
rect 5437 11169 5471 11203
rect 10425 11169 10459 11203
rect 13073 11169 13107 11203
rect 15025 11169 15059 11203
rect 15761 11169 15795 11203
rect 19349 11169 19383 11203
rect 26525 11169 26559 11203
rect 3157 11101 3191 11135
rect 5181 11101 5215 11135
rect 7389 11101 7423 11135
rect 10517 11101 10551 11135
rect 10609 11101 10643 11135
rect 12817 11101 12851 11135
rect 15945 11101 15979 11135
rect 16405 11101 16439 11135
rect 19441 11101 19475 11135
rect 19625 11101 19659 11135
rect 21925 11101 21959 11135
rect 1593 11033 1627 11067
rect 10057 11033 10091 11067
rect 15393 11033 15427 11067
rect 18889 11033 18923 11067
rect 26709 11033 26743 11067
rect 6929 10965 6963 10999
rect 8769 10965 8803 10999
rect 14197 10965 14231 10999
rect 18521 10965 18555 10999
rect 1593 10761 1627 10795
rect 2329 10761 2363 10795
rect 5273 10761 5307 10795
rect 6561 10761 6595 10795
rect 11069 10761 11103 10795
rect 12909 10761 12943 10795
rect 13737 10761 13771 10795
rect 14105 10761 14139 10795
rect 15945 10761 15979 10795
rect 18981 10761 19015 10795
rect 20821 10761 20855 10795
rect 22017 10761 22051 10795
rect 27353 10761 27387 10795
rect 5549 10693 5583 10727
rect 8493 10693 8527 10727
rect 9873 10693 9907 10727
rect 11805 10693 11839 10727
rect 15669 10693 15703 10727
rect 2421 10625 2455 10659
rect 7297 10625 7331 10659
rect 7389 10625 7423 10659
rect 9045 10625 9079 10659
rect 10517 10625 10551 10659
rect 10609 10625 10643 10659
rect 11437 10625 11471 10659
rect 13369 10625 13403 10659
rect 15117 10625 15151 10659
rect 16129 10625 16163 10659
rect 19625 10625 19659 10659
rect 8953 10557 8987 10591
rect 15025 10557 15059 10591
rect 19349 10557 19383 10591
rect 19993 10557 20027 10591
rect 26433 10557 26467 10591
rect 26985 10557 27019 10591
rect 27537 10557 27571 10591
rect 28089 10557 28123 10591
rect 2688 10489 2722 10523
rect 6285 10489 6319 10523
rect 7205 10489 7239 10523
rect 8861 10489 8895 10523
rect 10425 10489 10459 10523
rect 14933 10489 14967 10523
rect 18429 10489 18463 10523
rect 19441 10489 19475 10523
rect 22293 10489 22327 10523
rect 3801 10421 3835 10455
rect 6837 10421 6871 10455
rect 7849 10421 7883 10455
rect 8401 10421 8435 10455
rect 9505 10421 9539 10455
rect 10057 10421 10091 10455
rect 14381 10421 14415 10455
rect 14565 10421 14599 10455
rect 18889 10421 18923 10455
rect 20361 10421 20395 10455
rect 25237 10421 25271 10455
rect 26617 10421 26651 10455
rect 27721 10421 27755 10455
rect 3065 10217 3099 10251
rect 6377 10217 6411 10251
rect 7757 10217 7791 10251
rect 8585 10217 8619 10251
rect 8861 10217 8895 10251
rect 10057 10217 10091 10251
rect 10425 10217 10459 10251
rect 10609 10217 10643 10251
rect 11069 10217 11103 10251
rect 14013 10217 14047 10251
rect 14749 10217 14783 10251
rect 15117 10217 15151 10251
rect 15485 10217 15519 10251
rect 18981 10217 19015 10251
rect 25329 10217 25363 10251
rect 3525 10149 3559 10183
rect 10977 10149 11011 10183
rect 1409 10081 1443 10115
rect 2513 10081 2547 10115
rect 6745 10081 6779 10115
rect 8125 10081 8159 10115
rect 14105 10081 14139 10115
rect 18889 10081 18923 10115
rect 19349 10081 19383 10115
rect 25237 10081 25271 10115
rect 26525 10081 26559 10115
rect 6837 10013 6871 10047
rect 6929 10013 6963 10047
rect 11161 10013 11195 10047
rect 14197 10013 14231 10047
rect 19441 10013 19475 10047
rect 19625 10013 19659 10047
rect 25421 10013 25455 10047
rect 25881 10013 25915 10047
rect 1593 9877 1627 9911
rect 2697 9877 2731 9911
rect 7389 9877 7423 9911
rect 7941 9877 7975 9911
rect 12817 9877 12851 9911
rect 13645 9877 13679 9911
rect 18705 9877 18739 9911
rect 24685 9877 24719 9911
rect 24869 9877 24903 9911
rect 26709 9877 26743 9911
rect 2513 9673 2547 9707
rect 6009 9673 6043 9707
rect 8217 9673 8251 9707
rect 9781 9673 9815 9707
rect 10517 9673 10551 9707
rect 14197 9673 14231 9707
rect 14473 9673 14507 9707
rect 14841 9673 14875 9707
rect 18705 9673 18739 9707
rect 19809 9673 19843 9707
rect 22385 9673 22419 9707
rect 25421 9673 25455 9707
rect 26893 9673 26927 9707
rect 5549 9605 5583 9639
rect 6837 9605 6871 9639
rect 10609 9605 10643 9639
rect 2053 9537 2087 9571
rect 3525 9537 3559 9571
rect 7389 9537 7423 9571
rect 11161 9537 11195 9571
rect 11989 9537 12023 9571
rect 19441 9537 19475 9571
rect 26433 9537 26467 9571
rect 1409 9469 1443 9503
rect 3433 9469 3467 9503
rect 3792 9469 3826 9503
rect 6193 9469 6227 9503
rect 6653 9469 6687 9503
rect 7297 9469 7331 9503
rect 12817 9469 12851 9503
rect 15025 9469 15059 9503
rect 15281 9469 15315 9503
rect 21005 9469 21039 9503
rect 23673 9469 23707 9503
rect 25789 9469 25823 9503
rect 26249 9469 26283 9503
rect 5917 9401 5951 9435
rect 7205 9401 7239 9435
rect 7849 9401 7883 9435
rect 10149 9401 10183 9435
rect 11069 9401 11103 9435
rect 12725 9401 12759 9435
rect 13084 9401 13118 9435
rect 18981 9401 19015 9435
rect 20913 9401 20947 9435
rect 21250 9401 21284 9435
rect 23918 9401 23952 9435
rect 26341 9401 26375 9435
rect 1593 9333 1627 9367
rect 4905 9333 4939 9367
rect 10977 9333 11011 9367
rect 11621 9333 11655 9367
rect 16405 9333 16439 9367
rect 20453 9333 20487 9367
rect 23489 9333 23523 9367
rect 25053 9333 25087 9367
rect 25881 9333 25915 9367
rect 1685 9129 1719 9163
rect 3525 9129 3559 9163
rect 6101 9129 6135 9163
rect 6469 9129 6503 9163
rect 6837 9129 6871 9163
rect 11621 9129 11655 9163
rect 13737 9129 13771 9163
rect 14105 9129 14139 9163
rect 22477 9129 22511 9163
rect 22937 9129 22971 9163
rect 24225 9129 24259 9163
rect 24593 9129 24627 9163
rect 25237 9129 25271 9163
rect 2789 9061 2823 9095
rect 7297 9061 7331 9095
rect 10486 9061 10520 9095
rect 17386 9061 17420 9095
rect 21281 9061 21315 9095
rect 24685 9061 24719 9095
rect 7205 8993 7239 9027
rect 9137 8993 9171 9027
rect 15117 8993 15151 9027
rect 17141 8993 17175 9027
rect 19533 8993 19567 9027
rect 20729 8993 20763 9027
rect 22845 8993 22879 9027
rect 2329 8925 2363 8959
rect 2881 8925 2915 8959
rect 3065 8925 3099 8959
rect 7389 8925 7423 8959
rect 10241 8925 10275 8959
rect 21373 8925 21407 8959
rect 21465 8925 21499 8959
rect 23029 8925 23063 8959
rect 24777 8925 24811 8959
rect 25881 8925 25915 8959
rect 2421 8789 2455 8823
rect 4905 8789 4939 8823
rect 8953 8789 8987 8823
rect 12909 8789 12943 8823
rect 16497 8789 16531 8823
rect 18521 8789 18555 8823
rect 19349 8789 19383 8823
rect 20545 8789 20579 8823
rect 20913 8789 20947 8823
rect 23673 8789 23707 8823
rect 2513 8585 2547 8619
rect 3157 8585 3191 8619
rect 8585 8585 8619 8619
rect 10425 8585 10459 8619
rect 10701 8585 10735 8619
rect 10977 8585 11011 8619
rect 17417 8585 17451 8619
rect 17877 8585 17911 8619
rect 19349 8585 19383 8619
rect 21373 8585 21407 8619
rect 21649 8585 21683 8619
rect 24685 8585 24719 8619
rect 24961 8585 24995 8619
rect 26617 8585 26651 8619
rect 1593 8517 1627 8551
rect 3065 8517 3099 8551
rect 4813 8517 4847 8551
rect 2053 8449 2087 8483
rect 3617 8449 3651 8483
rect 3801 8449 3835 8483
rect 5365 8449 5399 8483
rect 6929 8449 6963 8483
rect 1409 8381 1443 8415
rect 3525 8381 3559 8415
rect 5181 8381 5215 8415
rect 9045 8381 9079 8415
rect 4629 8313 4663 8347
rect 6561 8313 6595 8347
rect 8953 8313 8987 8347
rect 9290 8313 9324 8347
rect 16865 8449 16899 8483
rect 17049 8449 17083 8483
rect 22845 8449 22879 8483
rect 19993 8381 20027 8415
rect 26433 8381 26467 8415
rect 26985 8381 27019 8415
rect 16313 8313 16347 8347
rect 16773 8313 16807 8347
rect 19901 8313 19935 8347
rect 20238 8313 20272 8347
rect 23213 8313 23247 8347
rect 4261 8245 4295 8279
rect 5273 8245 5307 8279
rect 7481 8245 7515 8279
rect 10977 8245 11011 8279
rect 11069 8245 11103 8279
rect 16405 8245 16439 8279
rect 22477 8245 22511 8279
rect 24225 8245 24259 8279
rect 3525 8041 3559 8075
rect 4905 8041 4939 8075
rect 6561 8041 6595 8075
rect 6929 8041 6963 8075
rect 16497 8041 16531 8075
rect 16957 8041 16991 8075
rect 18521 8041 18555 8075
rect 20545 8041 20579 8075
rect 21189 8041 21223 8075
rect 21557 8041 21591 8075
rect 22017 8041 22051 8075
rect 22477 8041 22511 8075
rect 23581 8041 23615 8075
rect 26709 8041 26743 8075
rect 2789 7973 2823 8007
rect 11406 7973 11440 8007
rect 17417 7973 17451 8007
rect 2881 7905 2915 7939
rect 5181 7905 5215 7939
rect 5448 7905 5482 7939
rect 17325 7905 17359 7939
rect 22385 7905 22419 7939
rect 23949 7905 23983 7939
rect 26525 7905 26559 7939
rect 3065 7837 3099 7871
rect 11161 7837 11195 7871
rect 13369 7837 13403 7871
rect 17509 7837 17543 7871
rect 22661 7837 22695 7871
rect 24041 7837 24075 7871
rect 24225 7837 24259 7871
rect 2329 7769 2363 7803
rect 23489 7769 23523 7803
rect 1685 7701 1719 7735
rect 2421 7701 2455 7735
rect 3893 7701 3927 7735
rect 9045 7701 9079 7735
rect 12541 7701 12575 7735
rect 18061 7701 18095 7735
rect 19993 7701 20027 7735
rect 25329 7701 25363 7735
rect 3065 7497 3099 7531
rect 4997 7497 5031 7531
rect 5181 7497 5215 7531
rect 16681 7497 16715 7531
rect 21833 7497 21867 7531
rect 22017 7497 22051 7531
rect 23121 7497 23155 7531
rect 24777 7497 24811 7531
rect 25145 7497 25179 7531
rect 26985 7497 27019 7531
rect 23673 7429 23707 7463
rect 26709 7429 26743 7463
rect 4169 7361 4203 7395
rect 4721 7361 4755 7395
rect 5825 7361 5859 7395
rect 12173 7361 12207 7395
rect 13093 7361 13127 7395
rect 14657 7361 14691 7395
rect 18613 7361 18647 7395
rect 21189 7361 21223 7395
rect 22477 7361 22511 7395
rect 22569 7361 22603 7395
rect 23489 7361 23523 7395
rect 24133 7361 24167 7395
rect 24317 7361 24351 7395
rect 1409 7293 1443 7327
rect 3985 7293 4019 7327
rect 6561 7293 6595 7327
rect 8309 7293 8343 7327
rect 14924 7293 14958 7327
rect 17785 7293 17819 7327
rect 18429 7293 18463 7327
rect 21557 7293 21591 7327
rect 24041 7293 24075 7327
rect 25329 7293 25363 7327
rect 25585 7293 25619 7327
rect 1676 7225 1710 7259
rect 5641 7225 5675 7259
rect 8217 7225 8251 7259
rect 8554 7225 8588 7259
rect 12909 7225 12943 7259
rect 14565 7225 14599 7259
rect 17325 7225 17359 7259
rect 18521 7225 18555 7259
rect 22385 7225 22419 7259
rect 2789 7157 2823 7191
rect 3433 7157 3467 7191
rect 3617 7157 3651 7191
rect 4077 7157 4111 7191
rect 5549 7157 5583 7191
rect 6285 7157 6319 7191
rect 6837 7157 6871 7191
rect 9689 7157 9723 7191
rect 10793 7157 10827 7191
rect 11253 7157 11287 7191
rect 11805 7157 11839 7191
rect 12449 7157 12483 7191
rect 12817 7157 12851 7191
rect 16037 7157 16071 7191
rect 16957 7157 16991 7191
rect 18061 7157 18095 7191
rect 1685 6953 1719 6987
rect 2329 6953 2363 6987
rect 2697 6953 2731 6987
rect 5733 6953 5767 6987
rect 13737 6953 13771 6987
rect 14657 6953 14691 6987
rect 22017 6953 22051 6987
rect 22477 6953 22511 6987
rect 23857 6953 23891 6987
rect 8401 6885 8435 6919
rect 12265 6885 12299 6919
rect 21281 6885 21315 6919
rect 22845 6885 22879 6919
rect 4353 6817 4387 6851
rect 5273 6817 5307 6851
rect 5825 6817 5859 6851
rect 12173 6817 12207 6851
rect 13829 6817 13863 6851
rect 16221 6817 16255 6851
rect 16865 6817 16899 6851
rect 16957 6817 16991 6851
rect 18429 6817 18463 6851
rect 18521 6817 18555 6851
rect 21373 6817 21407 6851
rect 26525 6817 26559 6851
rect 2789 6749 2823 6783
rect 2973 6749 3007 6783
rect 5917 6749 5951 6783
rect 6929 6749 6963 6783
rect 12357 6749 12391 6783
rect 14013 6749 14047 6783
rect 17141 6749 17175 6783
rect 18613 6749 18647 6783
rect 21557 6749 21591 6783
rect 23949 6749 23983 6783
rect 24133 6749 24167 6783
rect 5365 6681 5399 6715
rect 8861 6681 8895 6715
rect 11805 6681 11839 6715
rect 12909 6681 12943 6715
rect 18061 6681 18095 6715
rect 23489 6681 23523 6715
rect 26709 6681 26743 6715
rect 3617 6613 3651 6647
rect 10425 6613 10459 6647
rect 13369 6613 13403 6647
rect 16497 6613 16531 6647
rect 20913 6613 20947 6647
rect 24593 6613 24627 6647
rect 25329 6613 25363 6647
rect 1593 6409 1627 6443
rect 2053 6409 2087 6443
rect 2697 6409 2731 6443
rect 3065 6409 3099 6443
rect 5457 6409 5491 6443
rect 5825 6409 5859 6443
rect 6193 6409 6227 6443
rect 6561 6409 6595 6443
rect 10149 6409 10183 6443
rect 12265 6409 12299 6443
rect 12725 6409 12759 6443
rect 13829 6409 13863 6443
rect 18521 6409 18555 6443
rect 21741 6409 21775 6443
rect 22385 6409 22419 6443
rect 23489 6409 23523 6443
rect 26985 6409 27019 6443
rect 2329 6341 2363 6375
rect 8769 6341 8803 6375
rect 10333 6341 10367 6375
rect 11805 6341 11839 6375
rect 13461 6341 13495 6375
rect 17877 6341 17911 6375
rect 21373 6341 21407 6375
rect 23949 6341 23983 6375
rect 7297 6273 7331 6307
rect 7481 6273 7515 6307
rect 7849 6273 7883 6307
rect 9229 6273 9263 6307
rect 9321 6273 9355 6307
rect 10793 6273 10827 6307
rect 10885 6273 10919 6307
rect 16589 6273 16623 6307
rect 16681 6273 16715 6307
rect 18061 6273 18095 6307
rect 18889 6273 18923 6307
rect 21925 6273 21959 6307
rect 24317 6273 24351 6307
rect 1409 6205 1443 6239
rect 7205 6205 7239 6239
rect 8677 6205 8711 6239
rect 15853 6205 15887 6239
rect 17141 6205 17175 6239
rect 19717 6205 19751 6239
rect 26433 6205 26467 6239
rect 9137 6137 9171 6171
rect 9873 6137 9907 6171
rect 10701 6137 10735 6171
rect 15669 6137 15703 6171
rect 16497 6137 16531 6171
rect 19625 6137 19659 6171
rect 19984 6137 20018 6171
rect 26249 6137 26283 6171
rect 6837 6069 6871 6103
rect 14105 6069 14139 6103
rect 15853 6069 15887 6103
rect 15945 6069 15979 6103
rect 16129 6069 16163 6103
rect 21097 6069 21131 6103
rect 26617 6069 26651 6103
rect 6929 5865 6963 5899
rect 8861 5865 8895 5899
rect 10425 5865 10459 5899
rect 10885 5865 10919 5899
rect 11989 5865 12023 5899
rect 15945 5865 15979 5899
rect 16865 5865 16899 5899
rect 17049 5865 17083 5899
rect 17417 5865 17451 5899
rect 2044 5797 2078 5831
rect 5058 5797 5092 5831
rect 7389 5797 7423 5831
rect 10793 5797 10827 5831
rect 16589 5797 16623 5831
rect 19809 5797 19843 5831
rect 7481 5729 7515 5763
rect 12357 5729 12391 5763
rect 15853 5729 15887 5763
rect 21281 5729 21315 5763
rect 26525 5729 26559 5763
rect 1777 5661 1811 5695
rect 4813 5661 4847 5695
rect 7573 5661 7607 5695
rect 10977 5661 11011 5695
rect 12449 5661 12483 5695
rect 12633 5661 12667 5695
rect 16129 5661 16163 5695
rect 17509 5661 17543 5695
rect 17601 5661 17635 5695
rect 21373 5661 21407 5695
rect 21557 5661 21591 5695
rect 3157 5525 3191 5559
rect 6193 5525 6227 5559
rect 7021 5525 7055 5559
rect 11437 5525 11471 5559
rect 13001 5525 13035 5559
rect 13369 5525 13403 5559
rect 15485 5525 15519 5559
rect 20545 5525 20579 5559
rect 20913 5525 20947 5559
rect 23673 5525 23707 5559
rect 26709 5525 26743 5559
rect 1593 5321 1627 5355
rect 2329 5321 2363 5355
rect 2881 5321 2915 5355
rect 5181 5321 5215 5355
rect 6285 5321 6319 5355
rect 7941 5321 7975 5355
rect 9781 5321 9815 5355
rect 10701 5321 10735 5355
rect 12081 5321 12115 5355
rect 14013 5321 14047 5355
rect 16221 5321 16255 5355
rect 16589 5321 16623 5355
rect 17509 5321 17543 5355
rect 17785 5321 17819 5355
rect 21465 5321 21499 5355
rect 25053 5321 25087 5355
rect 26985 5321 27019 5355
rect 10425 5253 10459 5287
rect 17141 5253 17175 5287
rect 20269 5253 20303 5287
rect 2053 5185 2087 5219
rect 6653 5185 6687 5219
rect 7297 5185 7331 5219
rect 7389 5185 7423 5219
rect 10149 5185 10183 5219
rect 11345 5185 11379 5219
rect 14841 5185 14875 5219
rect 20913 5185 20947 5219
rect 21097 5185 21131 5219
rect 23673 5185 23707 5219
rect 1409 5117 1443 5151
rect 2973 5117 3007 5151
rect 7205 5117 7239 5151
rect 8217 5117 8251 5151
rect 12633 5117 12667 5151
rect 19993 5117 20027 5151
rect 20821 5117 20855 5151
rect 26433 5117 26467 5151
rect 3218 5049 3252 5083
rect 11069 5049 11103 5083
rect 12900 5049 12934 5083
rect 14749 5049 14783 5083
rect 15086 5049 15120 5083
rect 23918 5049 23952 5083
rect 26249 5049 26283 5083
rect 4353 4981 4387 5015
rect 4813 4981 4847 5015
rect 6837 4981 6871 5015
rect 11161 4981 11195 5015
rect 20453 4981 20487 5015
rect 23489 4981 23523 5015
rect 26617 4981 26651 5015
rect 1593 4777 1627 4811
rect 3157 4777 3191 4811
rect 3525 4777 3559 4811
rect 6377 4777 6411 4811
rect 7389 4777 7423 4811
rect 10793 4777 10827 4811
rect 11161 4777 11195 4811
rect 11345 4777 11379 4811
rect 12909 4777 12943 4811
rect 13277 4777 13311 4811
rect 13369 4777 13403 4811
rect 14841 4777 14875 4811
rect 15853 4777 15887 4811
rect 19625 4777 19659 4811
rect 20545 4777 20579 4811
rect 21925 4777 21959 4811
rect 2421 4709 2455 4743
rect 11805 4709 11839 4743
rect 15577 4709 15611 4743
rect 16304 4709 16338 4743
rect 22446 4709 22480 4743
rect 1409 4641 1443 4675
rect 2053 4641 2087 4675
rect 2513 4641 2547 4675
rect 4077 4641 4111 4675
rect 11713 4641 11747 4675
rect 16037 4641 16071 4675
rect 18061 4641 18095 4675
rect 21189 4641 21223 4675
rect 26525 4641 26559 4675
rect 6469 4573 6503 4607
rect 6561 4573 6595 4607
rect 7021 4573 7055 4607
rect 11989 4573 12023 4607
rect 12817 4573 12851 4607
rect 13553 4573 13587 4607
rect 19717 4573 19751 4607
rect 19901 4573 19935 4607
rect 22201 4573 22235 4607
rect 23581 4505 23615 4539
rect 2697 4437 2731 4471
rect 4261 4437 4295 4471
rect 6009 4437 6043 4471
rect 12449 4437 12483 4471
rect 17417 4437 17451 4471
rect 19257 4437 19291 4471
rect 26709 4437 26743 4471
rect 2329 4233 2363 4267
rect 5641 4233 5675 4267
rect 7481 4233 7515 4267
rect 11253 4233 11287 4267
rect 13277 4233 13311 4267
rect 13645 4233 13679 4267
rect 16405 4233 16439 4267
rect 17785 4233 17819 4267
rect 19809 4233 19843 4267
rect 21649 4233 21683 4267
rect 22845 4233 22879 4267
rect 27353 4233 27387 4267
rect 6101 4165 6135 4199
rect 11621 4165 11655 4199
rect 13001 4165 13035 4199
rect 16129 4165 16163 4199
rect 19441 4165 19475 4199
rect 21373 4165 21407 4199
rect 2697 4097 2731 4131
rect 3249 4097 3283 4131
rect 3341 4097 3375 4131
rect 4997 4097 5031 4131
rect 20177 4097 20211 4131
rect 20913 4097 20947 4131
rect 22293 4097 22327 4131
rect 22385 4097 22419 4131
rect 1409 4029 1443 4063
rect 4353 4029 4387 4063
rect 7205 4029 7239 4063
rect 7665 4029 7699 4063
rect 7921 4029 7955 4063
rect 9873 4029 9907 4063
rect 11897 4029 11931 4063
rect 18061 4029 18095 4063
rect 18317 4029 18351 4063
rect 20637 4029 20671 4063
rect 22201 4029 22235 4063
rect 26433 4029 26467 4063
rect 26985 4029 27019 4063
rect 27537 4029 27571 4063
rect 28089 4029 28123 4063
rect 10118 3961 10152 3995
rect 1593 3893 1627 3927
rect 2789 3893 2823 3927
rect 3157 3893 3191 3927
rect 4169 3893 4203 3927
rect 4537 3893 4571 3927
rect 6469 3893 6503 3927
rect 9045 3893 9079 3927
rect 9689 3893 9723 3927
rect 20269 3893 20303 3927
rect 20729 3893 20763 3927
rect 21833 3893 21867 3927
rect 26617 3893 26651 3927
rect 27721 3893 27755 3927
rect 1685 3689 1719 3723
rect 3341 3689 3375 3723
rect 5825 3689 5859 3723
rect 6929 3689 6963 3723
rect 9873 3689 9907 3723
rect 11437 3689 11471 3723
rect 19717 3689 19751 3723
rect 20361 3689 20395 3723
rect 21281 3689 21315 3723
rect 22293 3689 22327 3723
rect 2881 3621 2915 3655
rect 7297 3621 7331 3655
rect 21373 3621 21407 3655
rect 1961 3553 1995 3587
rect 4077 3553 4111 3587
rect 5733 3553 5767 3587
rect 15669 3553 15703 3587
rect 18061 3553 18095 3587
rect 26525 3553 26559 3587
rect 5917 3485 5951 3519
rect 7389 3485 7423 3519
rect 7481 3485 7515 3519
rect 15945 3485 15979 3519
rect 18153 3485 18187 3519
rect 18337 3485 18371 3519
rect 19349 3485 19383 3519
rect 21465 3485 21499 3519
rect 17693 3417 17727 3451
rect 20637 3417 20671 3451
rect 20913 3417 20947 3451
rect 2145 3349 2179 3383
rect 4261 3349 4295 3383
rect 5365 3349 5399 3383
rect 26709 3349 26743 3383
rect 2145 3145 2179 3179
rect 4445 3145 4479 3179
rect 4813 3145 4847 3179
rect 5825 3145 5859 3179
rect 6285 3145 6319 3179
rect 7573 3145 7607 3179
rect 13645 3145 13679 3179
rect 15301 3145 15335 3179
rect 15669 3145 15703 3179
rect 17325 3145 17359 3179
rect 21373 3145 21407 3179
rect 21741 3145 21775 3179
rect 27353 3145 27387 3179
rect 3341 3077 3375 3111
rect 5089 3077 5123 3111
rect 17785 3077 17819 3111
rect 21005 3077 21039 3111
rect 24961 3077 24995 3111
rect 3801 3009 3835 3043
rect 3893 3009 3927 3043
rect 6561 3009 6595 3043
rect 1409 2941 1443 2975
rect 4905 2941 4939 2975
rect 5457 2941 5491 2975
rect 6837 2941 6871 2975
rect 7941 2941 7975 2975
rect 12909 2941 12943 2975
rect 14473 2941 14507 2975
rect 18061 2941 18095 2975
rect 18797 2941 18831 2975
rect 23673 2941 23707 2975
rect 24317 2941 24351 2975
rect 24777 2941 24811 2975
rect 25329 2941 25363 2975
rect 26433 2941 26467 2975
rect 26985 2941 27019 2975
rect 27537 2941 27571 2975
rect 28089 2941 28123 2975
rect 1685 2873 1719 2907
rect 7113 2873 7147 2907
rect 13185 2873 13219 2907
rect 14749 2873 14783 2907
rect 18337 2873 18371 2907
rect 3249 2805 3283 2839
rect 3709 2805 3743 2839
rect 23857 2805 23891 2839
rect 26617 2805 26651 2839
rect 27721 2805 27755 2839
rect 1685 2601 1719 2635
rect 2973 2601 3007 2635
rect 5457 2601 5491 2635
rect 6285 2601 6319 2635
rect 7757 2601 7791 2635
rect 16865 2601 16899 2635
rect 17785 2601 17819 2635
rect 22569 2601 22603 2635
rect 3433 2533 3467 2567
rect 2145 2465 2179 2499
rect 3893 2465 3927 2499
rect 4353 2465 4387 2499
rect 5641 2465 5675 2499
rect 6929 2465 6963 2499
rect 8217 2465 8251 2499
rect 8953 2465 8987 2499
rect 9781 2465 9815 2499
rect 10517 2465 10551 2499
rect 12633 2465 12667 2499
rect 13369 2465 13403 2499
rect 16957 2465 16991 2499
rect 19165 2465 19199 2499
rect 19901 2465 19935 2499
rect 21833 2465 21867 2499
rect 24041 2465 24075 2499
rect 24777 2465 24811 2499
rect 25697 2465 25731 2499
rect 26249 2465 26283 2499
rect 2421 2397 2455 2431
rect 4629 2397 4663 2431
rect 7113 2397 7147 2431
rect 8493 2397 8527 2431
rect 10057 2397 10091 2431
rect 12817 2397 12851 2431
rect 17233 2397 17267 2431
rect 19441 2397 19475 2431
rect 22109 2397 22143 2431
rect 24225 2397 24259 2431
rect 5825 2261 5859 2295
rect 25881 2261 25915 2295
rect 27077 2261 27111 2295
<< metal1 >>
rect 3970 22176 3976 22228
rect 4028 22216 4034 22228
rect 12526 22216 12532 22228
rect 4028 22188 12532 22216
rect 4028 22176 4034 22188
rect 12526 22176 12532 22188
rect 12584 22176 12590 22228
rect 21450 22108 21456 22160
rect 21508 22148 21514 22160
rect 25774 22148 25780 22160
rect 21508 22120 25780 22148
rect 21508 22108 21514 22120
rect 25774 22108 25780 22120
rect 25832 22108 25838 22160
rect 1104 21786 28888 21808
rect 1104 21734 5982 21786
rect 6034 21734 6046 21786
rect 6098 21734 6110 21786
rect 6162 21734 6174 21786
rect 6226 21734 15982 21786
rect 16034 21734 16046 21786
rect 16098 21734 16110 21786
rect 16162 21734 16174 21786
rect 16226 21734 25982 21786
rect 26034 21734 26046 21786
rect 26098 21734 26110 21786
rect 26162 21734 26174 21786
rect 26226 21734 28888 21786
rect 1104 21712 28888 21734
rect 1104 21242 28888 21264
rect 1104 21190 10982 21242
rect 11034 21190 11046 21242
rect 11098 21190 11110 21242
rect 11162 21190 11174 21242
rect 11226 21190 20982 21242
rect 21034 21190 21046 21242
rect 21098 21190 21110 21242
rect 21162 21190 21174 21242
rect 21226 21190 28888 21242
rect 1104 21168 28888 21190
rect 10045 20995 10103 21001
rect 10045 20961 10057 20995
rect 10091 20992 10103 20995
rect 10502 20992 10508 21004
rect 10091 20964 10508 20992
rect 10091 20961 10103 20964
rect 10045 20955 10103 20961
rect 10502 20952 10508 20964
rect 10560 20952 10566 21004
rect 22370 20952 22376 21004
rect 22428 20992 22434 21004
rect 22537 20995 22595 21001
rect 22537 20992 22549 20995
rect 22428 20964 22549 20992
rect 22428 20952 22434 20964
rect 22537 20961 22549 20964
rect 22583 20961 22595 20995
rect 22537 20955 22595 20961
rect 10134 20924 10140 20936
rect 10095 20896 10140 20924
rect 10134 20884 10140 20896
rect 10192 20884 10198 20936
rect 10226 20884 10232 20936
rect 10284 20924 10290 20936
rect 10284 20896 10329 20924
rect 10284 20884 10290 20896
rect 19702 20884 19708 20936
rect 19760 20924 19766 20936
rect 19797 20927 19855 20933
rect 19797 20924 19809 20927
rect 19760 20896 19809 20924
rect 19760 20884 19766 20896
rect 19797 20893 19809 20896
rect 19843 20924 19855 20927
rect 22278 20924 22284 20936
rect 19843 20896 22284 20924
rect 19843 20893 19855 20896
rect 19797 20887 19855 20893
rect 22278 20884 22284 20896
rect 22336 20884 22342 20936
rect 4062 20816 4068 20868
rect 4120 20856 4126 20868
rect 9950 20856 9956 20868
rect 4120 20828 9956 20856
rect 4120 20816 4126 20828
rect 9950 20816 9956 20828
rect 10008 20816 10014 20868
rect 8754 20788 8760 20800
rect 8715 20760 8760 20788
rect 8754 20748 8760 20760
rect 8812 20748 8818 20800
rect 8846 20748 8852 20800
rect 8904 20788 8910 20800
rect 9677 20791 9735 20797
rect 9677 20788 9689 20791
rect 8904 20760 9689 20788
rect 8904 20748 8910 20760
rect 9677 20757 9689 20760
rect 9723 20757 9735 20791
rect 9677 20751 9735 20757
rect 22646 20748 22652 20800
rect 22704 20788 22710 20800
rect 23661 20791 23719 20797
rect 23661 20788 23673 20791
rect 22704 20760 23673 20788
rect 22704 20748 22710 20760
rect 23661 20757 23673 20760
rect 23707 20757 23719 20791
rect 23661 20751 23719 20757
rect 1104 20698 28888 20720
rect 1104 20646 5982 20698
rect 6034 20646 6046 20698
rect 6098 20646 6110 20698
rect 6162 20646 6174 20698
rect 6226 20646 15982 20698
rect 16034 20646 16046 20698
rect 16098 20646 16110 20698
rect 16162 20646 16174 20698
rect 16226 20646 25982 20698
rect 26034 20646 26046 20698
rect 26098 20646 26110 20698
rect 26162 20646 26174 20698
rect 26226 20646 28888 20698
rect 1104 20624 28888 20646
rect 7101 20587 7159 20593
rect 7101 20553 7113 20587
rect 7147 20584 7159 20587
rect 8202 20584 8208 20596
rect 7147 20556 8208 20584
rect 7147 20553 7159 20556
rect 7101 20547 7159 20553
rect 8202 20544 8208 20556
rect 8260 20544 8266 20596
rect 10134 20544 10140 20596
rect 10192 20584 10198 20596
rect 10781 20587 10839 20593
rect 10781 20584 10793 20587
rect 10192 20556 10793 20584
rect 10192 20544 10198 20556
rect 10781 20553 10793 20556
rect 10827 20553 10839 20587
rect 22370 20584 22376 20596
rect 22331 20556 22376 20584
rect 10781 20547 10839 20553
rect 22370 20544 22376 20556
rect 22428 20544 22434 20596
rect 27157 20587 27215 20593
rect 27157 20553 27169 20587
rect 27203 20584 27215 20587
rect 28258 20584 28264 20596
rect 27203 20556 28264 20584
rect 27203 20553 27215 20556
rect 27157 20547 27215 20553
rect 28258 20544 28264 20556
rect 28316 20544 28322 20596
rect 11606 20476 11612 20528
rect 11664 20516 11670 20528
rect 12161 20519 12219 20525
rect 12161 20516 12173 20519
rect 11664 20488 12173 20516
rect 11664 20476 11670 20488
rect 12161 20485 12173 20488
rect 12207 20485 12219 20519
rect 12161 20479 12219 20485
rect 8754 20448 8760 20460
rect 8715 20420 8760 20448
rect 8754 20408 8760 20420
rect 8812 20408 8818 20460
rect 10778 20340 10784 20392
rect 10836 20380 10842 20392
rect 10965 20383 11023 20389
rect 10965 20380 10977 20383
rect 10836 20352 10977 20380
rect 10836 20340 10842 20352
rect 10965 20349 10977 20352
rect 11011 20349 11023 20383
rect 10965 20343 11023 20349
rect 8665 20315 8723 20321
rect 8665 20281 8677 20315
rect 8711 20312 8723 20315
rect 9024 20315 9082 20321
rect 9024 20312 9036 20315
rect 8711 20284 9036 20312
rect 8711 20281 8723 20284
rect 8665 20275 8723 20281
rect 9024 20281 9036 20284
rect 9070 20312 9082 20315
rect 9306 20312 9312 20324
rect 9070 20284 9312 20312
rect 9070 20281 9082 20284
rect 9024 20275 9082 20281
rect 9306 20272 9312 20284
rect 9364 20272 9370 20324
rect 10502 20272 10508 20324
rect 10560 20312 10566 20324
rect 11425 20315 11483 20321
rect 11425 20312 11437 20315
rect 10560 20284 11437 20312
rect 10560 20272 10566 20284
rect 11425 20281 11437 20284
rect 11471 20281 11483 20315
rect 12176 20312 12204 20479
rect 22278 20476 22284 20528
rect 22336 20516 22342 20528
rect 22649 20519 22707 20525
rect 22649 20516 22661 20519
rect 22336 20488 22661 20516
rect 22336 20476 22342 20488
rect 22649 20485 22661 20488
rect 22695 20485 22707 20519
rect 22649 20479 22707 20485
rect 12434 20408 12440 20460
rect 12492 20448 12498 20460
rect 16114 20448 16120 20460
rect 12492 20420 12537 20448
rect 16075 20420 16120 20448
rect 12492 20408 12498 20420
rect 16114 20408 16120 20420
rect 16172 20408 16178 20460
rect 19702 20448 19708 20460
rect 19663 20420 19708 20448
rect 19702 20408 19708 20420
rect 19760 20408 19766 20460
rect 15838 20380 15844 20392
rect 15799 20352 15844 20380
rect 15838 20340 15844 20352
rect 15896 20380 15902 20392
rect 16577 20383 16635 20389
rect 16577 20380 16589 20383
rect 15896 20352 16589 20380
rect 15896 20340 15902 20352
rect 16577 20349 16589 20352
rect 16623 20349 16635 20383
rect 16577 20343 16635 20349
rect 25869 20383 25927 20389
rect 25869 20349 25881 20383
rect 25915 20380 25927 20383
rect 26973 20383 27031 20389
rect 25915 20352 26556 20380
rect 25915 20349 25927 20352
rect 25869 20343 25927 20349
rect 12704 20315 12762 20321
rect 12704 20312 12716 20315
rect 12176 20284 12716 20312
rect 11425 20275 11483 20281
rect 12704 20281 12716 20284
rect 12750 20281 12762 20315
rect 12704 20275 12762 20281
rect 19613 20315 19671 20321
rect 19613 20281 19625 20315
rect 19659 20312 19671 20315
rect 19950 20315 20008 20321
rect 19950 20312 19962 20315
rect 19659 20284 19962 20312
rect 19659 20281 19671 20284
rect 19613 20275 19671 20281
rect 19950 20281 19962 20284
rect 19996 20312 20008 20315
rect 20714 20312 20720 20324
rect 19996 20284 20720 20312
rect 19996 20281 20008 20284
rect 19950 20275 20008 20281
rect 20714 20272 20720 20284
rect 20772 20272 20778 20324
rect 9674 20204 9680 20256
rect 9732 20244 9738 20256
rect 10137 20247 10195 20253
rect 10137 20244 10149 20247
rect 9732 20216 10149 20244
rect 9732 20204 9738 20216
rect 10137 20213 10149 20216
rect 10183 20244 10195 20247
rect 10226 20244 10232 20256
rect 10183 20216 10232 20244
rect 10183 20213 10195 20216
rect 10137 20207 10195 20213
rect 10226 20204 10232 20216
rect 10284 20244 10290 20256
rect 10413 20247 10471 20253
rect 10413 20244 10425 20247
rect 10284 20216 10425 20244
rect 10284 20204 10290 20216
rect 10413 20213 10425 20216
rect 10459 20213 10471 20247
rect 13814 20244 13820 20256
rect 13775 20216 13820 20244
rect 10413 20207 10471 20213
rect 13814 20204 13820 20216
rect 13872 20204 13878 20256
rect 20806 20204 20812 20256
rect 20864 20244 20870 20256
rect 21085 20247 21143 20253
rect 21085 20244 21097 20247
rect 20864 20216 21097 20244
rect 20864 20204 20870 20216
rect 21085 20213 21097 20216
rect 21131 20213 21143 20247
rect 26050 20244 26056 20256
rect 26011 20216 26056 20244
rect 21085 20207 21143 20213
rect 26050 20204 26056 20216
rect 26108 20204 26114 20256
rect 26528 20253 26556 20352
rect 26973 20349 26985 20383
rect 27019 20380 27031 20383
rect 27019 20352 27476 20380
rect 27019 20349 27031 20352
rect 26973 20343 27031 20349
rect 27448 20256 27476 20352
rect 26513 20247 26571 20253
rect 26513 20213 26525 20247
rect 26559 20244 26571 20247
rect 27246 20244 27252 20256
rect 26559 20216 27252 20244
rect 26559 20213 26571 20216
rect 26513 20207 26571 20213
rect 27246 20204 27252 20216
rect 27304 20204 27310 20256
rect 27430 20204 27436 20256
rect 27488 20244 27494 20256
rect 27525 20247 27583 20253
rect 27525 20244 27537 20247
rect 27488 20216 27537 20244
rect 27488 20204 27494 20216
rect 27525 20213 27537 20216
rect 27571 20213 27583 20247
rect 27525 20207 27583 20213
rect 1104 20154 28888 20176
rect 1104 20102 10982 20154
rect 11034 20102 11046 20154
rect 11098 20102 11110 20154
rect 11162 20102 11174 20154
rect 11226 20102 20982 20154
rect 21034 20102 21046 20154
rect 21098 20102 21110 20154
rect 21162 20102 21174 20154
rect 21226 20102 28888 20154
rect 1104 20080 28888 20102
rect 8018 20040 8024 20052
rect 7979 20012 8024 20040
rect 8018 20000 8024 20012
rect 8076 20000 8082 20052
rect 8389 20043 8447 20049
rect 8389 20009 8401 20043
rect 8435 20040 8447 20043
rect 8478 20040 8484 20052
rect 8435 20012 8484 20040
rect 8435 20009 8447 20012
rect 8389 20003 8447 20009
rect 8478 20000 8484 20012
rect 8536 20040 8542 20052
rect 8846 20040 8852 20052
rect 8536 20012 8852 20040
rect 8536 20000 8542 20012
rect 8846 20000 8852 20012
rect 8904 20000 8910 20052
rect 10502 20040 10508 20052
rect 10463 20012 10508 20040
rect 10502 20000 10508 20012
rect 10560 20000 10566 20052
rect 12434 20040 12440 20052
rect 12395 20012 12440 20040
rect 12434 20000 12440 20012
rect 12492 20040 12498 20052
rect 12713 20043 12771 20049
rect 12713 20040 12725 20043
rect 12492 20012 12725 20040
rect 12492 20000 12498 20012
rect 12713 20009 12725 20012
rect 12759 20009 12771 20043
rect 12713 20003 12771 20009
rect 21085 20043 21143 20049
rect 21085 20009 21097 20043
rect 21131 20040 21143 20043
rect 21634 20040 21640 20052
rect 21131 20012 21640 20040
rect 21131 20009 21143 20012
rect 21085 20003 21143 20009
rect 21634 20000 21640 20012
rect 21692 20000 21698 20052
rect 5718 19864 5724 19916
rect 5776 19904 5782 19916
rect 5885 19907 5943 19913
rect 5885 19904 5897 19907
rect 5776 19876 5897 19904
rect 5776 19864 5782 19876
rect 5885 19873 5897 19876
rect 5931 19873 5943 19907
rect 5885 19867 5943 19873
rect 8481 19907 8539 19913
rect 8481 19873 8493 19907
rect 8527 19904 8539 19907
rect 8846 19904 8852 19916
rect 8527 19876 8852 19904
rect 8527 19873 8539 19876
rect 8481 19867 8539 19873
rect 8846 19864 8852 19876
rect 8904 19864 8910 19916
rect 10778 19864 10784 19916
rect 10836 19904 10842 19916
rect 10873 19907 10931 19913
rect 10873 19904 10885 19907
rect 10836 19876 10885 19904
rect 10836 19864 10842 19876
rect 10873 19873 10885 19876
rect 10919 19873 10931 19907
rect 10873 19867 10931 19873
rect 12434 19864 12440 19916
rect 12492 19904 12498 19916
rect 13061 19907 13119 19913
rect 13061 19904 13073 19907
rect 12492 19876 13073 19904
rect 12492 19864 12498 19876
rect 13061 19873 13073 19876
rect 13107 19904 13119 19907
rect 13814 19904 13820 19916
rect 13107 19876 13820 19904
rect 13107 19873 13119 19876
rect 13061 19867 13119 19873
rect 13814 19864 13820 19876
rect 13872 19864 13878 19916
rect 20806 19864 20812 19916
rect 20864 19904 20870 19916
rect 20901 19907 20959 19913
rect 20901 19904 20913 19907
rect 20864 19876 20913 19904
rect 20864 19864 20870 19876
rect 20901 19873 20913 19876
rect 20947 19873 20959 19907
rect 20901 19867 20959 19873
rect 22278 19864 22284 19916
rect 22336 19904 22342 19916
rect 22830 19904 22836 19916
rect 22336 19876 22836 19904
rect 22336 19864 22342 19876
rect 22830 19864 22836 19876
rect 22888 19864 22894 19916
rect 23106 19913 23112 19916
rect 23100 19904 23112 19913
rect 23067 19876 23112 19904
rect 23100 19867 23112 19876
rect 23106 19864 23112 19867
rect 23164 19864 23170 19916
rect 1670 19796 1676 19848
rect 1728 19836 1734 19848
rect 2682 19836 2688 19848
rect 1728 19808 2688 19836
rect 1728 19796 1734 19808
rect 2682 19796 2688 19808
rect 2740 19796 2746 19848
rect 5626 19836 5632 19848
rect 5587 19808 5632 19836
rect 5626 19796 5632 19808
rect 5684 19796 5690 19848
rect 8570 19836 8576 19848
rect 8531 19808 8576 19836
rect 8570 19796 8576 19808
rect 8628 19796 8634 19848
rect 10962 19836 10968 19848
rect 10923 19808 10968 19836
rect 10962 19796 10968 19808
rect 11020 19796 11026 19848
rect 11057 19839 11115 19845
rect 11057 19805 11069 19839
rect 11103 19805 11115 19839
rect 11057 19799 11115 19805
rect 10870 19728 10876 19780
rect 10928 19768 10934 19780
rect 11072 19768 11100 19799
rect 12618 19796 12624 19848
rect 12676 19836 12682 19848
rect 12713 19839 12771 19845
rect 12713 19836 12725 19839
rect 12676 19808 12725 19836
rect 12676 19796 12682 19808
rect 12713 19805 12725 19808
rect 12759 19836 12771 19839
rect 12805 19839 12863 19845
rect 12805 19836 12817 19839
rect 12759 19808 12817 19836
rect 12759 19805 12771 19808
rect 12713 19799 12771 19805
rect 12805 19805 12817 19808
rect 12851 19805 12863 19839
rect 12805 19799 12863 19805
rect 14182 19768 14188 19780
rect 10928 19740 11100 19768
rect 14143 19740 14188 19768
rect 10928 19728 10934 19740
rect 14182 19728 14188 19740
rect 14240 19728 14246 19780
rect 7009 19703 7067 19709
rect 7009 19669 7021 19703
rect 7055 19700 7067 19703
rect 7098 19700 7104 19712
rect 7055 19672 7104 19700
rect 7055 19669 7067 19672
rect 7009 19663 7067 19669
rect 7098 19660 7104 19672
rect 7156 19660 7162 19712
rect 10229 19703 10287 19709
rect 10229 19669 10241 19703
rect 10275 19700 10287 19703
rect 10594 19700 10600 19712
rect 10275 19672 10600 19700
rect 10275 19669 10287 19672
rect 10229 19663 10287 19669
rect 10594 19660 10600 19672
rect 10652 19660 10658 19712
rect 16209 19703 16267 19709
rect 16209 19669 16221 19703
rect 16255 19700 16267 19703
rect 16482 19700 16488 19712
rect 16255 19672 16488 19700
rect 16255 19669 16267 19672
rect 16209 19663 16267 19669
rect 16482 19660 16488 19672
rect 16540 19660 16546 19712
rect 19610 19700 19616 19712
rect 19571 19672 19616 19700
rect 19610 19660 19616 19672
rect 19668 19660 19674 19712
rect 22094 19660 22100 19712
rect 22152 19700 22158 19712
rect 24210 19700 24216 19712
rect 22152 19672 22197 19700
rect 24171 19672 24216 19700
rect 22152 19660 22158 19672
rect 24210 19660 24216 19672
rect 24268 19660 24274 19712
rect 25406 19660 25412 19712
rect 25464 19700 25470 19712
rect 25501 19703 25559 19709
rect 25501 19700 25513 19703
rect 25464 19672 25513 19700
rect 25464 19660 25470 19672
rect 25501 19669 25513 19672
rect 25547 19700 25559 19703
rect 27065 19703 27123 19709
rect 27065 19700 27077 19703
rect 25547 19672 27077 19700
rect 25547 19669 25559 19672
rect 25501 19663 25559 19669
rect 27065 19669 27077 19672
rect 27111 19669 27123 19703
rect 27065 19663 27123 19669
rect 1104 19610 28888 19632
rect 1104 19558 5982 19610
rect 6034 19558 6046 19610
rect 6098 19558 6110 19610
rect 6162 19558 6174 19610
rect 6226 19558 15982 19610
rect 16034 19558 16046 19610
rect 16098 19558 16110 19610
rect 16162 19558 16174 19610
rect 16226 19558 25982 19610
rect 26034 19558 26046 19610
rect 26098 19558 26110 19610
rect 26162 19558 26174 19610
rect 26226 19558 28888 19610
rect 1104 19536 28888 19558
rect 5718 19496 5724 19508
rect 5679 19468 5724 19496
rect 5718 19456 5724 19468
rect 5776 19456 5782 19508
rect 10134 19496 10140 19508
rect 10095 19468 10140 19496
rect 10134 19456 10140 19468
rect 10192 19456 10198 19508
rect 20806 19456 20812 19508
rect 20864 19496 20870 19508
rect 21269 19499 21327 19505
rect 21269 19496 21281 19499
rect 20864 19468 21281 19496
rect 20864 19456 20870 19468
rect 21269 19465 21281 19468
rect 21315 19465 21327 19499
rect 21269 19459 21327 19465
rect 22370 19456 22376 19508
rect 22428 19496 22434 19508
rect 23385 19499 23443 19505
rect 23385 19496 23397 19499
rect 22428 19468 23397 19496
rect 22428 19456 22434 19468
rect 23385 19465 23397 19468
rect 23431 19496 23443 19499
rect 23566 19496 23572 19508
rect 23431 19468 23572 19496
rect 23431 19465 23443 19468
rect 23385 19459 23443 19465
rect 23566 19456 23572 19468
rect 23624 19496 23630 19508
rect 24210 19496 24216 19508
rect 23624 19468 24216 19496
rect 23624 19456 23630 19468
rect 24210 19456 24216 19468
rect 24268 19456 24274 19508
rect 10042 19388 10048 19440
rect 10100 19428 10106 19440
rect 10962 19428 10968 19440
rect 10100 19400 10968 19428
rect 10100 19388 10106 19400
rect 10962 19388 10968 19400
rect 11020 19428 11026 19440
rect 11149 19431 11207 19437
rect 11149 19428 11161 19431
rect 11020 19400 11161 19428
rect 11020 19388 11026 19400
rect 11149 19397 11161 19400
rect 11195 19397 11207 19431
rect 11149 19391 11207 19397
rect 9306 19360 9312 19372
rect 6656 19332 6960 19360
rect 9219 19332 9312 19360
rect 6656 19301 6684 19332
rect 6641 19295 6699 19301
rect 6641 19261 6653 19295
rect 6687 19261 6699 19295
rect 6822 19292 6828 19304
rect 6783 19264 6828 19292
rect 6641 19255 6699 19261
rect 6822 19252 6828 19264
rect 6880 19252 6886 19304
rect 6932 19292 6960 19332
rect 9306 19320 9312 19332
rect 9364 19360 9370 19372
rect 9677 19363 9735 19369
rect 9677 19360 9689 19363
rect 9364 19332 9689 19360
rect 9364 19320 9370 19332
rect 9677 19329 9689 19332
rect 9723 19360 9735 19363
rect 10781 19363 10839 19369
rect 10781 19360 10793 19363
rect 9723 19332 10793 19360
rect 9723 19329 9735 19332
rect 9677 19323 9735 19329
rect 10781 19329 10793 19332
rect 10827 19360 10839 19363
rect 10870 19360 10876 19372
rect 10827 19332 10876 19360
rect 10827 19329 10839 19332
rect 10781 19323 10839 19329
rect 10870 19320 10876 19332
rect 10928 19320 10934 19372
rect 16669 19363 16727 19369
rect 16669 19360 16681 19363
rect 15580 19332 16681 19360
rect 9950 19292 9956 19304
rect 6932 19264 7144 19292
rect 9911 19264 9956 19292
rect 5718 19184 5724 19236
rect 5776 19224 5782 19236
rect 7116 19233 7144 19264
rect 9950 19252 9956 19264
rect 10008 19292 10014 19304
rect 10502 19292 10508 19304
rect 10008 19264 10508 19292
rect 10008 19252 10014 19264
rect 10502 19252 10508 19264
rect 10560 19252 10566 19304
rect 7092 19227 7150 19233
rect 5776 19196 7052 19224
rect 5776 19184 5782 19196
rect 5626 19116 5632 19168
rect 5684 19156 5690 19168
rect 6089 19159 6147 19165
rect 6089 19156 6101 19159
rect 5684 19128 6101 19156
rect 5684 19116 5690 19128
rect 6089 19125 6101 19128
rect 6135 19156 6147 19159
rect 6914 19156 6920 19168
rect 6135 19128 6920 19156
rect 6135 19125 6147 19128
rect 6089 19119 6147 19125
rect 6914 19116 6920 19128
rect 6972 19116 6978 19168
rect 7024 19156 7052 19196
rect 7092 19193 7104 19227
rect 7138 19224 7150 19227
rect 8018 19224 8024 19236
rect 7138 19196 8024 19224
rect 7138 19193 7150 19196
rect 7092 19187 7150 19193
rect 8018 19184 8024 19196
rect 8076 19184 8082 19236
rect 12618 19184 12624 19236
rect 12676 19224 12682 19236
rect 13173 19227 13231 19233
rect 13173 19224 13185 19227
rect 12676 19196 13185 19224
rect 12676 19184 12682 19196
rect 13173 19193 13185 19196
rect 13219 19193 13231 19227
rect 13173 19187 13231 19193
rect 8205 19159 8263 19165
rect 8205 19156 8217 19159
rect 7024 19128 8217 19156
rect 8205 19125 8217 19128
rect 8251 19156 8263 19159
rect 8481 19159 8539 19165
rect 8481 19156 8493 19159
rect 8251 19128 8493 19156
rect 8251 19125 8263 19128
rect 8205 19119 8263 19125
rect 8481 19125 8493 19128
rect 8527 19156 8539 19159
rect 8570 19156 8576 19168
rect 8527 19128 8576 19156
rect 8527 19125 8539 19128
rect 8481 19119 8539 19125
rect 8570 19116 8576 19128
rect 8628 19116 8634 19168
rect 8846 19156 8852 19168
rect 8807 19128 8852 19156
rect 8846 19116 8852 19128
rect 8904 19116 8910 19168
rect 10594 19156 10600 19168
rect 10555 19128 10600 19156
rect 10594 19116 10600 19128
rect 10652 19116 10658 19168
rect 12434 19116 12440 19168
rect 12492 19156 12498 19168
rect 12805 19159 12863 19165
rect 12805 19156 12817 19159
rect 12492 19128 12817 19156
rect 12492 19116 12498 19128
rect 12805 19125 12817 19128
rect 12851 19125 12863 19159
rect 12805 19119 12863 19125
rect 15194 19116 15200 19168
rect 15252 19156 15258 19168
rect 15580 19165 15608 19332
rect 16669 19329 16681 19332
rect 16715 19329 16727 19363
rect 19610 19360 19616 19372
rect 19571 19332 19616 19360
rect 16669 19323 16727 19329
rect 19610 19320 19616 19332
rect 19668 19320 19674 19372
rect 22646 19360 22652 19372
rect 22020 19332 22652 19360
rect 16485 19295 16543 19301
rect 16485 19292 16497 19295
rect 15764 19264 16497 19292
rect 15764 19168 15792 19264
rect 16485 19261 16497 19264
rect 16531 19261 16543 19295
rect 16485 19255 16543 19261
rect 20714 19252 20720 19304
rect 20772 19292 20778 19304
rect 21821 19295 21879 19301
rect 21821 19292 21833 19295
rect 20772 19264 21833 19292
rect 20772 19252 20778 19264
rect 21821 19261 21833 19264
rect 21867 19292 21879 19295
rect 22020 19292 22048 19332
rect 22646 19320 22652 19332
rect 22704 19320 22710 19372
rect 24228 19360 24256 19456
rect 25498 19428 25504 19440
rect 25459 19400 25504 19428
rect 25498 19388 25504 19400
rect 25556 19388 25562 19440
rect 24489 19363 24547 19369
rect 24489 19360 24501 19363
rect 24228 19332 24501 19360
rect 24489 19329 24501 19332
rect 24535 19329 24547 19363
rect 24489 19323 24547 19329
rect 24946 19320 24952 19372
rect 25004 19360 25010 19372
rect 25222 19360 25228 19372
rect 25004 19332 25228 19360
rect 25004 19320 25010 19332
rect 25222 19320 25228 19332
rect 25280 19320 25286 19372
rect 25406 19320 25412 19372
rect 25464 19360 25470 19372
rect 26053 19363 26111 19369
rect 26053 19360 26065 19363
rect 25464 19332 26065 19360
rect 25464 19320 25470 19332
rect 26053 19329 26065 19332
rect 26099 19360 26111 19363
rect 27617 19363 27675 19369
rect 27617 19360 27629 19363
rect 26099 19332 27629 19360
rect 26099 19329 26111 19332
rect 26053 19323 26111 19329
rect 27617 19329 27629 19332
rect 27663 19329 27675 19363
rect 27617 19323 27675 19329
rect 21867 19264 22048 19292
rect 21867 19261 21879 19264
rect 21821 19255 21879 19261
rect 22094 19252 22100 19304
rect 22152 19292 22158 19304
rect 22373 19295 22431 19301
rect 22373 19292 22385 19295
rect 22152 19264 22385 19292
rect 22152 19252 22158 19264
rect 22373 19261 22385 19264
rect 22419 19261 22431 19295
rect 22373 19255 22431 19261
rect 24305 19295 24363 19301
rect 24305 19261 24317 19295
rect 24351 19292 24363 19295
rect 24578 19292 24584 19304
rect 24351 19264 24584 19292
rect 24351 19261 24363 19264
rect 24305 19255 24363 19261
rect 15838 19184 15844 19236
rect 15896 19224 15902 19236
rect 19521 19227 19579 19233
rect 15896 19196 16160 19224
rect 15896 19184 15902 19196
rect 15565 19159 15623 19165
rect 15565 19156 15577 19159
rect 15252 19128 15577 19156
rect 15252 19116 15258 19128
rect 15565 19125 15577 19128
rect 15611 19125 15623 19159
rect 15565 19119 15623 19125
rect 15746 19116 15752 19168
rect 15804 19156 15810 19168
rect 16132 19165 16160 19196
rect 19521 19193 19533 19227
rect 19567 19224 19579 19227
rect 19858 19227 19916 19233
rect 19858 19224 19870 19227
rect 19567 19196 19870 19224
rect 19567 19193 19579 19196
rect 19521 19187 19579 19193
rect 19858 19193 19870 19196
rect 19904 19224 19916 19227
rect 19978 19224 19984 19236
rect 19904 19196 19984 19224
rect 19904 19193 19916 19196
rect 19858 19187 19916 19193
rect 19978 19184 19984 19196
rect 20036 19184 20042 19236
rect 22388 19224 22416 19255
rect 24578 19252 24584 19264
rect 24636 19292 24642 19304
rect 27522 19292 27528 19304
rect 24636 19264 26832 19292
rect 27483 19264 27528 19292
rect 24636 19252 24642 19264
rect 22388 19196 23980 19224
rect 15933 19159 15991 19165
rect 15933 19156 15945 19159
rect 15804 19128 15945 19156
rect 15804 19116 15810 19128
rect 15933 19125 15945 19128
rect 15979 19125 15991 19159
rect 15933 19119 15991 19125
rect 16117 19159 16175 19165
rect 16117 19125 16129 19159
rect 16163 19125 16175 19159
rect 16117 19119 16175 19125
rect 16482 19116 16488 19168
rect 16540 19156 16546 19168
rect 16577 19159 16635 19165
rect 16577 19156 16589 19159
rect 16540 19128 16589 19156
rect 16540 19116 16546 19128
rect 16577 19125 16589 19128
rect 16623 19156 16635 19159
rect 16850 19156 16856 19168
rect 16623 19128 16856 19156
rect 16623 19125 16635 19128
rect 16577 19119 16635 19125
rect 16850 19116 16856 19128
rect 16908 19116 16914 19168
rect 20993 19159 21051 19165
rect 20993 19125 21005 19159
rect 21039 19156 21051 19159
rect 21266 19156 21272 19168
rect 21039 19128 21272 19156
rect 21039 19125 21051 19128
rect 20993 19119 21051 19125
rect 21266 19116 21272 19128
rect 21324 19116 21330 19168
rect 21726 19116 21732 19168
rect 21784 19156 21790 19168
rect 22005 19159 22063 19165
rect 22005 19156 22017 19159
rect 21784 19128 22017 19156
rect 21784 19116 21790 19128
rect 22005 19125 22017 19128
rect 22051 19125 22063 19159
rect 22462 19156 22468 19168
rect 22423 19128 22468 19156
rect 22005 19119 22063 19125
rect 22462 19116 22468 19128
rect 22520 19116 22526 19168
rect 23106 19156 23112 19168
rect 23067 19128 23112 19156
rect 23106 19116 23112 19128
rect 23164 19116 23170 19168
rect 23952 19165 23980 19196
rect 24118 19184 24124 19236
rect 24176 19224 24182 19236
rect 24397 19227 24455 19233
rect 24397 19224 24409 19227
rect 24176 19196 24409 19224
rect 24176 19184 24182 19196
rect 24397 19193 24409 19196
rect 24443 19224 24455 19227
rect 25498 19224 25504 19236
rect 24443 19196 25504 19224
rect 24443 19193 24455 19196
rect 24397 19187 24455 19193
rect 25498 19184 25504 19196
rect 25556 19184 25562 19236
rect 25682 19184 25688 19236
rect 25740 19224 25746 19236
rect 25961 19227 26019 19233
rect 25961 19224 25973 19227
rect 25740 19196 25973 19224
rect 25740 19184 25746 19196
rect 25961 19193 25973 19196
rect 26007 19193 26019 19227
rect 25961 19187 26019 19193
rect 23937 19159 23995 19165
rect 23937 19125 23949 19159
rect 23983 19125 23995 19159
rect 25314 19156 25320 19168
rect 25275 19128 25320 19156
rect 23937 19119 23995 19125
rect 25314 19116 25320 19128
rect 25372 19156 25378 19168
rect 25869 19159 25927 19165
rect 25869 19156 25881 19159
rect 25372 19128 25881 19156
rect 25372 19116 25378 19128
rect 25869 19125 25881 19128
rect 25915 19156 25927 19159
rect 26418 19156 26424 19168
rect 25915 19128 26424 19156
rect 25915 19125 25927 19128
rect 25869 19119 25927 19125
rect 26418 19116 26424 19128
rect 26476 19116 26482 19168
rect 26804 19156 26832 19264
rect 27522 19252 27528 19264
rect 27580 19252 27586 19304
rect 26970 19224 26976 19236
rect 26883 19196 26976 19224
rect 26970 19184 26976 19196
rect 27028 19224 27034 19236
rect 27540 19224 27568 19252
rect 27028 19196 27568 19224
rect 27028 19184 27034 19196
rect 27065 19159 27123 19165
rect 27065 19156 27077 19159
rect 26804 19128 27077 19156
rect 27065 19125 27077 19128
rect 27111 19125 27123 19159
rect 27065 19119 27123 19125
rect 27154 19116 27160 19168
rect 27212 19156 27218 19168
rect 27433 19159 27491 19165
rect 27433 19156 27445 19159
rect 27212 19128 27445 19156
rect 27212 19116 27218 19128
rect 27433 19125 27445 19128
rect 27479 19125 27491 19159
rect 27433 19119 27491 19125
rect 1104 19066 28888 19088
rect 1104 19014 10982 19066
rect 11034 19014 11046 19066
rect 11098 19014 11110 19066
rect 11162 19014 11174 19066
rect 11226 19014 20982 19066
rect 21034 19014 21046 19066
rect 21098 19014 21110 19066
rect 21162 19014 21174 19066
rect 21226 19014 28888 19066
rect 1104 18992 28888 19014
rect 8478 18952 8484 18964
rect 8439 18924 8484 18952
rect 8478 18912 8484 18924
rect 8536 18912 8542 18964
rect 10778 18952 10784 18964
rect 10739 18924 10784 18952
rect 10778 18912 10784 18924
rect 10836 18912 10842 18964
rect 22097 18955 22155 18961
rect 22097 18921 22109 18955
rect 22143 18952 22155 18955
rect 22462 18952 22468 18964
rect 22143 18924 22468 18952
rect 22143 18921 22155 18924
rect 22097 18915 22155 18921
rect 22462 18912 22468 18924
rect 22520 18952 22526 18964
rect 23017 18955 23075 18961
rect 23017 18952 23029 18955
rect 22520 18924 23029 18952
rect 22520 18912 22526 18924
rect 23017 18921 23029 18924
rect 23063 18921 23075 18955
rect 24118 18952 24124 18964
rect 24079 18924 24124 18952
rect 23017 18915 23075 18921
rect 24118 18912 24124 18924
rect 24176 18912 24182 18964
rect 24489 18955 24547 18961
rect 24489 18921 24501 18955
rect 24535 18952 24547 18955
rect 24578 18952 24584 18964
rect 24535 18924 24584 18952
rect 24535 18921 24547 18924
rect 24489 18915 24547 18921
rect 24578 18912 24584 18924
rect 24636 18912 24642 18964
rect 26513 18955 26571 18961
rect 26513 18921 26525 18955
rect 26559 18952 26571 18955
rect 27154 18952 27160 18964
rect 26559 18924 27160 18952
rect 26559 18921 26571 18924
rect 26513 18915 26571 18921
rect 27154 18912 27160 18924
rect 27212 18912 27218 18964
rect 22830 18884 22836 18896
rect 22791 18856 22836 18884
rect 22830 18844 22836 18856
rect 22888 18844 22894 18896
rect 4246 18776 4252 18828
rect 4304 18816 4310 18828
rect 4433 18819 4491 18825
rect 4433 18816 4445 18819
rect 4304 18788 4445 18816
rect 4304 18776 4310 18788
rect 4433 18785 4445 18788
rect 4479 18785 4491 18819
rect 4433 18779 4491 18785
rect 9766 18776 9772 18828
rect 9824 18816 9830 18828
rect 10045 18819 10103 18825
rect 10045 18816 10057 18819
rect 9824 18788 10057 18816
rect 9824 18776 9830 18788
rect 10045 18785 10057 18788
rect 10091 18785 10103 18819
rect 10045 18779 10103 18785
rect 15194 18776 15200 18828
rect 15252 18816 15258 18828
rect 15545 18819 15603 18825
rect 15545 18816 15557 18819
rect 15252 18788 15557 18816
rect 15252 18776 15258 18788
rect 15545 18785 15557 18788
rect 15591 18785 15603 18819
rect 15545 18779 15603 18785
rect 23290 18776 23296 18828
rect 23348 18816 23354 18828
rect 23385 18819 23443 18825
rect 23385 18816 23397 18819
rect 23348 18788 23397 18816
rect 23348 18776 23354 18788
rect 23385 18785 23397 18788
rect 23431 18785 23443 18819
rect 23385 18779 23443 18785
rect 23474 18776 23480 18828
rect 23532 18816 23538 18828
rect 23532 18788 23577 18816
rect 23532 18776 23538 18788
rect 4522 18748 4528 18760
rect 4483 18720 4528 18748
rect 4522 18708 4528 18720
rect 4580 18708 4586 18760
rect 4709 18751 4767 18757
rect 4709 18717 4721 18751
rect 4755 18748 4767 18751
rect 4798 18748 4804 18760
rect 4755 18720 4804 18748
rect 4755 18717 4767 18720
rect 4709 18711 4767 18717
rect 4798 18708 4804 18720
rect 4856 18708 4862 18760
rect 10134 18748 10140 18760
rect 10095 18720 10140 18748
rect 10134 18708 10140 18720
rect 10192 18708 10198 18760
rect 10321 18751 10379 18757
rect 10321 18717 10333 18751
rect 10367 18748 10379 18751
rect 10870 18748 10876 18760
rect 10367 18720 10876 18748
rect 10367 18717 10379 18720
rect 10321 18711 10379 18717
rect 10870 18708 10876 18720
rect 10928 18708 10934 18760
rect 15286 18748 15292 18760
rect 15247 18720 15292 18748
rect 15286 18708 15292 18720
rect 15344 18708 15350 18760
rect 19429 18751 19487 18757
rect 19429 18717 19441 18751
rect 19475 18748 19487 18751
rect 20438 18748 20444 18760
rect 19475 18720 20444 18748
rect 19475 18717 19487 18720
rect 19429 18711 19487 18717
rect 20438 18708 20444 18720
rect 20496 18708 20502 18760
rect 23566 18748 23572 18760
rect 23527 18720 23572 18748
rect 23566 18708 23572 18720
rect 23624 18708 23630 18760
rect 8205 18683 8263 18689
rect 8205 18649 8217 18683
rect 8251 18680 8263 18683
rect 8386 18680 8392 18692
rect 8251 18652 8392 18680
rect 8251 18649 8263 18652
rect 8205 18643 8263 18649
rect 8386 18640 8392 18652
rect 8444 18680 8450 18692
rect 9677 18683 9735 18689
rect 9677 18680 9689 18683
rect 8444 18652 9689 18680
rect 8444 18640 8450 18652
rect 9677 18649 9689 18652
rect 9723 18649 9735 18683
rect 9677 18643 9735 18649
rect 4065 18615 4123 18621
rect 4065 18581 4077 18615
rect 4111 18612 4123 18615
rect 4154 18612 4160 18624
rect 4111 18584 4160 18612
rect 4111 18581 4123 18584
rect 4065 18575 4123 18581
rect 4154 18572 4160 18584
rect 4212 18572 4218 18624
rect 5074 18612 5080 18624
rect 5035 18584 5080 18612
rect 5074 18572 5080 18584
rect 5132 18572 5138 18624
rect 6914 18612 6920 18624
rect 6827 18584 6920 18612
rect 6914 18572 6920 18584
rect 6972 18612 6978 18624
rect 7190 18612 7196 18624
rect 6972 18584 7196 18612
rect 6972 18572 6978 18584
rect 7190 18572 7196 18584
rect 7248 18572 7254 18624
rect 12618 18572 12624 18624
rect 12676 18612 12682 18624
rect 12805 18615 12863 18621
rect 12805 18612 12817 18615
rect 12676 18584 12817 18612
rect 12676 18572 12682 18584
rect 12805 18581 12817 18584
rect 12851 18581 12863 18615
rect 16666 18612 16672 18624
rect 16627 18584 16672 18612
rect 12805 18575 12863 18581
rect 16666 18572 16672 18584
rect 16724 18572 16730 18624
rect 25593 18615 25651 18621
rect 25593 18581 25605 18615
rect 25639 18612 25651 18615
rect 25682 18612 25688 18624
rect 25639 18584 25688 18612
rect 25639 18581 25651 18584
rect 25593 18575 25651 18581
rect 25682 18572 25688 18584
rect 25740 18572 25746 18624
rect 1104 18522 28888 18544
rect 1104 18470 5982 18522
rect 6034 18470 6046 18522
rect 6098 18470 6110 18522
rect 6162 18470 6174 18522
rect 6226 18470 15982 18522
rect 16034 18470 16046 18522
rect 16098 18470 16110 18522
rect 16162 18470 16174 18522
rect 16226 18470 25982 18522
rect 26034 18470 26046 18522
rect 26098 18470 26110 18522
rect 26162 18470 26174 18522
rect 26226 18470 28888 18522
rect 1104 18448 28888 18470
rect 4522 18368 4528 18420
rect 4580 18408 4586 18420
rect 5350 18408 5356 18420
rect 4580 18380 5356 18408
rect 4580 18368 4586 18380
rect 5350 18368 5356 18380
rect 5408 18368 5414 18420
rect 8113 18411 8171 18417
rect 8113 18377 8125 18411
rect 8159 18408 8171 18411
rect 8846 18408 8852 18420
rect 8159 18380 8852 18408
rect 8159 18377 8171 18380
rect 8113 18371 8171 18377
rect 8846 18368 8852 18380
rect 8904 18368 8910 18420
rect 9217 18411 9275 18417
rect 9217 18377 9229 18411
rect 9263 18408 9275 18411
rect 10781 18411 10839 18417
rect 10781 18408 10793 18411
rect 9263 18380 10793 18408
rect 9263 18377 9275 18380
rect 9217 18371 9275 18377
rect 9677 18343 9735 18349
rect 9677 18340 9689 18343
rect 8588 18312 9689 18340
rect 3970 18232 3976 18284
rect 4028 18272 4034 18284
rect 4798 18272 4804 18284
rect 4028 18244 4804 18272
rect 4028 18232 4034 18244
rect 4798 18232 4804 18244
rect 4856 18272 4862 18284
rect 4985 18275 5043 18281
rect 4985 18272 4997 18275
rect 4856 18244 4997 18272
rect 4856 18232 4862 18244
rect 4985 18241 4997 18244
rect 5031 18272 5043 18275
rect 5721 18275 5779 18281
rect 5721 18272 5733 18275
rect 5031 18244 5733 18272
rect 5031 18241 5043 18244
rect 4985 18235 5043 18241
rect 5721 18241 5733 18244
rect 5767 18241 5779 18275
rect 5721 18235 5779 18241
rect 8202 18232 8208 18284
rect 8260 18272 8266 18284
rect 8588 18281 8616 18312
rect 9677 18309 9689 18312
rect 9723 18309 9735 18343
rect 9677 18303 9735 18309
rect 8573 18275 8631 18281
rect 8573 18272 8585 18275
rect 8260 18244 8585 18272
rect 8260 18232 8266 18244
rect 8573 18241 8585 18244
rect 8619 18241 8631 18275
rect 8573 18235 8631 18241
rect 8757 18275 8815 18281
rect 8757 18241 8769 18275
rect 8803 18272 8815 18275
rect 9582 18272 9588 18284
rect 8803 18244 9588 18272
rect 8803 18241 8815 18244
rect 8757 18235 8815 18241
rect 2133 18207 2191 18213
rect 2133 18173 2145 18207
rect 2179 18204 2191 18207
rect 2222 18204 2228 18216
rect 2179 18176 2228 18204
rect 2179 18173 2191 18176
rect 2133 18167 2191 18173
rect 2222 18164 2228 18176
rect 2280 18164 2286 18216
rect 4062 18164 4068 18216
rect 4120 18204 4126 18216
rect 4709 18207 4767 18213
rect 4709 18204 4721 18207
rect 4120 18176 4721 18204
rect 4120 18164 4126 18176
rect 4709 18173 4721 18176
rect 4755 18204 4767 18207
rect 5074 18204 5080 18216
rect 4755 18176 5080 18204
rect 4755 18173 4767 18176
rect 4709 18167 4767 18173
rect 5074 18164 5080 18176
rect 5132 18164 5138 18216
rect 8386 18164 8392 18216
rect 8444 18204 8450 18216
rect 8481 18207 8539 18213
rect 8481 18204 8493 18207
rect 8444 18176 8493 18204
rect 8444 18164 8450 18176
rect 8481 18173 8493 18176
rect 8527 18173 8539 18207
rect 8481 18167 8539 18173
rect 2041 18139 2099 18145
rect 2041 18105 2053 18139
rect 2087 18136 2099 18139
rect 2378 18139 2436 18145
rect 2378 18136 2390 18139
rect 2087 18108 2390 18136
rect 2087 18105 2099 18108
rect 2041 18099 2099 18105
rect 2378 18105 2390 18108
rect 2424 18136 2436 18139
rect 2774 18136 2780 18148
rect 2424 18108 2780 18136
rect 2424 18105 2436 18108
rect 2378 18099 2436 18105
rect 2774 18096 2780 18108
rect 2832 18096 2838 18148
rect 4157 18139 4215 18145
rect 4157 18105 4169 18139
rect 4203 18136 4215 18139
rect 4246 18136 4252 18148
rect 4203 18108 4252 18136
rect 4203 18105 4215 18108
rect 4157 18099 4215 18105
rect 4246 18096 4252 18108
rect 4304 18096 4310 18148
rect 8018 18136 8024 18148
rect 7931 18108 8024 18136
rect 8018 18096 8024 18108
rect 8076 18136 8082 18148
rect 8772 18136 8800 18235
rect 9582 18232 9588 18244
rect 9640 18232 9646 18284
rect 10244 18281 10272 18380
rect 10781 18377 10793 18380
rect 10827 18408 10839 18411
rect 10870 18408 10876 18420
rect 10827 18380 10876 18408
rect 10827 18377 10839 18380
rect 10781 18371 10839 18377
rect 10870 18368 10876 18380
rect 10928 18368 10934 18420
rect 18874 18408 18880 18420
rect 18835 18380 18880 18408
rect 18874 18368 18880 18380
rect 18932 18408 18938 18420
rect 20438 18408 20444 18420
rect 18932 18380 19932 18408
rect 20399 18380 20444 18408
rect 18932 18368 18938 18380
rect 10229 18275 10287 18281
rect 10229 18241 10241 18275
rect 10275 18241 10287 18275
rect 10229 18235 10287 18241
rect 14553 18275 14611 18281
rect 14553 18241 14565 18275
rect 14599 18272 14611 18275
rect 15838 18272 15844 18284
rect 14599 18244 15844 18272
rect 14599 18241 14611 18244
rect 14553 18235 14611 18241
rect 15838 18232 15844 18244
rect 15896 18232 15902 18284
rect 16025 18275 16083 18281
rect 16025 18241 16037 18275
rect 16071 18272 16083 18275
rect 16666 18272 16672 18284
rect 16071 18244 16672 18272
rect 16071 18241 16083 18244
rect 16025 18235 16083 18241
rect 10137 18207 10195 18213
rect 10137 18173 10149 18207
rect 10183 18204 10195 18207
rect 10318 18204 10324 18216
rect 10183 18176 10324 18204
rect 10183 18173 10195 18176
rect 10137 18167 10195 18173
rect 10318 18164 10324 18176
rect 10376 18204 10382 18216
rect 11057 18207 11115 18213
rect 11057 18204 11069 18207
rect 10376 18176 11069 18204
rect 10376 18164 10382 18176
rect 11057 18173 11069 18176
rect 11103 18173 11115 18207
rect 11057 18167 11115 18173
rect 12618 18164 12624 18216
rect 12676 18204 12682 18216
rect 12805 18207 12863 18213
rect 12805 18204 12817 18207
rect 12676 18176 12817 18204
rect 12676 18164 12682 18176
rect 12805 18173 12817 18176
rect 12851 18173 12863 18207
rect 13072 18207 13130 18213
rect 13072 18204 13084 18207
rect 12805 18167 12863 18173
rect 13004 18176 13084 18204
rect 8076 18108 8800 18136
rect 10045 18139 10103 18145
rect 8076 18096 8082 18108
rect 10045 18105 10057 18139
rect 10091 18136 10103 18139
rect 10226 18136 10232 18148
rect 10091 18108 10232 18136
rect 10091 18105 10103 18108
rect 10045 18099 10103 18105
rect 10226 18096 10232 18108
rect 10284 18136 10290 18148
rect 11425 18139 11483 18145
rect 11425 18136 11437 18139
rect 10284 18108 11437 18136
rect 10284 18096 10290 18108
rect 11425 18105 11437 18108
rect 11471 18105 11483 18139
rect 11425 18099 11483 18105
rect 12713 18139 12771 18145
rect 12713 18105 12725 18139
rect 12759 18136 12771 18139
rect 13004 18136 13032 18176
rect 13072 18173 13084 18176
rect 13118 18204 13130 18207
rect 14458 18204 14464 18216
rect 13118 18176 14464 18204
rect 13118 18173 13130 18176
rect 13072 18167 13130 18173
rect 14458 18164 14464 18176
rect 14516 18204 14522 18216
rect 14921 18207 14979 18213
rect 14921 18204 14933 18207
rect 14516 18176 14933 18204
rect 14516 18164 14522 18176
rect 14921 18173 14933 18176
rect 14967 18204 14979 18207
rect 16040 18204 16068 18235
rect 16666 18232 16672 18244
rect 16724 18232 16730 18284
rect 19904 18281 19932 18380
rect 20438 18368 20444 18380
rect 20496 18368 20502 18420
rect 23109 18411 23167 18417
rect 23109 18377 23121 18411
rect 23155 18408 23167 18411
rect 23566 18408 23572 18420
rect 23155 18380 23572 18408
rect 23155 18377 23167 18380
rect 23109 18371 23167 18377
rect 23566 18368 23572 18380
rect 23624 18368 23630 18420
rect 20714 18300 20720 18352
rect 20772 18340 20778 18352
rect 20993 18343 21051 18349
rect 20993 18340 21005 18343
rect 20772 18312 21005 18340
rect 20772 18300 20778 18312
rect 20993 18309 21005 18312
rect 21039 18309 21051 18343
rect 20993 18303 21051 18309
rect 19889 18275 19947 18281
rect 19889 18241 19901 18275
rect 19935 18241 19947 18275
rect 19889 18235 19947 18241
rect 19978 18232 19984 18284
rect 20036 18272 20042 18284
rect 20806 18272 20812 18284
rect 20036 18244 20812 18272
rect 20036 18232 20042 18244
rect 20806 18232 20812 18244
rect 20864 18272 20870 18284
rect 21545 18275 21603 18281
rect 21545 18272 21557 18275
rect 20864 18244 21557 18272
rect 20864 18232 20870 18244
rect 21545 18241 21557 18244
rect 21591 18241 21603 18275
rect 21545 18235 21603 18241
rect 19334 18204 19340 18216
rect 14967 18176 16068 18204
rect 19295 18176 19340 18204
rect 14967 18173 14979 18176
rect 14921 18167 14979 18173
rect 19334 18164 19340 18176
rect 19392 18204 19398 18216
rect 19797 18207 19855 18213
rect 19797 18204 19809 18207
rect 19392 18176 19809 18204
rect 19392 18164 19398 18176
rect 19797 18173 19809 18176
rect 19843 18173 19855 18207
rect 19797 18167 19855 18173
rect 12759 18108 13032 18136
rect 15749 18139 15807 18145
rect 12759 18105 12771 18108
rect 12713 18099 12771 18105
rect 15749 18105 15761 18139
rect 15795 18136 15807 18139
rect 18598 18136 18604 18148
rect 15795 18108 16252 18136
rect 18511 18108 18604 18136
rect 15795 18105 15807 18108
rect 15749 18099 15807 18105
rect 16224 18080 16252 18108
rect 18598 18096 18604 18108
rect 18656 18136 18662 18148
rect 19996 18136 20024 18232
rect 20438 18164 20444 18216
rect 20496 18204 20502 18216
rect 21361 18207 21419 18213
rect 21361 18204 21373 18207
rect 20496 18176 21373 18204
rect 20496 18164 20502 18176
rect 21361 18173 21373 18176
rect 21407 18173 21419 18207
rect 21361 18167 21419 18173
rect 18656 18108 20024 18136
rect 18656 18096 18662 18108
rect 23290 18096 23296 18148
rect 23348 18136 23354 18148
rect 23845 18139 23903 18145
rect 23845 18136 23857 18139
rect 23348 18108 23857 18136
rect 23348 18096 23354 18108
rect 23845 18105 23857 18108
rect 23891 18105 23903 18139
rect 23845 18099 23903 18105
rect 3510 18068 3516 18080
rect 3471 18040 3516 18068
rect 3510 18028 3516 18040
rect 3568 18028 3574 18080
rect 4341 18071 4399 18077
rect 4341 18037 4353 18071
rect 4387 18068 4399 18071
rect 4430 18068 4436 18080
rect 4387 18040 4436 18068
rect 4387 18037 4399 18040
rect 4341 18031 4399 18037
rect 4430 18028 4436 18040
rect 4488 18028 4494 18080
rect 4801 18071 4859 18077
rect 4801 18037 4813 18071
rect 4847 18068 4859 18071
rect 5166 18068 5172 18080
rect 4847 18040 5172 18068
rect 4847 18037 4859 18040
rect 4801 18031 4859 18037
rect 5166 18028 5172 18040
rect 5224 18028 5230 18080
rect 9585 18071 9643 18077
rect 9585 18037 9597 18071
rect 9631 18068 9643 18071
rect 9674 18068 9680 18080
rect 9631 18040 9680 18068
rect 9631 18037 9643 18040
rect 9585 18031 9643 18037
rect 9674 18028 9680 18040
rect 9732 18028 9738 18080
rect 13814 18028 13820 18080
rect 13872 18068 13878 18080
rect 14185 18071 14243 18077
rect 14185 18068 14197 18071
rect 13872 18040 14197 18068
rect 13872 18028 13878 18040
rect 14185 18037 14197 18040
rect 14231 18037 14243 18071
rect 15194 18068 15200 18080
rect 15155 18040 15200 18068
rect 14185 18031 14243 18037
rect 15194 18028 15200 18040
rect 15252 18028 15258 18080
rect 15378 18068 15384 18080
rect 15339 18040 15384 18068
rect 15378 18028 15384 18040
rect 15436 18028 15442 18080
rect 16206 18028 16212 18080
rect 16264 18068 16270 18080
rect 16393 18071 16451 18077
rect 16393 18068 16405 18071
rect 16264 18040 16405 18068
rect 16264 18028 16270 18040
rect 16393 18037 16405 18040
rect 16439 18037 16451 18071
rect 16942 18068 16948 18080
rect 16903 18040 16948 18068
rect 16393 18031 16451 18037
rect 16942 18028 16948 18040
rect 17000 18028 17006 18080
rect 19429 18071 19487 18077
rect 19429 18037 19441 18071
rect 19475 18068 19487 18071
rect 19702 18068 19708 18080
rect 19475 18040 19708 18068
rect 19475 18037 19487 18040
rect 19429 18031 19487 18037
rect 19702 18028 19708 18040
rect 19760 18028 19766 18080
rect 20901 18071 20959 18077
rect 20901 18037 20913 18071
rect 20947 18068 20959 18071
rect 21358 18068 21364 18080
rect 20947 18040 21364 18068
rect 20947 18037 20959 18040
rect 20901 18031 20959 18037
rect 21358 18028 21364 18040
rect 21416 18068 21422 18080
rect 21453 18071 21511 18077
rect 21453 18068 21465 18071
rect 21416 18040 21465 18068
rect 21416 18028 21422 18040
rect 21453 18037 21465 18040
rect 21499 18037 21511 18071
rect 23474 18068 23480 18080
rect 23387 18040 23480 18068
rect 21453 18031 21511 18037
rect 23474 18028 23480 18040
rect 23532 18068 23538 18080
rect 24762 18068 24768 18080
rect 23532 18040 24768 18068
rect 23532 18028 23538 18040
rect 24762 18028 24768 18040
rect 24820 18028 24826 18080
rect 1104 17978 28888 18000
rect 1104 17926 10982 17978
rect 11034 17926 11046 17978
rect 11098 17926 11110 17978
rect 11162 17926 11174 17978
rect 11226 17926 20982 17978
rect 21034 17926 21046 17978
rect 21098 17926 21110 17978
rect 21162 17926 21174 17978
rect 21226 17926 28888 17978
rect 1104 17904 28888 17926
rect 2961 17867 3019 17873
rect 2961 17833 2973 17867
rect 3007 17864 3019 17867
rect 4062 17864 4068 17876
rect 3007 17836 4068 17864
rect 3007 17833 3019 17836
rect 2961 17827 3019 17833
rect 4062 17824 4068 17836
rect 4120 17824 4126 17876
rect 4154 17824 4160 17876
rect 4212 17864 4218 17876
rect 4525 17867 4583 17873
rect 4525 17864 4537 17867
rect 4212 17836 4537 17864
rect 4212 17824 4218 17836
rect 4525 17833 4537 17836
rect 4571 17864 4583 17867
rect 4614 17864 4620 17876
rect 4571 17836 4620 17864
rect 4571 17833 4583 17836
rect 4525 17827 4583 17833
rect 4614 17824 4620 17836
rect 4672 17824 4678 17876
rect 8202 17864 8208 17876
rect 8163 17836 8208 17864
rect 8202 17824 8208 17836
rect 8260 17824 8266 17876
rect 10226 17864 10232 17876
rect 10187 17836 10232 17864
rect 10226 17824 10232 17836
rect 10284 17824 10290 17876
rect 13262 17864 13268 17876
rect 13223 17836 13268 17864
rect 13262 17824 13268 17836
rect 13320 17824 13326 17876
rect 16206 17864 16212 17876
rect 16167 17836 16212 17864
rect 16206 17824 16212 17836
rect 16264 17824 16270 17876
rect 19702 17864 19708 17876
rect 19663 17836 19708 17864
rect 19702 17824 19708 17836
rect 19760 17824 19766 17876
rect 20806 17824 20812 17876
rect 20864 17864 20870 17876
rect 21085 17867 21143 17873
rect 21085 17864 21097 17867
rect 20864 17836 21097 17864
rect 20864 17824 20870 17836
rect 21085 17833 21097 17836
rect 21131 17833 21143 17867
rect 21085 17827 21143 17833
rect 23017 17867 23075 17873
rect 23017 17833 23029 17867
rect 23063 17864 23075 17867
rect 23290 17864 23296 17876
rect 23063 17836 23296 17864
rect 23063 17833 23075 17836
rect 23017 17827 23075 17833
rect 23290 17824 23296 17836
rect 23348 17824 23354 17876
rect 24854 17864 24860 17876
rect 24815 17836 24860 17864
rect 24854 17824 24860 17836
rect 24912 17824 24918 17876
rect 2774 17756 2780 17808
rect 2832 17796 2838 17808
rect 3881 17799 3939 17805
rect 3881 17796 3893 17799
rect 2832 17768 3893 17796
rect 2832 17756 2838 17768
rect 3881 17765 3893 17768
rect 3927 17796 3939 17799
rect 3970 17796 3976 17808
rect 3927 17768 3976 17796
rect 3927 17765 3939 17768
rect 3881 17759 3939 17765
rect 3970 17756 3976 17768
rect 4028 17756 4034 17808
rect 16666 17796 16672 17808
rect 16627 17768 16672 17796
rect 16666 17756 16672 17768
rect 16724 17756 16730 17808
rect 24670 17756 24676 17808
rect 24728 17796 24734 17808
rect 25317 17799 25375 17805
rect 25317 17796 25329 17799
rect 24728 17768 25329 17796
rect 24728 17756 24734 17768
rect 25317 17765 25329 17768
rect 25363 17765 25375 17799
rect 25317 17759 25375 17765
rect 1394 17728 1400 17740
rect 1355 17700 1400 17728
rect 1394 17688 1400 17700
rect 1452 17688 1458 17740
rect 4430 17728 4436 17740
rect 4391 17700 4436 17728
rect 4430 17688 4436 17700
rect 4488 17688 4494 17740
rect 6362 17737 6368 17740
rect 6356 17728 6368 17737
rect 4724 17700 6368 17728
rect 3510 17620 3516 17672
rect 3568 17660 3574 17672
rect 4338 17660 4344 17672
rect 3568 17632 4344 17660
rect 3568 17620 3574 17632
rect 4338 17620 4344 17632
rect 4396 17660 4402 17672
rect 4724 17669 4752 17700
rect 6356 17691 6368 17700
rect 6420 17728 6426 17740
rect 9493 17731 9551 17737
rect 6420 17700 6456 17728
rect 6362 17688 6368 17691
rect 6420 17688 6426 17700
rect 9493 17697 9505 17731
rect 9539 17728 9551 17731
rect 10134 17728 10140 17740
rect 9539 17700 10140 17728
rect 9539 17697 9551 17700
rect 9493 17691 9551 17697
rect 10134 17688 10140 17700
rect 10192 17688 10198 17740
rect 10594 17728 10600 17740
rect 10555 17700 10600 17728
rect 10594 17688 10600 17700
rect 10652 17688 10658 17740
rect 10689 17731 10747 17737
rect 10689 17697 10701 17731
rect 10735 17728 10747 17731
rect 10778 17728 10784 17740
rect 10735 17700 10784 17728
rect 10735 17697 10747 17700
rect 10689 17691 10747 17697
rect 10778 17688 10784 17700
rect 10836 17688 10842 17740
rect 16577 17731 16635 17737
rect 16577 17697 16589 17731
rect 16623 17728 16635 17731
rect 16942 17728 16948 17740
rect 16623 17700 16948 17728
rect 16623 17697 16635 17700
rect 16577 17691 16635 17697
rect 16942 17688 16948 17700
rect 17000 17688 17006 17740
rect 19613 17731 19671 17737
rect 19613 17697 19625 17731
rect 19659 17728 19671 17731
rect 20622 17728 20628 17740
rect 19659 17700 20628 17728
rect 19659 17697 19671 17700
rect 19613 17691 19671 17697
rect 20622 17688 20628 17700
rect 20680 17688 20686 17740
rect 23198 17688 23204 17740
rect 23256 17728 23262 17740
rect 23385 17731 23443 17737
rect 23385 17728 23397 17731
rect 23256 17700 23397 17728
rect 23256 17688 23262 17700
rect 23385 17697 23397 17700
rect 23431 17697 23443 17731
rect 23385 17691 23443 17697
rect 24765 17731 24823 17737
rect 24765 17697 24777 17731
rect 24811 17728 24823 17731
rect 24854 17728 24860 17740
rect 24811 17700 24860 17728
rect 24811 17697 24823 17700
rect 24765 17691 24823 17697
rect 24854 17688 24860 17700
rect 24912 17728 24918 17740
rect 25225 17731 25283 17737
rect 25225 17728 25237 17731
rect 24912 17700 25237 17728
rect 24912 17688 24918 17700
rect 25225 17697 25237 17700
rect 25271 17697 25283 17731
rect 25225 17691 25283 17697
rect 4709 17663 4767 17669
rect 4709 17660 4721 17663
rect 4396 17632 4721 17660
rect 4396 17620 4402 17632
rect 4709 17629 4721 17632
rect 4755 17629 4767 17663
rect 5166 17660 5172 17672
rect 5127 17632 5172 17660
rect 4709 17623 4767 17629
rect 5166 17620 5172 17632
rect 5224 17620 5230 17672
rect 5718 17620 5724 17672
rect 5776 17660 5782 17672
rect 6089 17663 6147 17669
rect 6089 17660 6101 17663
rect 5776 17632 6101 17660
rect 5776 17620 5782 17632
rect 6089 17629 6101 17632
rect 6135 17629 6147 17663
rect 10870 17660 10876 17672
rect 10831 17632 10876 17660
rect 6089 17623 6147 17629
rect 10870 17620 10876 17632
rect 10928 17620 10934 17672
rect 13354 17660 13360 17672
rect 13315 17632 13360 17660
rect 13354 17620 13360 17632
rect 13412 17620 13418 17672
rect 13541 17663 13599 17669
rect 13541 17629 13553 17663
rect 13587 17660 13599 17663
rect 13722 17660 13728 17672
rect 13587 17632 13728 17660
rect 13587 17629 13599 17632
rect 13541 17623 13599 17629
rect 13722 17620 13728 17632
rect 13780 17620 13786 17672
rect 16758 17620 16764 17672
rect 16816 17660 16822 17672
rect 16816 17632 16861 17660
rect 16816 17620 16822 17632
rect 19794 17620 19800 17672
rect 19852 17660 19858 17672
rect 19889 17663 19947 17669
rect 19889 17660 19901 17663
rect 19852 17632 19901 17660
rect 19852 17620 19858 17632
rect 19889 17629 19901 17632
rect 19935 17660 19947 17663
rect 21266 17660 21272 17672
rect 19935 17632 21272 17660
rect 19935 17629 19947 17632
rect 19889 17623 19947 17629
rect 21266 17620 21272 17632
rect 21324 17620 21330 17672
rect 22925 17663 22983 17669
rect 22925 17629 22937 17663
rect 22971 17660 22983 17663
rect 23474 17660 23480 17672
rect 22971 17632 23480 17660
rect 22971 17629 22983 17632
rect 22925 17623 22983 17629
rect 23474 17620 23480 17632
rect 23532 17620 23538 17672
rect 23569 17663 23627 17669
rect 23569 17629 23581 17663
rect 23615 17629 23627 17663
rect 25406 17660 25412 17672
rect 25367 17632 25412 17660
rect 23569 17623 23627 17629
rect 15657 17595 15715 17601
rect 15657 17561 15669 17595
rect 15703 17592 15715 17595
rect 16390 17592 16396 17604
rect 15703 17564 16396 17592
rect 15703 17561 15715 17564
rect 15657 17555 15715 17561
rect 16390 17552 16396 17564
rect 16448 17552 16454 17604
rect 23106 17552 23112 17604
rect 23164 17592 23170 17604
rect 23584 17592 23612 17623
rect 25406 17620 25412 17632
rect 25464 17620 25470 17672
rect 23164 17564 23612 17592
rect 23164 17552 23170 17564
rect 1394 17484 1400 17536
rect 1452 17524 1458 17536
rect 1581 17527 1639 17533
rect 1581 17524 1593 17527
rect 1452 17496 1593 17524
rect 1452 17484 1458 17496
rect 1581 17493 1593 17496
rect 1627 17493 1639 17527
rect 1581 17487 1639 17493
rect 2225 17527 2283 17533
rect 2225 17493 2237 17527
rect 2271 17524 2283 17527
rect 2314 17524 2320 17536
rect 2271 17496 2320 17524
rect 2271 17493 2283 17496
rect 2225 17487 2283 17493
rect 2314 17484 2320 17496
rect 2372 17484 2378 17536
rect 4062 17524 4068 17536
rect 4023 17496 4068 17524
rect 4062 17484 4068 17496
rect 4120 17484 4126 17536
rect 7466 17524 7472 17536
rect 7427 17496 7472 17524
rect 7466 17484 7472 17496
rect 7524 17484 7530 17536
rect 10137 17527 10195 17533
rect 10137 17493 10149 17527
rect 10183 17524 10195 17527
rect 10410 17524 10416 17536
rect 10183 17496 10416 17524
rect 10183 17493 10195 17496
rect 10137 17487 10195 17493
rect 10410 17484 10416 17496
rect 10468 17484 10474 17536
rect 12710 17484 12716 17536
rect 12768 17524 12774 17536
rect 12897 17527 12955 17533
rect 12897 17524 12909 17527
rect 12768 17496 12909 17524
rect 12768 17484 12774 17496
rect 12897 17493 12909 17496
rect 12943 17493 12955 17527
rect 12897 17487 12955 17493
rect 13814 17484 13820 17536
rect 13872 17524 13878 17536
rect 13909 17527 13967 17533
rect 13909 17524 13921 17527
rect 13872 17496 13921 17524
rect 13872 17484 13878 17496
rect 13909 17493 13921 17496
rect 13955 17493 13967 17527
rect 13909 17487 13967 17493
rect 15286 17484 15292 17536
rect 15344 17524 15350 17536
rect 16025 17527 16083 17533
rect 16025 17524 16037 17527
rect 15344 17496 16037 17524
rect 15344 17484 15350 17496
rect 16025 17493 16037 17496
rect 16071 17524 16083 17527
rect 16298 17524 16304 17536
rect 16071 17496 16304 17524
rect 16071 17493 16083 17496
rect 16025 17487 16083 17493
rect 16298 17484 16304 17496
rect 16356 17484 16362 17536
rect 19153 17527 19211 17533
rect 19153 17493 19165 17527
rect 19199 17524 19211 17527
rect 19245 17527 19303 17533
rect 19245 17524 19257 17527
rect 19199 17496 19257 17524
rect 19199 17493 19211 17496
rect 19153 17487 19211 17493
rect 19245 17493 19257 17496
rect 19291 17524 19303 17527
rect 19518 17524 19524 17536
rect 19291 17496 19524 17524
rect 19291 17493 19303 17496
rect 19245 17487 19303 17493
rect 19518 17484 19524 17496
rect 19576 17484 19582 17536
rect 25774 17484 25780 17536
rect 25832 17524 25838 17536
rect 25869 17527 25927 17533
rect 25869 17524 25881 17527
rect 25832 17496 25881 17524
rect 25832 17484 25838 17496
rect 25869 17493 25881 17496
rect 25915 17493 25927 17527
rect 25869 17487 25927 17493
rect 1104 17434 28888 17456
rect 1104 17382 5982 17434
rect 6034 17382 6046 17434
rect 6098 17382 6110 17434
rect 6162 17382 6174 17434
rect 6226 17382 15982 17434
rect 16034 17382 16046 17434
rect 16098 17382 16110 17434
rect 16162 17382 16174 17434
rect 16226 17382 25982 17434
rect 26034 17382 26046 17434
rect 26098 17382 26110 17434
rect 26162 17382 26174 17434
rect 26226 17382 28888 17434
rect 1104 17360 28888 17382
rect 2038 17320 2044 17332
rect 1999 17292 2044 17320
rect 2038 17280 2044 17292
rect 2096 17280 2102 17332
rect 4338 17320 4344 17332
rect 4299 17292 4344 17320
rect 4338 17280 4344 17292
rect 4396 17280 4402 17332
rect 4430 17280 4436 17332
rect 4488 17320 4494 17332
rect 4985 17323 5043 17329
rect 4985 17320 4997 17323
rect 4488 17292 4997 17320
rect 4488 17280 4494 17292
rect 4985 17289 4997 17292
rect 5031 17289 5043 17323
rect 4985 17283 5043 17289
rect 6181 17323 6239 17329
rect 6181 17289 6193 17323
rect 6227 17320 6239 17323
rect 6362 17320 6368 17332
rect 6227 17292 6368 17320
rect 6227 17289 6239 17292
rect 6181 17283 6239 17289
rect 6362 17280 6368 17292
rect 6420 17280 6426 17332
rect 10045 17323 10103 17329
rect 10045 17289 10057 17323
rect 10091 17320 10103 17323
rect 10134 17320 10140 17332
rect 10091 17292 10140 17320
rect 10091 17289 10103 17292
rect 10045 17283 10103 17289
rect 10134 17280 10140 17292
rect 10192 17280 10198 17332
rect 13354 17320 13360 17332
rect 13315 17292 13360 17320
rect 13354 17280 13360 17292
rect 13412 17280 13418 17332
rect 14458 17320 14464 17332
rect 14419 17292 14464 17320
rect 14458 17280 14464 17292
rect 14516 17280 14522 17332
rect 16666 17320 16672 17332
rect 16627 17292 16672 17320
rect 16666 17280 16672 17292
rect 16724 17280 16730 17332
rect 16942 17320 16948 17332
rect 16903 17292 16948 17320
rect 16942 17280 16948 17292
rect 17000 17280 17006 17332
rect 19702 17280 19708 17332
rect 19760 17320 19766 17332
rect 20165 17323 20223 17329
rect 20165 17320 20177 17323
rect 19760 17292 20177 17320
rect 19760 17280 19766 17292
rect 20165 17289 20177 17292
rect 20211 17289 20223 17323
rect 22738 17320 22744 17332
rect 20165 17283 20223 17289
rect 20272 17292 22744 17320
rect 1581 17255 1639 17261
rect 1581 17221 1593 17255
rect 1627 17252 1639 17255
rect 3786 17252 3792 17264
rect 1627 17224 3792 17252
rect 1627 17221 1639 17224
rect 1581 17215 1639 17221
rect 3786 17212 3792 17224
rect 3844 17212 3850 17264
rect 3145 17187 3203 17193
rect 3145 17153 3157 17187
rect 3191 17184 3203 17187
rect 3881 17187 3939 17193
rect 3881 17184 3893 17187
rect 3191 17156 3893 17184
rect 3191 17153 3203 17156
rect 3145 17147 3203 17153
rect 3881 17153 3893 17156
rect 3927 17184 3939 17187
rect 4356 17184 4384 17280
rect 4614 17252 4620 17264
rect 4575 17224 4620 17252
rect 4614 17212 4620 17224
rect 4672 17212 4678 17264
rect 9582 17252 9588 17264
rect 9495 17224 9588 17252
rect 9582 17212 9588 17224
rect 9640 17252 9646 17264
rect 10594 17252 10600 17264
rect 9640 17224 10600 17252
rect 9640 17212 9646 17224
rect 10594 17212 10600 17224
rect 10652 17212 10658 17264
rect 10870 17252 10876 17264
rect 10704 17224 10876 17252
rect 10704 17193 10732 17224
rect 10870 17212 10876 17224
rect 10928 17252 10934 17264
rect 11517 17255 11575 17261
rect 11517 17252 11529 17255
rect 10928 17224 11529 17252
rect 10928 17212 10934 17224
rect 11517 17221 11529 17224
rect 11563 17252 11575 17255
rect 12342 17252 12348 17264
rect 11563 17224 12348 17252
rect 11563 17221 11575 17224
rect 11517 17215 11575 17221
rect 12342 17212 12348 17224
rect 12400 17212 12406 17264
rect 12989 17255 13047 17261
rect 12989 17221 13001 17255
rect 13035 17252 13047 17255
rect 13722 17252 13728 17264
rect 13035 17224 13728 17252
rect 13035 17221 13047 17224
rect 12989 17215 13047 17221
rect 13722 17212 13728 17224
rect 13780 17212 13786 17264
rect 3927 17156 4384 17184
rect 9217 17187 9275 17193
rect 3927 17153 3939 17156
rect 3881 17147 3939 17153
rect 9217 17153 9229 17187
rect 9263 17184 9275 17187
rect 10689 17187 10747 17193
rect 10689 17184 10701 17187
rect 9263 17156 10701 17184
rect 9263 17153 9275 17156
rect 9217 17147 9275 17153
rect 10689 17153 10701 17156
rect 10735 17153 10747 17187
rect 10689 17147 10747 17153
rect 12253 17187 12311 17193
rect 12253 17153 12265 17187
rect 12299 17184 12311 17187
rect 13262 17184 13268 17196
rect 12299 17156 13268 17184
rect 12299 17153 12311 17156
rect 12253 17147 12311 17153
rect 13262 17144 13268 17156
rect 13320 17144 13326 17196
rect 14001 17187 14059 17193
rect 14001 17153 14013 17187
rect 14047 17184 14059 17187
rect 14476 17184 14504 17280
rect 16758 17212 16764 17264
rect 16816 17252 16822 17264
rect 17313 17255 17371 17261
rect 17313 17252 17325 17255
rect 16816 17224 17325 17252
rect 16816 17212 16822 17224
rect 17313 17221 17325 17224
rect 17359 17252 17371 17255
rect 17494 17252 17500 17264
rect 17359 17224 17500 17252
rect 17359 17221 17371 17224
rect 17313 17215 17371 17221
rect 17494 17212 17500 17224
rect 17552 17212 17558 17264
rect 18230 17212 18236 17264
rect 18288 17252 18294 17264
rect 19153 17255 19211 17261
rect 19153 17252 19165 17255
rect 18288 17224 19165 17252
rect 18288 17212 18294 17224
rect 19153 17221 19165 17224
rect 19199 17221 19211 17255
rect 19153 17215 19211 17221
rect 14047 17156 14504 17184
rect 16209 17187 16267 17193
rect 14047 17153 14059 17156
rect 14001 17147 14059 17153
rect 16209 17153 16221 17187
rect 16255 17184 16267 17187
rect 16390 17184 16396 17196
rect 16255 17156 16396 17184
rect 16255 17153 16267 17156
rect 16209 17147 16267 17153
rect 16390 17144 16396 17156
rect 16448 17144 16454 17196
rect 19061 17187 19119 17193
rect 19061 17153 19073 17187
rect 19107 17184 19119 17187
rect 19797 17187 19855 17193
rect 19797 17184 19809 17187
rect 19107 17156 19809 17184
rect 19107 17153 19119 17156
rect 19061 17147 19119 17153
rect 19797 17153 19809 17156
rect 19843 17184 19855 17187
rect 20272 17184 20300 17292
rect 22738 17280 22744 17292
rect 22796 17280 22802 17332
rect 23474 17280 23480 17332
rect 23532 17320 23538 17332
rect 23661 17323 23719 17329
rect 23661 17320 23673 17323
rect 23532 17292 23673 17320
rect 23532 17280 23538 17292
rect 23661 17289 23673 17292
rect 23707 17289 23719 17323
rect 23661 17283 23719 17289
rect 25406 17280 25412 17332
rect 25464 17320 25470 17332
rect 27065 17323 27123 17329
rect 27065 17320 27077 17323
rect 25464 17292 27077 17320
rect 25464 17280 25470 17292
rect 27065 17289 27077 17292
rect 27111 17289 27123 17323
rect 27065 17283 27123 17289
rect 20622 17252 20628 17264
rect 20583 17224 20628 17252
rect 20622 17212 20628 17224
rect 20680 17212 20686 17264
rect 21266 17252 21272 17264
rect 21227 17224 21272 17252
rect 21266 17212 21272 17224
rect 21324 17212 21330 17264
rect 23106 17212 23112 17264
rect 23164 17252 23170 17264
rect 24857 17255 24915 17261
rect 24857 17252 24869 17255
rect 23164 17224 24869 17252
rect 23164 17212 23170 17224
rect 24857 17221 24869 17224
rect 24903 17252 24915 17255
rect 25424 17252 25452 17280
rect 24903 17224 25452 17252
rect 24903 17221 24915 17224
rect 24857 17215 24915 17221
rect 19843 17156 20300 17184
rect 21284 17184 21312 17212
rect 24210 17184 24216 17196
rect 21284 17156 21496 17184
rect 24171 17156 24216 17184
rect 19843 17153 19855 17156
rect 19797 17147 19855 17153
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17116 1455 17119
rect 2038 17116 2044 17128
rect 1443 17088 2044 17116
rect 1443 17085 1455 17088
rect 1397 17079 1455 17085
rect 2038 17076 2044 17088
rect 2096 17076 2102 17128
rect 7190 17116 7196 17128
rect 6472 17088 7196 17116
rect 2777 17051 2835 17057
rect 2777 17017 2789 17051
rect 2823 17048 2835 17051
rect 3605 17051 3663 17057
rect 3605 17048 3617 17051
rect 2823 17020 3617 17048
rect 2823 17017 2835 17020
rect 2777 17011 2835 17017
rect 3605 17017 3617 17020
rect 3651 17048 3663 17051
rect 4062 17048 4068 17060
rect 3651 17020 4068 17048
rect 3651 17017 3663 17020
rect 3605 17011 3663 17017
rect 4062 17008 4068 17020
rect 4120 17008 4126 17060
rect 3234 16980 3240 16992
rect 3195 16952 3240 16980
rect 3234 16940 3240 16952
rect 3292 16940 3298 16992
rect 3694 16980 3700 16992
rect 3655 16952 3700 16980
rect 3694 16940 3700 16952
rect 3752 16940 3758 16992
rect 5718 16940 5724 16992
rect 5776 16980 5782 16992
rect 6472 16989 6500 17088
rect 7190 17076 7196 17088
rect 7248 17076 7254 17128
rect 19518 17116 19524 17128
rect 19479 17088 19524 17116
rect 19518 17076 19524 17088
rect 19576 17076 19582 17128
rect 21358 17116 21364 17128
rect 21319 17088 21364 17116
rect 21358 17076 21364 17088
rect 21416 17076 21422 17128
rect 21468 17116 21496 17156
rect 24210 17144 24216 17156
rect 24268 17184 24274 17196
rect 25406 17184 25412 17196
rect 24268 17156 25412 17184
rect 24268 17144 24274 17156
rect 25406 17144 25412 17156
rect 25464 17184 25470 17196
rect 25501 17187 25559 17193
rect 25501 17184 25513 17187
rect 25464 17156 25513 17184
rect 25464 17144 25470 17156
rect 25501 17153 25513 17156
rect 25547 17184 25559 17187
rect 25547 17156 25820 17184
rect 25547 17153 25559 17156
rect 25501 17147 25559 17153
rect 21617 17119 21675 17125
rect 21617 17116 21629 17119
rect 21468 17088 21629 17116
rect 21617 17085 21629 17088
rect 21663 17085 21675 17119
rect 21617 17079 21675 17085
rect 24762 17076 24768 17128
rect 24820 17116 24826 17128
rect 25685 17119 25743 17125
rect 25685 17116 25697 17119
rect 24820 17088 25697 17116
rect 24820 17076 24826 17088
rect 25685 17085 25697 17088
rect 25731 17085 25743 17119
rect 25792 17116 25820 17156
rect 25941 17119 25999 17125
rect 25941 17116 25953 17119
rect 25792 17088 25953 17116
rect 25685 17079 25743 17085
rect 25941 17085 25953 17088
rect 25987 17085 25999 17119
rect 25941 17079 25999 17085
rect 7466 17057 7472 17060
rect 7438 17051 7472 17057
rect 7438 17048 7450 17051
rect 7024 17020 7450 17048
rect 7024 16992 7052 17020
rect 7438 17017 7450 17020
rect 7524 17048 7530 17060
rect 10505 17051 10563 17057
rect 10505 17048 10517 17051
rect 7524 17020 7586 17048
rect 9876 17020 10517 17048
rect 7438 17011 7472 17017
rect 7466 17008 7472 17011
rect 7524 17008 7530 17020
rect 9876 16992 9904 17020
rect 10505 17017 10517 17020
rect 10551 17048 10563 17051
rect 11606 17048 11612 17060
rect 10551 17020 11612 17048
rect 10551 17017 10563 17020
rect 10505 17011 10563 17017
rect 11606 17008 11612 17020
rect 11664 17008 11670 17060
rect 13446 17008 13452 17060
rect 13504 17048 13510 17060
rect 13725 17051 13783 17057
rect 13725 17048 13737 17051
rect 13504 17020 13737 17048
rect 13504 17008 13510 17020
rect 13725 17017 13737 17020
rect 13771 17048 13783 17051
rect 14737 17051 14795 17057
rect 14737 17048 14749 17051
rect 13771 17020 14749 17048
rect 13771 17017 13783 17020
rect 13725 17011 13783 17017
rect 14737 17017 14749 17020
rect 14783 17017 14795 17051
rect 16025 17051 16083 17057
rect 16025 17048 16037 17051
rect 14737 17011 14795 17017
rect 15396 17020 16037 17048
rect 15396 16992 15424 17020
rect 16025 17017 16037 17020
rect 16071 17017 16083 17051
rect 16025 17011 16083 17017
rect 18693 17051 18751 17057
rect 18693 17017 18705 17051
rect 18739 17048 18751 17051
rect 19794 17048 19800 17060
rect 18739 17020 19800 17048
rect 18739 17017 18751 17020
rect 18693 17011 18751 17017
rect 19794 17008 19800 17020
rect 19852 17008 19858 17060
rect 23474 17048 23480 17060
rect 23435 17020 23480 17048
rect 23474 17008 23480 17020
rect 23532 17048 23538 17060
rect 24121 17051 24179 17057
rect 24121 17048 24133 17051
rect 23532 17020 24133 17048
rect 23532 17008 23538 17020
rect 24121 17017 24133 17020
rect 24167 17017 24179 17051
rect 25700 17048 25728 17079
rect 25774 17048 25780 17060
rect 25700 17020 25780 17048
rect 24121 17011 24179 17017
rect 25774 17008 25780 17020
rect 25832 17008 25838 17060
rect 6457 16983 6515 16989
rect 6457 16980 6469 16983
rect 5776 16952 6469 16980
rect 5776 16940 5782 16952
rect 6457 16949 6469 16952
rect 6503 16949 6515 16983
rect 7006 16980 7012 16992
rect 6967 16952 7012 16980
rect 6457 16943 6515 16949
rect 7006 16940 7012 16952
rect 7064 16940 7070 16992
rect 8570 16980 8576 16992
rect 8531 16952 8576 16980
rect 8570 16940 8576 16952
rect 8628 16940 8634 16992
rect 9858 16980 9864 16992
rect 9819 16952 9864 16980
rect 9858 16940 9864 16952
rect 9916 16940 9922 16992
rect 10410 16980 10416 16992
rect 10371 16952 10416 16980
rect 10410 16940 10416 16952
rect 10468 16940 10474 16992
rect 10778 16940 10784 16992
rect 10836 16980 10842 16992
rect 11057 16983 11115 16989
rect 11057 16980 11069 16983
rect 10836 16952 11069 16980
rect 10836 16940 10842 16952
rect 11057 16949 11069 16952
rect 11103 16949 11115 16983
rect 13814 16980 13820 16992
rect 13775 16952 13820 16980
rect 11057 16943 11115 16949
rect 13814 16940 13820 16952
rect 13872 16940 13878 16992
rect 15378 16980 15384 16992
rect 15339 16952 15384 16980
rect 15378 16940 15384 16952
rect 15436 16940 15442 16992
rect 15470 16940 15476 16992
rect 15528 16980 15534 16992
rect 15565 16983 15623 16989
rect 15565 16980 15577 16983
rect 15528 16952 15577 16980
rect 15528 16940 15534 16952
rect 15565 16949 15577 16952
rect 15611 16949 15623 16983
rect 15565 16943 15623 16949
rect 15838 16940 15844 16992
rect 15896 16980 15902 16992
rect 15933 16983 15991 16989
rect 15933 16980 15945 16983
rect 15896 16952 15945 16980
rect 15896 16940 15902 16952
rect 15933 16949 15945 16952
rect 15979 16949 15991 16983
rect 18322 16980 18328 16992
rect 18283 16952 18328 16980
rect 15933 16943 15991 16949
rect 18322 16940 18328 16952
rect 18380 16940 18386 16992
rect 19610 16980 19616 16992
rect 19571 16952 19616 16980
rect 19610 16940 19616 16952
rect 19668 16940 19674 16992
rect 23109 16983 23167 16989
rect 23109 16949 23121 16983
rect 23155 16980 23167 16983
rect 23198 16980 23204 16992
rect 23155 16952 23204 16980
rect 23155 16949 23167 16952
rect 23109 16943 23167 16949
rect 23198 16940 23204 16952
rect 23256 16940 23262 16992
rect 23658 16940 23664 16992
rect 23716 16980 23722 16992
rect 24029 16983 24087 16989
rect 24029 16980 24041 16983
rect 23716 16952 24041 16980
rect 23716 16940 23722 16952
rect 24029 16949 24041 16952
rect 24075 16949 24087 16983
rect 24029 16943 24087 16949
rect 1104 16890 28888 16912
rect 1104 16838 10982 16890
rect 11034 16838 11046 16890
rect 11098 16838 11110 16890
rect 11162 16838 11174 16890
rect 11226 16838 20982 16890
rect 21034 16838 21046 16890
rect 21098 16838 21110 16890
rect 21162 16838 21174 16890
rect 21226 16838 28888 16890
rect 1104 16816 28888 16838
rect 1486 16736 1492 16788
rect 1544 16776 1550 16788
rect 1581 16779 1639 16785
rect 1581 16776 1593 16779
rect 1544 16748 1593 16776
rect 1544 16736 1550 16748
rect 1581 16745 1593 16748
rect 1627 16745 1639 16779
rect 1581 16739 1639 16745
rect 3329 16779 3387 16785
rect 3329 16745 3341 16779
rect 3375 16776 3387 16779
rect 3694 16776 3700 16788
rect 3375 16748 3700 16776
rect 3375 16745 3387 16748
rect 3329 16739 3387 16745
rect 3694 16736 3700 16748
rect 3752 16736 3758 16788
rect 4062 16776 4068 16788
rect 4023 16748 4068 16776
rect 4062 16736 4068 16748
rect 4120 16736 4126 16788
rect 4433 16779 4491 16785
rect 4433 16745 4445 16779
rect 4479 16776 4491 16779
rect 4706 16776 4712 16788
rect 4479 16748 4712 16776
rect 4479 16745 4491 16748
rect 4433 16739 4491 16745
rect 4706 16736 4712 16748
rect 4764 16736 4770 16788
rect 6822 16776 6828 16788
rect 6783 16748 6828 16776
rect 6822 16736 6828 16748
rect 6880 16736 6886 16788
rect 7190 16736 7196 16788
rect 7248 16776 7254 16788
rect 7377 16779 7435 16785
rect 7377 16776 7389 16779
rect 7248 16748 7389 16776
rect 7248 16736 7254 16748
rect 7377 16745 7389 16748
rect 7423 16745 7435 16779
rect 7377 16739 7435 16745
rect 10137 16779 10195 16785
rect 10137 16745 10149 16779
rect 10183 16776 10195 16779
rect 10318 16776 10324 16788
rect 10183 16748 10324 16776
rect 10183 16745 10195 16748
rect 10137 16739 10195 16745
rect 10318 16736 10324 16748
rect 10376 16736 10382 16788
rect 13446 16776 13452 16788
rect 13407 16748 13452 16776
rect 13446 16736 13452 16748
rect 13504 16736 13510 16788
rect 17494 16776 17500 16788
rect 17455 16748 17500 16776
rect 17494 16736 17500 16748
rect 17552 16736 17558 16788
rect 18322 16736 18328 16788
rect 18380 16776 18386 16788
rect 19153 16779 19211 16785
rect 19153 16776 19165 16779
rect 18380 16748 19165 16776
rect 18380 16736 18386 16748
rect 19153 16745 19165 16748
rect 19199 16776 19211 16779
rect 19610 16776 19616 16788
rect 19199 16748 19616 16776
rect 19199 16745 19211 16748
rect 19153 16739 19211 16745
rect 19610 16736 19616 16748
rect 19668 16736 19674 16788
rect 21358 16776 21364 16788
rect 21319 16748 21364 16776
rect 21358 16736 21364 16748
rect 21416 16736 21422 16788
rect 23106 16776 23112 16788
rect 23067 16748 23112 16776
rect 23106 16736 23112 16748
rect 23164 16736 23170 16788
rect 24121 16779 24179 16785
rect 24121 16745 24133 16779
rect 24167 16776 24179 16779
rect 24210 16776 24216 16788
rect 24167 16748 24216 16776
rect 24167 16745 24179 16748
rect 24121 16739 24179 16745
rect 24210 16736 24216 16748
rect 24268 16736 24274 16788
rect 24854 16776 24860 16788
rect 24815 16748 24860 16776
rect 24854 16736 24860 16748
rect 24912 16736 24918 16788
rect 25774 16736 25780 16788
rect 25832 16776 25838 16788
rect 26697 16779 26755 16785
rect 26697 16776 26709 16779
rect 25832 16748 26709 16776
rect 25832 16736 25838 16748
rect 26697 16745 26709 16748
rect 26743 16745 26755 16779
rect 26697 16739 26755 16745
rect 5810 16668 5816 16720
rect 5868 16708 5874 16720
rect 6733 16711 6791 16717
rect 6733 16708 6745 16711
rect 5868 16680 6745 16708
rect 5868 16668 5874 16680
rect 6733 16677 6745 16680
rect 6779 16677 6791 16711
rect 6733 16671 6791 16677
rect 12989 16711 13047 16717
rect 12989 16677 13001 16711
rect 13035 16708 13047 16711
rect 13354 16708 13360 16720
rect 13035 16680 13360 16708
rect 13035 16677 13047 16680
rect 12989 16671 13047 16677
rect 13354 16668 13360 16680
rect 13412 16668 13418 16720
rect 13630 16668 13636 16720
rect 13688 16708 13694 16720
rect 13817 16711 13875 16717
rect 13817 16708 13829 16711
rect 13688 16680 13829 16708
rect 13688 16668 13694 16680
rect 13817 16677 13829 16680
rect 13863 16708 13875 16711
rect 13906 16708 13912 16720
rect 13863 16680 13912 16708
rect 13863 16677 13875 16680
rect 13817 16671 13875 16677
rect 13906 16668 13912 16680
rect 13964 16708 13970 16720
rect 14458 16708 14464 16720
rect 13964 16680 14464 16708
rect 13964 16668 13970 16680
rect 14458 16668 14464 16680
rect 14516 16668 14522 16720
rect 19061 16711 19119 16717
rect 19061 16677 19073 16711
rect 19107 16708 19119 16711
rect 25317 16711 25375 16717
rect 19107 16680 19656 16708
rect 19107 16677 19119 16680
rect 19061 16671 19119 16677
rect 4525 16643 4583 16649
rect 4525 16609 4537 16643
rect 4571 16640 4583 16643
rect 5074 16640 5080 16652
rect 4571 16612 5080 16640
rect 4571 16609 4583 16612
rect 4525 16603 4583 16609
rect 5074 16600 5080 16612
rect 5132 16600 5138 16652
rect 7006 16640 7012 16652
rect 6932 16612 7012 16640
rect 6932 16581 6960 16612
rect 7006 16600 7012 16612
rect 7064 16600 7070 16652
rect 10502 16640 10508 16652
rect 10415 16612 10508 16640
rect 10502 16600 10508 16612
rect 10560 16640 10566 16652
rect 15838 16640 15844 16652
rect 10560 16612 15844 16640
rect 10560 16600 10566 16612
rect 15838 16600 15844 16612
rect 15896 16600 15902 16652
rect 16117 16643 16175 16649
rect 16117 16609 16129 16643
rect 16163 16640 16175 16643
rect 16206 16640 16212 16652
rect 16163 16612 16212 16640
rect 16163 16609 16175 16612
rect 16117 16603 16175 16609
rect 16206 16600 16212 16612
rect 16264 16600 16270 16652
rect 16390 16649 16396 16652
rect 16384 16640 16396 16649
rect 16351 16612 16396 16640
rect 16384 16603 16396 16612
rect 16390 16600 16396 16603
rect 16448 16600 16454 16652
rect 19426 16600 19432 16652
rect 19484 16640 19490 16652
rect 19628 16649 19656 16680
rect 25317 16677 25329 16711
rect 25363 16677 25375 16711
rect 25317 16671 25375 16677
rect 19521 16643 19579 16649
rect 19521 16640 19533 16643
rect 19484 16612 19533 16640
rect 19484 16600 19490 16612
rect 19521 16609 19533 16612
rect 19567 16609 19579 16643
rect 19521 16603 19579 16609
rect 19613 16643 19671 16649
rect 19613 16609 19625 16643
rect 19659 16640 19671 16643
rect 23658 16640 23664 16652
rect 19659 16612 20668 16640
rect 23619 16612 23664 16640
rect 19659 16609 19671 16612
rect 19613 16603 19671 16609
rect 4617 16575 4675 16581
rect 4617 16541 4629 16575
rect 4663 16541 4675 16575
rect 4617 16535 4675 16541
rect 6917 16575 6975 16581
rect 6917 16541 6929 16575
rect 6963 16541 6975 16575
rect 10594 16572 10600 16584
rect 10555 16544 10600 16572
rect 6917 16535 6975 16541
rect 3970 16464 3976 16516
rect 4028 16504 4034 16516
rect 4632 16504 4660 16535
rect 4028 16476 4660 16504
rect 4028 16464 4034 16476
rect 6454 16464 6460 16516
rect 6512 16504 6518 16516
rect 6932 16504 6960 16535
rect 10594 16532 10600 16544
rect 10652 16532 10658 16584
rect 10781 16575 10839 16581
rect 10781 16541 10793 16575
rect 10827 16572 10839 16575
rect 10870 16572 10876 16584
rect 10827 16544 10876 16572
rect 10827 16541 10839 16544
rect 10781 16535 10839 16541
rect 10870 16532 10876 16544
rect 10928 16532 10934 16584
rect 13354 16532 13360 16584
rect 13412 16572 13418 16584
rect 13909 16575 13967 16581
rect 13909 16572 13921 16575
rect 13412 16544 13921 16572
rect 13412 16532 13418 16544
rect 13909 16541 13921 16544
rect 13955 16541 13967 16575
rect 13909 16535 13967 16541
rect 13998 16532 14004 16584
rect 14056 16572 14062 16584
rect 19794 16572 19800 16584
rect 14056 16544 14101 16572
rect 19755 16544 19800 16572
rect 14056 16532 14062 16544
rect 19794 16532 19800 16544
rect 19852 16532 19858 16584
rect 20640 16572 20668 16612
rect 23658 16600 23664 16612
rect 23716 16600 23722 16652
rect 24394 16600 24400 16652
rect 24452 16640 24458 16652
rect 25225 16643 25283 16649
rect 25225 16640 25237 16643
rect 24452 16612 25237 16640
rect 24452 16600 24458 16612
rect 25225 16609 25237 16612
rect 25271 16609 25283 16643
rect 25225 16603 25283 16609
rect 25332 16584 25360 16671
rect 26510 16640 26516 16652
rect 26471 16612 26516 16640
rect 26510 16600 26516 16612
rect 26568 16600 26574 16652
rect 20990 16572 20996 16584
rect 20640 16544 20996 16572
rect 20990 16532 20996 16544
rect 21048 16532 21054 16584
rect 25314 16532 25320 16584
rect 25372 16532 25378 16584
rect 25501 16575 25559 16581
rect 25501 16541 25513 16575
rect 25547 16541 25559 16575
rect 25501 16535 25559 16541
rect 6512 16476 6960 16504
rect 6512 16464 6518 16476
rect 25406 16464 25412 16516
rect 25464 16504 25470 16516
rect 25516 16504 25544 16535
rect 25869 16507 25927 16513
rect 25869 16504 25881 16507
rect 25464 16476 25881 16504
rect 25464 16464 25470 16476
rect 25869 16473 25881 16476
rect 25915 16473 25927 16507
rect 25869 16467 25927 16473
rect 2041 16439 2099 16445
rect 2041 16405 2053 16439
rect 2087 16436 2099 16439
rect 2314 16436 2320 16448
rect 2087 16408 2320 16436
rect 2087 16405 2099 16408
rect 2041 16399 2099 16405
rect 2314 16396 2320 16408
rect 2372 16396 2378 16448
rect 3694 16436 3700 16448
rect 3655 16408 3700 16436
rect 3694 16396 3700 16408
rect 3752 16396 3758 16448
rect 6362 16436 6368 16448
rect 6323 16408 6368 16436
rect 6362 16396 6368 16408
rect 6420 16396 6426 16448
rect 15105 16439 15163 16445
rect 15105 16405 15117 16439
rect 15151 16436 15163 16439
rect 15378 16436 15384 16448
rect 15151 16408 15384 16436
rect 15151 16405 15163 16408
rect 15105 16399 15163 16405
rect 15378 16396 15384 16408
rect 15436 16396 15442 16448
rect 15657 16439 15715 16445
rect 15657 16405 15669 16439
rect 15703 16436 15715 16439
rect 15838 16436 15844 16448
rect 15703 16408 15844 16436
rect 15703 16405 15715 16408
rect 15657 16399 15715 16405
rect 15838 16396 15844 16408
rect 15896 16436 15902 16448
rect 18782 16436 18788 16448
rect 15896 16408 18788 16436
rect 15896 16396 15902 16408
rect 18782 16396 18788 16408
rect 18840 16396 18846 16448
rect 24670 16436 24676 16448
rect 24631 16408 24676 16436
rect 24670 16396 24676 16408
rect 24728 16396 24734 16448
rect 1104 16346 28888 16368
rect 1104 16294 5982 16346
rect 6034 16294 6046 16346
rect 6098 16294 6110 16346
rect 6162 16294 6174 16346
rect 6226 16294 15982 16346
rect 16034 16294 16046 16346
rect 16098 16294 16110 16346
rect 16162 16294 16174 16346
rect 16226 16294 25982 16346
rect 26034 16294 26046 16346
rect 26098 16294 26110 16346
rect 26162 16294 26174 16346
rect 26226 16294 28888 16346
rect 1104 16272 28888 16294
rect 3602 16232 3608 16244
rect 3563 16204 3608 16232
rect 3602 16192 3608 16204
rect 3660 16192 3666 16244
rect 4706 16232 4712 16244
rect 4667 16204 4712 16232
rect 4706 16192 4712 16204
rect 4764 16192 4770 16244
rect 5074 16232 5080 16244
rect 5035 16204 5080 16232
rect 5074 16192 5080 16204
rect 5132 16192 5138 16244
rect 5810 16192 5816 16244
rect 5868 16232 5874 16244
rect 5997 16235 6055 16241
rect 5997 16232 6009 16235
rect 5868 16204 6009 16232
rect 5868 16192 5874 16204
rect 5997 16201 6009 16204
rect 6043 16201 6055 16235
rect 6454 16232 6460 16244
rect 6415 16204 6460 16232
rect 5997 16195 6055 16201
rect 6454 16192 6460 16204
rect 6512 16192 6518 16244
rect 6914 16192 6920 16244
rect 6972 16232 6978 16244
rect 7009 16235 7067 16241
rect 7009 16232 7021 16235
rect 6972 16204 7021 16232
rect 6972 16192 6978 16204
rect 7009 16201 7021 16204
rect 7055 16201 7067 16235
rect 10502 16232 10508 16244
rect 10463 16204 10508 16232
rect 7009 16195 7067 16201
rect 10502 16192 10508 16204
rect 10560 16192 10566 16244
rect 10870 16232 10876 16244
rect 10831 16204 10876 16232
rect 10870 16192 10876 16204
rect 10928 16192 10934 16244
rect 13265 16235 13323 16241
rect 13265 16201 13277 16235
rect 13311 16232 13323 16235
rect 13630 16232 13636 16244
rect 13311 16204 13636 16232
rect 13311 16201 13323 16204
rect 13265 16195 13323 16201
rect 13630 16192 13636 16204
rect 13688 16192 13694 16244
rect 13814 16192 13820 16244
rect 13872 16232 13878 16244
rect 15013 16235 15071 16241
rect 15013 16232 15025 16235
rect 13872 16204 15025 16232
rect 13872 16192 13878 16204
rect 15013 16201 15025 16204
rect 15059 16201 15071 16235
rect 18598 16232 18604 16244
rect 18559 16204 18604 16232
rect 15013 16195 15071 16201
rect 18598 16192 18604 16204
rect 18656 16232 18662 16244
rect 20441 16235 20499 16241
rect 20441 16232 20453 16235
rect 18656 16204 20453 16232
rect 18656 16192 18662 16204
rect 2777 16167 2835 16173
rect 2777 16133 2789 16167
rect 2823 16164 2835 16167
rect 3970 16164 3976 16176
rect 2823 16136 3976 16164
rect 2823 16133 2835 16136
rect 2777 16127 2835 16133
rect 3970 16124 3976 16136
rect 4028 16164 4034 16176
rect 5353 16167 5411 16173
rect 5353 16164 5365 16167
rect 4028 16136 5365 16164
rect 4028 16124 4034 16136
rect 3694 16056 3700 16108
rect 3752 16096 3758 16108
rect 4062 16096 4068 16108
rect 3752 16068 4068 16096
rect 3752 16056 3758 16068
rect 4062 16056 4068 16068
rect 4120 16056 4126 16108
rect 4264 16105 4292 16136
rect 5353 16133 5365 16136
rect 5399 16133 5411 16167
rect 5353 16127 5411 16133
rect 10229 16167 10287 16173
rect 10229 16133 10241 16167
rect 10275 16164 10287 16167
rect 10594 16164 10600 16176
rect 10275 16136 10600 16164
rect 10275 16133 10287 16136
rect 10229 16127 10287 16133
rect 10594 16124 10600 16136
rect 10652 16124 10658 16176
rect 16114 16164 16120 16176
rect 14384 16136 16120 16164
rect 4249 16099 4307 16105
rect 4249 16065 4261 16099
rect 4295 16096 4307 16099
rect 4295 16068 4329 16096
rect 4295 16065 4307 16068
rect 4249 16059 4307 16065
rect 13262 16056 13268 16108
rect 13320 16096 13326 16108
rect 14384 16105 14412 16136
rect 16114 16124 16120 16136
rect 16172 16164 16178 16176
rect 16390 16164 16396 16176
rect 16172 16136 16396 16164
rect 16172 16124 16178 16136
rect 16390 16124 16396 16136
rect 16448 16124 16454 16176
rect 19334 16164 19340 16176
rect 19295 16136 19340 16164
rect 19334 16124 19340 16136
rect 19392 16124 19398 16176
rect 13909 16099 13967 16105
rect 13909 16096 13921 16099
rect 13320 16068 13921 16096
rect 13320 16056 13326 16068
rect 13909 16065 13921 16068
rect 13955 16096 13967 16099
rect 14369 16099 14427 16105
rect 14369 16096 14381 16099
rect 13955 16068 14381 16096
rect 13955 16065 13967 16068
rect 13909 16059 13967 16065
rect 14369 16065 14381 16068
rect 14415 16065 14427 16099
rect 15470 16096 15476 16108
rect 15431 16068 15476 16096
rect 14369 16059 14427 16065
rect 15470 16056 15476 16068
rect 15528 16056 15534 16108
rect 15565 16099 15623 16105
rect 15565 16065 15577 16099
rect 15611 16065 15623 16099
rect 15565 16059 15623 16065
rect 1397 16031 1455 16037
rect 1397 15997 1409 16031
rect 1443 16028 1455 16031
rect 1443 16000 2360 16028
rect 1443 15997 1455 16000
rect 1397 15991 1455 15997
rect 2332 15972 2360 16000
rect 8202 15988 8208 16040
rect 8260 16028 8266 16040
rect 9309 16031 9367 16037
rect 9309 16028 9321 16031
rect 8260 16000 9321 16028
rect 8260 15988 8266 16000
rect 9309 15997 9321 16000
rect 9355 16028 9367 16031
rect 9585 16031 9643 16037
rect 9585 16028 9597 16031
rect 9355 16000 9597 16028
rect 9355 15997 9367 16000
rect 9309 15991 9367 15997
rect 9585 15997 9597 16000
rect 9631 15997 9643 16031
rect 9585 15991 9643 15997
rect 13998 15988 14004 16040
rect 14056 16028 14062 16040
rect 14829 16031 14887 16037
rect 14829 16028 14841 16031
rect 14056 16000 14841 16028
rect 14056 15988 14062 16000
rect 14829 15997 14841 16000
rect 14875 15997 14887 16031
rect 15378 16028 15384 16040
rect 15339 16000 15384 16028
rect 14829 15991 14887 15997
rect 1670 15969 1676 15972
rect 1664 15960 1676 15969
rect 1631 15932 1676 15960
rect 1664 15923 1676 15932
rect 1670 15920 1676 15923
rect 1728 15920 1734 15972
rect 2314 15920 2320 15972
rect 2372 15920 2378 15972
rect 2682 15920 2688 15972
rect 2740 15960 2746 15972
rect 8754 15960 8760 15972
rect 2740 15932 8760 15960
rect 2740 15920 2746 15932
rect 8754 15920 8760 15932
rect 8812 15920 8818 15972
rect 13817 15963 13875 15969
rect 13817 15960 13829 15963
rect 12820 15932 13829 15960
rect 12820 15904 12848 15932
rect 13817 15929 13829 15932
rect 13863 15929 13875 15963
rect 14844 15960 14872 15991
rect 15378 15988 15384 16000
rect 15436 15988 15442 16040
rect 15580 16028 15608 16059
rect 15488 16000 15608 16028
rect 19352 16028 19380 16124
rect 20088 16105 20116 16204
rect 20441 16201 20453 16204
rect 20487 16201 20499 16235
rect 20990 16232 20996 16244
rect 20951 16204 20996 16232
rect 20441 16195 20499 16201
rect 20990 16192 20996 16204
rect 21048 16192 21054 16244
rect 22646 16192 22652 16244
rect 22704 16232 22710 16244
rect 22830 16232 22836 16244
rect 22704 16204 22836 16232
rect 22704 16192 22710 16204
rect 22830 16192 22836 16204
rect 22888 16232 22894 16244
rect 23017 16235 23075 16241
rect 23017 16232 23029 16235
rect 22888 16204 23029 16232
rect 22888 16192 22894 16204
rect 23017 16201 23029 16204
rect 23063 16201 23075 16235
rect 24762 16232 24768 16244
rect 23017 16195 23075 16201
rect 23676 16204 24768 16232
rect 20073 16099 20131 16105
rect 20073 16065 20085 16099
rect 20119 16096 20131 16099
rect 20714 16096 20720 16108
rect 20119 16068 20720 16096
rect 20119 16065 20131 16068
rect 20073 16059 20131 16065
rect 20714 16056 20720 16068
rect 20772 16096 20778 16108
rect 21545 16099 21603 16105
rect 21545 16096 21557 16099
rect 20772 16068 21557 16096
rect 20772 16056 20778 16068
rect 21545 16065 21557 16068
rect 21591 16065 21603 16099
rect 23032 16096 23060 16195
rect 23676 16105 23704 16204
rect 24762 16192 24768 16204
rect 24820 16192 24826 16244
rect 25041 16235 25099 16241
rect 25041 16201 25053 16235
rect 25087 16232 25099 16235
rect 25406 16232 25412 16244
rect 25087 16204 25412 16232
rect 25087 16201 25099 16204
rect 25041 16195 25099 16201
rect 25406 16192 25412 16204
rect 25464 16192 25470 16244
rect 25682 16232 25688 16244
rect 25643 16204 25688 16232
rect 25682 16192 25688 16204
rect 25740 16232 25746 16244
rect 25740 16204 26372 16232
rect 25740 16192 25746 16204
rect 24670 16124 24676 16176
rect 24728 16164 24734 16176
rect 25869 16167 25927 16173
rect 25869 16164 25881 16167
rect 24728 16136 25881 16164
rect 24728 16124 24734 16136
rect 25869 16133 25881 16136
rect 25915 16133 25927 16167
rect 25869 16127 25927 16133
rect 26344 16105 26372 16204
rect 26510 16192 26516 16244
rect 26568 16232 26574 16244
rect 26881 16235 26939 16241
rect 26881 16232 26893 16235
rect 26568 16204 26893 16232
rect 26568 16192 26574 16204
rect 26881 16201 26893 16204
rect 26927 16201 26939 16235
rect 26881 16195 26939 16201
rect 23661 16099 23719 16105
rect 23661 16096 23673 16099
rect 23032 16068 23673 16096
rect 21545 16059 21603 16065
rect 23661 16065 23673 16068
rect 23707 16065 23719 16099
rect 23661 16059 23719 16065
rect 26329 16099 26387 16105
rect 26329 16065 26341 16099
rect 26375 16065 26387 16099
rect 26329 16059 26387 16065
rect 26421 16099 26479 16105
rect 26421 16065 26433 16099
rect 26467 16065 26479 16099
rect 26421 16059 26479 16065
rect 19797 16031 19855 16037
rect 19797 16028 19809 16031
rect 19352 16000 19809 16028
rect 15194 15960 15200 15972
rect 14844 15932 15200 15960
rect 13817 15923 13875 15929
rect 15194 15920 15200 15932
rect 15252 15960 15258 15972
rect 15488 15960 15516 16000
rect 19797 15997 19809 16000
rect 19843 15997 19855 16031
rect 25314 16028 25320 16040
rect 19797 15991 19855 15997
rect 21376 16000 25320 16028
rect 19886 15960 19892 15972
rect 15252 15932 15516 15960
rect 18892 15932 19892 15960
rect 15252 15920 15258 15932
rect 18892 15904 18920 15932
rect 19886 15920 19892 15932
rect 19944 15920 19950 15972
rect 3513 15895 3571 15901
rect 3513 15861 3525 15895
rect 3559 15892 3571 15895
rect 3602 15892 3608 15904
rect 3559 15864 3608 15892
rect 3559 15861 3571 15864
rect 3513 15855 3571 15861
rect 3602 15852 3608 15864
rect 3660 15892 3666 15904
rect 3973 15895 4031 15901
rect 3973 15892 3985 15895
rect 3660 15864 3985 15892
rect 3660 15852 3666 15864
rect 3973 15861 3985 15864
rect 4019 15861 4031 15895
rect 3973 15855 4031 15861
rect 8386 15852 8392 15904
rect 8444 15892 8450 15904
rect 9401 15895 9459 15901
rect 9401 15892 9413 15895
rect 8444 15864 9413 15892
rect 8444 15852 8450 15864
rect 9401 15861 9413 15864
rect 9447 15892 9459 15895
rect 9674 15892 9680 15904
rect 9447 15864 9680 15892
rect 9447 15861 9459 15864
rect 9401 15855 9459 15861
rect 9674 15852 9680 15864
rect 9732 15852 9738 15904
rect 12802 15892 12808 15904
rect 12763 15864 12808 15892
rect 12802 15852 12808 15864
rect 12860 15852 12866 15904
rect 13354 15892 13360 15904
rect 13315 15864 13360 15892
rect 13354 15852 13360 15864
rect 13412 15852 13418 15904
rect 13630 15852 13636 15904
rect 13688 15892 13694 15904
rect 13725 15895 13783 15901
rect 13725 15892 13737 15895
rect 13688 15864 13737 15892
rect 13688 15852 13694 15864
rect 13725 15861 13737 15864
rect 13771 15861 13783 15895
rect 13725 15855 13783 15861
rect 16298 15852 16304 15904
rect 16356 15892 16362 15904
rect 16577 15895 16635 15901
rect 16577 15892 16589 15895
rect 16356 15864 16589 15892
rect 16356 15852 16362 15864
rect 16577 15861 16589 15864
rect 16623 15892 16635 15895
rect 17770 15892 17776 15904
rect 16623 15864 17776 15892
rect 16623 15861 16635 15864
rect 16577 15855 16635 15861
rect 17770 15852 17776 15864
rect 17828 15852 17834 15904
rect 18874 15892 18880 15904
rect 18835 15864 18880 15892
rect 18874 15852 18880 15864
rect 18932 15852 18938 15904
rect 19426 15892 19432 15904
rect 19387 15864 19432 15892
rect 19426 15852 19432 15864
rect 19484 15852 19490 15904
rect 19610 15852 19616 15904
rect 19668 15892 19674 15904
rect 21376 15901 21404 16000
rect 25314 15988 25320 16000
rect 25372 15988 25378 16040
rect 25406 15988 25412 16040
rect 25464 16028 25470 16040
rect 26436 16028 26464 16059
rect 25464 16000 26464 16028
rect 25464 15988 25470 16000
rect 23906 15963 23964 15969
rect 23906 15960 23918 15963
rect 23768 15932 23918 15960
rect 23768 15904 23796 15932
rect 23906 15929 23918 15932
rect 23952 15929 23964 15963
rect 23906 15923 23964 15929
rect 20809 15895 20867 15901
rect 20809 15892 20821 15895
rect 19668 15864 20821 15892
rect 19668 15852 19674 15864
rect 20809 15861 20821 15864
rect 20855 15892 20867 15895
rect 21361 15895 21419 15901
rect 21361 15892 21373 15895
rect 20855 15864 21373 15892
rect 20855 15861 20867 15864
rect 20809 15855 20867 15861
rect 21361 15861 21373 15864
rect 21407 15861 21419 15895
rect 21361 15855 21419 15861
rect 21450 15852 21456 15904
rect 21508 15892 21514 15904
rect 23477 15895 23535 15901
rect 21508 15864 21553 15892
rect 21508 15852 21514 15864
rect 23477 15861 23489 15895
rect 23523 15892 23535 15895
rect 23750 15892 23756 15904
rect 23523 15864 23756 15892
rect 23523 15861 23535 15864
rect 23477 15855 23535 15861
rect 23750 15852 23756 15864
rect 23808 15852 23814 15904
rect 26234 15892 26240 15904
rect 26195 15864 26240 15892
rect 26234 15852 26240 15864
rect 26292 15852 26298 15904
rect 1104 15802 28888 15824
rect 1104 15750 10982 15802
rect 11034 15750 11046 15802
rect 11098 15750 11110 15802
rect 11162 15750 11174 15802
rect 11226 15750 20982 15802
rect 21034 15750 21046 15802
rect 21098 15750 21110 15802
rect 21162 15750 21174 15802
rect 21226 15750 28888 15802
rect 1104 15728 28888 15750
rect 4062 15688 4068 15700
rect 4023 15660 4068 15688
rect 4062 15648 4068 15660
rect 4120 15648 4126 15700
rect 4430 15688 4436 15700
rect 4391 15660 4436 15688
rect 4430 15648 4436 15660
rect 4488 15648 4494 15700
rect 4522 15648 4528 15700
rect 4580 15688 4586 15700
rect 13262 15688 13268 15700
rect 4580 15660 4625 15688
rect 13223 15660 13268 15688
rect 4580 15648 4586 15660
rect 13262 15648 13268 15660
rect 13320 15648 13326 15700
rect 13354 15648 13360 15700
rect 13412 15688 13418 15700
rect 14277 15691 14335 15697
rect 14277 15688 14289 15691
rect 13412 15660 14289 15688
rect 13412 15648 13418 15660
rect 14277 15657 14289 15660
rect 14323 15657 14335 15691
rect 14277 15651 14335 15657
rect 15378 15648 15384 15700
rect 15436 15688 15442 15700
rect 15565 15691 15623 15697
rect 15565 15688 15577 15691
rect 15436 15660 15577 15688
rect 15436 15648 15442 15660
rect 15565 15657 15577 15660
rect 15611 15657 15623 15691
rect 15565 15651 15623 15657
rect 15746 15648 15752 15700
rect 15804 15688 15810 15700
rect 15933 15691 15991 15697
rect 15933 15688 15945 15691
rect 15804 15660 15945 15688
rect 15804 15648 15810 15660
rect 15933 15657 15945 15660
rect 15979 15657 15991 15691
rect 15933 15651 15991 15657
rect 16022 15648 16028 15700
rect 16080 15688 16086 15700
rect 18785 15691 18843 15697
rect 16080 15660 16125 15688
rect 16080 15648 16086 15660
rect 18785 15657 18797 15691
rect 18831 15688 18843 15691
rect 19426 15688 19432 15700
rect 18831 15660 19432 15688
rect 18831 15657 18843 15660
rect 18785 15651 18843 15657
rect 19426 15648 19432 15660
rect 19484 15648 19490 15700
rect 19518 15648 19524 15700
rect 19576 15688 19582 15700
rect 19705 15691 19763 15697
rect 19705 15688 19717 15691
rect 19576 15660 19717 15688
rect 19576 15648 19582 15660
rect 19705 15657 19717 15660
rect 19751 15657 19763 15691
rect 19705 15651 19763 15657
rect 21358 15648 21364 15700
rect 21416 15688 21422 15700
rect 21637 15691 21695 15697
rect 21637 15688 21649 15691
rect 21416 15660 21649 15688
rect 21416 15648 21422 15660
rect 21637 15657 21649 15660
rect 21683 15657 21695 15691
rect 21637 15651 21695 15657
rect 21910 15648 21916 15700
rect 21968 15688 21974 15700
rect 25130 15688 25136 15700
rect 21968 15660 25136 15688
rect 21968 15648 21974 15660
rect 25130 15648 25136 15660
rect 25188 15648 25194 15700
rect 25317 15691 25375 15697
rect 25317 15657 25329 15691
rect 25363 15688 25375 15691
rect 25406 15688 25412 15700
rect 25363 15660 25412 15688
rect 25363 15657 25375 15660
rect 25317 15651 25375 15657
rect 25406 15648 25412 15660
rect 25464 15648 25470 15700
rect 3697 15623 3755 15629
rect 3697 15589 3709 15623
rect 3743 15620 3755 15623
rect 3970 15620 3976 15632
rect 3743 15592 3976 15620
rect 3743 15589 3755 15592
rect 3697 15583 3755 15589
rect 3970 15580 3976 15592
rect 4028 15580 4034 15632
rect 11882 15580 11888 15632
rect 11940 15620 11946 15632
rect 12130 15623 12188 15629
rect 12130 15620 12142 15623
rect 11940 15592 12142 15620
rect 11940 15580 11946 15592
rect 12130 15589 12142 15592
rect 12176 15589 12188 15623
rect 13998 15620 14004 15632
rect 13959 15592 14004 15620
rect 12130 15583 12188 15589
rect 13998 15580 14004 15592
rect 14056 15580 14062 15632
rect 15105 15623 15163 15629
rect 15105 15589 15117 15623
rect 15151 15620 15163 15623
rect 15470 15620 15476 15632
rect 15151 15592 15476 15620
rect 15151 15589 15163 15592
rect 15105 15583 15163 15589
rect 15470 15580 15476 15592
rect 15528 15580 15534 15632
rect 19153 15623 19211 15629
rect 19153 15589 19165 15623
rect 19199 15620 19211 15623
rect 19794 15620 19800 15632
rect 19199 15592 19800 15620
rect 19199 15589 19211 15592
rect 19153 15583 19211 15589
rect 19794 15580 19800 15592
rect 19852 15580 19858 15632
rect 22738 15580 22744 15632
rect 22796 15620 22802 15632
rect 22894 15623 22952 15629
rect 22894 15620 22906 15623
rect 22796 15592 22906 15620
rect 22796 15580 22802 15592
rect 22894 15589 22906 15592
rect 22940 15589 22952 15623
rect 22894 15583 22952 15589
rect 5810 15512 5816 15564
rect 5868 15552 5874 15564
rect 5905 15555 5963 15561
rect 5905 15552 5917 15555
rect 5868 15524 5917 15552
rect 5868 15512 5874 15524
rect 5905 15521 5917 15524
rect 5951 15521 5963 15555
rect 5905 15515 5963 15521
rect 6264 15555 6322 15561
rect 6264 15521 6276 15555
rect 6310 15552 6322 15555
rect 6546 15552 6552 15564
rect 6310 15524 6552 15552
rect 6310 15521 6322 15524
rect 6264 15515 6322 15521
rect 6546 15512 6552 15524
rect 6604 15512 6610 15564
rect 9674 15552 9680 15564
rect 9635 15524 9680 15552
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 9950 15561 9956 15564
rect 9944 15552 9956 15561
rect 9911 15524 9956 15552
rect 9944 15515 9956 15524
rect 9950 15512 9956 15515
rect 10008 15512 10014 15564
rect 13170 15512 13176 15564
rect 13228 15552 13234 15564
rect 13630 15552 13636 15564
rect 13228 15524 13636 15552
rect 13228 15512 13234 15524
rect 13630 15512 13636 15524
rect 13688 15512 13694 15564
rect 17954 15512 17960 15564
rect 18012 15552 18018 15564
rect 18049 15555 18107 15561
rect 18049 15552 18061 15555
rect 18012 15524 18061 15552
rect 18012 15512 18018 15524
rect 18049 15521 18061 15524
rect 18095 15552 18107 15555
rect 19242 15552 19248 15564
rect 18095 15524 19248 15552
rect 18095 15521 18107 15524
rect 18049 15515 18107 15521
rect 19242 15512 19248 15524
rect 19300 15512 19306 15564
rect 19610 15552 19616 15564
rect 19352 15524 19616 15552
rect 1854 15484 1860 15496
rect 1815 15456 1860 15484
rect 1854 15444 1860 15456
rect 1912 15444 1918 15496
rect 4709 15487 4767 15493
rect 4709 15453 4721 15487
rect 4755 15453 4767 15487
rect 4709 15447 4767 15453
rect 1670 15416 1676 15428
rect 1583 15388 1676 15416
rect 1670 15376 1676 15388
rect 1728 15416 1734 15428
rect 4724 15416 4752 15447
rect 5718 15444 5724 15496
rect 5776 15484 5782 15496
rect 5997 15487 6055 15493
rect 5997 15484 6009 15487
rect 5776 15456 6009 15484
rect 5776 15444 5782 15456
rect 5997 15453 6009 15456
rect 6043 15453 6055 15487
rect 5997 15447 6055 15453
rect 10686 15444 10692 15496
rect 10744 15484 10750 15496
rect 11790 15484 11796 15496
rect 10744 15456 11796 15484
rect 10744 15444 10750 15456
rect 11790 15444 11796 15456
rect 11848 15484 11854 15496
rect 11885 15487 11943 15493
rect 11885 15484 11897 15487
rect 11848 15456 11897 15484
rect 11848 15444 11854 15456
rect 11885 15453 11897 15456
rect 11931 15453 11943 15487
rect 11885 15447 11943 15453
rect 16114 15444 16120 15496
rect 16172 15484 16178 15496
rect 16298 15484 16304 15496
rect 16172 15456 16304 15484
rect 16172 15444 16178 15456
rect 16298 15444 16304 15456
rect 16356 15444 16362 15496
rect 18874 15444 18880 15496
rect 18932 15484 18938 15496
rect 19352 15484 19380 15524
rect 19610 15512 19616 15524
rect 19668 15512 19674 15564
rect 21818 15552 21824 15564
rect 21779 15524 21824 15552
rect 21818 15512 21824 15524
rect 21876 15512 21882 15564
rect 22646 15552 22652 15564
rect 22607 15524 22652 15552
rect 22646 15512 22652 15524
rect 22704 15512 22710 15564
rect 26326 15512 26332 15564
rect 26384 15552 26390 15564
rect 26513 15555 26571 15561
rect 26513 15552 26525 15555
rect 26384 15524 26525 15552
rect 26384 15512 26390 15524
rect 26513 15521 26525 15524
rect 26559 15552 26571 15555
rect 27338 15552 27344 15564
rect 26559 15524 27344 15552
rect 26559 15521 26571 15524
rect 26513 15515 26571 15521
rect 27338 15512 27344 15524
rect 27396 15512 27402 15564
rect 18932 15456 19380 15484
rect 18932 15444 18938 15456
rect 19794 15444 19800 15496
rect 19852 15484 19858 15496
rect 19852 15456 19897 15484
rect 19852 15444 19858 15456
rect 4890 15416 4896 15428
rect 1728 15388 4896 15416
rect 1728 15376 1734 15388
rect 4890 15376 4896 15388
rect 4948 15416 4954 15428
rect 19245 15419 19303 15425
rect 4948 15388 5856 15416
rect 4948 15376 4954 15388
rect 2314 15308 2320 15360
rect 2372 15348 2378 15360
rect 2409 15351 2467 15357
rect 2409 15348 2421 15351
rect 2372 15320 2421 15348
rect 2372 15308 2378 15320
rect 2409 15317 2421 15320
rect 2455 15348 2467 15351
rect 5718 15348 5724 15360
rect 2455 15320 5724 15348
rect 2455 15317 2467 15320
rect 2409 15311 2467 15317
rect 5718 15308 5724 15320
rect 5776 15308 5782 15360
rect 5828 15348 5856 15388
rect 19245 15385 19257 15419
rect 19291 15416 19303 15419
rect 21085 15419 21143 15425
rect 21085 15416 21097 15419
rect 19291 15388 21097 15416
rect 19291 15385 19303 15388
rect 19245 15379 19303 15385
rect 21085 15385 21097 15388
rect 21131 15416 21143 15419
rect 21450 15416 21456 15428
rect 21131 15388 21456 15416
rect 21131 15385 21143 15388
rect 21085 15379 21143 15385
rect 21450 15376 21456 15388
rect 21508 15376 21514 15428
rect 24394 15376 24400 15428
rect 24452 15416 24458 15428
rect 24857 15419 24915 15425
rect 24857 15416 24869 15419
rect 24452 15388 24869 15416
rect 24452 15376 24458 15388
rect 24857 15385 24869 15388
rect 24903 15385 24915 15419
rect 24857 15379 24915 15385
rect 7377 15351 7435 15357
rect 7377 15348 7389 15351
rect 5828 15320 7389 15348
rect 7377 15317 7389 15320
rect 7423 15317 7435 15351
rect 8386 15348 8392 15360
rect 8347 15320 8392 15348
rect 7377 15311 7435 15317
rect 8386 15308 8392 15320
rect 8444 15308 8450 15360
rect 11054 15348 11060 15360
rect 11015 15320 11060 15348
rect 11054 15308 11060 15320
rect 11112 15308 11118 15360
rect 17770 15308 17776 15360
rect 17828 15348 17834 15360
rect 17865 15351 17923 15357
rect 17865 15348 17877 15351
rect 17828 15320 17877 15348
rect 17828 15308 17834 15320
rect 17865 15317 17877 15320
rect 17911 15317 17923 15351
rect 17865 15311 17923 15317
rect 21358 15308 21364 15360
rect 21416 15348 21422 15360
rect 22646 15348 22652 15360
rect 21416 15320 22652 15348
rect 21416 15308 21422 15320
rect 22646 15308 22652 15320
rect 22704 15308 22710 15360
rect 24029 15351 24087 15357
rect 24029 15317 24041 15351
rect 24075 15348 24087 15351
rect 24762 15348 24768 15360
rect 24075 15320 24768 15348
rect 24075 15317 24087 15320
rect 24029 15311 24087 15317
rect 24762 15308 24768 15320
rect 24820 15308 24826 15360
rect 25406 15308 25412 15360
rect 25464 15348 25470 15360
rect 25961 15351 26019 15357
rect 25961 15348 25973 15351
rect 25464 15320 25973 15348
rect 25464 15308 25470 15320
rect 25961 15317 25973 15320
rect 26007 15348 26019 15351
rect 26326 15348 26332 15360
rect 26007 15320 26332 15348
rect 26007 15317 26019 15320
rect 25961 15311 26019 15317
rect 26326 15308 26332 15320
rect 26384 15308 26390 15360
rect 26697 15351 26755 15357
rect 26697 15317 26709 15351
rect 26743 15348 26755 15351
rect 26786 15348 26792 15360
rect 26743 15320 26792 15348
rect 26743 15317 26755 15320
rect 26697 15311 26755 15317
rect 26786 15308 26792 15320
rect 26844 15308 26850 15360
rect 1104 15258 28888 15280
rect 1104 15206 5982 15258
rect 6034 15206 6046 15258
rect 6098 15206 6110 15258
rect 6162 15206 6174 15258
rect 6226 15206 15982 15258
rect 16034 15206 16046 15258
rect 16098 15206 16110 15258
rect 16162 15206 16174 15258
rect 16226 15206 25982 15258
rect 26034 15206 26046 15258
rect 26098 15206 26110 15258
rect 26162 15206 26174 15258
rect 26226 15206 28888 15258
rect 1104 15184 28888 15206
rect 4154 15104 4160 15156
rect 4212 15144 4218 15156
rect 4430 15144 4436 15156
rect 4212 15116 4436 15144
rect 4212 15104 4218 15116
rect 4430 15104 4436 15116
rect 4488 15104 4494 15156
rect 4890 15144 4896 15156
rect 4851 15116 4896 15144
rect 4890 15104 4896 15116
rect 4948 15104 4954 15156
rect 5718 15144 5724 15156
rect 5679 15116 5724 15144
rect 5718 15104 5724 15116
rect 5776 15104 5782 15156
rect 5810 15104 5816 15156
rect 5868 15144 5874 15156
rect 6457 15147 6515 15153
rect 6457 15144 6469 15147
rect 5868 15116 6469 15144
rect 5868 15104 5874 15116
rect 6457 15113 6469 15116
rect 6503 15144 6515 15147
rect 8202 15144 8208 15156
rect 6503 15116 8208 15144
rect 6503 15113 6515 15116
rect 6457 15107 6515 15113
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 8297 15147 8355 15153
rect 8297 15113 8309 15147
rect 8343 15144 8355 15147
rect 8570 15144 8576 15156
rect 8343 15116 8576 15144
rect 8343 15113 8355 15116
rect 8297 15107 8355 15113
rect 8570 15104 8576 15116
rect 8628 15104 8634 15156
rect 9674 15104 9680 15156
rect 9732 15144 9738 15156
rect 10413 15147 10471 15153
rect 10413 15144 10425 15147
rect 9732 15116 10425 15144
rect 9732 15104 9738 15116
rect 10413 15113 10425 15116
rect 10459 15144 10471 15147
rect 10594 15144 10600 15156
rect 10459 15116 10600 15144
rect 10459 15113 10471 15116
rect 10413 15107 10471 15113
rect 10594 15104 10600 15116
rect 10652 15104 10658 15156
rect 11790 15104 11796 15156
rect 11848 15144 11854 15156
rect 12618 15144 12624 15156
rect 11848 15116 12624 15144
rect 11848 15104 11854 15116
rect 12618 15104 12624 15116
rect 12676 15104 12682 15156
rect 13449 15147 13507 15153
rect 13449 15113 13461 15147
rect 13495 15144 13507 15147
rect 13814 15144 13820 15156
rect 13495 15116 13820 15144
rect 13495 15113 13507 15116
rect 13449 15107 13507 15113
rect 13814 15104 13820 15116
rect 13872 15104 13878 15156
rect 15746 15104 15752 15156
rect 15804 15144 15810 15156
rect 15933 15147 15991 15153
rect 15933 15144 15945 15147
rect 15804 15116 15945 15144
rect 15804 15104 15810 15116
rect 15933 15113 15945 15116
rect 15979 15113 15991 15147
rect 16298 15144 16304 15156
rect 16259 15116 16304 15144
rect 15933 15107 15991 15113
rect 16298 15104 16304 15116
rect 16356 15104 16362 15156
rect 17862 15144 17868 15156
rect 17823 15116 17868 15144
rect 17862 15104 17868 15116
rect 17920 15104 17926 15156
rect 18874 15144 18880 15156
rect 18835 15116 18880 15144
rect 18874 15104 18880 15116
rect 18932 15104 18938 15156
rect 19150 15144 19156 15156
rect 19111 15116 19156 15144
rect 19150 15104 19156 15116
rect 19208 15104 19214 15156
rect 19702 15144 19708 15156
rect 19352 15116 19708 15144
rect 15286 15036 15292 15088
rect 15344 15076 15350 15088
rect 15657 15079 15715 15085
rect 15657 15076 15669 15079
rect 15344 15048 15669 15076
rect 15344 15036 15350 15048
rect 15657 15045 15669 15048
rect 15703 15076 15715 15079
rect 15838 15076 15844 15088
rect 15703 15048 15844 15076
rect 15703 15045 15715 15048
rect 15657 15039 15715 15045
rect 15838 15036 15844 15048
rect 15896 15036 15902 15088
rect 17954 15036 17960 15088
rect 18012 15076 18018 15088
rect 19168 15076 19196 15104
rect 18012 15048 19196 15076
rect 18012 15036 18018 15048
rect 2314 15008 2320 15020
rect 2275 14980 2320 15008
rect 2314 14968 2320 14980
rect 2372 14968 2378 15020
rect 4157 15011 4215 15017
rect 4157 14977 4169 15011
rect 4203 15008 4215 15011
rect 4338 15008 4344 15020
rect 4203 14980 4344 15008
rect 4203 14977 4215 14980
rect 4157 14971 4215 14977
rect 4338 14968 4344 14980
rect 4396 15008 4402 15020
rect 4522 15008 4528 15020
rect 4396 14980 4528 15008
rect 4396 14968 4402 14980
rect 4522 14968 4528 14980
rect 4580 14968 4586 15020
rect 8386 15008 8392 15020
rect 8347 14980 8392 15008
rect 8386 14968 8392 14980
rect 8444 14968 8450 15020
rect 17770 14968 17776 15020
rect 17828 15008 17834 15020
rect 18874 15008 18880 15020
rect 17828 14980 18880 15008
rect 17828 14968 17834 14980
rect 18874 14968 18880 14980
rect 18932 15008 18938 15020
rect 19352 15017 19380 15116
rect 19702 15104 19708 15116
rect 19760 15144 19766 15156
rect 20714 15144 20720 15156
rect 19760 15116 20300 15144
rect 20675 15116 20720 15144
rect 19760 15104 19766 15116
rect 20272 15076 20300 15116
rect 20714 15104 20720 15116
rect 20772 15104 20778 15156
rect 21729 15147 21787 15153
rect 21729 15113 21741 15147
rect 21775 15144 21787 15147
rect 21818 15144 21824 15156
rect 21775 15116 21824 15144
rect 21775 15113 21787 15116
rect 21729 15107 21787 15113
rect 21818 15104 21824 15116
rect 21876 15104 21882 15156
rect 22738 15144 22744 15156
rect 22699 15116 22744 15144
rect 22738 15104 22744 15116
rect 22796 15104 22802 15156
rect 24486 15104 24492 15156
rect 24544 15144 24550 15156
rect 25866 15144 25872 15156
rect 24544 15116 25872 15144
rect 24544 15104 24550 15116
rect 25866 15104 25872 15116
rect 25924 15104 25930 15156
rect 27338 15144 27344 15156
rect 27299 15116 27344 15144
rect 27338 15104 27344 15116
rect 27396 15104 27402 15156
rect 20993 15079 21051 15085
rect 20993 15076 21005 15079
rect 20272 15048 21005 15076
rect 20993 15045 21005 15048
rect 21039 15045 21051 15079
rect 20993 15039 21051 15045
rect 22646 15036 22652 15088
rect 22704 15076 22710 15088
rect 23017 15079 23075 15085
rect 23017 15076 23029 15079
rect 22704 15048 23029 15076
rect 22704 15036 22710 15048
rect 23017 15045 23029 15048
rect 23063 15076 23075 15079
rect 25133 15079 25191 15085
rect 25133 15076 25145 15079
rect 23063 15048 25145 15076
rect 23063 15045 23075 15048
rect 23017 15039 23075 15045
rect 25133 15045 25145 15048
rect 25179 15045 25191 15079
rect 25133 15039 25191 15045
rect 19337 15011 19395 15017
rect 19337 15008 19349 15011
rect 18932 14980 19349 15008
rect 18932 14968 18938 14980
rect 19337 14977 19349 14980
rect 19383 14977 19395 15011
rect 25148 15008 25176 15039
rect 25406 15008 25412 15020
rect 25148 14980 25412 15008
rect 19337 14971 19395 14977
rect 25406 14968 25412 14980
rect 25464 15008 25470 15020
rect 25685 15011 25743 15017
rect 25685 15008 25697 15011
rect 25464 14980 25697 15008
rect 25464 14968 25470 14980
rect 25685 14977 25697 14980
rect 25731 14977 25743 15011
rect 25685 14971 25743 14977
rect 13814 14949 13820 14952
rect 13541 14943 13599 14949
rect 13541 14909 13553 14943
rect 13587 14909 13599 14943
rect 13808 14940 13820 14949
rect 13775 14912 13820 14940
rect 13541 14903 13599 14909
rect 13808 14903 13820 14912
rect 2225 14875 2283 14881
rect 2225 14841 2237 14875
rect 2271 14872 2283 14875
rect 2498 14872 2504 14884
rect 2271 14844 2504 14872
rect 2271 14841 2283 14844
rect 2225 14835 2283 14841
rect 2498 14832 2504 14844
rect 2556 14881 2562 14884
rect 2556 14875 2620 14881
rect 2556 14841 2574 14875
rect 2608 14841 2620 14875
rect 2556 14835 2620 14841
rect 6089 14875 6147 14881
rect 6089 14841 6101 14875
rect 6135 14872 6147 14875
rect 6546 14872 6552 14884
rect 6135 14844 6552 14872
rect 6135 14841 6147 14844
rect 6089 14835 6147 14841
rect 2556 14832 2562 14835
rect 6546 14832 6552 14844
rect 6604 14832 6610 14884
rect 8570 14832 8576 14884
rect 8628 14881 8634 14884
rect 8628 14875 8692 14881
rect 8628 14841 8646 14875
rect 8680 14841 8692 14875
rect 13556 14872 13584 14903
rect 13814 14900 13820 14903
rect 13872 14900 13878 14952
rect 13722 14872 13728 14884
rect 13556 14844 13728 14872
rect 8628 14835 8692 14841
rect 8628 14832 8634 14835
rect 13722 14832 13728 14844
rect 13780 14832 13786 14884
rect 18509 14875 18567 14881
rect 18509 14841 18521 14875
rect 18555 14872 18567 14875
rect 19582 14875 19640 14881
rect 19582 14872 19594 14875
rect 18555 14844 19594 14872
rect 18555 14841 18567 14844
rect 18509 14835 18567 14841
rect 19582 14841 19594 14844
rect 19628 14872 19640 14875
rect 19794 14872 19800 14884
rect 19628 14844 19800 14872
rect 19628 14841 19640 14844
rect 19582 14835 19640 14841
rect 19794 14832 19800 14844
rect 19852 14832 19858 14884
rect 25498 14832 25504 14884
rect 25556 14872 25562 14884
rect 25593 14875 25651 14881
rect 25593 14872 25605 14875
rect 25556 14844 25605 14872
rect 25556 14832 25562 14844
rect 25593 14841 25605 14844
rect 25639 14872 25651 14875
rect 25930 14875 25988 14881
rect 25930 14872 25942 14875
rect 25639 14844 25942 14872
rect 25639 14841 25651 14844
rect 25593 14835 25651 14841
rect 25930 14841 25942 14844
rect 25976 14841 25988 14875
rect 25930 14835 25988 14841
rect 1670 14804 1676 14816
rect 1631 14776 1676 14804
rect 1670 14764 1676 14776
rect 1728 14764 1734 14816
rect 1762 14764 1768 14816
rect 1820 14804 1826 14816
rect 3694 14804 3700 14816
rect 1820 14776 3700 14804
rect 1820 14764 1826 14776
rect 3694 14764 3700 14776
rect 3752 14764 3758 14816
rect 9214 14764 9220 14816
rect 9272 14804 9278 14816
rect 9769 14807 9827 14813
rect 9769 14804 9781 14807
rect 9272 14776 9781 14804
rect 9272 14764 9278 14776
rect 9769 14773 9781 14776
rect 9815 14804 9827 14807
rect 9950 14804 9956 14816
rect 9815 14776 9956 14804
rect 9815 14773 9827 14776
rect 9769 14767 9827 14773
rect 9950 14764 9956 14776
rect 10008 14804 10014 14816
rect 10045 14807 10103 14813
rect 10045 14804 10057 14807
rect 10008 14776 10057 14804
rect 10008 14764 10014 14776
rect 10045 14773 10057 14776
rect 10091 14773 10103 14807
rect 11882 14804 11888 14816
rect 11843 14776 11888 14804
rect 10045 14767 10103 14773
rect 11882 14764 11888 14776
rect 11940 14764 11946 14816
rect 14918 14804 14924 14816
rect 14879 14776 14924 14804
rect 14918 14764 14924 14776
rect 14976 14764 14982 14816
rect 24578 14764 24584 14816
rect 24636 14804 24642 14816
rect 27065 14807 27123 14813
rect 27065 14804 27077 14807
rect 24636 14776 27077 14804
rect 24636 14764 24642 14776
rect 27065 14773 27077 14776
rect 27111 14773 27123 14807
rect 27065 14767 27123 14773
rect 1104 14714 28888 14736
rect 1104 14662 10982 14714
rect 11034 14662 11046 14714
rect 11098 14662 11110 14714
rect 11162 14662 11174 14714
rect 11226 14662 20982 14714
rect 21034 14662 21046 14714
rect 21098 14662 21110 14714
rect 21162 14662 21174 14714
rect 21226 14662 28888 14714
rect 1104 14640 28888 14662
rect 1673 14603 1731 14609
rect 1673 14569 1685 14603
rect 1719 14600 1731 14603
rect 1762 14600 1768 14612
rect 1719 14572 1768 14600
rect 1719 14569 1731 14572
rect 1673 14563 1731 14569
rect 1762 14560 1768 14572
rect 1820 14560 1826 14612
rect 1854 14560 1860 14612
rect 1912 14600 1918 14612
rect 2225 14603 2283 14609
rect 2225 14600 2237 14603
rect 1912 14572 2237 14600
rect 1912 14560 1918 14572
rect 2225 14569 2237 14572
rect 2271 14600 2283 14603
rect 2958 14600 2964 14612
rect 2271 14572 2964 14600
rect 2271 14569 2283 14572
rect 2225 14563 2283 14569
rect 2958 14560 2964 14572
rect 3016 14560 3022 14612
rect 8113 14603 8171 14609
rect 8113 14569 8125 14603
rect 8159 14600 8171 14603
rect 8202 14600 8208 14612
rect 8159 14572 8208 14600
rect 8159 14569 8171 14572
rect 8113 14563 8171 14569
rect 8202 14560 8208 14572
rect 8260 14560 8266 14612
rect 19794 14600 19800 14612
rect 19755 14572 19800 14600
rect 19794 14560 19800 14572
rect 19852 14600 19858 14612
rect 20073 14603 20131 14609
rect 20073 14600 20085 14603
rect 19852 14572 20085 14600
rect 19852 14560 19858 14572
rect 20073 14569 20085 14572
rect 20119 14569 20131 14603
rect 20073 14563 20131 14569
rect 25406 14560 25412 14612
rect 25464 14600 25470 14612
rect 25501 14603 25559 14609
rect 25501 14600 25513 14603
rect 25464 14572 25513 14600
rect 25464 14560 25470 14572
rect 25501 14569 25513 14572
rect 25547 14569 25559 14603
rect 25501 14563 25559 14569
rect 2317 14535 2375 14541
rect 2317 14501 2329 14535
rect 2363 14532 2375 14535
rect 2590 14532 2596 14544
rect 2363 14504 2596 14532
rect 2363 14501 2375 14504
rect 2317 14495 2375 14501
rect 2590 14492 2596 14504
rect 2648 14532 2654 14544
rect 3234 14532 3240 14544
rect 2648 14504 3240 14532
rect 2648 14492 2654 14504
rect 3234 14492 3240 14504
rect 3292 14492 3298 14544
rect 5810 14541 5816 14544
rect 5804 14532 5816 14541
rect 5723 14504 5816 14532
rect 5804 14495 5816 14504
rect 5868 14532 5874 14544
rect 6822 14532 6828 14544
rect 5868 14504 6828 14532
rect 5810 14492 5816 14495
rect 5868 14492 5874 14504
rect 6822 14492 6828 14504
rect 6880 14492 6886 14544
rect 10778 14492 10784 14544
rect 10836 14541 10842 14544
rect 10836 14535 10900 14541
rect 10836 14501 10854 14535
rect 10888 14501 10900 14535
rect 10836 14495 10900 14501
rect 10836 14492 10842 14495
rect 15194 14492 15200 14544
rect 15252 14532 15258 14544
rect 15749 14535 15807 14541
rect 15749 14532 15761 14535
rect 15252 14504 15761 14532
rect 15252 14492 15258 14504
rect 15749 14501 15761 14504
rect 15795 14501 15807 14535
rect 22646 14532 22652 14544
rect 15749 14495 15807 14501
rect 22296 14504 22652 14532
rect 5537 14467 5595 14473
rect 5537 14433 5549 14467
rect 5583 14464 5595 14467
rect 5626 14464 5632 14476
rect 5583 14436 5632 14464
rect 5583 14433 5595 14436
rect 5537 14427 5595 14433
rect 5626 14424 5632 14436
rect 5684 14424 5690 14476
rect 8294 14464 8300 14476
rect 8255 14436 8300 14464
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 10594 14464 10600 14476
rect 10555 14436 10600 14464
rect 10594 14424 10600 14436
rect 10652 14424 10658 14476
rect 15657 14467 15715 14473
rect 15657 14433 15669 14467
rect 15703 14464 15715 14467
rect 16298 14464 16304 14476
rect 15703 14436 16304 14464
rect 15703 14433 15715 14436
rect 15657 14427 15715 14433
rect 16298 14424 16304 14436
rect 16356 14424 16362 14476
rect 18138 14424 18144 14476
rect 18196 14464 18202 14476
rect 22296 14473 22324 14504
rect 22646 14492 22652 14504
rect 22704 14492 22710 14544
rect 18673 14467 18731 14473
rect 18673 14464 18685 14467
rect 18196 14436 18685 14464
rect 18196 14424 18202 14436
rect 18673 14433 18685 14436
rect 18719 14433 18731 14467
rect 18673 14427 18731 14433
rect 22281 14467 22339 14473
rect 22281 14433 22293 14467
rect 22327 14433 22339 14467
rect 22281 14427 22339 14433
rect 22370 14424 22376 14476
rect 22428 14464 22434 14476
rect 22548 14467 22606 14473
rect 22548 14464 22560 14467
rect 22428 14436 22560 14464
rect 22428 14424 22434 14436
rect 22548 14433 22560 14436
rect 22594 14464 22606 14467
rect 24578 14464 24584 14476
rect 22594 14436 24584 14464
rect 22594 14433 22606 14436
rect 22548 14427 22606 14433
rect 24578 14424 24584 14436
rect 24636 14424 24642 14476
rect 2498 14396 2504 14408
rect 2459 14368 2504 14396
rect 2498 14356 2504 14368
rect 2556 14356 2562 14408
rect 15838 14396 15844 14408
rect 15799 14368 15844 14396
rect 15838 14356 15844 14368
rect 15896 14356 15902 14408
rect 18417 14399 18475 14405
rect 18417 14365 18429 14399
rect 18463 14365 18475 14399
rect 18417 14359 18475 14365
rect 1857 14263 1915 14269
rect 1857 14229 1869 14263
rect 1903 14260 1915 14263
rect 1946 14260 1952 14272
rect 1903 14232 1952 14260
rect 1903 14229 1915 14232
rect 1857 14223 1915 14229
rect 1946 14220 1952 14232
rect 2004 14220 2010 14272
rect 5074 14260 5080 14272
rect 5035 14232 5080 14260
rect 5074 14220 5080 14232
rect 5132 14220 5138 14272
rect 6914 14260 6920 14272
rect 6875 14232 6920 14260
rect 6914 14220 6920 14232
rect 6972 14220 6978 14272
rect 8665 14263 8723 14269
rect 8665 14229 8677 14263
rect 8711 14260 8723 14263
rect 9214 14260 9220 14272
rect 8711 14232 9220 14260
rect 8711 14229 8723 14232
rect 8665 14223 8723 14229
rect 9214 14220 9220 14232
rect 9272 14220 9278 14272
rect 10870 14220 10876 14272
rect 10928 14260 10934 14272
rect 11882 14260 11888 14272
rect 10928 14232 11888 14260
rect 10928 14220 10934 14232
rect 11882 14220 11888 14232
rect 11940 14260 11946 14272
rect 11977 14263 12035 14269
rect 11977 14260 11989 14263
rect 11940 14232 11989 14260
rect 11940 14220 11946 14232
rect 11977 14229 11989 14232
rect 12023 14229 12035 14263
rect 11977 14223 12035 14229
rect 13633 14263 13691 14269
rect 13633 14229 13645 14263
rect 13679 14260 13691 14263
rect 13722 14260 13728 14272
rect 13679 14232 13728 14260
rect 13679 14229 13691 14232
rect 13633 14223 13691 14229
rect 13722 14220 13728 14232
rect 13780 14220 13786 14272
rect 15102 14220 15108 14272
rect 15160 14260 15166 14272
rect 15289 14263 15347 14269
rect 15289 14260 15301 14263
rect 15160 14232 15301 14260
rect 15160 14220 15166 14232
rect 15289 14229 15301 14232
rect 15335 14229 15347 14263
rect 18432 14260 18460 14359
rect 18782 14260 18788 14272
rect 18432 14232 18788 14260
rect 15289 14223 15347 14229
rect 18782 14220 18788 14232
rect 18840 14220 18846 14272
rect 23661 14263 23719 14269
rect 23661 14229 23673 14263
rect 23707 14260 23719 14263
rect 23750 14260 23756 14272
rect 23707 14232 23756 14260
rect 23707 14229 23719 14232
rect 23661 14223 23719 14229
rect 23750 14220 23756 14232
rect 23808 14220 23814 14272
rect 1104 14170 28888 14192
rect 1104 14118 5982 14170
rect 6034 14118 6046 14170
rect 6098 14118 6110 14170
rect 6162 14118 6174 14170
rect 6226 14118 15982 14170
rect 16034 14118 16046 14170
rect 16098 14118 16110 14170
rect 16162 14118 16174 14170
rect 16226 14118 25982 14170
rect 26034 14118 26046 14170
rect 26098 14118 26110 14170
rect 26162 14118 26174 14170
rect 26226 14118 28888 14170
rect 1104 14096 28888 14118
rect 2590 14056 2596 14068
rect 2551 14028 2596 14056
rect 2590 14016 2596 14028
rect 2648 14016 2654 14068
rect 2958 14056 2964 14068
rect 2919 14028 2964 14056
rect 2958 14016 2964 14028
rect 3016 14016 3022 14068
rect 5810 14016 5816 14068
rect 5868 14056 5874 14068
rect 5997 14059 6055 14065
rect 5997 14056 6009 14059
rect 5868 14028 6009 14056
rect 5868 14016 5874 14028
rect 5997 14025 6009 14028
rect 6043 14025 6055 14059
rect 5997 14019 6055 14025
rect 10594 14016 10600 14068
rect 10652 14056 10658 14068
rect 10965 14059 11023 14065
rect 10965 14056 10977 14059
rect 10652 14028 10977 14056
rect 10652 14016 10658 14028
rect 10965 14025 10977 14028
rect 11011 14025 11023 14059
rect 10965 14019 11023 14025
rect 14829 14059 14887 14065
rect 14829 14025 14841 14059
rect 14875 14056 14887 14059
rect 16298 14056 16304 14068
rect 14875 14028 16304 14056
rect 14875 14025 14887 14028
rect 14829 14019 14887 14025
rect 16298 14016 16304 14028
rect 16356 14016 16362 14068
rect 18874 14056 18880 14068
rect 18835 14028 18880 14056
rect 18874 14016 18880 14028
rect 18932 14016 18938 14068
rect 19242 14016 19248 14068
rect 19300 14056 19306 14068
rect 19521 14059 19579 14065
rect 19521 14056 19533 14059
rect 19300 14028 19533 14056
rect 19300 14016 19306 14028
rect 19521 14025 19533 14028
rect 19567 14056 19579 14059
rect 21818 14056 21824 14068
rect 19567 14028 21824 14056
rect 19567 14025 19579 14028
rect 19521 14019 19579 14025
rect 21818 14016 21824 14028
rect 21876 14016 21882 14068
rect 22370 14056 22376 14068
rect 22331 14028 22376 14056
rect 22370 14016 22376 14028
rect 22428 14016 22434 14068
rect 22646 14056 22652 14068
rect 22607 14028 22652 14056
rect 22646 14016 22652 14028
rect 22704 14016 22710 14068
rect 24854 14016 24860 14068
rect 24912 14056 24918 14068
rect 25317 14059 25375 14065
rect 25317 14056 25329 14059
rect 24912 14028 25329 14056
rect 24912 14016 24918 14028
rect 25317 14025 25329 14028
rect 25363 14025 25375 14059
rect 25317 14019 25375 14025
rect 1762 13948 1768 14000
rect 1820 13988 1826 14000
rect 1820 13960 2176 13988
rect 1820 13948 1826 13960
rect 1670 13880 1676 13932
rect 1728 13920 1734 13932
rect 2148 13929 2176 13960
rect 4062 13948 4068 14000
rect 4120 13988 4126 14000
rect 4985 13991 5043 13997
rect 4985 13988 4997 13991
rect 4120 13960 4997 13988
rect 4120 13948 4126 13960
rect 4985 13957 4997 13960
rect 5031 13957 5043 13991
rect 4985 13951 5043 13957
rect 5718 13948 5724 14000
rect 5776 13988 5782 14000
rect 6365 13991 6423 13997
rect 6365 13988 6377 13991
rect 5776 13960 6377 13988
rect 5776 13948 5782 13960
rect 6365 13957 6377 13960
rect 6411 13957 6423 13991
rect 6365 13951 6423 13957
rect 16574 13948 16580 14000
rect 16632 13988 16638 14000
rect 16669 13991 16727 13997
rect 16669 13988 16681 13991
rect 16632 13960 16681 13988
rect 16632 13948 16638 13960
rect 16669 13957 16681 13960
rect 16715 13957 16727 13991
rect 16669 13951 16727 13957
rect 2041 13923 2099 13929
rect 2041 13920 2053 13923
rect 1728 13892 2053 13920
rect 1728 13880 1734 13892
rect 2041 13889 2053 13892
rect 2087 13889 2099 13923
rect 2041 13883 2099 13889
rect 2133 13923 2191 13929
rect 2133 13889 2145 13923
rect 2179 13889 2191 13923
rect 2133 13883 2191 13889
rect 5074 13880 5080 13932
rect 5132 13920 5138 13932
rect 5350 13920 5356 13932
rect 5132 13892 5356 13920
rect 5132 13880 5138 13892
rect 5350 13880 5356 13892
rect 5408 13920 5414 13932
rect 5445 13923 5503 13929
rect 5445 13920 5457 13923
rect 5408 13892 5457 13920
rect 5408 13880 5414 13892
rect 5445 13889 5457 13892
rect 5491 13889 5503 13923
rect 5445 13883 5503 13889
rect 5629 13923 5687 13929
rect 5629 13889 5641 13923
rect 5675 13920 5687 13923
rect 6914 13920 6920 13932
rect 5675 13892 6920 13920
rect 5675 13889 5687 13892
rect 5629 13883 5687 13889
rect 2498 13812 2504 13864
rect 2556 13852 2562 13864
rect 3421 13855 3479 13861
rect 3421 13852 3433 13855
rect 2556 13824 3433 13852
rect 2556 13812 2562 13824
rect 3421 13821 3433 13824
rect 3467 13852 3479 13855
rect 4893 13855 4951 13861
rect 4893 13852 4905 13855
rect 3467 13824 4905 13852
rect 3467 13821 3479 13824
rect 3421 13815 3479 13821
rect 4893 13821 4905 13824
rect 4939 13852 4951 13855
rect 4982 13852 4988 13864
rect 4939 13824 4988 13852
rect 4939 13821 4951 13824
rect 4893 13815 4951 13821
rect 4982 13812 4988 13824
rect 5040 13852 5046 13864
rect 5644 13852 5672 13883
rect 6914 13880 6920 13892
rect 6972 13880 6978 13932
rect 7745 13923 7803 13929
rect 7745 13889 7757 13923
rect 7791 13920 7803 13923
rect 8294 13920 8300 13932
rect 7791 13892 8300 13920
rect 7791 13889 7803 13892
rect 7745 13883 7803 13889
rect 8294 13880 8300 13892
rect 8352 13880 8358 13932
rect 9214 13920 9220 13932
rect 9175 13892 9220 13920
rect 9214 13880 9220 13892
rect 9272 13880 9278 13932
rect 24854 13880 24860 13932
rect 24912 13920 24918 13932
rect 25222 13920 25228 13932
rect 24912 13892 25228 13920
rect 24912 13880 24918 13892
rect 25222 13880 25228 13892
rect 25280 13880 25286 13932
rect 25332 13920 25360 14019
rect 25332 13892 25636 13920
rect 5040 13824 5672 13852
rect 5040 13812 5046 13824
rect 8018 13812 8024 13864
rect 8076 13852 8082 13864
rect 8113 13855 8171 13861
rect 8113 13852 8125 13855
rect 8076 13824 8125 13852
rect 8076 13812 8082 13824
rect 8113 13821 8125 13824
rect 8159 13852 8171 13855
rect 9033 13855 9091 13861
rect 9033 13852 9045 13855
rect 8159 13824 9045 13852
rect 8159 13821 8171 13824
rect 8113 13815 8171 13821
rect 9033 13821 9045 13824
rect 9079 13821 9091 13855
rect 9033 13815 9091 13821
rect 10689 13855 10747 13861
rect 10689 13821 10701 13855
rect 10735 13852 10747 13855
rect 10778 13852 10784 13864
rect 10735 13824 10784 13852
rect 10735 13821 10747 13824
rect 10689 13815 10747 13821
rect 10778 13812 10784 13824
rect 10836 13812 10842 13864
rect 15194 13852 15200 13864
rect 15155 13824 15200 13852
rect 15194 13812 15200 13824
rect 15252 13812 15258 13864
rect 15289 13855 15347 13861
rect 15289 13821 15301 13855
rect 15335 13852 15347 13855
rect 15378 13852 15384 13864
rect 15335 13824 15384 13852
rect 15335 13821 15347 13824
rect 15289 13815 15347 13821
rect 15378 13812 15384 13824
rect 15436 13812 15442 13864
rect 16945 13855 17003 13861
rect 16945 13852 16957 13855
rect 15856 13824 16957 13852
rect 15856 13796 15884 13824
rect 16945 13821 16957 13824
rect 16991 13821 17003 13855
rect 19702 13852 19708 13864
rect 19663 13824 19708 13852
rect 16945 13815 17003 13821
rect 19702 13812 19708 13824
rect 19760 13852 19766 13864
rect 19981 13855 20039 13861
rect 19981 13852 19993 13855
rect 19760 13824 19993 13852
rect 19760 13812 19766 13824
rect 19981 13821 19993 13824
rect 20027 13821 20039 13855
rect 19981 13815 20039 13821
rect 25406 13812 25412 13864
rect 25464 13852 25470 13864
rect 25501 13855 25559 13861
rect 25501 13852 25513 13855
rect 25464 13824 25513 13852
rect 25464 13812 25470 13824
rect 25501 13821 25513 13824
rect 25547 13821 25559 13855
rect 25608 13852 25636 13892
rect 25774 13861 25780 13864
rect 25757 13855 25780 13861
rect 25757 13852 25769 13855
rect 25608 13824 25769 13852
rect 25501 13815 25559 13821
rect 25757 13821 25769 13824
rect 25832 13852 25838 13864
rect 25832 13824 25905 13852
rect 25757 13815 25780 13821
rect 25774 13812 25780 13815
rect 25832 13812 25838 13824
rect 4525 13787 4583 13793
rect 4525 13753 4537 13787
rect 4571 13784 4583 13787
rect 5166 13784 5172 13796
rect 4571 13756 5172 13784
rect 4571 13753 4583 13756
rect 4525 13747 4583 13753
rect 5166 13744 5172 13756
rect 5224 13784 5230 13796
rect 5353 13787 5411 13793
rect 5353 13784 5365 13787
rect 5224 13756 5365 13784
rect 5224 13744 5230 13756
rect 5353 13753 5365 13756
rect 5399 13753 5411 13787
rect 8389 13787 8447 13793
rect 8389 13784 8401 13787
rect 5353 13747 5411 13753
rect 5644 13756 8401 13784
rect 1578 13716 1584 13728
rect 1539 13688 1584 13716
rect 1578 13676 1584 13688
rect 1636 13676 1642 13728
rect 1946 13716 1952 13728
rect 1907 13688 1952 13716
rect 1946 13676 1952 13688
rect 2004 13676 2010 13728
rect 4798 13676 4804 13728
rect 4856 13716 4862 13728
rect 5644 13716 5672 13756
rect 8389 13753 8401 13756
rect 8435 13784 8447 13787
rect 8941 13787 8999 13793
rect 8941 13784 8953 13787
rect 8435 13756 8953 13784
rect 8435 13753 8447 13756
rect 8389 13747 8447 13753
rect 8941 13753 8953 13756
rect 8987 13784 8999 13787
rect 9398 13784 9404 13796
rect 8987 13756 9404 13784
rect 8987 13753 8999 13756
rect 8941 13747 8999 13753
rect 9398 13744 9404 13756
rect 9456 13744 9462 13796
rect 14918 13784 14924 13796
rect 14384 13756 14924 13784
rect 4856 13688 5672 13716
rect 4856 13676 4862 13688
rect 5718 13676 5724 13728
rect 5776 13716 5782 13728
rect 6362 13716 6368 13728
rect 5776 13688 6368 13716
rect 5776 13676 5782 13688
rect 6362 13676 6368 13688
rect 6420 13676 6426 13728
rect 8570 13716 8576 13728
rect 8531 13688 8576 13716
rect 8570 13676 8576 13688
rect 8628 13676 8634 13728
rect 14182 13676 14188 13728
rect 14240 13716 14246 13728
rect 14384 13725 14412 13756
rect 14918 13744 14924 13756
rect 14976 13784 14982 13796
rect 15534 13787 15592 13793
rect 15534 13784 15546 13787
rect 14976 13756 15546 13784
rect 14976 13744 14982 13756
rect 15534 13753 15546 13756
rect 15580 13784 15592 13787
rect 15838 13784 15844 13796
rect 15580 13756 15844 13784
rect 15580 13753 15592 13756
rect 15534 13747 15592 13753
rect 15838 13744 15844 13756
rect 15896 13744 15902 13796
rect 14369 13719 14427 13725
rect 14369 13716 14381 13719
rect 14240 13688 14381 13716
rect 14240 13676 14246 13688
rect 14369 13685 14381 13688
rect 14415 13685 14427 13719
rect 14369 13679 14427 13685
rect 18138 13676 18144 13728
rect 18196 13716 18202 13728
rect 18417 13719 18475 13725
rect 18417 13716 18429 13719
rect 18196 13688 18429 13716
rect 18196 13676 18202 13688
rect 18417 13685 18429 13688
rect 18463 13685 18475 13719
rect 18417 13679 18475 13685
rect 26510 13676 26516 13728
rect 26568 13716 26574 13728
rect 26881 13719 26939 13725
rect 26881 13716 26893 13719
rect 26568 13688 26893 13716
rect 26568 13676 26574 13688
rect 26881 13685 26893 13688
rect 26927 13685 26939 13719
rect 26881 13679 26939 13685
rect 1104 13626 28888 13648
rect 1104 13574 10982 13626
rect 11034 13574 11046 13626
rect 11098 13574 11110 13626
rect 11162 13574 11174 13626
rect 11226 13574 20982 13626
rect 21034 13574 21046 13626
rect 21098 13574 21110 13626
rect 21162 13574 21174 13626
rect 21226 13574 28888 13626
rect 1104 13552 28888 13574
rect 1670 13472 1676 13524
rect 1728 13512 1734 13524
rect 1857 13515 1915 13521
rect 1857 13512 1869 13515
rect 1728 13484 1869 13512
rect 1728 13472 1734 13484
rect 1857 13481 1869 13484
rect 1903 13481 1915 13515
rect 1857 13475 1915 13481
rect 1946 13472 1952 13524
rect 2004 13512 2010 13524
rect 2869 13515 2927 13521
rect 2869 13512 2881 13515
rect 2004 13484 2881 13512
rect 2004 13472 2010 13484
rect 2869 13481 2881 13484
rect 2915 13481 2927 13515
rect 2869 13475 2927 13481
rect 3513 13515 3571 13521
rect 3513 13481 3525 13515
rect 3559 13512 3571 13515
rect 4062 13512 4068 13524
rect 3559 13484 4068 13512
rect 3559 13481 3571 13484
rect 3513 13475 3571 13481
rect 4062 13472 4068 13484
rect 4120 13472 4126 13524
rect 4433 13515 4491 13521
rect 4433 13481 4445 13515
rect 4479 13512 4491 13515
rect 4985 13515 5043 13521
rect 4985 13512 4997 13515
rect 4479 13484 4997 13512
rect 4479 13481 4491 13484
rect 4433 13475 4491 13481
rect 4985 13481 4997 13484
rect 5031 13512 5043 13515
rect 6089 13515 6147 13521
rect 6089 13512 6101 13515
rect 5031 13484 6101 13512
rect 5031 13481 5043 13484
rect 4985 13475 5043 13481
rect 6089 13481 6101 13484
rect 6135 13481 6147 13515
rect 6089 13475 6147 13481
rect 6457 13515 6515 13521
rect 6457 13481 6469 13515
rect 6503 13512 6515 13515
rect 6638 13512 6644 13524
rect 6503 13484 6644 13512
rect 6503 13481 6515 13484
rect 6457 13475 6515 13481
rect 6638 13472 6644 13484
rect 6696 13472 6702 13524
rect 8018 13512 8024 13524
rect 7979 13484 8024 13512
rect 8018 13472 8024 13484
rect 8076 13472 8082 13524
rect 15010 13512 15016 13524
rect 14971 13484 15016 13512
rect 15010 13472 15016 13484
rect 15068 13472 15074 13524
rect 18138 13472 18144 13524
rect 18196 13512 18202 13524
rect 19153 13515 19211 13521
rect 19153 13512 19165 13515
rect 18196 13484 19165 13512
rect 18196 13472 18202 13484
rect 19153 13481 19165 13484
rect 19199 13481 19211 13515
rect 19153 13475 19211 13481
rect 4890 13444 4896 13456
rect 4851 13416 4896 13444
rect 4890 13404 4896 13416
rect 4948 13404 4954 13456
rect 5629 13447 5687 13453
rect 5629 13413 5641 13447
rect 5675 13444 5687 13447
rect 5810 13444 5816 13456
rect 5675 13416 5816 13444
rect 5675 13413 5687 13416
rect 5629 13407 5687 13413
rect 5810 13404 5816 13416
rect 5868 13444 5874 13456
rect 11241 13447 11299 13453
rect 5868 13416 6592 13444
rect 5868 13404 5874 13416
rect 2222 13376 2228 13388
rect 2183 13348 2228 13376
rect 2222 13336 2228 13348
rect 2280 13336 2286 13388
rect 2317 13379 2375 13385
rect 2317 13345 2329 13379
rect 2363 13376 2375 13379
rect 2866 13376 2872 13388
rect 2363 13348 2872 13376
rect 2363 13345 2375 13348
rect 2317 13339 2375 13345
rect 2866 13336 2872 13348
rect 2924 13336 2930 13388
rect 6564 13376 6592 13416
rect 11241 13413 11253 13447
rect 11287 13444 11299 13447
rect 11330 13444 11336 13456
rect 11287 13416 11336 13444
rect 11287 13413 11299 13416
rect 11241 13407 11299 13413
rect 11330 13404 11336 13416
rect 11388 13404 11394 13456
rect 15746 13444 15752 13456
rect 15707 13416 15752 13444
rect 15746 13404 15752 13416
rect 15804 13404 15810 13456
rect 22922 13404 22928 13456
rect 22980 13444 22986 13456
rect 23658 13444 23664 13456
rect 22980 13416 23664 13444
rect 22980 13404 22986 13416
rect 23658 13404 23664 13416
rect 23716 13404 23722 13456
rect 8386 13376 8392 13388
rect 6564 13348 6684 13376
rect 8347 13348 8392 13376
rect 2498 13308 2504 13320
rect 2459 13280 2504 13308
rect 2498 13268 2504 13280
rect 2556 13268 2562 13320
rect 4982 13268 4988 13320
rect 5040 13308 5046 13320
rect 5077 13311 5135 13317
rect 5077 13308 5089 13311
rect 5040 13280 5089 13308
rect 5040 13268 5046 13280
rect 5077 13277 5089 13280
rect 5123 13277 5135 13311
rect 5077 13271 5135 13277
rect 5534 13268 5540 13320
rect 5592 13308 5598 13320
rect 6362 13308 6368 13320
rect 5592 13280 6368 13308
rect 5592 13268 5598 13280
rect 6362 13268 6368 13280
rect 6420 13308 6426 13320
rect 6656 13317 6684 13348
rect 8386 13336 8392 13348
rect 8444 13336 8450 13388
rect 10778 13336 10784 13388
rect 10836 13376 10842 13388
rect 11146 13376 11152 13388
rect 10836 13348 11152 13376
rect 10836 13336 10842 13348
rect 11146 13336 11152 13348
rect 11204 13376 11210 13388
rect 11204 13348 11468 13376
rect 11204 13336 11210 13348
rect 6549 13311 6607 13317
rect 6549 13308 6561 13311
rect 6420 13280 6561 13308
rect 6420 13268 6426 13280
rect 6549 13277 6561 13280
rect 6595 13277 6607 13311
rect 6549 13271 6607 13277
rect 6641 13311 6699 13317
rect 6641 13277 6653 13311
rect 6687 13308 6699 13311
rect 7006 13308 7012 13320
rect 6687 13280 7012 13308
rect 6687 13277 6699 13280
rect 6641 13271 6699 13277
rect 7006 13268 7012 13280
rect 7064 13268 7070 13320
rect 8018 13268 8024 13320
rect 8076 13308 8082 13320
rect 8481 13311 8539 13317
rect 8481 13308 8493 13311
rect 8076 13280 8493 13308
rect 8076 13268 8082 13280
rect 8481 13277 8493 13280
rect 8527 13277 8539 13311
rect 8662 13308 8668 13320
rect 8623 13280 8668 13308
rect 8481 13271 8539 13277
rect 1765 13243 1823 13249
rect 1765 13209 1777 13243
rect 1811 13240 1823 13243
rect 2516 13240 2544 13268
rect 1811 13212 2544 13240
rect 8496 13240 8524 13271
rect 8662 13268 8668 13280
rect 8720 13268 8726 13320
rect 11440 13317 11468 13348
rect 13906 13336 13912 13388
rect 13964 13376 13970 13388
rect 14001 13379 14059 13385
rect 14001 13376 14013 13379
rect 13964 13348 14013 13376
rect 13964 13336 13970 13348
rect 14001 13345 14013 13348
rect 14047 13345 14059 13379
rect 14001 13339 14059 13345
rect 14090 13336 14096 13388
rect 14148 13376 14154 13388
rect 15657 13379 15715 13385
rect 14148 13348 14193 13376
rect 14148 13336 14154 13348
rect 15657 13345 15669 13379
rect 15703 13376 15715 13379
rect 16390 13376 16396 13388
rect 15703 13348 16396 13376
rect 15703 13345 15715 13348
rect 15657 13339 15715 13345
rect 16390 13336 16396 13348
rect 16448 13336 16454 13388
rect 17770 13376 17776 13388
rect 17731 13348 17776 13376
rect 17770 13336 17776 13348
rect 17828 13336 17834 13388
rect 18046 13385 18052 13388
rect 18040 13376 18052 13385
rect 18007 13348 18052 13376
rect 18040 13339 18052 13348
rect 18046 13336 18052 13339
rect 18104 13336 18110 13388
rect 21266 13376 21272 13388
rect 21227 13348 21272 13376
rect 21266 13336 21272 13348
rect 21324 13336 21330 13388
rect 23566 13376 23572 13388
rect 23527 13348 23572 13376
rect 23566 13336 23572 13348
rect 23624 13336 23630 13388
rect 25130 13336 25136 13388
rect 25188 13376 25194 13388
rect 25225 13379 25283 13385
rect 25225 13376 25237 13379
rect 25188 13348 25237 13376
rect 25188 13336 25194 13348
rect 25225 13345 25237 13348
rect 25271 13345 25283 13379
rect 25225 13339 25283 13345
rect 11333 13311 11391 13317
rect 11333 13277 11345 13311
rect 11379 13277 11391 13311
rect 11333 13271 11391 13277
rect 11425 13311 11483 13317
rect 11425 13277 11437 13311
rect 11471 13277 11483 13311
rect 11425 13271 11483 13277
rect 9490 13240 9496 13252
rect 8496 13212 9496 13240
rect 1811 13209 1823 13212
rect 1765 13203 1823 13209
rect 9490 13200 9496 13212
rect 9548 13200 9554 13252
rect 11348 13240 11376 13271
rect 12342 13268 12348 13320
rect 12400 13308 12406 13320
rect 12437 13311 12495 13317
rect 12437 13308 12449 13311
rect 12400 13280 12449 13308
rect 12400 13268 12406 13280
rect 12437 13277 12449 13280
rect 12483 13277 12495 13311
rect 14182 13308 14188 13320
rect 14143 13280 14188 13308
rect 12437 13271 12495 13277
rect 14182 13268 14188 13280
rect 14240 13268 14246 13320
rect 15838 13308 15844 13320
rect 15799 13280 15844 13308
rect 15838 13268 15844 13280
rect 15896 13268 15902 13320
rect 21358 13308 21364 13320
rect 21319 13280 21364 13308
rect 21358 13268 21364 13280
rect 21416 13268 21422 13320
rect 21450 13268 21456 13320
rect 21508 13308 21514 13320
rect 23750 13308 23756 13320
rect 21508 13280 21553 13308
rect 23711 13280 23756 13308
rect 21508 13268 21514 13280
rect 23750 13268 23756 13280
rect 23808 13268 23814 13320
rect 24765 13311 24823 13317
rect 24765 13277 24777 13311
rect 24811 13308 24823 13311
rect 25314 13308 25320 13320
rect 24811 13280 25320 13308
rect 24811 13277 24823 13280
rect 24765 13271 24823 13277
rect 25314 13268 25320 13280
rect 25372 13268 25378 13320
rect 25498 13308 25504 13320
rect 25459 13280 25504 13308
rect 25498 13268 25504 13280
rect 25556 13308 25562 13320
rect 26510 13308 26516 13320
rect 25556 13280 26516 13308
rect 25556 13268 25562 13280
rect 26510 13268 26516 13280
rect 26568 13308 26574 13320
rect 27065 13311 27123 13317
rect 27065 13308 27077 13311
rect 26568 13280 27077 13308
rect 26568 13268 26574 13280
rect 27065 13277 27077 13280
rect 27111 13277 27123 13311
rect 27065 13271 27123 13277
rect 11514 13240 11520 13252
rect 11348 13212 11520 13240
rect 11514 13200 11520 13212
rect 11572 13200 11578 13252
rect 4522 13172 4528 13184
rect 4483 13144 4528 13172
rect 4522 13132 4528 13144
rect 4580 13132 4586 13184
rect 9122 13172 9128 13184
rect 9083 13144 9128 13172
rect 9122 13132 9128 13144
rect 9180 13132 9186 13184
rect 10042 13132 10048 13184
rect 10100 13172 10106 13184
rect 10137 13175 10195 13181
rect 10137 13172 10149 13175
rect 10100 13144 10149 13172
rect 10100 13132 10106 13144
rect 10137 13141 10149 13144
rect 10183 13141 10195 13175
rect 10137 13135 10195 13141
rect 10502 13132 10508 13184
rect 10560 13172 10566 13184
rect 10873 13175 10931 13181
rect 10873 13172 10885 13175
rect 10560 13144 10885 13172
rect 10560 13132 10566 13144
rect 10873 13141 10885 13144
rect 10919 13141 10931 13175
rect 10873 13135 10931 13141
rect 13633 13175 13691 13181
rect 13633 13141 13645 13175
rect 13679 13172 13691 13175
rect 13814 13172 13820 13184
rect 13679 13144 13820 13172
rect 13679 13141 13691 13144
rect 13633 13135 13691 13141
rect 13814 13132 13820 13144
rect 13872 13132 13878 13184
rect 15289 13175 15347 13181
rect 15289 13141 15301 13175
rect 15335 13172 15347 13175
rect 15654 13172 15660 13184
rect 15335 13144 15660 13172
rect 15335 13141 15347 13144
rect 15289 13135 15347 13141
rect 15654 13132 15660 13144
rect 15712 13132 15718 13184
rect 20898 13172 20904 13184
rect 20859 13144 20904 13172
rect 20898 13132 20904 13144
rect 20956 13132 20962 13184
rect 22554 13132 22560 13184
rect 22612 13172 22618 13184
rect 23201 13175 23259 13181
rect 23201 13172 23213 13175
rect 22612 13144 23213 13172
rect 22612 13132 22618 13144
rect 23201 13141 23213 13144
rect 23247 13141 23259 13175
rect 24302 13172 24308 13184
rect 24263 13144 24308 13172
rect 23201 13135 23259 13141
rect 24302 13132 24308 13144
rect 24360 13132 24366 13184
rect 24854 13172 24860 13184
rect 24815 13144 24860 13172
rect 24854 13132 24860 13144
rect 24912 13132 24918 13184
rect 25038 13132 25044 13184
rect 25096 13172 25102 13184
rect 25498 13172 25504 13184
rect 25096 13144 25504 13172
rect 25096 13132 25102 13144
rect 25498 13132 25504 13144
rect 25556 13132 25562 13184
rect 1104 13082 28888 13104
rect 1104 13030 5982 13082
rect 6034 13030 6046 13082
rect 6098 13030 6110 13082
rect 6162 13030 6174 13082
rect 6226 13030 15982 13082
rect 16034 13030 16046 13082
rect 16098 13030 16110 13082
rect 16162 13030 16174 13082
rect 16226 13030 25982 13082
rect 26034 13030 26046 13082
rect 26098 13030 26110 13082
rect 26162 13030 26174 13082
rect 26226 13030 28888 13082
rect 1104 13008 28888 13030
rect 4617 12971 4675 12977
rect 4617 12937 4629 12971
rect 4663 12968 4675 12971
rect 4890 12968 4896 12980
rect 4663 12940 4896 12968
rect 4663 12937 4675 12940
rect 4617 12931 4675 12937
rect 4890 12928 4896 12940
rect 4948 12928 4954 12980
rect 5166 12968 5172 12980
rect 5127 12940 5172 12968
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 6273 12971 6331 12977
rect 6273 12937 6285 12971
rect 6319 12968 6331 12971
rect 6362 12968 6368 12980
rect 6319 12940 6368 12968
rect 6319 12937 6331 12940
rect 6273 12931 6331 12937
rect 6362 12928 6368 12940
rect 6420 12928 6426 12980
rect 7006 12968 7012 12980
rect 6967 12940 7012 12968
rect 7006 12928 7012 12940
rect 7064 12928 7070 12980
rect 8573 12971 8631 12977
rect 8573 12937 8585 12971
rect 8619 12968 8631 12971
rect 10042 12968 10048 12980
rect 8619 12940 10048 12968
rect 8619 12937 8631 12940
rect 8573 12931 8631 12937
rect 10042 12928 10048 12940
rect 10100 12968 10106 12980
rect 11514 12968 11520 12980
rect 10100 12940 10640 12968
rect 11475 12940 11520 12968
rect 10100 12928 10106 12940
rect 3421 12903 3479 12909
rect 3421 12900 3433 12903
rect 2240 12872 3433 12900
rect 2038 12792 2044 12844
rect 2096 12832 2102 12844
rect 2240 12841 2268 12872
rect 3421 12869 3433 12872
rect 3467 12869 3479 12903
rect 3421 12863 3479 12869
rect 4798 12860 4804 12912
rect 4856 12900 4862 12912
rect 4985 12903 5043 12909
rect 4985 12900 4997 12903
rect 4856 12872 4997 12900
rect 4856 12860 4862 12872
rect 4985 12869 4997 12872
rect 5031 12900 5043 12903
rect 7745 12903 7803 12909
rect 5031 12872 5672 12900
rect 5031 12869 5043 12872
rect 4985 12863 5043 12869
rect 2225 12835 2283 12841
rect 2225 12832 2237 12835
rect 2096 12804 2237 12832
rect 2096 12792 2102 12804
rect 2225 12801 2237 12804
rect 2271 12801 2283 12835
rect 2225 12795 2283 12801
rect 2409 12835 2467 12841
rect 2409 12801 2421 12835
rect 2455 12832 2467 12835
rect 3050 12832 3056 12844
rect 2455 12804 3056 12832
rect 2455 12801 2467 12804
rect 2409 12795 2467 12801
rect 3050 12792 3056 12804
rect 3108 12832 3114 12844
rect 3145 12835 3203 12841
rect 3145 12832 3157 12835
rect 3108 12804 3157 12832
rect 3108 12792 3114 12804
rect 3145 12801 3157 12804
rect 3191 12801 3203 12835
rect 3145 12795 3203 12801
rect 3694 12792 3700 12844
rect 3752 12832 3758 12844
rect 5644 12841 5672 12872
rect 7745 12869 7757 12903
rect 7791 12900 7803 12903
rect 8662 12900 8668 12912
rect 7791 12872 8668 12900
rect 7791 12869 7803 12872
rect 7745 12863 7803 12869
rect 8662 12860 8668 12872
rect 8720 12860 8726 12912
rect 8754 12860 8760 12912
rect 8812 12900 8818 12912
rect 8812 12872 9628 12900
rect 8812 12860 8818 12872
rect 9600 12844 9628 12872
rect 9766 12860 9772 12912
rect 9824 12900 9830 12912
rect 10137 12903 10195 12909
rect 10137 12900 10149 12903
rect 9824 12872 10149 12900
rect 9824 12860 9830 12872
rect 10137 12869 10149 12872
rect 10183 12869 10195 12903
rect 10137 12863 10195 12869
rect 3973 12835 4031 12841
rect 3973 12832 3985 12835
rect 3752 12804 3985 12832
rect 3752 12792 3758 12804
rect 3973 12801 3985 12804
rect 4019 12801 4031 12835
rect 3973 12795 4031 12801
rect 5629 12835 5687 12841
rect 5629 12801 5641 12835
rect 5675 12801 5687 12835
rect 5810 12832 5816 12844
rect 5771 12804 5816 12832
rect 5629 12795 5687 12801
rect 5810 12792 5816 12804
rect 5868 12792 5874 12844
rect 8570 12792 8576 12844
rect 8628 12832 8634 12844
rect 8846 12832 8852 12844
rect 8628 12804 8852 12832
rect 8628 12792 8634 12804
rect 8846 12792 8852 12804
rect 8904 12832 8910 12844
rect 9033 12835 9091 12841
rect 9033 12832 9045 12835
rect 8904 12804 9045 12832
rect 8904 12792 8910 12804
rect 9033 12801 9045 12804
rect 9079 12801 9091 12835
rect 9033 12795 9091 12801
rect 9125 12835 9183 12841
rect 9125 12801 9137 12835
rect 9171 12801 9183 12835
rect 9125 12795 9183 12801
rect 1578 12724 1584 12776
rect 1636 12764 1642 12776
rect 2133 12767 2191 12773
rect 2133 12764 2145 12767
rect 1636 12736 2145 12764
rect 1636 12724 1642 12736
rect 2133 12733 2145 12736
rect 2179 12764 2191 12767
rect 2590 12764 2596 12776
rect 2179 12736 2596 12764
rect 2179 12733 2191 12736
rect 2133 12727 2191 12733
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 3789 12767 3847 12773
rect 3789 12733 3801 12767
rect 3835 12764 3847 12767
rect 3878 12764 3884 12776
rect 3835 12736 3884 12764
rect 3835 12733 3847 12736
rect 3789 12727 3847 12733
rect 3878 12724 3884 12736
rect 3936 12764 3942 12776
rect 4522 12764 4528 12776
rect 3936 12736 4528 12764
rect 3936 12724 3942 12736
rect 4522 12724 4528 12736
rect 4580 12724 4586 12776
rect 8662 12724 8668 12776
rect 8720 12764 8726 12776
rect 9140 12764 9168 12795
rect 9582 12792 9588 12844
rect 9640 12792 9646 12844
rect 10612 12841 10640 12940
rect 11514 12928 11520 12940
rect 11572 12968 11578 12980
rect 12434 12968 12440 12980
rect 11572 12940 12440 12968
rect 11572 12928 11578 12940
rect 12434 12928 12440 12940
rect 12492 12928 12498 12980
rect 14826 12968 14832 12980
rect 14787 12940 14832 12968
rect 14826 12928 14832 12940
rect 14884 12928 14890 12980
rect 15562 12928 15568 12980
rect 15620 12968 15626 12980
rect 15657 12971 15715 12977
rect 15657 12968 15669 12971
rect 15620 12940 15669 12968
rect 15620 12928 15626 12940
rect 15657 12937 15669 12940
rect 15703 12968 15715 12971
rect 15746 12968 15752 12980
rect 15703 12940 15752 12968
rect 15703 12937 15715 12940
rect 15657 12931 15715 12937
rect 15746 12928 15752 12940
rect 15804 12928 15810 12980
rect 15838 12928 15844 12980
rect 15896 12968 15902 12980
rect 16301 12971 16359 12977
rect 16301 12968 16313 12971
rect 15896 12940 16313 12968
rect 15896 12928 15902 12940
rect 16301 12937 16313 12940
rect 16347 12937 16359 12971
rect 16301 12931 16359 12937
rect 21266 12928 21272 12980
rect 21324 12968 21330 12980
rect 22373 12971 22431 12977
rect 22373 12968 22385 12971
rect 21324 12940 22385 12968
rect 21324 12928 21330 12940
rect 22373 12937 22385 12940
rect 22419 12937 22431 12971
rect 22922 12968 22928 12980
rect 22883 12940 22928 12968
rect 22373 12931 22431 12937
rect 22922 12928 22928 12940
rect 22980 12928 22986 12980
rect 23566 12928 23572 12980
rect 23624 12968 23630 12980
rect 23937 12971 23995 12977
rect 23937 12968 23949 12971
rect 23624 12940 23949 12968
rect 23624 12928 23630 12940
rect 23937 12937 23949 12940
rect 23983 12937 23995 12971
rect 23937 12931 23995 12937
rect 25314 12928 25320 12980
rect 25372 12968 25378 12980
rect 25501 12971 25559 12977
rect 25501 12968 25513 12971
rect 25372 12940 25513 12968
rect 25372 12928 25378 12940
rect 25501 12937 25513 12940
rect 25547 12937 25559 12971
rect 26510 12968 26516 12980
rect 26471 12940 26516 12968
rect 25501 12931 25559 12937
rect 26510 12928 26516 12940
rect 26568 12968 26574 12980
rect 27338 12968 27344 12980
rect 26568 12940 27344 12968
rect 26568 12928 26574 12940
rect 27338 12928 27344 12940
rect 27396 12968 27402 12980
rect 27396 12940 27568 12968
rect 27396 12928 27402 12940
rect 10778 12860 10784 12912
rect 10836 12900 10842 12912
rect 12989 12903 13047 12909
rect 12989 12900 13001 12903
rect 10836 12872 13001 12900
rect 10836 12860 10842 12872
rect 12989 12869 13001 12872
rect 13035 12869 13047 12903
rect 12989 12863 13047 12869
rect 16025 12903 16083 12909
rect 16025 12869 16037 12903
rect 16071 12900 16083 12903
rect 16390 12900 16396 12912
rect 16071 12872 16396 12900
rect 16071 12869 16083 12872
rect 16025 12863 16083 12869
rect 10597 12835 10655 12841
rect 10597 12801 10609 12835
rect 10643 12801 10655 12835
rect 10597 12795 10655 12801
rect 10689 12835 10747 12841
rect 10689 12801 10701 12835
rect 10735 12832 10747 12835
rect 10870 12832 10876 12844
rect 10735 12804 10876 12832
rect 10735 12801 10747 12804
rect 10689 12795 10747 12801
rect 9490 12764 9496 12776
rect 8720 12736 9496 12764
rect 8720 12724 8726 12736
rect 9490 12724 9496 12736
rect 9548 12724 9554 12776
rect 9677 12767 9735 12773
rect 9677 12733 9689 12767
rect 9723 12764 9735 12767
rect 10502 12764 10508 12776
rect 9723 12736 10508 12764
rect 9723 12733 9735 12736
rect 9677 12727 9735 12733
rect 10502 12724 10508 12736
rect 10560 12724 10566 12776
rect 10704 12764 10732 12795
rect 10870 12792 10876 12804
rect 10928 12792 10934 12844
rect 11146 12764 11152 12776
rect 10612 12736 10732 12764
rect 11107 12736 11152 12764
rect 1673 12699 1731 12705
rect 1673 12665 1685 12699
rect 1719 12696 1731 12699
rect 2222 12696 2228 12708
rect 1719 12668 2228 12696
rect 1719 12665 1731 12668
rect 1673 12659 1731 12665
rect 2222 12656 2228 12668
rect 2280 12696 2286 12708
rect 2958 12696 2964 12708
rect 2280 12668 2964 12696
rect 2280 12656 2286 12668
rect 2958 12656 2964 12668
rect 3016 12656 3022 12708
rect 8941 12699 8999 12705
rect 8941 12665 8953 12699
rect 8987 12696 8999 12699
rect 9122 12696 9128 12708
rect 8987 12668 9128 12696
rect 8987 12665 8999 12668
rect 8941 12659 8999 12665
rect 9122 12656 9128 12668
rect 9180 12696 9186 12708
rect 9582 12696 9588 12708
rect 9180 12668 9588 12696
rect 9180 12656 9186 12668
rect 9582 12656 9588 12668
rect 9640 12656 9646 12708
rect 10045 12699 10103 12705
rect 10045 12665 10057 12699
rect 10091 12696 10103 12699
rect 10612 12696 10640 12736
rect 11146 12724 11152 12736
rect 11204 12724 11210 12776
rect 13004 12764 13032 12863
rect 13541 12767 13599 12773
rect 13541 12764 13553 12767
rect 13004 12736 13553 12764
rect 13541 12733 13553 12736
rect 13587 12733 13599 12767
rect 13541 12727 13599 12733
rect 15654 12724 15660 12776
rect 15712 12764 15718 12776
rect 16040 12764 16068 12863
rect 16390 12860 16396 12872
rect 16448 12860 16454 12912
rect 21358 12860 21364 12912
rect 21416 12900 21422 12912
rect 22005 12903 22063 12909
rect 22005 12900 22017 12903
rect 21416 12872 22017 12900
rect 21416 12860 21422 12872
rect 22005 12869 22017 12872
rect 22051 12869 22063 12903
rect 22005 12863 22063 12869
rect 23293 12903 23351 12909
rect 23293 12869 23305 12903
rect 23339 12900 23351 12903
rect 23750 12900 23756 12912
rect 23339 12872 23756 12900
rect 23339 12869 23351 12872
rect 23293 12863 23351 12869
rect 23750 12860 23756 12872
rect 23808 12860 23814 12912
rect 23860 12872 25360 12900
rect 17497 12835 17555 12841
rect 17497 12801 17509 12835
rect 17543 12832 17555 12835
rect 17865 12835 17923 12841
rect 17865 12832 17877 12835
rect 17543 12804 17877 12832
rect 17543 12801 17555 12804
rect 17497 12795 17555 12801
rect 17865 12801 17877 12804
rect 17911 12832 17923 12835
rect 18046 12832 18052 12844
rect 17911 12804 18052 12832
rect 17911 12801 17923 12804
rect 17865 12795 17923 12801
rect 18046 12792 18052 12804
rect 18104 12832 18110 12844
rect 18782 12832 18788 12844
rect 18104 12804 18788 12832
rect 18104 12792 18110 12804
rect 18782 12792 18788 12804
rect 18840 12792 18846 12844
rect 20346 12832 20352 12844
rect 20307 12804 20352 12832
rect 20346 12792 20352 12804
rect 20404 12792 20410 12844
rect 15712 12736 16068 12764
rect 15712 12724 15718 12736
rect 20438 12724 20444 12776
rect 20496 12764 20502 12776
rect 23860 12764 23888 12872
rect 24578 12832 24584 12844
rect 24539 12804 24584 12832
rect 24578 12792 24584 12804
rect 24636 12792 24642 12844
rect 20496 12736 23888 12764
rect 24305 12767 24363 12773
rect 20496 12724 20502 12736
rect 24305 12733 24317 12767
rect 24351 12764 24363 12767
rect 24394 12764 24400 12776
rect 24351 12736 24400 12764
rect 24351 12733 24363 12736
rect 24305 12727 24363 12733
rect 24394 12724 24400 12736
rect 24452 12724 24458 12776
rect 24762 12724 24768 12776
rect 24820 12764 24826 12776
rect 24820 12736 25268 12764
rect 24820 12724 24826 12736
rect 25240 12708 25268 12736
rect 10091 12668 10640 12696
rect 10091 12665 10103 12668
rect 10045 12659 10103 12665
rect 10778 12656 10784 12708
rect 10836 12696 10842 12708
rect 14274 12696 14280 12708
rect 10836 12668 14280 12696
rect 10836 12656 10842 12668
rect 14274 12656 14280 12668
rect 14332 12656 14338 12708
rect 18506 12696 18512 12708
rect 18419 12668 18512 12696
rect 18506 12656 18512 12668
rect 18564 12696 18570 12708
rect 19521 12699 19579 12705
rect 19521 12696 19533 12699
rect 18564 12668 19533 12696
rect 18564 12656 18570 12668
rect 19521 12665 19533 12668
rect 19567 12665 19579 12699
rect 19521 12659 19579 12665
rect 19610 12656 19616 12708
rect 19668 12696 19674 12708
rect 20257 12699 20315 12705
rect 20257 12696 20269 12699
rect 19668 12668 20269 12696
rect 19668 12656 19674 12668
rect 20257 12665 20269 12668
rect 20303 12696 20315 12699
rect 20616 12699 20674 12705
rect 20616 12696 20628 12699
rect 20303 12668 20628 12696
rect 20303 12665 20315 12668
rect 20257 12659 20315 12665
rect 20616 12665 20628 12668
rect 20662 12696 20674 12699
rect 22094 12696 22100 12708
rect 20662 12668 22100 12696
rect 20662 12665 20674 12668
rect 20616 12659 20674 12665
rect 22094 12656 22100 12668
rect 22152 12656 22158 12708
rect 25038 12696 25044 12708
rect 24412 12668 25044 12696
rect 1765 12631 1823 12637
rect 1765 12597 1777 12631
rect 1811 12628 1823 12631
rect 1946 12628 1952 12640
rect 1811 12600 1952 12628
rect 1811 12597 1823 12600
rect 1765 12591 1823 12597
rect 1946 12588 1952 12600
rect 2004 12588 2010 12640
rect 2866 12628 2872 12640
rect 2827 12600 2872 12628
rect 2866 12588 2872 12600
rect 2924 12588 2930 12640
rect 3881 12631 3939 12637
rect 3881 12597 3893 12631
rect 3927 12628 3939 12631
rect 4062 12628 4068 12640
rect 3927 12600 4068 12628
rect 3927 12597 3939 12600
rect 3881 12591 3939 12597
rect 4062 12588 4068 12600
rect 4120 12588 4126 12640
rect 5258 12588 5264 12640
rect 5316 12628 5322 12640
rect 5537 12631 5595 12637
rect 5537 12628 5549 12631
rect 5316 12600 5549 12628
rect 5316 12588 5322 12600
rect 5537 12597 5549 12600
rect 5583 12597 5595 12631
rect 6638 12628 6644 12640
rect 6599 12600 6644 12628
rect 5537 12591 5595 12597
rect 6638 12588 6644 12600
rect 6696 12588 6702 12640
rect 8018 12628 8024 12640
rect 7979 12600 8024 12628
rect 8018 12588 8024 12600
rect 8076 12588 8082 12640
rect 8386 12588 8392 12640
rect 8444 12628 8450 12640
rect 8481 12631 8539 12637
rect 8481 12628 8493 12631
rect 8444 12600 8493 12628
rect 8444 12588 8450 12600
rect 8481 12597 8493 12600
rect 8527 12628 8539 12631
rect 9490 12628 9496 12640
rect 8527 12600 9496 12628
rect 8527 12597 8539 12600
rect 8481 12591 8539 12597
rect 9490 12588 9496 12600
rect 9548 12588 9554 12640
rect 10594 12588 10600 12640
rect 10652 12628 10658 12640
rect 11422 12628 11428 12640
rect 10652 12600 11428 12628
rect 10652 12588 10658 12600
rect 11422 12588 11428 12600
rect 11480 12588 11486 12640
rect 13446 12628 13452 12640
rect 13407 12600 13452 12628
rect 13446 12588 13452 12600
rect 13504 12588 13510 12640
rect 17402 12588 17408 12640
rect 17460 12628 17466 12640
rect 18141 12631 18199 12637
rect 18141 12628 18153 12631
rect 17460 12600 18153 12628
rect 17460 12588 17466 12600
rect 18141 12597 18153 12600
rect 18187 12597 18199 12631
rect 18141 12591 18199 12597
rect 18598 12588 18604 12640
rect 18656 12628 18662 12640
rect 19153 12631 19211 12637
rect 19153 12628 19165 12631
rect 18656 12600 19165 12628
rect 18656 12588 18662 12600
rect 19153 12597 19165 12600
rect 19199 12597 19211 12631
rect 19153 12591 19211 12597
rect 20806 12588 20812 12640
rect 20864 12628 20870 12640
rect 21450 12628 21456 12640
rect 20864 12600 21456 12628
rect 20864 12588 20870 12600
rect 21450 12588 21456 12600
rect 21508 12628 21514 12640
rect 21729 12631 21787 12637
rect 21729 12628 21741 12631
rect 21508 12600 21741 12628
rect 21508 12588 21514 12600
rect 21729 12597 21741 12600
rect 21775 12597 21787 12631
rect 21729 12591 21787 12597
rect 24302 12588 24308 12640
rect 24360 12628 24366 12640
rect 24412 12637 24440 12668
rect 25038 12656 25044 12668
rect 25096 12656 25102 12708
rect 25222 12656 25228 12708
rect 25280 12656 25286 12708
rect 24397 12631 24455 12637
rect 24397 12628 24409 12631
rect 24360 12600 24409 12628
rect 24360 12588 24366 12600
rect 24397 12597 24409 12600
rect 24443 12597 24455 12631
rect 24397 12591 24455 12597
rect 24949 12631 25007 12637
rect 24949 12597 24961 12631
rect 24995 12628 25007 12631
rect 25130 12628 25136 12640
rect 24995 12600 25136 12628
rect 24995 12597 25007 12600
rect 24949 12591 25007 12597
rect 25130 12588 25136 12600
rect 25188 12588 25194 12640
rect 25332 12628 25360 12872
rect 26142 12860 26148 12912
rect 26200 12900 26206 12912
rect 27065 12903 27123 12909
rect 27065 12900 27077 12903
rect 26200 12872 27077 12900
rect 26200 12860 26206 12872
rect 27065 12869 27077 12872
rect 27111 12869 27123 12903
rect 27065 12863 27123 12869
rect 25774 12792 25780 12844
rect 25832 12832 25838 12844
rect 26053 12835 26111 12841
rect 26053 12832 26065 12835
rect 25832 12804 26065 12832
rect 25832 12792 25838 12804
rect 26053 12801 26065 12804
rect 26099 12801 26111 12835
rect 27540 12832 27568 12940
rect 27617 12835 27675 12841
rect 27617 12832 27629 12835
rect 27540 12804 27629 12832
rect 26053 12795 26111 12801
rect 27617 12801 27629 12804
rect 27663 12801 27675 12835
rect 27617 12795 27675 12801
rect 25406 12724 25412 12776
rect 25464 12764 25470 12776
rect 25869 12767 25927 12773
rect 25869 12764 25881 12767
rect 25464 12736 25881 12764
rect 25464 12724 25470 12736
rect 25869 12733 25881 12736
rect 25915 12764 25927 12767
rect 25958 12764 25964 12776
rect 25915 12736 25964 12764
rect 25915 12733 25927 12736
rect 25869 12727 25927 12733
rect 25958 12724 25964 12736
rect 26016 12724 26022 12776
rect 27522 12764 27528 12776
rect 27483 12736 27528 12764
rect 27522 12724 27528 12736
rect 27580 12724 27586 12776
rect 25590 12656 25596 12708
rect 25648 12696 25654 12708
rect 26418 12696 26424 12708
rect 25648 12668 26424 12696
rect 25648 12656 25654 12668
rect 26418 12656 26424 12668
rect 26476 12656 26482 12708
rect 25409 12631 25467 12637
rect 25409 12628 25421 12631
rect 25332 12600 25421 12628
rect 25409 12597 25421 12600
rect 25455 12628 25467 12631
rect 25961 12631 26019 12637
rect 25961 12628 25973 12631
rect 25455 12600 25973 12628
rect 25455 12597 25467 12600
rect 25409 12591 25467 12597
rect 25961 12597 25973 12600
rect 26007 12597 26019 12631
rect 26878 12628 26884 12640
rect 26839 12600 26884 12628
rect 25961 12591 26019 12597
rect 26878 12588 26884 12600
rect 26936 12628 26942 12640
rect 27433 12631 27491 12637
rect 27433 12628 27445 12631
rect 26936 12600 27445 12628
rect 26936 12588 26942 12600
rect 27433 12597 27445 12600
rect 27479 12597 27491 12631
rect 27433 12591 27491 12597
rect 1104 12538 28888 12560
rect 1104 12486 10982 12538
rect 11034 12486 11046 12538
rect 11098 12486 11110 12538
rect 11162 12486 11174 12538
rect 11226 12486 20982 12538
rect 21034 12486 21046 12538
rect 21098 12486 21110 12538
rect 21162 12486 21174 12538
rect 21226 12486 28888 12538
rect 1104 12464 28888 12486
rect 3878 12424 3884 12436
rect 3839 12396 3884 12424
rect 3878 12384 3884 12396
rect 3936 12384 3942 12436
rect 4617 12427 4675 12433
rect 4617 12393 4629 12427
rect 4663 12424 4675 12427
rect 4982 12424 4988 12436
rect 4663 12396 4988 12424
rect 4663 12393 4675 12396
rect 4617 12387 4675 12393
rect 4982 12384 4988 12396
rect 5040 12384 5046 12436
rect 5534 12384 5540 12436
rect 5592 12424 5598 12436
rect 5629 12427 5687 12433
rect 5629 12424 5641 12427
rect 5592 12396 5641 12424
rect 5592 12384 5598 12396
rect 5629 12393 5641 12396
rect 5675 12393 5687 12427
rect 8662 12424 8668 12436
rect 8623 12396 8668 12424
rect 5629 12387 5687 12393
rect 8662 12384 8668 12396
rect 8720 12384 8726 12436
rect 8846 12384 8852 12436
rect 8904 12424 8910 12436
rect 8941 12427 8999 12433
rect 8941 12424 8953 12427
rect 8904 12396 8953 12424
rect 8904 12384 8910 12396
rect 8941 12393 8953 12396
rect 8987 12393 8999 12427
rect 9674 12424 9680 12436
rect 9635 12396 9680 12424
rect 8941 12387 8999 12393
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 10778 12424 10784 12436
rect 10739 12396 10784 12424
rect 10778 12384 10784 12396
rect 10836 12384 10842 12436
rect 11149 12427 11207 12433
rect 11149 12393 11161 12427
rect 11195 12424 11207 12427
rect 11330 12424 11336 12436
rect 11195 12396 11336 12424
rect 11195 12393 11207 12396
rect 11149 12387 11207 12393
rect 11330 12384 11336 12396
rect 11388 12424 11394 12436
rect 11425 12427 11483 12433
rect 11425 12424 11437 12427
rect 11388 12396 11437 12424
rect 11388 12384 11394 12396
rect 11425 12393 11437 12396
rect 11471 12393 11483 12427
rect 11425 12387 11483 12393
rect 11793 12427 11851 12433
rect 11793 12393 11805 12427
rect 11839 12424 11851 12427
rect 11882 12424 11888 12436
rect 11839 12396 11888 12424
rect 11839 12393 11851 12396
rect 11793 12387 11851 12393
rect 11882 12384 11888 12396
rect 11940 12424 11946 12436
rect 12342 12424 12348 12436
rect 11940 12396 12348 12424
rect 11940 12384 11946 12396
rect 12342 12384 12348 12396
rect 12400 12384 12406 12436
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 14093 12427 14151 12433
rect 12492 12396 12537 12424
rect 12492 12384 12498 12396
rect 14093 12393 14105 12427
rect 14139 12424 14151 12427
rect 14182 12424 14188 12436
rect 14139 12396 14188 12424
rect 14139 12393 14151 12396
rect 14093 12387 14151 12393
rect 14182 12384 14188 12396
rect 14240 12384 14246 12436
rect 17402 12424 17408 12436
rect 17363 12396 17408 12424
rect 17402 12384 17408 12396
rect 17460 12384 17466 12436
rect 17770 12384 17776 12436
rect 17828 12424 17834 12436
rect 17957 12427 18015 12433
rect 17957 12424 17969 12427
rect 17828 12396 17969 12424
rect 17828 12384 17834 12396
rect 17957 12393 17969 12396
rect 18003 12393 18015 12427
rect 18506 12424 18512 12436
rect 18467 12396 18512 12424
rect 17957 12387 18015 12393
rect 18506 12384 18512 12396
rect 18564 12384 18570 12436
rect 20346 12424 20352 12436
rect 20307 12396 20352 12424
rect 20346 12384 20352 12396
rect 20404 12384 20410 12436
rect 20806 12384 20812 12436
rect 20864 12424 20870 12436
rect 21085 12427 21143 12433
rect 21085 12424 21097 12427
rect 20864 12396 21097 12424
rect 20864 12384 20870 12396
rect 21085 12393 21097 12396
rect 21131 12393 21143 12427
rect 21085 12387 21143 12393
rect 21358 12384 21364 12436
rect 21416 12424 21422 12436
rect 21453 12427 21511 12433
rect 21453 12424 21465 12427
rect 21416 12396 21465 12424
rect 21416 12384 21422 12396
rect 21453 12393 21465 12396
rect 21499 12393 21511 12427
rect 21453 12387 21511 12393
rect 21634 12384 21640 12436
rect 21692 12424 21698 12436
rect 21818 12424 21824 12436
rect 21692 12396 21824 12424
rect 21692 12384 21698 12396
rect 21818 12384 21824 12396
rect 21876 12424 21882 12436
rect 21913 12427 21971 12433
rect 21913 12424 21925 12427
rect 21876 12396 21925 12424
rect 21876 12384 21882 12396
rect 21913 12393 21925 12396
rect 21959 12393 21971 12427
rect 23566 12424 23572 12436
rect 23527 12396 23572 12424
rect 21913 12387 21971 12393
rect 23566 12384 23572 12396
rect 23624 12384 23630 12436
rect 23658 12384 23664 12436
rect 23716 12424 23722 12436
rect 24489 12427 24547 12433
rect 24489 12424 24501 12427
rect 23716 12396 24501 12424
rect 23716 12384 23722 12396
rect 24489 12393 24501 12396
rect 24535 12393 24547 12427
rect 24762 12424 24768 12436
rect 24489 12387 24547 12393
rect 24688 12396 24768 12424
rect 1762 12316 1768 12368
rect 1820 12365 1826 12368
rect 1820 12359 1884 12365
rect 1820 12325 1838 12359
rect 1872 12325 1884 12359
rect 1820 12319 1884 12325
rect 3513 12359 3571 12365
rect 3513 12325 3525 12359
rect 3559 12356 3571 12359
rect 3694 12356 3700 12368
rect 3559 12328 3700 12356
rect 3559 12325 3571 12328
rect 3513 12319 3571 12325
rect 1820 12316 1826 12319
rect 3694 12316 3700 12328
rect 3752 12316 3758 12368
rect 6089 12359 6147 12365
rect 6089 12356 6101 12359
rect 5644 12328 6101 12356
rect 5644 12300 5672 12328
rect 6089 12325 6101 12328
rect 6135 12356 6147 12359
rect 8018 12356 8024 12368
rect 6135 12328 8024 12356
rect 6135 12325 6147 12328
rect 6089 12319 6147 12325
rect 8018 12316 8024 12328
rect 8076 12316 8082 12368
rect 15657 12359 15715 12365
rect 15657 12325 15669 12359
rect 15703 12356 15715 12359
rect 15838 12356 15844 12368
rect 15703 12328 15844 12356
rect 15703 12325 15715 12328
rect 15657 12319 15715 12325
rect 15838 12316 15844 12328
rect 15896 12316 15902 12368
rect 18414 12316 18420 12368
rect 18472 12356 18478 12368
rect 18877 12359 18935 12365
rect 18877 12356 18889 12359
rect 18472 12328 18889 12356
rect 18472 12316 18478 12328
rect 18877 12325 18889 12328
rect 18923 12325 18935 12359
rect 18877 12319 18935 12325
rect 24029 12359 24087 12365
rect 24029 12325 24041 12359
rect 24075 12356 24087 12359
rect 24118 12356 24124 12368
rect 24075 12328 24124 12356
rect 24075 12325 24087 12328
rect 24029 12319 24087 12325
rect 24118 12316 24124 12328
rect 24176 12356 24182 12368
rect 24578 12356 24584 12368
rect 24176 12328 24584 12356
rect 24176 12316 24182 12328
rect 1581 12291 1639 12297
rect 1581 12257 1593 12291
rect 1627 12288 1639 12291
rect 2222 12288 2228 12300
rect 1627 12260 2228 12288
rect 1627 12257 1639 12260
rect 1581 12251 1639 12257
rect 2222 12248 2228 12260
rect 2280 12248 2286 12300
rect 5626 12248 5632 12300
rect 5684 12248 5690 12300
rect 5994 12288 6000 12300
rect 5955 12260 6000 12288
rect 5994 12248 6000 12260
rect 6052 12248 6058 12300
rect 10042 12288 10048 12300
rect 10003 12260 10048 12288
rect 10042 12248 10048 12260
rect 10100 12248 10106 12300
rect 12526 12248 12532 12300
rect 12584 12288 12590 12300
rect 12802 12288 12808 12300
rect 12584 12260 12808 12288
rect 12584 12248 12590 12260
rect 12802 12248 12808 12260
rect 12860 12248 12866 12300
rect 13630 12288 13636 12300
rect 13591 12260 13636 12288
rect 13630 12248 13636 12260
rect 13688 12248 13694 12300
rect 13814 12248 13820 12300
rect 13872 12288 13878 12300
rect 14090 12288 14096 12300
rect 13872 12260 14096 12288
rect 13872 12248 13878 12260
rect 14090 12248 14096 12260
rect 14148 12288 14154 12300
rect 14645 12291 14703 12297
rect 14645 12288 14657 12291
rect 14148 12260 14657 12288
rect 14148 12248 14154 12260
rect 14645 12257 14657 12260
rect 14691 12257 14703 12291
rect 15102 12288 15108 12300
rect 14645 12251 14703 12257
rect 14752 12260 15108 12288
rect 5810 12180 5816 12232
rect 5868 12220 5874 12232
rect 6181 12223 6239 12229
rect 6181 12220 6193 12223
rect 5868 12192 6193 12220
rect 5868 12180 5874 12192
rect 6181 12189 6193 12192
rect 6227 12220 6239 12223
rect 6362 12220 6368 12232
rect 6227 12192 6368 12220
rect 6227 12189 6239 12192
rect 6181 12183 6239 12189
rect 6362 12180 6368 12192
rect 6420 12180 6426 12232
rect 9674 12180 9680 12232
rect 9732 12220 9738 12232
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 9732 12192 10149 12220
rect 9732 12180 9738 12192
rect 10137 12189 10149 12192
rect 10183 12189 10195 12223
rect 10137 12183 10195 12189
rect 10226 12180 10232 12232
rect 10284 12220 10290 12232
rect 10284 12192 10329 12220
rect 10284 12180 10290 12192
rect 11422 12180 11428 12232
rect 11480 12220 11486 12232
rect 11885 12223 11943 12229
rect 11885 12220 11897 12223
rect 11480 12192 11897 12220
rect 11480 12180 11486 12192
rect 11885 12189 11897 12192
rect 11931 12189 11943 12223
rect 11885 12183 11943 12189
rect 11977 12223 12035 12229
rect 11977 12189 11989 12223
rect 12023 12189 12035 12223
rect 12894 12220 12900 12232
rect 12855 12192 12900 12220
rect 11977 12183 12035 12189
rect 10244 12152 10272 12180
rect 11992 12152 12020 12183
rect 12894 12180 12900 12192
rect 12952 12180 12958 12232
rect 12989 12223 13047 12229
rect 12989 12189 13001 12223
rect 13035 12189 13047 12223
rect 12989 12183 13047 12189
rect 12434 12152 12440 12164
rect 10244 12124 12440 12152
rect 12434 12112 12440 12124
rect 12492 12152 12498 12164
rect 13004 12152 13032 12183
rect 14550 12180 14556 12232
rect 14608 12220 14614 12232
rect 14752 12229 14780 12260
rect 15102 12248 15108 12260
rect 15160 12248 15166 12300
rect 15746 12248 15752 12300
rect 15804 12288 15810 12300
rect 16669 12291 16727 12297
rect 16669 12288 16681 12291
rect 15804 12260 16681 12288
rect 15804 12248 15810 12260
rect 16669 12257 16681 12260
rect 16715 12257 16727 12291
rect 16669 12251 16727 12257
rect 17034 12248 17040 12300
rect 17092 12288 17098 12300
rect 17310 12288 17316 12300
rect 17092 12260 17316 12288
rect 17092 12248 17098 12260
rect 17310 12248 17316 12260
rect 17368 12248 17374 12300
rect 21634 12248 21640 12300
rect 21692 12288 21698 12300
rect 21821 12291 21879 12297
rect 21821 12288 21833 12291
rect 21692 12260 21833 12288
rect 21692 12248 21698 12260
rect 21821 12257 21833 12260
rect 21867 12257 21879 12291
rect 21821 12251 21879 12257
rect 14737 12223 14795 12229
rect 14737 12220 14749 12223
rect 14608 12192 14749 12220
rect 14608 12180 14614 12192
rect 14737 12189 14749 12192
rect 14783 12189 14795 12223
rect 14918 12220 14924 12232
rect 14879 12192 14924 12220
rect 14737 12183 14795 12189
rect 14918 12180 14924 12192
rect 14976 12220 14982 12232
rect 15841 12223 15899 12229
rect 15841 12220 15853 12223
rect 14976 12192 15853 12220
rect 14976 12180 14982 12192
rect 15841 12189 15853 12192
rect 15887 12220 15899 12223
rect 16574 12220 16580 12232
rect 15887 12192 16580 12220
rect 15887 12189 15899 12192
rect 15841 12183 15899 12189
rect 16574 12180 16580 12192
rect 16632 12180 16638 12232
rect 17126 12180 17132 12232
rect 17184 12220 17190 12232
rect 17589 12223 17647 12229
rect 17589 12220 17601 12223
rect 17184 12192 17601 12220
rect 17184 12180 17190 12192
rect 17589 12189 17601 12192
rect 17635 12220 17647 12223
rect 18138 12220 18144 12232
rect 17635 12192 18144 12220
rect 17635 12189 17647 12192
rect 17589 12183 17647 12189
rect 18138 12180 18144 12192
rect 18196 12180 18202 12232
rect 18417 12223 18475 12229
rect 18417 12189 18429 12223
rect 18463 12220 18475 12223
rect 18966 12220 18972 12232
rect 18463 12192 18972 12220
rect 18463 12189 18475 12192
rect 18417 12183 18475 12189
rect 18966 12180 18972 12192
rect 19024 12180 19030 12232
rect 19150 12220 19156 12232
rect 19111 12192 19156 12220
rect 19150 12180 19156 12192
rect 19208 12180 19214 12232
rect 22094 12220 22100 12232
rect 22055 12192 22100 12220
rect 22094 12180 22100 12192
rect 22152 12180 22158 12232
rect 23014 12220 23020 12232
rect 22975 12192 23020 12220
rect 23014 12180 23020 12192
rect 23072 12180 23078 12232
rect 12492 12124 13032 12152
rect 24504 12152 24532 12328
rect 24578 12316 24584 12328
rect 24636 12316 24642 12368
rect 24578 12180 24584 12232
rect 24636 12220 24642 12232
rect 24688 12220 24716 12396
rect 24762 12384 24768 12396
rect 24820 12424 24826 12436
rect 24949 12427 25007 12433
rect 24949 12424 24961 12427
rect 24820 12396 24961 12424
rect 24820 12384 24826 12396
rect 24949 12393 24961 12396
rect 24995 12393 25007 12427
rect 24949 12387 25007 12393
rect 25774 12384 25780 12436
rect 25832 12424 25838 12436
rect 25869 12427 25927 12433
rect 25869 12424 25881 12427
rect 25832 12396 25881 12424
rect 25832 12384 25838 12396
rect 25869 12393 25881 12396
rect 25915 12393 25927 12427
rect 25869 12387 25927 12393
rect 27157 12427 27215 12433
rect 27157 12393 27169 12427
rect 27203 12424 27215 12427
rect 27522 12424 27528 12436
rect 27203 12396 27528 12424
rect 27203 12393 27215 12396
rect 27157 12387 27215 12393
rect 27522 12384 27528 12396
rect 27580 12384 27586 12436
rect 24857 12359 24915 12365
rect 24857 12325 24869 12359
rect 24903 12356 24915 12359
rect 26142 12356 26148 12368
rect 24903 12328 26148 12356
rect 24903 12325 24915 12328
rect 24857 12319 24915 12325
rect 24636 12192 24716 12220
rect 25041 12223 25099 12229
rect 24636 12180 24642 12192
rect 25041 12189 25053 12223
rect 25087 12189 25099 12223
rect 25041 12183 25099 12189
rect 25056 12152 25084 12183
rect 24504 12124 25084 12152
rect 12492 12112 12498 12124
rect 2961 12087 3019 12093
rect 2961 12053 2973 12087
rect 3007 12084 3019 12087
rect 3050 12084 3056 12096
rect 3007 12056 3056 12084
rect 3007 12053 3019 12056
rect 2961 12047 3019 12053
rect 3050 12044 3056 12056
rect 3108 12044 3114 12096
rect 5258 12084 5264 12096
rect 5171 12056 5264 12084
rect 5258 12044 5264 12056
rect 5316 12084 5322 12096
rect 5442 12084 5448 12096
rect 5316 12056 5448 12084
rect 5316 12044 5322 12056
rect 5442 12044 5448 12056
rect 5500 12044 5506 12096
rect 14274 12084 14280 12096
rect 14235 12056 14280 12084
rect 14274 12044 14280 12056
rect 14332 12044 14338 12096
rect 14366 12044 14372 12096
rect 14424 12084 14430 12096
rect 15289 12087 15347 12093
rect 15289 12084 15301 12087
rect 14424 12056 15301 12084
rect 14424 12044 14430 12056
rect 15289 12053 15301 12056
rect 15335 12053 15347 12087
rect 16390 12084 16396 12096
rect 16351 12056 16396 12084
rect 15289 12047 15347 12053
rect 16390 12044 16396 12056
rect 16448 12044 16454 12096
rect 16945 12087 17003 12093
rect 16945 12053 16957 12087
rect 16991 12084 17003 12087
rect 17678 12084 17684 12096
rect 16991 12056 17684 12084
rect 16991 12053 17003 12056
rect 16945 12047 17003 12053
rect 17678 12044 17684 12056
rect 17736 12044 17742 12096
rect 24302 12084 24308 12096
rect 24263 12056 24308 12084
rect 24302 12044 24308 12056
rect 24360 12044 24366 12096
rect 24946 12044 24952 12096
rect 25004 12084 25010 12096
rect 25148 12084 25176 12328
rect 26142 12316 26148 12328
rect 26200 12316 26206 12368
rect 26513 12291 26571 12297
rect 26513 12257 26525 12291
rect 26559 12288 26571 12291
rect 26878 12288 26884 12300
rect 26559 12260 26884 12288
rect 26559 12257 26571 12260
rect 26513 12251 26571 12257
rect 26878 12248 26884 12260
rect 26936 12248 26942 12300
rect 25004 12056 25176 12084
rect 25004 12044 25010 12056
rect 25406 12044 25412 12096
rect 25464 12084 25470 12096
rect 25501 12087 25559 12093
rect 25501 12084 25513 12087
rect 25464 12056 25513 12084
rect 25464 12044 25470 12056
rect 25501 12053 25513 12056
rect 25547 12053 25559 12087
rect 25501 12047 25559 12053
rect 25774 12044 25780 12096
rect 25832 12084 25838 12096
rect 26697 12087 26755 12093
rect 26697 12084 26709 12087
rect 25832 12056 26709 12084
rect 25832 12044 25838 12056
rect 26697 12053 26709 12056
rect 26743 12053 26755 12087
rect 26697 12047 26755 12053
rect 1104 11994 28888 12016
rect 1104 11942 5982 11994
rect 6034 11942 6046 11994
rect 6098 11942 6110 11994
rect 6162 11942 6174 11994
rect 6226 11942 15982 11994
rect 16034 11942 16046 11994
rect 16098 11942 16110 11994
rect 16162 11942 16174 11994
rect 16226 11942 25982 11994
rect 26034 11942 26046 11994
rect 26098 11942 26110 11994
rect 26162 11942 26174 11994
rect 26226 11942 28888 11994
rect 1104 11920 28888 11942
rect 1762 11840 1768 11892
rect 1820 11880 1826 11892
rect 2409 11883 2467 11889
rect 2409 11880 2421 11883
rect 1820 11852 2421 11880
rect 1820 11840 1826 11852
rect 2409 11849 2421 11852
rect 2455 11849 2467 11883
rect 2409 11843 2467 11849
rect 2590 11840 2596 11892
rect 2648 11880 2654 11892
rect 2777 11883 2835 11889
rect 2777 11880 2789 11883
rect 2648 11852 2789 11880
rect 2648 11840 2654 11852
rect 2777 11849 2789 11852
rect 2823 11849 2835 11883
rect 2777 11843 2835 11849
rect 3234 11840 3240 11892
rect 3292 11880 3298 11892
rect 5626 11880 5632 11892
rect 3292 11852 5632 11880
rect 3292 11840 3298 11852
rect 5626 11840 5632 11852
rect 5684 11840 5690 11892
rect 6362 11880 6368 11892
rect 6323 11852 6368 11880
rect 6362 11840 6368 11852
rect 6420 11840 6426 11892
rect 9769 11883 9827 11889
rect 9769 11849 9781 11883
rect 9815 11880 9827 11883
rect 10042 11880 10048 11892
rect 9815 11852 10048 11880
rect 9815 11849 9827 11852
rect 9769 11843 9827 11849
rect 10042 11840 10048 11852
rect 10100 11840 10106 11892
rect 11882 11880 11888 11892
rect 11843 11852 11888 11880
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 12894 11840 12900 11892
rect 12952 11880 12958 11892
rect 12989 11883 13047 11889
rect 12989 11880 13001 11883
rect 12952 11852 13001 11880
rect 12952 11840 12958 11852
rect 12989 11849 13001 11852
rect 13035 11849 13047 11883
rect 15378 11880 15384 11892
rect 15291 11852 15384 11880
rect 12989 11843 13047 11849
rect 15378 11840 15384 11852
rect 15436 11880 15442 11892
rect 15838 11880 15844 11892
rect 15436 11852 15844 11880
rect 15436 11840 15442 11852
rect 15838 11840 15844 11852
rect 15896 11840 15902 11892
rect 17037 11883 17095 11889
rect 17037 11849 17049 11883
rect 17083 11880 17095 11883
rect 17126 11880 17132 11892
rect 17083 11852 17132 11880
rect 17083 11849 17095 11852
rect 17037 11843 17095 11849
rect 17126 11840 17132 11852
rect 17184 11840 17190 11892
rect 17402 11880 17408 11892
rect 17363 11852 17408 11880
rect 17402 11840 17408 11852
rect 17460 11840 17466 11892
rect 18509 11883 18567 11889
rect 18509 11849 18521 11883
rect 18555 11880 18567 11883
rect 18598 11880 18604 11892
rect 18555 11852 18604 11880
rect 18555 11849 18567 11852
rect 18509 11843 18567 11849
rect 18598 11840 18604 11852
rect 18656 11840 18662 11892
rect 20530 11840 20536 11892
rect 20588 11880 20594 11892
rect 20901 11883 20959 11889
rect 20901 11880 20913 11883
rect 20588 11852 20913 11880
rect 20588 11840 20594 11852
rect 20901 11849 20913 11852
rect 20947 11849 20959 11883
rect 20901 11843 20959 11849
rect 2041 11815 2099 11821
rect 2041 11781 2053 11815
rect 2087 11812 2099 11815
rect 2498 11812 2504 11824
rect 2087 11784 2504 11812
rect 2087 11781 2099 11784
rect 2041 11775 2099 11781
rect 1397 11679 1455 11685
rect 1397 11645 1409 11679
rect 1443 11676 1455 11679
rect 2056 11676 2084 11775
rect 2498 11772 2504 11784
rect 2556 11772 2562 11824
rect 6089 11815 6147 11821
rect 6089 11781 6101 11815
rect 6135 11812 6147 11815
rect 6270 11812 6276 11824
rect 6135 11784 6276 11812
rect 6135 11781 6147 11784
rect 6089 11775 6147 11781
rect 6270 11772 6276 11784
rect 6328 11772 6334 11824
rect 12713 11815 12771 11821
rect 12713 11781 12725 11815
rect 12759 11812 12771 11815
rect 12802 11812 12808 11824
rect 12759 11784 12808 11812
rect 12759 11781 12771 11784
rect 12713 11775 12771 11781
rect 12802 11772 12808 11784
rect 12860 11812 12866 11824
rect 16666 11812 16672 11824
rect 12860 11784 16672 11812
rect 12860 11772 12866 11784
rect 9033 11747 9091 11753
rect 9033 11713 9045 11747
rect 9079 11744 9091 11747
rect 10410 11744 10416 11756
rect 9079 11716 10416 11744
rect 9079 11713 9091 11716
rect 9033 11707 9091 11713
rect 10410 11704 10416 11716
rect 10468 11744 10474 11756
rect 10689 11747 10747 11753
rect 10689 11744 10701 11747
rect 10468 11716 10701 11744
rect 10468 11704 10474 11716
rect 10689 11713 10701 11716
rect 10735 11713 10747 11747
rect 10689 11707 10747 11713
rect 14182 11704 14188 11756
rect 14240 11744 14246 11756
rect 14553 11747 14611 11753
rect 14553 11744 14565 11747
rect 14240 11716 14565 11744
rect 14240 11704 14246 11716
rect 14553 11713 14565 11716
rect 14599 11713 14611 11747
rect 14553 11707 14611 11713
rect 1443 11648 2084 11676
rect 10505 11679 10563 11685
rect 1443 11645 1455 11648
rect 1397 11639 1455 11645
rect 10505 11645 10517 11679
rect 10551 11676 10563 11679
rect 10778 11676 10784 11688
rect 10551 11648 10784 11676
rect 10551 11645 10563 11648
rect 10505 11639 10563 11645
rect 10778 11636 10784 11648
rect 10836 11636 10842 11688
rect 13814 11636 13820 11688
rect 13872 11676 13878 11688
rect 14274 11676 14280 11688
rect 13872 11648 14280 11676
rect 13872 11636 13878 11648
rect 14274 11636 14280 11648
rect 14332 11676 14338 11688
rect 15948 11685 15976 11784
rect 16666 11772 16672 11784
rect 16724 11772 16730 11824
rect 19610 11812 19616 11824
rect 19571 11784 19616 11812
rect 19610 11772 19616 11784
rect 19668 11772 19674 11824
rect 16114 11744 16120 11756
rect 16075 11716 16120 11744
rect 16114 11704 16120 11716
rect 16172 11704 16178 11756
rect 17773 11747 17831 11753
rect 17773 11713 17785 11747
rect 17819 11744 17831 11747
rect 19150 11744 19156 11756
rect 17819 11716 19156 11744
rect 17819 11713 17831 11716
rect 17773 11707 17831 11713
rect 19150 11704 19156 11716
rect 19208 11744 19214 11756
rect 19628 11744 19656 11772
rect 19208 11716 19656 11744
rect 20916 11744 20944 11843
rect 21266 11840 21272 11892
rect 21324 11880 21330 11892
rect 21453 11883 21511 11889
rect 21453 11880 21465 11883
rect 21324 11852 21465 11880
rect 21324 11840 21330 11852
rect 21453 11849 21465 11852
rect 21499 11849 21511 11883
rect 24118 11880 24124 11892
rect 24079 11852 24124 11880
rect 21453 11843 21511 11849
rect 24118 11840 24124 11852
rect 24176 11840 24182 11892
rect 25038 11840 25044 11892
rect 25096 11880 25102 11892
rect 25317 11883 25375 11889
rect 25317 11880 25329 11883
rect 25096 11852 25329 11880
rect 25096 11840 25102 11852
rect 25317 11849 25329 11852
rect 25363 11849 25375 11883
rect 25317 11843 25375 11849
rect 26605 11883 26663 11889
rect 26605 11849 26617 11883
rect 26651 11880 26663 11883
rect 26878 11880 26884 11892
rect 26651 11852 26884 11880
rect 26651 11849 26663 11852
rect 26605 11843 26663 11849
rect 26878 11840 26884 11852
rect 26936 11840 26942 11892
rect 24857 11815 24915 11821
rect 24857 11781 24869 11815
rect 24903 11812 24915 11815
rect 25222 11812 25228 11824
rect 24903 11784 25228 11812
rect 24903 11781 24915 11784
rect 24857 11775 24915 11781
rect 25222 11772 25228 11784
rect 25280 11812 25286 11824
rect 25280 11784 25820 11812
rect 25280 11772 25286 11784
rect 21913 11747 21971 11753
rect 21913 11744 21925 11747
rect 20916 11716 21925 11744
rect 19208 11704 19214 11716
rect 21913 11713 21925 11716
rect 21959 11713 21971 11747
rect 22094 11744 22100 11756
rect 22007 11716 22100 11744
rect 21913 11707 21971 11713
rect 22094 11704 22100 11716
rect 22152 11744 22158 11756
rect 22281 11747 22339 11753
rect 22281 11744 22293 11747
rect 22152 11716 22293 11744
rect 22152 11704 22158 11716
rect 22281 11713 22293 11716
rect 22327 11713 22339 11747
rect 25130 11744 25136 11756
rect 25091 11716 25136 11744
rect 22281 11707 22339 11713
rect 25130 11704 25136 11716
rect 25188 11744 25194 11756
rect 25792 11753 25820 11784
rect 25777 11747 25835 11753
rect 25188 11716 25728 11744
rect 25188 11704 25194 11716
rect 25700 11688 25728 11716
rect 25777 11713 25789 11747
rect 25823 11713 25835 11747
rect 25777 11707 25835 11713
rect 25869 11747 25927 11753
rect 25869 11713 25881 11747
rect 25915 11744 25927 11747
rect 27430 11744 27436 11756
rect 25915 11716 27436 11744
rect 25915 11713 25927 11716
rect 25869 11707 25927 11713
rect 14461 11679 14519 11685
rect 14461 11676 14473 11679
rect 14332 11648 14473 11676
rect 14332 11636 14338 11648
rect 14461 11645 14473 11648
rect 14507 11645 14519 11679
rect 14461 11639 14519 11645
rect 15933 11679 15991 11685
rect 15933 11645 15945 11679
rect 15979 11645 15991 11679
rect 25682 11676 25688 11688
rect 25595 11648 25688 11676
rect 15933 11639 15991 11645
rect 25682 11636 25688 11648
rect 25740 11636 25746 11688
rect 9306 11568 9312 11620
rect 9364 11608 9370 11620
rect 9401 11611 9459 11617
rect 9401 11608 9413 11611
rect 9364 11580 9413 11608
rect 9364 11568 9370 11580
rect 9401 11577 9413 11580
rect 9447 11608 9459 11611
rect 9447 11580 10640 11608
rect 9447 11577 9459 11580
rect 9401 11571 9459 11577
rect 1578 11540 1584 11552
rect 1539 11512 1584 11540
rect 1578 11500 1584 11512
rect 1636 11500 1642 11552
rect 10134 11540 10140 11552
rect 10095 11512 10140 11540
rect 10134 11500 10140 11512
rect 10192 11500 10198 11552
rect 10612 11549 10640 11580
rect 13906 11568 13912 11620
rect 13964 11608 13970 11620
rect 14366 11608 14372 11620
rect 13964 11580 14372 11608
rect 13964 11568 13970 11580
rect 14366 11568 14372 11580
rect 14424 11568 14430 11620
rect 15286 11568 15292 11620
rect 15344 11608 15350 11620
rect 16025 11611 16083 11617
rect 16025 11608 16037 11611
rect 15344 11580 16037 11608
rect 15344 11568 15350 11580
rect 16025 11577 16037 11580
rect 16071 11608 16083 11611
rect 16390 11608 16396 11620
rect 16071 11580 16396 11608
rect 16071 11577 16083 11580
rect 16025 11571 16083 11577
rect 16390 11568 16396 11580
rect 16448 11568 16454 11620
rect 18969 11611 19027 11617
rect 18969 11577 18981 11611
rect 19015 11608 19027 11611
rect 19058 11608 19064 11620
rect 19015 11580 19064 11608
rect 19015 11577 19027 11580
rect 18969 11571 19027 11577
rect 19058 11568 19064 11580
rect 19116 11608 19122 11620
rect 19889 11611 19947 11617
rect 19889 11608 19901 11611
rect 19116 11580 19901 11608
rect 19116 11568 19122 11580
rect 19889 11577 19901 11580
rect 19935 11577 19947 11611
rect 19889 11571 19947 11577
rect 20625 11611 20683 11617
rect 20625 11577 20637 11611
rect 20671 11608 20683 11611
rect 21821 11611 21879 11617
rect 21821 11608 21833 11611
rect 20671 11580 21833 11608
rect 20671 11577 20683 11580
rect 20625 11571 20683 11577
rect 21821 11577 21833 11580
rect 21867 11608 21879 11611
rect 23014 11608 23020 11620
rect 21867 11580 23020 11608
rect 21867 11577 21879 11580
rect 21821 11571 21879 11577
rect 23014 11568 23020 11580
rect 23072 11568 23078 11620
rect 24489 11611 24547 11617
rect 24489 11577 24501 11611
rect 24535 11608 24547 11611
rect 25884 11608 25912 11707
rect 27430 11704 27436 11716
rect 27488 11704 27494 11756
rect 27062 11636 27068 11688
rect 27120 11676 27126 11688
rect 27341 11679 27399 11685
rect 27341 11676 27353 11679
rect 27120 11648 27353 11676
rect 27120 11636 27126 11648
rect 27341 11645 27353 11648
rect 27387 11645 27399 11679
rect 27341 11639 27399 11645
rect 27893 11611 27951 11617
rect 27893 11608 27905 11611
rect 24535 11580 25912 11608
rect 27264 11580 27905 11608
rect 24535 11577 24547 11580
rect 24489 11571 24547 11577
rect 27264 11552 27292 11580
rect 27893 11577 27905 11580
rect 27939 11577 27951 11611
rect 27893 11571 27951 11577
rect 10597 11543 10655 11549
rect 10597 11509 10609 11543
rect 10643 11540 10655 11543
rect 10778 11540 10784 11552
rect 10643 11512 10784 11540
rect 10643 11509 10655 11512
rect 10597 11503 10655 11509
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 11422 11540 11428 11552
rect 11383 11512 11428 11540
rect 11422 11500 11428 11512
rect 11480 11500 11486 11552
rect 12253 11543 12311 11549
rect 12253 11509 12265 11543
rect 12299 11540 12311 11543
rect 12434 11540 12440 11552
rect 12299 11512 12440 11540
rect 12299 11509 12311 11512
rect 12253 11503 12311 11509
rect 12434 11500 12440 11512
rect 12492 11500 12498 11552
rect 13538 11540 13544 11552
rect 13499 11512 13544 11540
rect 13538 11500 13544 11512
rect 13596 11500 13602 11552
rect 13814 11540 13820 11552
rect 13775 11512 13820 11540
rect 13814 11500 13820 11512
rect 13872 11500 13878 11552
rect 13998 11540 14004 11552
rect 13959 11512 14004 11540
rect 13998 11500 14004 11512
rect 14056 11500 14062 11552
rect 15378 11500 15384 11552
rect 15436 11540 15442 11552
rect 15565 11543 15623 11549
rect 15565 11540 15577 11543
rect 15436 11512 15577 11540
rect 15436 11500 15442 11512
rect 15565 11509 15577 11512
rect 15611 11509 15623 11543
rect 18414 11540 18420 11552
rect 18375 11512 18420 11540
rect 15565 11503 15623 11509
rect 18414 11500 18420 11512
rect 18472 11500 18478 11552
rect 18506 11500 18512 11552
rect 18564 11540 18570 11552
rect 18877 11543 18935 11549
rect 18877 11540 18889 11543
rect 18564 11512 18889 11540
rect 18564 11500 18570 11512
rect 18877 11509 18889 11512
rect 18923 11509 18935 11543
rect 18877 11503 18935 11509
rect 20806 11500 20812 11552
rect 20864 11540 20870 11552
rect 21269 11543 21327 11549
rect 21269 11540 21281 11543
rect 20864 11512 21281 11540
rect 20864 11500 20870 11512
rect 21269 11509 21281 11512
rect 21315 11540 21327 11543
rect 21634 11540 21640 11552
rect 21315 11512 21640 11540
rect 21315 11509 21327 11512
rect 21269 11503 21327 11509
rect 21634 11500 21640 11512
rect 21692 11500 21698 11552
rect 22281 11543 22339 11549
rect 22281 11509 22293 11543
rect 22327 11540 22339 11543
rect 22557 11543 22615 11549
rect 22557 11540 22569 11543
rect 22327 11512 22569 11540
rect 22327 11509 22339 11512
rect 22281 11503 22339 11509
rect 22557 11509 22569 11512
rect 22603 11540 22615 11543
rect 22922 11540 22928 11552
rect 22603 11512 22928 11540
rect 22603 11509 22615 11512
rect 22557 11503 22615 11509
rect 22922 11500 22928 11512
rect 22980 11500 22986 11552
rect 26234 11500 26240 11552
rect 26292 11540 26298 11552
rect 26881 11543 26939 11549
rect 26881 11540 26893 11543
rect 26292 11512 26893 11540
rect 26292 11500 26298 11512
rect 26881 11509 26893 11512
rect 26927 11509 26939 11543
rect 27246 11540 27252 11552
rect 27207 11512 27252 11540
rect 26881 11503 26939 11509
rect 27246 11500 27252 11512
rect 27304 11500 27310 11552
rect 1104 11450 28888 11472
rect 1104 11398 10982 11450
rect 11034 11398 11046 11450
rect 11098 11398 11110 11450
rect 11162 11398 11174 11450
rect 11226 11398 20982 11450
rect 21034 11398 21046 11450
rect 21098 11398 21110 11450
rect 21162 11398 21174 11450
rect 21226 11398 28888 11450
rect 1104 11376 28888 11398
rect 2038 11336 2044 11348
rect 1999 11308 2044 11336
rect 2038 11296 2044 11308
rect 2096 11296 2102 11348
rect 2222 11296 2228 11348
rect 2280 11336 2286 11348
rect 2317 11339 2375 11345
rect 2317 11336 2329 11339
rect 2280 11308 2329 11336
rect 2280 11296 2286 11308
rect 2317 11305 2329 11308
rect 2363 11305 2375 11339
rect 2682 11336 2688 11348
rect 2643 11308 2688 11336
rect 2317 11299 2375 11305
rect 2332 11268 2360 11299
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 6546 11336 6552 11348
rect 6507 11308 6552 11336
rect 6546 11296 6552 11308
rect 6604 11296 6610 11348
rect 9214 11296 9220 11348
rect 9272 11336 9278 11348
rect 9493 11339 9551 11345
rect 9493 11336 9505 11339
rect 9272 11308 9505 11336
rect 9272 11296 9278 11308
rect 9493 11305 9505 11308
rect 9539 11336 9551 11339
rect 10226 11336 10232 11348
rect 9539 11308 10232 11336
rect 9539 11305 9551 11308
rect 9493 11299 9551 11305
rect 10226 11296 10232 11308
rect 10284 11296 10290 11348
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 14550 11336 14556 11348
rect 12492 11308 12537 11336
rect 14511 11308 14556 11336
rect 12492 11296 12498 11308
rect 14550 11296 14556 11308
rect 14608 11296 14614 11348
rect 17034 11336 17040 11348
rect 16995 11308 17040 11336
rect 17034 11296 17040 11308
rect 17092 11296 17098 11348
rect 18966 11336 18972 11348
rect 18927 11308 18972 11336
rect 18966 11296 18972 11308
rect 19024 11296 19030 11348
rect 21545 11339 21603 11345
rect 21545 11305 21557 11339
rect 21591 11336 21603 11339
rect 21818 11336 21824 11348
rect 21591 11308 21824 11336
rect 21591 11305 21603 11308
rect 21545 11299 21603 11305
rect 21818 11296 21824 11308
rect 21876 11296 21882 11348
rect 22922 11296 22928 11348
rect 22980 11336 22986 11348
rect 23293 11339 23351 11345
rect 23293 11336 23305 11339
rect 22980 11308 23305 11336
rect 22980 11296 22986 11308
rect 23293 11305 23305 11308
rect 23339 11305 23351 11339
rect 24578 11336 24584 11348
rect 24539 11308 24584 11336
rect 23293 11299 23351 11305
rect 24578 11296 24584 11308
rect 24636 11296 24642 11348
rect 24946 11336 24952 11348
rect 24907 11308 24952 11336
rect 24946 11296 24952 11308
rect 25004 11296 25010 11348
rect 25409 11339 25467 11345
rect 25409 11305 25421 11339
rect 25455 11336 25467 11339
rect 27246 11336 27252 11348
rect 25455 11308 27252 11336
rect 25455 11305 25467 11308
rect 25409 11299 25467 11305
rect 27246 11296 27252 11308
rect 27304 11296 27310 11348
rect 27430 11336 27436 11348
rect 27391 11308 27436 11336
rect 27430 11296 27436 11308
rect 27488 11296 27494 11348
rect 2332 11240 3188 11268
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 1486 11200 1492 11212
rect 1443 11172 1492 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 1486 11160 1492 11172
rect 1544 11160 1550 11212
rect 2501 11203 2559 11209
rect 2501 11169 2513 11203
rect 2547 11200 2559 11203
rect 2682 11200 2688 11212
rect 2547 11172 2688 11200
rect 2547 11169 2559 11172
rect 2501 11163 2559 11169
rect 2682 11160 2688 11172
rect 2740 11160 2746 11212
rect 3160 11141 3188 11240
rect 7374 11228 7380 11280
rect 7432 11268 7438 11280
rect 7622 11271 7680 11277
rect 7622 11268 7634 11271
rect 7432 11240 7634 11268
rect 7432 11228 7438 11240
rect 7622 11237 7634 11240
rect 7668 11237 7680 11271
rect 7622 11231 7680 11237
rect 9674 11228 9680 11280
rect 9732 11268 9738 11280
rect 9861 11271 9919 11277
rect 9861 11268 9873 11271
rect 9732 11240 9873 11268
rect 9732 11228 9738 11240
rect 9861 11237 9873 11240
rect 9907 11237 9919 11271
rect 9861 11231 9919 11237
rect 15841 11271 15899 11277
rect 15841 11237 15853 11271
rect 15887 11268 15899 11271
rect 15930 11268 15936 11280
rect 15887 11240 15936 11268
rect 15887 11237 15899 11240
rect 15841 11231 15899 11237
rect 15930 11228 15936 11240
rect 15988 11228 15994 11280
rect 22094 11228 22100 11280
rect 22152 11277 22158 11280
rect 22152 11271 22216 11277
rect 22152 11237 22170 11271
rect 22204 11237 22216 11271
rect 22152 11231 22216 11237
rect 22152 11228 22158 11231
rect 26418 11228 26424 11280
rect 26476 11268 26482 11280
rect 27062 11268 27068 11280
rect 26476 11240 27068 11268
rect 26476 11228 26482 11240
rect 27062 11228 27068 11240
rect 27120 11228 27126 11280
rect 5258 11160 5264 11212
rect 5316 11200 5322 11212
rect 5425 11203 5483 11209
rect 5425 11200 5437 11203
rect 5316 11172 5437 11200
rect 5316 11160 5322 11172
rect 5425 11169 5437 11172
rect 5471 11169 5483 11203
rect 5425 11163 5483 11169
rect 10413 11203 10471 11209
rect 10413 11169 10425 11203
rect 10459 11200 10471 11203
rect 10962 11200 10968 11212
rect 10459 11172 10968 11200
rect 10459 11169 10471 11172
rect 10413 11163 10471 11169
rect 10962 11160 10968 11172
rect 11020 11160 11026 11212
rect 12894 11160 12900 11212
rect 12952 11200 12958 11212
rect 13061 11203 13119 11209
rect 13061 11200 13073 11203
rect 12952 11172 13073 11200
rect 12952 11160 12958 11172
rect 13061 11169 13073 11172
rect 13107 11200 13119 11203
rect 13814 11200 13820 11212
rect 13107 11172 13820 11200
rect 13107 11169 13119 11172
rect 13061 11163 13119 11169
rect 13814 11160 13820 11172
rect 13872 11200 13878 11212
rect 14918 11200 14924 11212
rect 13872 11172 14924 11200
rect 13872 11160 13878 11172
rect 14918 11160 14924 11172
rect 14976 11200 14982 11212
rect 15013 11203 15071 11209
rect 15013 11200 15025 11203
rect 14976 11172 15025 11200
rect 14976 11160 14982 11172
rect 15013 11169 15025 11172
rect 15059 11200 15071 11203
rect 15470 11200 15476 11212
rect 15059 11172 15476 11200
rect 15059 11169 15071 11172
rect 15013 11163 15071 11169
rect 15470 11160 15476 11172
rect 15528 11160 15534 11212
rect 15746 11200 15752 11212
rect 15707 11172 15752 11200
rect 15746 11160 15752 11172
rect 15804 11160 15810 11212
rect 19337 11203 19395 11209
rect 19337 11169 19349 11203
rect 19383 11200 19395 11203
rect 20070 11200 20076 11212
rect 19383 11172 20076 11200
rect 19383 11169 19395 11172
rect 19337 11163 19395 11169
rect 20070 11160 20076 11172
rect 20128 11200 20134 11212
rect 20254 11200 20260 11212
rect 20128 11172 20260 11200
rect 20128 11160 20134 11172
rect 20254 11160 20260 11172
rect 20312 11160 20318 11212
rect 25682 11160 25688 11212
rect 25740 11200 25746 11212
rect 26513 11203 26571 11209
rect 26513 11200 26525 11203
rect 25740 11172 26525 11200
rect 25740 11160 25746 11172
rect 26513 11169 26525 11172
rect 26559 11200 26571 11203
rect 27246 11200 27252 11212
rect 26559 11172 27252 11200
rect 26559 11169 26571 11172
rect 26513 11163 26571 11169
rect 27246 11160 27252 11172
rect 27304 11160 27310 11212
rect 3145 11135 3203 11141
rect 3145 11101 3157 11135
rect 3191 11132 3203 11135
rect 5166 11132 5172 11144
rect 3191 11104 5172 11132
rect 3191 11101 3203 11104
rect 3145 11095 3203 11101
rect 5166 11092 5172 11104
rect 5224 11092 5230 11144
rect 7377 11135 7435 11141
rect 7377 11101 7389 11135
rect 7423 11101 7435 11135
rect 7377 11095 7435 11101
rect 1581 11067 1639 11073
rect 1581 11033 1593 11067
rect 1627 11064 1639 11067
rect 1762 11064 1768 11076
rect 1627 11036 1768 11064
rect 1627 11033 1639 11036
rect 1581 11027 1639 11033
rect 1762 11024 1768 11036
rect 1820 11024 1826 11076
rect 6917 10999 6975 11005
rect 6917 10965 6929 10999
rect 6963 10996 6975 10999
rect 7282 10996 7288 11008
rect 6963 10968 7288 10996
rect 6963 10965 6975 10968
rect 6917 10959 6975 10965
rect 7282 10956 7288 10968
rect 7340 10956 7346 11008
rect 7392 10996 7420 11095
rect 9858 11092 9864 11144
rect 9916 11132 9922 11144
rect 10226 11132 10232 11144
rect 9916 11104 10232 11132
rect 9916 11092 9922 11104
rect 10226 11092 10232 11104
rect 10284 11092 10290 11144
rect 10502 11132 10508 11144
rect 10463 11104 10508 11132
rect 10502 11092 10508 11104
rect 10560 11092 10566 11144
rect 10594 11092 10600 11144
rect 10652 11132 10658 11144
rect 12802 11132 12808 11144
rect 10652 11104 10697 11132
rect 12763 11104 12808 11132
rect 10652 11092 10658 11104
rect 12802 11092 12808 11104
rect 12860 11092 12866 11144
rect 15488 11132 15516 11160
rect 15933 11135 15991 11141
rect 15933 11132 15945 11135
rect 15488 11104 15945 11132
rect 15933 11101 15945 11104
rect 15979 11132 15991 11135
rect 16114 11132 16120 11144
rect 15979 11104 16120 11132
rect 15979 11101 15991 11104
rect 15933 11095 15991 11101
rect 16114 11092 16120 11104
rect 16172 11132 16178 11144
rect 16393 11135 16451 11141
rect 16393 11132 16405 11135
rect 16172 11104 16405 11132
rect 16172 11092 16178 11104
rect 16393 11101 16405 11104
rect 16439 11101 16451 11135
rect 16393 11095 16451 11101
rect 19429 11135 19487 11141
rect 19429 11101 19441 11135
rect 19475 11132 19487 11135
rect 19518 11132 19524 11144
rect 19475 11104 19524 11132
rect 19475 11101 19487 11104
rect 19429 11095 19487 11101
rect 19518 11092 19524 11104
rect 19576 11092 19582 11144
rect 19613 11135 19671 11141
rect 19613 11101 19625 11135
rect 19659 11101 19671 11135
rect 21910 11132 21916 11144
rect 21871 11104 21916 11132
rect 19613 11095 19671 11101
rect 10045 11067 10103 11073
rect 10045 11064 10057 11067
rect 9600 11036 10057 11064
rect 9600 11008 9628 11036
rect 10045 11033 10057 11036
rect 10091 11033 10103 11067
rect 15381 11067 15439 11073
rect 15381 11064 15393 11067
rect 10045 11027 10103 11033
rect 15120 11036 15393 11064
rect 15120 11008 15148 11036
rect 15381 11033 15393 11036
rect 15427 11033 15439 11067
rect 15381 11027 15439 11033
rect 18877 11067 18935 11073
rect 18877 11033 18889 11067
rect 18923 11064 18935 11067
rect 18923 11036 19380 11064
rect 18923 11033 18935 11036
rect 18877 11027 18935 11033
rect 7742 10996 7748 11008
rect 7392 10968 7748 10996
rect 7742 10956 7748 10968
rect 7800 10956 7806 11008
rect 8386 10956 8392 11008
rect 8444 10996 8450 11008
rect 8757 10999 8815 11005
rect 8757 10996 8769 10999
rect 8444 10968 8769 10996
rect 8444 10956 8450 10968
rect 8757 10965 8769 10968
rect 8803 10965 8815 10999
rect 8757 10959 8815 10965
rect 9582 10956 9588 11008
rect 9640 10956 9646 11008
rect 14182 10996 14188 11008
rect 14143 10968 14188 10996
rect 14182 10956 14188 10968
rect 14240 10956 14246 11008
rect 15102 10956 15108 11008
rect 15160 10956 15166 11008
rect 18506 10996 18512 11008
rect 18467 10968 18512 10996
rect 18506 10956 18512 10968
rect 18564 10956 18570 11008
rect 19352 10996 19380 11036
rect 19628 11008 19656 11095
rect 21910 11092 21916 11104
rect 21968 11092 21974 11144
rect 26694 11064 26700 11076
rect 26655 11036 26700 11064
rect 26694 11024 26700 11036
rect 26752 11024 26758 11076
rect 19610 10996 19616 11008
rect 19352 10968 19616 10996
rect 19610 10956 19616 10968
rect 19668 10956 19674 11008
rect 1104 10906 28888 10928
rect 1104 10854 5982 10906
rect 6034 10854 6046 10906
rect 6098 10854 6110 10906
rect 6162 10854 6174 10906
rect 6226 10854 15982 10906
rect 16034 10854 16046 10906
rect 16098 10854 16110 10906
rect 16162 10854 16174 10906
rect 16226 10854 25982 10906
rect 26034 10854 26046 10906
rect 26098 10854 26110 10906
rect 26162 10854 26174 10906
rect 26226 10854 28888 10906
rect 1104 10832 28888 10854
rect 1486 10752 1492 10804
rect 1544 10792 1550 10804
rect 1581 10795 1639 10801
rect 1581 10792 1593 10795
rect 1544 10764 1593 10792
rect 1544 10752 1550 10764
rect 1581 10761 1593 10764
rect 1627 10761 1639 10795
rect 1581 10755 1639 10761
rect 2317 10795 2375 10801
rect 2317 10761 2329 10795
rect 2363 10792 2375 10795
rect 2682 10792 2688 10804
rect 2363 10764 2688 10792
rect 2363 10761 2375 10764
rect 2317 10755 2375 10761
rect 2682 10752 2688 10764
rect 2740 10752 2746 10804
rect 5258 10792 5264 10804
rect 5219 10764 5264 10792
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 6546 10792 6552 10804
rect 6507 10764 6552 10792
rect 6546 10752 6552 10764
rect 6604 10752 6610 10804
rect 7742 10792 7748 10804
rect 6656 10764 7748 10792
rect 5166 10684 5172 10736
rect 5224 10724 5230 10736
rect 5537 10727 5595 10733
rect 5537 10724 5549 10727
rect 5224 10696 5549 10724
rect 5224 10684 5230 10696
rect 5537 10693 5549 10696
rect 5583 10724 5595 10727
rect 5810 10724 5816 10736
rect 5583 10696 5816 10724
rect 5583 10693 5595 10696
rect 5537 10687 5595 10693
rect 5810 10684 5816 10696
rect 5868 10724 5874 10736
rect 6656 10724 6684 10764
rect 7742 10752 7748 10764
rect 7800 10752 7806 10804
rect 10502 10752 10508 10804
rect 10560 10792 10566 10804
rect 11057 10795 11115 10801
rect 11057 10792 11069 10795
rect 10560 10764 11069 10792
rect 10560 10752 10566 10764
rect 11057 10761 11069 10764
rect 11103 10761 11115 10795
rect 12894 10792 12900 10804
rect 12855 10764 12900 10792
rect 11057 10755 11115 10761
rect 12894 10752 12900 10764
rect 12952 10752 12958 10804
rect 13722 10792 13728 10804
rect 13683 10764 13728 10792
rect 13722 10752 13728 10764
rect 13780 10752 13786 10804
rect 14090 10792 14096 10804
rect 14051 10764 14096 10792
rect 14090 10752 14096 10764
rect 14148 10752 14154 10804
rect 15746 10752 15752 10804
rect 15804 10792 15810 10804
rect 15933 10795 15991 10801
rect 15933 10792 15945 10795
rect 15804 10764 15945 10792
rect 15804 10752 15810 10764
rect 15933 10761 15945 10764
rect 15979 10792 15991 10795
rect 18969 10795 19027 10801
rect 15979 10764 16160 10792
rect 15979 10761 15991 10764
rect 15933 10755 15991 10761
rect 8481 10727 8539 10733
rect 8481 10724 8493 10727
rect 5868 10696 6684 10724
rect 7300 10696 8493 10724
rect 5868 10684 5874 10696
rect 7300 10668 7328 10696
rect 8481 10693 8493 10696
rect 8527 10693 8539 10727
rect 9858 10724 9864 10736
rect 9819 10696 9864 10724
rect 8481 10687 8539 10693
rect 9858 10684 9864 10696
rect 9916 10724 9922 10736
rect 10318 10724 10324 10736
rect 9916 10696 10324 10724
rect 9916 10684 9922 10696
rect 10318 10684 10324 10696
rect 10376 10684 10382 10736
rect 11793 10727 11851 10733
rect 11793 10724 11805 10727
rect 10520 10696 11805 10724
rect 2222 10616 2228 10668
rect 2280 10656 2286 10668
rect 2409 10659 2467 10665
rect 2409 10656 2421 10659
rect 2280 10628 2421 10656
rect 2280 10616 2286 10628
rect 2409 10625 2421 10628
rect 2455 10625 2467 10659
rect 2409 10619 2467 10625
rect 5626 10616 5632 10668
rect 5684 10656 5690 10668
rect 6638 10656 6644 10668
rect 5684 10628 6644 10656
rect 5684 10616 5690 10628
rect 6638 10616 6644 10628
rect 6696 10616 6702 10668
rect 7282 10656 7288 10668
rect 7243 10628 7288 10656
rect 7282 10616 7288 10628
rect 7340 10616 7346 10668
rect 7377 10659 7435 10665
rect 7377 10625 7389 10659
rect 7423 10625 7435 10659
rect 7377 10619 7435 10625
rect 6546 10548 6552 10600
rect 6604 10588 6610 10600
rect 7392 10588 7420 10619
rect 8386 10616 8392 10668
rect 8444 10656 8450 10668
rect 9033 10659 9091 10665
rect 9033 10656 9045 10659
rect 8444 10628 9045 10656
rect 8444 10616 8450 10628
rect 9033 10625 9045 10628
rect 9079 10625 9091 10659
rect 9033 10619 9091 10625
rect 9490 10616 9496 10668
rect 9548 10656 9554 10668
rect 9548 10628 9904 10656
rect 9548 10616 9554 10628
rect 9876 10600 9904 10628
rect 10134 10616 10140 10668
rect 10192 10656 10198 10668
rect 10520 10665 10548 10696
rect 11793 10693 11805 10696
rect 11839 10693 11851 10727
rect 11793 10687 11851 10693
rect 15657 10727 15715 10733
rect 15657 10693 15669 10727
rect 15703 10724 15715 10727
rect 15838 10724 15844 10736
rect 15703 10696 15844 10724
rect 15703 10693 15715 10696
rect 15657 10687 15715 10693
rect 15838 10684 15844 10696
rect 15896 10684 15902 10736
rect 10505 10659 10563 10665
rect 10505 10656 10517 10659
rect 10192 10628 10517 10656
rect 10192 10616 10198 10628
rect 10505 10625 10517 10628
rect 10551 10625 10563 10659
rect 10505 10619 10563 10625
rect 10594 10616 10600 10668
rect 10652 10656 10658 10668
rect 10652 10628 10745 10656
rect 10652 10616 10658 10628
rect 11054 10616 11060 10668
rect 11112 10656 11118 10668
rect 11425 10659 11483 10665
rect 11425 10656 11437 10659
rect 11112 10628 11437 10656
rect 11112 10616 11118 10628
rect 11425 10625 11437 10628
rect 11471 10625 11483 10659
rect 11425 10619 11483 10625
rect 13357 10659 13415 10665
rect 13357 10625 13369 10659
rect 13403 10656 13415 10659
rect 13722 10656 13728 10668
rect 13403 10628 13728 10656
rect 13403 10625 13415 10628
rect 13357 10619 13415 10625
rect 13722 10616 13728 10628
rect 13780 10616 13786 10668
rect 14182 10616 14188 10668
rect 14240 10656 14246 10668
rect 16132 10665 16160 10764
rect 18969 10761 18981 10795
rect 19015 10792 19027 10795
rect 19058 10792 19064 10804
rect 19015 10764 19064 10792
rect 19015 10761 19027 10764
rect 18969 10755 19027 10761
rect 19058 10752 19064 10764
rect 19116 10752 19122 10804
rect 20809 10795 20867 10801
rect 20809 10761 20821 10795
rect 20855 10792 20867 10795
rect 22002 10792 22008 10804
rect 20855 10764 22008 10792
rect 20855 10761 20867 10764
rect 20809 10755 20867 10761
rect 22002 10752 22008 10764
rect 22060 10752 22066 10804
rect 27246 10752 27252 10804
rect 27304 10792 27310 10804
rect 27341 10795 27399 10801
rect 27341 10792 27353 10795
rect 27304 10764 27353 10792
rect 27304 10752 27310 10764
rect 27341 10761 27353 10764
rect 27387 10761 27399 10795
rect 27341 10755 27399 10761
rect 15105 10659 15163 10665
rect 15105 10656 15117 10659
rect 14240 10628 15117 10656
rect 14240 10616 14246 10628
rect 15105 10625 15117 10628
rect 15151 10625 15163 10659
rect 15105 10619 15163 10625
rect 16117 10659 16175 10665
rect 16117 10625 16129 10659
rect 16163 10625 16175 10659
rect 19610 10656 19616 10668
rect 19571 10628 19616 10656
rect 16117 10619 16175 10625
rect 19610 10616 19616 10628
rect 19668 10616 19674 10668
rect 6604 10560 7420 10588
rect 6604 10548 6610 10560
rect 8570 10548 8576 10600
rect 8628 10588 8634 10600
rect 8941 10591 8999 10597
rect 8941 10588 8953 10591
rect 8628 10560 8953 10588
rect 8628 10548 8634 10560
rect 8941 10557 8953 10560
rect 8987 10588 8999 10591
rect 9582 10588 9588 10600
rect 8987 10560 9588 10588
rect 8987 10557 8999 10560
rect 8941 10551 8999 10557
rect 9582 10548 9588 10560
rect 9640 10548 9646 10600
rect 9858 10548 9864 10600
rect 9916 10548 9922 10600
rect 10042 10548 10048 10600
rect 10100 10588 10106 10600
rect 10612 10588 10640 10616
rect 11330 10588 11336 10600
rect 10100 10560 11336 10588
rect 10100 10548 10106 10560
rect 11330 10548 11336 10560
rect 11388 10548 11394 10600
rect 14734 10548 14740 10600
rect 14792 10588 14798 10600
rect 15013 10591 15071 10597
rect 15013 10588 15025 10591
rect 14792 10560 15025 10588
rect 14792 10548 14798 10560
rect 15013 10557 15025 10560
rect 15059 10588 15071 10591
rect 15378 10588 15384 10600
rect 15059 10560 15384 10588
rect 15059 10557 15071 10560
rect 15013 10551 15071 10557
rect 15378 10548 15384 10560
rect 15436 10548 15442 10600
rect 19334 10588 19340 10600
rect 19295 10560 19340 10588
rect 19334 10548 19340 10560
rect 19392 10588 19398 10600
rect 19981 10591 20039 10597
rect 19981 10588 19993 10591
rect 19392 10560 19993 10588
rect 19392 10548 19398 10560
rect 19981 10557 19993 10560
rect 20027 10557 20039 10591
rect 26418 10588 26424 10600
rect 26379 10560 26424 10588
rect 19981 10551 20039 10557
rect 26418 10548 26424 10560
rect 26476 10588 26482 10600
rect 26973 10591 27031 10597
rect 26973 10588 26985 10591
rect 26476 10560 26985 10588
rect 26476 10548 26482 10560
rect 26973 10557 26985 10560
rect 27019 10557 27031 10591
rect 27522 10588 27528 10600
rect 27483 10560 27528 10588
rect 26973 10551 27031 10557
rect 27522 10548 27528 10560
rect 27580 10588 27586 10600
rect 28077 10591 28135 10597
rect 28077 10588 28089 10591
rect 27580 10560 28089 10588
rect 27580 10548 27586 10560
rect 28077 10557 28089 10560
rect 28123 10557 28135 10591
rect 28077 10551 28135 10557
rect 2676 10523 2734 10529
rect 2676 10489 2688 10523
rect 2722 10520 2734 10523
rect 3050 10520 3056 10532
rect 2722 10492 3056 10520
rect 2722 10489 2734 10492
rect 2676 10483 2734 10489
rect 3050 10480 3056 10492
rect 3108 10480 3114 10532
rect 3878 10480 3884 10532
rect 3936 10520 3942 10532
rect 4798 10520 4804 10532
rect 3936 10492 4804 10520
rect 3936 10480 3942 10492
rect 4798 10480 4804 10492
rect 4856 10480 4862 10532
rect 6273 10523 6331 10529
rect 6273 10489 6285 10523
rect 6319 10520 6331 10523
rect 6362 10520 6368 10532
rect 6319 10492 6368 10520
rect 6319 10489 6331 10492
rect 6273 10483 6331 10489
rect 6362 10480 6368 10492
rect 6420 10520 6426 10532
rect 7193 10523 7251 10529
rect 7193 10520 7205 10523
rect 6420 10492 7205 10520
rect 6420 10480 6426 10492
rect 7193 10489 7205 10492
rect 7239 10489 7251 10523
rect 8846 10520 8852 10532
rect 7193 10483 7251 10489
rect 7852 10492 8708 10520
rect 8759 10492 8852 10520
rect 3786 10452 3792 10464
rect 3747 10424 3792 10452
rect 3786 10412 3792 10424
rect 3844 10412 3850 10464
rect 6638 10412 6644 10464
rect 6696 10452 6702 10464
rect 6825 10455 6883 10461
rect 6825 10452 6837 10455
rect 6696 10424 6837 10452
rect 6696 10412 6702 10424
rect 6825 10421 6837 10424
rect 6871 10421 6883 10455
rect 6825 10415 6883 10421
rect 7374 10412 7380 10464
rect 7432 10452 7438 10464
rect 7852 10461 7880 10492
rect 7837 10455 7895 10461
rect 7837 10452 7849 10455
rect 7432 10424 7849 10452
rect 7432 10412 7438 10424
rect 7837 10421 7849 10424
rect 7883 10421 7895 10455
rect 8386 10452 8392 10464
rect 8347 10424 8392 10452
rect 7837 10415 7895 10421
rect 8386 10412 8392 10424
rect 8444 10412 8450 10464
rect 8680 10452 8708 10492
rect 8846 10480 8852 10492
rect 8904 10520 8910 10532
rect 8904 10492 10088 10520
rect 8904 10480 8910 10492
rect 9490 10452 9496 10464
rect 8680 10424 9496 10452
rect 9490 10412 9496 10424
rect 9548 10412 9554 10464
rect 10060 10461 10088 10492
rect 10318 10480 10324 10532
rect 10376 10520 10382 10532
rect 10413 10523 10471 10529
rect 10413 10520 10425 10523
rect 10376 10492 10425 10520
rect 10376 10480 10382 10492
rect 10413 10489 10425 10492
rect 10459 10489 10471 10523
rect 10413 10483 10471 10489
rect 14921 10523 14979 10529
rect 14921 10489 14933 10523
rect 14967 10520 14979 10523
rect 15102 10520 15108 10532
rect 14967 10492 15108 10520
rect 14967 10489 14979 10492
rect 14921 10483 14979 10489
rect 15102 10480 15108 10492
rect 15160 10480 15166 10532
rect 18414 10520 18420 10532
rect 18375 10492 18420 10520
rect 18414 10480 18420 10492
rect 18472 10480 18478 10532
rect 19429 10523 19487 10529
rect 19429 10489 19441 10523
rect 19475 10520 19487 10523
rect 20438 10520 20444 10532
rect 19475 10492 20444 10520
rect 19475 10489 19487 10492
rect 19429 10483 19487 10489
rect 10045 10455 10103 10461
rect 10045 10421 10057 10455
rect 10091 10421 10103 10455
rect 10045 10415 10103 10421
rect 13814 10412 13820 10464
rect 13872 10452 13878 10464
rect 14182 10452 14188 10464
rect 13872 10424 14188 10452
rect 13872 10412 13878 10424
rect 14182 10412 14188 10424
rect 14240 10452 14246 10464
rect 14369 10455 14427 10461
rect 14369 10452 14381 10455
rect 14240 10424 14381 10452
rect 14240 10412 14246 10424
rect 14369 10421 14381 10424
rect 14415 10421 14427 10455
rect 14550 10452 14556 10464
rect 14511 10424 14556 10452
rect 14369 10415 14427 10421
rect 14550 10412 14556 10424
rect 14608 10412 14614 10464
rect 18874 10452 18880 10464
rect 18835 10424 18880 10452
rect 18874 10412 18880 10424
rect 18932 10452 18938 10464
rect 19444 10452 19472 10483
rect 20438 10480 20444 10492
rect 20496 10480 20502 10532
rect 21910 10480 21916 10532
rect 21968 10520 21974 10532
rect 22094 10520 22100 10532
rect 21968 10492 22100 10520
rect 21968 10480 21974 10492
rect 22094 10480 22100 10492
rect 22152 10520 22158 10532
rect 22281 10523 22339 10529
rect 22281 10520 22293 10523
rect 22152 10492 22293 10520
rect 22152 10480 22158 10492
rect 22281 10489 22293 10492
rect 22327 10489 22339 10523
rect 22281 10483 22339 10489
rect 18932 10424 19472 10452
rect 18932 10412 18938 10424
rect 20254 10412 20260 10464
rect 20312 10452 20318 10464
rect 20349 10455 20407 10461
rect 20349 10452 20361 10455
rect 20312 10424 20361 10452
rect 20312 10412 20318 10424
rect 20349 10421 20361 10424
rect 20395 10421 20407 10455
rect 25222 10452 25228 10464
rect 25183 10424 25228 10452
rect 20349 10415 20407 10421
rect 25222 10412 25228 10424
rect 25280 10412 25286 10464
rect 26602 10452 26608 10464
rect 26563 10424 26608 10452
rect 26602 10412 26608 10424
rect 26660 10412 26666 10464
rect 27706 10452 27712 10464
rect 27667 10424 27712 10452
rect 27706 10412 27712 10424
rect 27764 10412 27770 10464
rect 1104 10362 28888 10384
rect 1104 10310 10982 10362
rect 11034 10310 11046 10362
rect 11098 10310 11110 10362
rect 11162 10310 11174 10362
rect 11226 10310 20982 10362
rect 21034 10310 21046 10362
rect 21098 10310 21110 10362
rect 21162 10310 21174 10362
rect 21226 10310 28888 10362
rect 1104 10288 28888 10310
rect 3050 10248 3056 10260
rect 3011 10220 3056 10248
rect 3050 10208 3056 10220
rect 3108 10208 3114 10260
rect 6362 10248 6368 10260
rect 6323 10220 6368 10248
rect 6362 10208 6368 10220
rect 6420 10208 6426 10260
rect 7742 10248 7748 10260
rect 7703 10220 7748 10248
rect 7742 10208 7748 10220
rect 7800 10208 7806 10260
rect 8570 10248 8576 10260
rect 8531 10220 8576 10248
rect 8570 10208 8576 10220
rect 8628 10208 8634 10260
rect 8846 10248 8852 10260
rect 8807 10220 8852 10248
rect 8846 10208 8852 10220
rect 8904 10208 8910 10260
rect 9490 10208 9496 10260
rect 9548 10248 9554 10260
rect 10042 10248 10048 10260
rect 9548 10220 10048 10248
rect 9548 10208 9554 10220
rect 10042 10208 10048 10220
rect 10100 10208 10106 10260
rect 10410 10248 10416 10260
rect 10371 10220 10416 10248
rect 10410 10208 10416 10220
rect 10468 10208 10474 10260
rect 10502 10208 10508 10260
rect 10560 10248 10566 10260
rect 10597 10251 10655 10257
rect 10597 10248 10609 10251
rect 10560 10220 10609 10248
rect 10560 10208 10566 10220
rect 10597 10217 10609 10220
rect 10643 10217 10655 10251
rect 10597 10211 10655 10217
rect 10686 10208 10692 10260
rect 10744 10248 10750 10260
rect 11057 10251 11115 10257
rect 11057 10248 11069 10251
rect 10744 10220 11069 10248
rect 10744 10208 10750 10220
rect 11057 10217 11069 10220
rect 11103 10217 11115 10251
rect 11057 10211 11115 10217
rect 14001 10251 14059 10257
rect 14001 10217 14013 10251
rect 14047 10248 14059 10251
rect 14090 10248 14096 10260
rect 14047 10220 14096 10248
rect 14047 10217 14059 10220
rect 14001 10211 14059 10217
rect 14090 10208 14096 10220
rect 14148 10248 14154 10260
rect 14550 10248 14556 10260
rect 14148 10220 14556 10248
rect 14148 10208 14154 10220
rect 14550 10208 14556 10220
rect 14608 10208 14614 10260
rect 14734 10248 14740 10260
rect 14695 10220 14740 10248
rect 14734 10208 14740 10220
rect 14792 10208 14798 10260
rect 15102 10248 15108 10260
rect 15063 10220 15108 10248
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 15470 10248 15476 10260
rect 15431 10220 15476 10248
rect 15470 10208 15476 10220
rect 15528 10208 15534 10260
rect 18506 10208 18512 10260
rect 18564 10248 18570 10260
rect 18969 10251 19027 10257
rect 18969 10248 18981 10251
rect 18564 10220 18981 10248
rect 18564 10208 18570 10220
rect 18969 10217 18981 10220
rect 19015 10217 19027 10251
rect 18969 10211 19027 10217
rect 25317 10251 25375 10257
rect 25317 10217 25329 10251
rect 25363 10248 25375 10251
rect 25498 10248 25504 10260
rect 25363 10220 25504 10248
rect 25363 10217 25375 10220
rect 25317 10211 25375 10217
rect 25498 10208 25504 10220
rect 25556 10208 25562 10260
rect 2222 10140 2228 10192
rect 2280 10180 2286 10192
rect 3510 10180 3516 10192
rect 2280 10152 3516 10180
rect 2280 10140 2286 10152
rect 3510 10140 3516 10152
rect 3568 10140 3574 10192
rect 9858 10140 9864 10192
rect 9916 10180 9922 10192
rect 10965 10183 11023 10189
rect 10965 10180 10977 10183
rect 9916 10152 10977 10180
rect 9916 10140 9922 10152
rect 10965 10149 10977 10152
rect 11011 10180 11023 10183
rect 11514 10180 11520 10192
rect 11011 10152 11520 10180
rect 11011 10149 11023 10152
rect 10965 10143 11023 10149
rect 11514 10140 11520 10152
rect 11572 10140 11578 10192
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10112 1455 10115
rect 1670 10112 1676 10124
rect 1443 10084 1676 10112
rect 1443 10081 1455 10084
rect 1397 10075 1455 10081
rect 1670 10072 1676 10084
rect 1728 10072 1734 10124
rect 2498 10112 2504 10124
rect 2459 10084 2504 10112
rect 2498 10072 2504 10084
rect 2556 10072 2562 10124
rect 6730 10112 6736 10124
rect 6691 10084 6736 10112
rect 6730 10072 6736 10084
rect 6788 10072 6794 10124
rect 8113 10115 8171 10121
rect 8113 10081 8125 10115
rect 8159 10112 8171 10115
rect 8202 10112 8208 10124
rect 8159 10084 8208 10112
rect 8159 10081 8171 10084
rect 8113 10075 8171 10081
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 13722 10072 13728 10124
rect 13780 10112 13786 10124
rect 13998 10112 14004 10124
rect 13780 10084 14004 10112
rect 13780 10072 13786 10084
rect 13998 10072 14004 10084
rect 14056 10112 14062 10124
rect 14093 10115 14151 10121
rect 14093 10112 14105 10115
rect 14056 10084 14105 10112
rect 14056 10072 14062 10084
rect 14093 10081 14105 10084
rect 14139 10081 14151 10115
rect 14093 10075 14151 10081
rect 18690 10072 18696 10124
rect 18748 10112 18754 10124
rect 18877 10115 18935 10121
rect 18877 10112 18889 10115
rect 18748 10084 18889 10112
rect 18748 10072 18754 10084
rect 18877 10081 18889 10084
rect 18923 10081 18935 10115
rect 19334 10112 19340 10124
rect 19295 10084 19340 10112
rect 18877 10075 18935 10081
rect 19334 10072 19340 10084
rect 19392 10112 19398 10124
rect 19702 10112 19708 10124
rect 19392 10084 19708 10112
rect 19392 10072 19398 10084
rect 19702 10072 19708 10084
rect 19760 10072 19766 10124
rect 25222 10112 25228 10124
rect 25183 10084 25228 10112
rect 25222 10072 25228 10084
rect 25280 10072 25286 10124
rect 26510 10112 26516 10124
rect 26471 10084 26516 10112
rect 26510 10072 26516 10084
rect 26568 10072 26574 10124
rect 6822 10044 6828 10056
rect 6783 10016 6828 10044
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 6917 10047 6975 10053
rect 6917 10013 6929 10047
rect 6963 10013 6975 10047
rect 6917 10007 6975 10013
rect 5258 9936 5264 9988
rect 5316 9976 5322 9988
rect 6454 9976 6460 9988
rect 5316 9948 6460 9976
rect 5316 9936 5322 9948
rect 6454 9936 6460 9948
rect 6512 9976 6518 9988
rect 6932 9976 6960 10007
rect 10410 10004 10416 10056
rect 10468 10044 10474 10056
rect 11149 10047 11207 10053
rect 11149 10044 11161 10047
rect 10468 10016 11161 10044
rect 10468 10004 10474 10016
rect 10980 9988 11008 10016
rect 11149 10013 11161 10016
rect 11195 10013 11207 10047
rect 14182 10044 14188 10056
rect 14143 10016 14188 10044
rect 11149 10007 11207 10013
rect 14182 10004 14188 10016
rect 14240 10004 14246 10056
rect 19426 10044 19432 10056
rect 19387 10016 19432 10044
rect 19426 10004 19432 10016
rect 19484 10004 19490 10056
rect 19610 10044 19616 10056
rect 19571 10016 19616 10044
rect 19610 10004 19616 10016
rect 19668 10004 19674 10056
rect 25409 10047 25467 10053
rect 25409 10044 25421 10047
rect 24688 10016 25421 10044
rect 6512 9948 6960 9976
rect 6512 9936 6518 9948
rect 10962 9936 10968 9988
rect 11020 9936 11026 9988
rect 19444 9976 19472 10004
rect 20162 9976 20168 9988
rect 19444 9948 20168 9976
rect 20162 9936 20168 9948
rect 20220 9936 20226 9988
rect 24688 9920 24716 10016
rect 25409 10013 25421 10016
rect 25455 10044 25467 10047
rect 25866 10044 25872 10056
rect 25455 10016 25872 10044
rect 25455 10013 25467 10016
rect 25409 10007 25467 10013
rect 25866 10004 25872 10016
rect 25924 10004 25930 10056
rect 1578 9908 1584 9920
rect 1539 9880 1584 9908
rect 1578 9868 1584 9880
rect 1636 9868 1642 9920
rect 2682 9908 2688 9920
rect 2643 9880 2688 9908
rect 2682 9868 2688 9880
rect 2740 9868 2746 9920
rect 7374 9908 7380 9920
rect 7335 9880 7380 9908
rect 7374 9868 7380 9880
rect 7432 9868 7438 9920
rect 7929 9911 7987 9917
rect 7929 9877 7941 9911
rect 7975 9908 7987 9911
rect 8110 9908 8116 9920
rect 7975 9880 8116 9908
rect 7975 9877 7987 9880
rect 7929 9871 7987 9877
rect 8110 9868 8116 9880
rect 8168 9868 8174 9920
rect 12802 9908 12808 9920
rect 12763 9880 12808 9908
rect 12802 9868 12808 9880
rect 12860 9868 12866 9920
rect 13630 9908 13636 9920
rect 13591 9880 13636 9908
rect 13630 9868 13636 9880
rect 13688 9868 13694 9920
rect 18693 9911 18751 9917
rect 18693 9877 18705 9911
rect 18739 9908 18751 9911
rect 19242 9908 19248 9920
rect 18739 9880 19248 9908
rect 18739 9877 18751 9880
rect 18693 9871 18751 9877
rect 19242 9868 19248 9880
rect 19300 9868 19306 9920
rect 24670 9908 24676 9920
rect 24631 9880 24676 9908
rect 24670 9868 24676 9880
rect 24728 9868 24734 9920
rect 24854 9908 24860 9920
rect 24815 9880 24860 9908
rect 24854 9868 24860 9880
rect 24912 9868 24918 9920
rect 26694 9908 26700 9920
rect 26655 9880 26700 9908
rect 26694 9868 26700 9880
rect 26752 9868 26758 9920
rect 1104 9818 28888 9840
rect 1104 9766 5982 9818
rect 6034 9766 6046 9818
rect 6098 9766 6110 9818
rect 6162 9766 6174 9818
rect 6226 9766 15982 9818
rect 16034 9766 16046 9818
rect 16098 9766 16110 9818
rect 16162 9766 16174 9818
rect 16226 9766 25982 9818
rect 26034 9766 26046 9818
rect 26098 9766 26110 9818
rect 26162 9766 26174 9818
rect 26226 9766 28888 9818
rect 1104 9744 28888 9766
rect 2498 9704 2504 9716
rect 2459 9676 2504 9704
rect 2498 9664 2504 9676
rect 2556 9664 2562 9716
rect 5810 9664 5816 9716
rect 5868 9704 5874 9716
rect 5997 9707 6055 9713
rect 5997 9704 6009 9707
rect 5868 9676 6009 9704
rect 5868 9664 5874 9676
rect 5997 9673 6009 9676
rect 6043 9673 6055 9707
rect 8018 9704 8024 9716
rect 5997 9667 6055 9673
rect 6932 9676 8024 9704
rect 5537 9639 5595 9645
rect 5537 9605 5549 9639
rect 5583 9636 5595 9639
rect 6730 9636 6736 9648
rect 5583 9608 6736 9636
rect 5583 9605 5595 9608
rect 5537 9599 5595 9605
rect 6730 9596 6736 9608
rect 6788 9636 6794 9648
rect 6825 9639 6883 9645
rect 6825 9636 6837 9639
rect 6788 9608 6837 9636
rect 6788 9596 6794 9608
rect 6825 9605 6837 9608
rect 6871 9605 6883 9639
rect 6825 9599 6883 9605
rect 2038 9568 2044 9580
rect 1412 9540 2044 9568
rect 1412 9509 1440 9540
rect 2038 9528 2044 9540
rect 2096 9528 2102 9580
rect 3510 9568 3516 9580
rect 3471 9540 3516 9568
rect 3510 9528 3516 9540
rect 3568 9528 3574 9580
rect 6932 9568 6960 9676
rect 8018 9664 8024 9676
rect 8076 9664 8082 9716
rect 8202 9704 8208 9716
rect 8163 9676 8208 9704
rect 8202 9664 8208 9676
rect 8260 9664 8266 9716
rect 9769 9707 9827 9713
rect 9769 9673 9781 9707
rect 9815 9704 9827 9707
rect 9858 9704 9864 9716
rect 9815 9676 9864 9704
rect 9815 9673 9827 9676
rect 9769 9667 9827 9673
rect 9858 9664 9864 9676
rect 9916 9664 9922 9716
rect 10505 9707 10563 9713
rect 10505 9673 10517 9707
rect 10551 9704 10563 9707
rect 10686 9704 10692 9716
rect 10551 9676 10692 9704
rect 10551 9673 10563 9676
rect 10505 9667 10563 9673
rect 10686 9664 10692 9676
rect 10744 9664 10750 9716
rect 13170 9664 13176 9716
rect 13228 9704 13234 9716
rect 13446 9704 13452 9716
rect 13228 9676 13452 9704
rect 13228 9664 13234 9676
rect 13446 9664 13452 9676
rect 13504 9664 13510 9716
rect 14182 9704 14188 9716
rect 14143 9676 14188 9704
rect 14182 9664 14188 9676
rect 14240 9704 14246 9716
rect 14461 9707 14519 9713
rect 14461 9704 14473 9707
rect 14240 9676 14473 9704
rect 14240 9664 14246 9676
rect 14461 9673 14473 9676
rect 14507 9704 14519 9707
rect 14829 9707 14887 9713
rect 14829 9704 14841 9707
rect 14507 9676 14841 9704
rect 14507 9673 14519 9676
rect 14461 9667 14519 9673
rect 14829 9673 14841 9676
rect 14875 9673 14887 9707
rect 16850 9704 16856 9716
rect 14829 9667 14887 9673
rect 16500 9676 16856 9704
rect 7282 9596 7288 9648
rect 7340 9636 7346 9648
rect 7466 9636 7472 9648
rect 7340 9608 7472 9636
rect 7340 9596 7346 9608
rect 7466 9596 7472 9608
rect 7524 9596 7530 9648
rect 10597 9639 10655 9645
rect 10597 9605 10609 9639
rect 10643 9636 10655 9639
rect 10870 9636 10876 9648
rect 10643 9608 10876 9636
rect 10643 9605 10655 9608
rect 10597 9599 10655 9605
rect 10870 9596 10876 9608
rect 10928 9596 10934 9648
rect 7374 9568 7380 9580
rect 6196 9540 6960 9568
rect 7335 9540 7380 9568
rect 3786 9509 3792 9512
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9469 1455 9503
rect 1397 9463 1455 9469
rect 3421 9503 3479 9509
rect 3421 9469 3433 9503
rect 3467 9500 3479 9503
rect 3780 9500 3792 9509
rect 3467 9472 3792 9500
rect 3467 9469 3479 9472
rect 3421 9463 3479 9469
rect 3780 9463 3792 9472
rect 3786 9460 3792 9463
rect 3844 9460 3850 9512
rect 6086 9460 6092 9512
rect 6144 9500 6150 9512
rect 6196 9509 6224 9540
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 10962 9528 10968 9580
rect 11020 9568 11026 9580
rect 11149 9571 11207 9577
rect 11149 9568 11161 9571
rect 11020 9540 11161 9568
rect 11020 9528 11026 9540
rect 11149 9537 11161 9540
rect 11195 9568 11207 9571
rect 11977 9571 12035 9577
rect 11977 9568 11989 9571
rect 11195 9540 11989 9568
rect 11195 9537 11207 9540
rect 11149 9531 11207 9537
rect 11977 9537 11989 9540
rect 12023 9537 12035 9571
rect 14844 9568 14872 9667
rect 14844 9540 15148 9568
rect 11977 9531 12035 9537
rect 6181 9503 6239 9509
rect 6181 9500 6193 9503
rect 6144 9472 6193 9500
rect 6144 9460 6150 9472
rect 6181 9469 6193 9472
rect 6227 9469 6239 9503
rect 6181 9463 6239 9469
rect 6546 9460 6552 9512
rect 6604 9500 6610 9512
rect 6641 9503 6699 9509
rect 6641 9500 6653 9503
rect 6604 9472 6653 9500
rect 6604 9460 6610 9472
rect 6641 9469 6653 9472
rect 6687 9500 6699 9503
rect 7285 9503 7343 9509
rect 7285 9500 7297 9503
rect 6687 9472 7297 9500
rect 6687 9469 6699 9472
rect 6641 9463 6699 9469
rect 7285 9469 7297 9472
rect 7331 9500 7343 9503
rect 7742 9500 7748 9512
rect 7331 9472 7748 9500
rect 7331 9469 7343 9472
rect 7285 9463 7343 9469
rect 7742 9460 7748 9472
rect 7800 9460 7806 9512
rect 9674 9460 9680 9512
rect 9732 9500 9738 9512
rect 12802 9500 12808 9512
rect 9732 9472 10088 9500
rect 12763 9472 12808 9500
rect 9732 9460 9738 9472
rect 5905 9435 5963 9441
rect 5905 9401 5917 9435
rect 5951 9432 5963 9435
rect 6822 9432 6828 9444
rect 5951 9404 6828 9432
rect 5951 9401 5963 9404
rect 5905 9395 5963 9401
rect 6822 9392 6828 9404
rect 6880 9392 6886 9444
rect 6914 9392 6920 9444
rect 6972 9432 6978 9444
rect 7193 9435 7251 9441
rect 7193 9432 7205 9435
rect 6972 9404 7205 9432
rect 6972 9392 6978 9404
rect 7193 9401 7205 9404
rect 7239 9432 7251 9435
rect 7837 9435 7895 9441
rect 7837 9432 7849 9435
rect 7239 9404 7849 9432
rect 7239 9401 7251 9404
rect 7193 9395 7251 9401
rect 7837 9401 7849 9404
rect 7883 9401 7895 9435
rect 7837 9395 7895 9401
rect 1394 9324 1400 9376
rect 1452 9364 1458 9376
rect 1581 9367 1639 9373
rect 1581 9364 1593 9367
rect 1452 9336 1593 9364
rect 1452 9324 1458 9336
rect 1581 9333 1593 9336
rect 1627 9333 1639 9367
rect 1581 9327 1639 9333
rect 4246 9324 4252 9376
rect 4304 9364 4310 9376
rect 4893 9367 4951 9373
rect 4893 9364 4905 9367
rect 4304 9336 4905 9364
rect 4304 9324 4310 9336
rect 4893 9333 4905 9336
rect 4939 9333 4951 9367
rect 4893 9327 4951 9333
rect 5534 9324 5540 9376
rect 5592 9364 5598 9376
rect 6730 9364 6736 9376
rect 5592 9336 6736 9364
rect 5592 9324 5598 9336
rect 6730 9324 6736 9336
rect 6788 9324 6794 9376
rect 10060 9364 10088 9472
rect 12802 9460 12808 9472
rect 12860 9460 12866 9512
rect 12894 9460 12900 9512
rect 12952 9500 12958 9512
rect 13446 9500 13452 9512
rect 12952 9472 13452 9500
rect 12952 9460 12958 9472
rect 13446 9460 13452 9472
rect 13504 9460 13510 9512
rect 15010 9500 15016 9512
rect 14971 9472 15016 9500
rect 15010 9460 15016 9472
rect 15068 9460 15074 9512
rect 15120 9500 15148 9540
rect 16298 9528 16304 9580
rect 16356 9568 16362 9580
rect 16500 9568 16528 9676
rect 16850 9664 16856 9676
rect 16908 9664 16914 9716
rect 18690 9704 18696 9716
rect 18651 9676 18696 9704
rect 18690 9664 18696 9676
rect 18748 9664 18754 9716
rect 19610 9664 19616 9716
rect 19668 9704 19674 9716
rect 19797 9707 19855 9713
rect 19797 9704 19809 9707
rect 19668 9676 19809 9704
rect 19668 9664 19674 9676
rect 19797 9673 19809 9676
rect 19843 9704 19855 9707
rect 22002 9704 22008 9716
rect 19843 9676 22008 9704
rect 19843 9673 19855 9676
rect 19797 9667 19855 9673
rect 22002 9664 22008 9676
rect 22060 9704 22066 9716
rect 22373 9707 22431 9713
rect 22373 9704 22385 9707
rect 22060 9676 22385 9704
rect 22060 9664 22066 9676
rect 22373 9673 22385 9676
rect 22419 9673 22431 9707
rect 22373 9667 22431 9673
rect 25409 9707 25467 9713
rect 25409 9673 25421 9707
rect 25455 9704 25467 9707
rect 25498 9704 25504 9716
rect 25455 9676 25504 9704
rect 25455 9673 25467 9676
rect 25409 9667 25467 9673
rect 25498 9664 25504 9676
rect 25556 9664 25562 9716
rect 26510 9664 26516 9716
rect 26568 9704 26574 9716
rect 26881 9707 26939 9713
rect 26881 9704 26893 9707
rect 26568 9676 26893 9704
rect 26568 9664 26574 9676
rect 26881 9673 26893 9676
rect 26927 9673 26939 9707
rect 26881 9667 26939 9673
rect 16356 9540 16528 9568
rect 16356 9528 16362 9540
rect 19334 9528 19340 9580
rect 19392 9568 19398 9580
rect 19429 9571 19487 9577
rect 19429 9568 19441 9571
rect 19392 9540 19441 9568
rect 19392 9528 19398 9540
rect 19429 9537 19441 9540
rect 19475 9568 19487 9571
rect 20622 9568 20628 9580
rect 19475 9540 20628 9568
rect 19475 9537 19487 9540
rect 19429 9531 19487 9537
rect 20622 9528 20628 9540
rect 20680 9528 20686 9580
rect 25866 9528 25872 9580
rect 25924 9568 25930 9580
rect 26326 9568 26332 9580
rect 25924 9540 26332 9568
rect 25924 9528 25930 9540
rect 26326 9528 26332 9540
rect 26384 9568 26390 9580
rect 26421 9571 26479 9577
rect 26421 9568 26433 9571
rect 26384 9540 26433 9568
rect 26384 9528 26390 9540
rect 26421 9537 26433 9540
rect 26467 9537 26479 9571
rect 26421 9531 26479 9537
rect 15269 9503 15327 9509
rect 15269 9500 15281 9503
rect 15120 9472 15281 9500
rect 15269 9469 15281 9472
rect 15315 9469 15327 9503
rect 20993 9503 21051 9509
rect 20993 9500 21005 9503
rect 15269 9463 15327 9469
rect 20456 9472 21005 9500
rect 10137 9435 10195 9441
rect 10137 9401 10149 9435
rect 10183 9432 10195 9435
rect 11057 9435 11115 9441
rect 11057 9432 11069 9435
rect 10183 9404 11069 9432
rect 10183 9401 10195 9404
rect 10137 9395 10195 9401
rect 11057 9401 11069 9404
rect 11103 9432 11115 9435
rect 12713 9435 12771 9441
rect 11103 9404 12388 9432
rect 11103 9401 11115 9404
rect 11057 9395 11115 9401
rect 10965 9367 11023 9373
rect 10965 9364 10977 9367
rect 10060 9336 10977 9364
rect 10965 9333 10977 9336
rect 11011 9364 11023 9367
rect 11609 9367 11667 9373
rect 11609 9364 11621 9367
rect 11011 9336 11621 9364
rect 11011 9333 11023 9336
rect 10965 9327 11023 9333
rect 11609 9333 11621 9336
rect 11655 9333 11667 9367
rect 12360 9364 12388 9404
rect 12713 9401 12725 9435
rect 12759 9432 12771 9435
rect 13072 9435 13130 9441
rect 13072 9432 13084 9435
rect 12759 9404 13084 9432
rect 12759 9401 12771 9404
rect 12713 9395 12771 9401
rect 13072 9401 13084 9404
rect 13118 9432 13130 9435
rect 13538 9432 13544 9444
rect 13118 9404 13544 9432
rect 13118 9401 13130 9404
rect 13072 9395 13130 9401
rect 13538 9392 13544 9404
rect 13596 9392 13602 9444
rect 18969 9435 19027 9441
rect 18969 9432 18981 9435
rect 16224 9404 18981 9432
rect 16224 9364 16252 9404
rect 18969 9401 18981 9404
rect 19015 9432 19027 9435
rect 19426 9432 19432 9444
rect 19015 9404 19432 9432
rect 19015 9401 19027 9404
rect 18969 9395 19027 9401
rect 19426 9392 19432 9404
rect 19484 9392 19490 9444
rect 20456 9376 20484 9472
rect 20993 9469 21005 9472
rect 21039 9500 21051 9503
rect 22094 9500 22100 9512
rect 21039 9472 22100 9500
rect 21039 9469 21051 9472
rect 20993 9463 21051 9469
rect 22094 9460 22100 9472
rect 22152 9460 22158 9512
rect 23658 9500 23664 9512
rect 23619 9472 23664 9500
rect 23658 9460 23664 9472
rect 23716 9460 23722 9512
rect 25777 9503 25835 9509
rect 25777 9469 25789 9503
rect 25823 9500 25835 9503
rect 26237 9503 26295 9509
rect 26237 9500 26249 9503
rect 25823 9472 26249 9500
rect 25823 9469 25835 9472
rect 25777 9463 25835 9469
rect 26237 9469 26249 9472
rect 26283 9500 26295 9503
rect 26510 9500 26516 9512
rect 26283 9472 26516 9500
rect 26283 9469 26295 9472
rect 26237 9463 26295 9469
rect 26510 9460 26516 9472
rect 26568 9460 26574 9512
rect 20901 9435 20959 9441
rect 20901 9401 20913 9435
rect 20947 9432 20959 9435
rect 21238 9435 21296 9441
rect 21238 9432 21250 9435
rect 20947 9404 21250 9432
rect 20947 9401 20959 9404
rect 20901 9395 20959 9401
rect 21238 9401 21250 9404
rect 21284 9432 21296 9435
rect 21450 9432 21456 9444
rect 21284 9404 21456 9432
rect 21284 9401 21296 9404
rect 21238 9395 21296 9401
rect 21450 9392 21456 9404
rect 21508 9392 21514 9444
rect 23906 9435 23964 9441
rect 23906 9432 23918 9435
rect 23492 9404 23918 9432
rect 23492 9376 23520 9404
rect 23906 9401 23918 9404
rect 23952 9432 23964 9435
rect 24670 9432 24676 9444
rect 23952 9404 24676 9432
rect 23952 9401 23964 9404
rect 23906 9395 23964 9401
rect 24670 9392 24676 9404
rect 24728 9392 24734 9444
rect 25958 9392 25964 9444
rect 26016 9432 26022 9444
rect 26329 9435 26387 9441
rect 26329 9432 26341 9435
rect 26016 9404 26341 9432
rect 26016 9392 26022 9404
rect 26329 9401 26341 9404
rect 26375 9401 26387 9435
rect 26329 9395 26387 9401
rect 16390 9364 16396 9376
rect 12360 9336 16252 9364
rect 16351 9336 16396 9364
rect 11609 9327 11667 9333
rect 16390 9324 16396 9336
rect 16448 9324 16454 9376
rect 20438 9364 20444 9376
rect 20399 9336 20444 9364
rect 20438 9324 20444 9336
rect 20496 9324 20502 9376
rect 23474 9364 23480 9376
rect 23435 9336 23480 9364
rect 23474 9324 23480 9336
rect 23532 9324 23538 9376
rect 25038 9364 25044 9376
rect 24999 9336 25044 9364
rect 25038 9324 25044 9336
rect 25096 9324 25102 9376
rect 25866 9364 25872 9376
rect 25827 9336 25872 9364
rect 25866 9324 25872 9336
rect 25924 9324 25930 9376
rect 1104 9274 28888 9296
rect 1104 9222 10982 9274
rect 11034 9222 11046 9274
rect 11098 9222 11110 9274
rect 11162 9222 11174 9274
rect 11226 9222 20982 9274
rect 21034 9222 21046 9274
rect 21098 9222 21110 9274
rect 21162 9222 21174 9274
rect 21226 9222 28888 9274
rect 1104 9200 28888 9222
rect 1670 9160 1676 9172
rect 1631 9132 1676 9160
rect 1670 9120 1676 9132
rect 1728 9120 1734 9172
rect 3513 9163 3571 9169
rect 3513 9129 3525 9163
rect 3559 9160 3571 9163
rect 3786 9160 3792 9172
rect 3559 9132 3792 9160
rect 3559 9129 3571 9132
rect 3513 9123 3571 9129
rect 3786 9120 3792 9132
rect 3844 9120 3850 9172
rect 6086 9160 6092 9172
rect 6047 9132 6092 9160
rect 6086 9120 6092 9132
rect 6144 9120 6150 9172
rect 6454 9160 6460 9172
rect 6415 9132 6460 9160
rect 6454 9120 6460 9132
rect 6512 9120 6518 9172
rect 6822 9160 6828 9172
rect 6783 9132 6828 9160
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 11330 9120 11336 9172
rect 11388 9160 11394 9172
rect 11609 9163 11667 9169
rect 11609 9160 11621 9163
rect 11388 9132 11621 9160
rect 11388 9120 11394 9132
rect 11609 9129 11621 9132
rect 11655 9129 11667 9163
rect 13722 9160 13728 9172
rect 13683 9132 13728 9160
rect 11609 9123 11667 9129
rect 13722 9120 13728 9132
rect 13780 9120 13786 9172
rect 14090 9160 14096 9172
rect 14051 9132 14096 9160
rect 14090 9120 14096 9132
rect 14148 9120 14154 9172
rect 21358 9120 21364 9172
rect 21416 9160 21422 9172
rect 22465 9163 22523 9169
rect 22465 9160 22477 9163
rect 21416 9132 22477 9160
rect 21416 9120 21422 9132
rect 22465 9129 22477 9132
rect 22511 9129 22523 9163
rect 22465 9123 22523 9129
rect 22738 9120 22744 9172
rect 22796 9160 22802 9172
rect 22925 9163 22983 9169
rect 22925 9160 22937 9163
rect 22796 9132 22937 9160
rect 22796 9120 22802 9132
rect 22925 9129 22937 9132
rect 22971 9129 22983 9163
rect 22925 9123 22983 9129
rect 24213 9163 24271 9169
rect 24213 9129 24225 9163
rect 24259 9129 24271 9163
rect 24213 9123 24271 9129
rect 24581 9163 24639 9169
rect 24581 9129 24593 9163
rect 24627 9160 24639 9163
rect 24854 9160 24860 9172
rect 24627 9132 24860 9160
rect 24627 9129 24639 9132
rect 24581 9123 24639 9129
rect 2498 9052 2504 9104
rect 2556 9092 2562 9104
rect 2777 9095 2835 9101
rect 2777 9092 2789 9095
rect 2556 9064 2789 9092
rect 2556 9052 2562 9064
rect 2777 9061 2789 9064
rect 2823 9092 2835 9095
rect 3602 9092 3608 9104
rect 2823 9064 3608 9092
rect 2823 9061 2835 9064
rect 2777 9055 2835 9061
rect 3602 9052 3608 9064
rect 3660 9052 3666 9104
rect 7282 9092 7288 9104
rect 6472 9064 7288 9092
rect 6472 9036 6500 9064
rect 7282 9052 7288 9064
rect 7340 9052 7346 9104
rect 10410 9052 10416 9104
rect 10468 9101 10474 9104
rect 10468 9095 10532 9101
rect 10468 9061 10486 9095
rect 10520 9061 10532 9095
rect 10468 9055 10532 9061
rect 10468 9052 10474 9055
rect 16390 9052 16396 9104
rect 16448 9092 16454 9104
rect 17402 9101 17408 9104
rect 17374 9095 17408 9101
rect 17374 9092 17386 9095
rect 16448 9064 17386 9092
rect 16448 9052 16454 9064
rect 17374 9061 17386 9064
rect 17460 9092 17466 9104
rect 21269 9095 21327 9101
rect 17460 9064 17522 9092
rect 17374 9055 17408 9061
rect 17402 9052 17408 9055
rect 17460 9052 17466 9064
rect 21269 9061 21281 9095
rect 21315 9092 21327 9095
rect 21542 9092 21548 9104
rect 21315 9064 21548 9092
rect 21315 9061 21327 9064
rect 21269 9055 21327 9061
rect 21542 9052 21548 9064
rect 21600 9092 21606 9104
rect 24228 9092 24256 9123
rect 24854 9120 24860 9132
rect 24912 9120 24918 9172
rect 25222 9160 25228 9172
rect 25183 9132 25228 9160
rect 25222 9120 25228 9132
rect 25280 9120 25286 9172
rect 24670 9092 24676 9104
rect 21600 9064 24256 9092
rect 24583 9064 24676 9092
rect 21600 9052 21606 9064
rect 24670 9052 24676 9064
rect 24728 9092 24734 9104
rect 25866 9092 25872 9104
rect 24728 9064 25872 9092
rect 24728 9052 24734 9064
rect 25866 9052 25872 9064
rect 25924 9052 25930 9104
rect 6454 8984 6460 9036
rect 6512 8984 6518 9036
rect 7193 9027 7251 9033
rect 7193 8993 7205 9027
rect 7239 9024 7251 9027
rect 7466 9024 7472 9036
rect 7239 8996 7472 9024
rect 7239 8993 7251 8996
rect 7193 8987 7251 8993
rect 7466 8984 7472 8996
rect 7524 8984 7530 9036
rect 8110 8984 8116 9036
rect 8168 9024 8174 9036
rect 8570 9024 8576 9036
rect 8168 8996 8576 9024
rect 8168 8984 8174 8996
rect 8570 8984 8576 8996
rect 8628 9024 8634 9036
rect 9125 9027 9183 9033
rect 9125 9024 9137 9027
rect 8628 8996 9137 9024
rect 8628 8984 8634 8996
rect 9125 8993 9137 8996
rect 9171 8993 9183 9027
rect 9125 8987 9183 8993
rect 15010 8984 15016 9036
rect 15068 9024 15074 9036
rect 15105 9027 15163 9033
rect 15105 9024 15117 9027
rect 15068 8996 15117 9024
rect 15068 8984 15074 8996
rect 15105 8993 15117 8996
rect 15151 9024 15163 9027
rect 17129 9027 17187 9033
rect 17129 9024 17141 9027
rect 15151 8996 17141 9024
rect 15151 8993 15163 8996
rect 15105 8987 15163 8993
rect 17129 8993 17141 8996
rect 17175 9024 17187 9027
rect 17862 9024 17868 9036
rect 17175 8996 17868 9024
rect 17175 8993 17187 8996
rect 17129 8987 17187 8993
rect 17862 8984 17868 8996
rect 17920 8984 17926 9036
rect 19334 8984 19340 9036
rect 19392 9024 19398 9036
rect 19521 9027 19579 9033
rect 19521 9024 19533 9027
rect 19392 8996 19533 9024
rect 19392 8984 19398 8996
rect 19521 8993 19533 8996
rect 19567 9024 19579 9027
rect 20530 9024 20536 9036
rect 19567 8996 20536 9024
rect 19567 8993 19579 8996
rect 19521 8987 19579 8993
rect 20530 8984 20536 8996
rect 20588 9024 20594 9036
rect 20717 9027 20775 9033
rect 20717 9024 20729 9027
rect 20588 8996 20729 9024
rect 20588 8984 20594 8996
rect 20717 8993 20729 8996
rect 20763 8993 20775 9027
rect 22830 9024 22836 9036
rect 22791 8996 22836 9024
rect 20717 8987 20775 8993
rect 22830 8984 22836 8996
rect 22888 8984 22894 9036
rect 2317 8959 2375 8965
rect 2317 8925 2329 8959
rect 2363 8956 2375 8959
rect 2866 8956 2872 8968
rect 2363 8928 2872 8956
rect 2363 8925 2375 8928
rect 2317 8919 2375 8925
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 3053 8959 3111 8965
rect 3053 8925 3065 8959
rect 3099 8956 3111 8959
rect 4246 8956 4252 8968
rect 3099 8928 4252 8956
rect 3099 8925 3111 8928
rect 3053 8919 3111 8925
rect 4246 8916 4252 8928
rect 4304 8916 4310 8968
rect 7374 8956 7380 8968
rect 7335 8928 7380 8956
rect 7374 8916 7380 8928
rect 7432 8916 7438 8968
rect 10229 8959 10287 8965
rect 10229 8956 10241 8959
rect 9048 8928 10241 8956
rect 9048 8832 9076 8928
rect 10229 8925 10241 8928
rect 10275 8925 10287 8959
rect 21358 8956 21364 8968
rect 21319 8928 21364 8956
rect 10229 8919 10287 8925
rect 21358 8916 21364 8928
rect 21416 8916 21422 8968
rect 21450 8916 21456 8968
rect 21508 8956 21514 8968
rect 23014 8956 23020 8968
rect 21508 8928 21553 8956
rect 22975 8928 23020 8956
rect 21508 8916 21514 8928
rect 23014 8916 23020 8928
rect 23072 8956 23078 8968
rect 24765 8959 24823 8965
rect 24765 8956 24777 8959
rect 23072 8928 24777 8956
rect 23072 8916 23078 8928
rect 24765 8925 24777 8928
rect 24811 8956 24823 8959
rect 25038 8956 25044 8968
rect 24811 8928 25044 8956
rect 24811 8925 24823 8928
rect 24765 8919 24823 8925
rect 25038 8916 25044 8928
rect 25096 8916 25102 8968
rect 25866 8956 25872 8968
rect 25827 8928 25872 8956
rect 25866 8916 25872 8928
rect 25924 8916 25930 8968
rect 2409 8823 2467 8829
rect 2409 8789 2421 8823
rect 2455 8820 2467 8823
rect 2590 8820 2596 8832
rect 2455 8792 2596 8820
rect 2455 8789 2467 8792
rect 2409 8783 2467 8789
rect 2590 8780 2596 8792
rect 2648 8780 2654 8832
rect 4890 8820 4896 8832
rect 4851 8792 4896 8820
rect 4890 8780 4896 8792
rect 4948 8780 4954 8832
rect 8941 8823 8999 8829
rect 8941 8789 8953 8823
rect 8987 8820 8999 8823
rect 9030 8820 9036 8832
rect 8987 8792 9036 8820
rect 8987 8789 8999 8792
rect 8941 8783 8999 8789
rect 9030 8780 9036 8792
rect 9088 8780 9094 8832
rect 12802 8780 12808 8832
rect 12860 8820 12866 8832
rect 12897 8823 12955 8829
rect 12897 8820 12909 8823
rect 12860 8792 12909 8820
rect 12860 8780 12866 8792
rect 12897 8789 12909 8792
rect 12943 8820 12955 8823
rect 13262 8820 13268 8832
rect 12943 8792 13268 8820
rect 12943 8789 12955 8792
rect 12897 8783 12955 8789
rect 13262 8780 13268 8792
rect 13320 8780 13326 8832
rect 16482 8820 16488 8832
rect 16443 8792 16488 8820
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 18506 8820 18512 8832
rect 18467 8792 18512 8820
rect 18506 8780 18512 8792
rect 18564 8780 18570 8832
rect 19337 8823 19395 8829
rect 19337 8789 19349 8823
rect 19383 8820 19395 8823
rect 19426 8820 19432 8832
rect 19383 8792 19432 8820
rect 19383 8789 19395 8792
rect 19337 8783 19395 8789
rect 19426 8780 19432 8792
rect 19484 8780 19490 8832
rect 19702 8780 19708 8832
rect 19760 8820 19766 8832
rect 20438 8820 20444 8832
rect 19760 8792 20444 8820
rect 19760 8780 19766 8792
rect 20438 8780 20444 8792
rect 20496 8820 20502 8832
rect 20533 8823 20591 8829
rect 20533 8820 20545 8823
rect 20496 8792 20545 8820
rect 20496 8780 20502 8792
rect 20533 8789 20545 8792
rect 20579 8789 20591 8823
rect 20533 8783 20591 8789
rect 20806 8780 20812 8832
rect 20864 8820 20870 8832
rect 20901 8823 20959 8829
rect 20901 8820 20913 8823
rect 20864 8792 20913 8820
rect 20864 8780 20870 8792
rect 20901 8789 20913 8792
rect 20947 8789 20959 8823
rect 23658 8820 23664 8832
rect 23619 8792 23664 8820
rect 20901 8783 20959 8789
rect 23658 8780 23664 8792
rect 23716 8780 23722 8832
rect 1104 8730 28888 8752
rect 1104 8678 5982 8730
rect 6034 8678 6046 8730
rect 6098 8678 6110 8730
rect 6162 8678 6174 8730
rect 6226 8678 15982 8730
rect 16034 8678 16046 8730
rect 16098 8678 16110 8730
rect 16162 8678 16174 8730
rect 16226 8678 25982 8730
rect 26034 8678 26046 8730
rect 26098 8678 26110 8730
rect 26162 8678 26174 8730
rect 26226 8678 28888 8730
rect 1104 8656 28888 8678
rect 2498 8616 2504 8628
rect 2459 8588 2504 8616
rect 2498 8576 2504 8588
rect 2556 8576 2562 8628
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 3145 8619 3203 8625
rect 3145 8616 3157 8619
rect 2924 8588 3157 8616
rect 2924 8576 2930 8588
rect 3145 8585 3157 8588
rect 3191 8585 3203 8619
rect 8570 8616 8576 8628
rect 8531 8588 8576 8616
rect 3145 8579 3203 8585
rect 8570 8576 8576 8588
rect 8628 8576 8634 8628
rect 10410 8616 10416 8628
rect 10371 8588 10416 8616
rect 10410 8576 10416 8588
rect 10468 8616 10474 8628
rect 10689 8619 10747 8625
rect 10689 8616 10701 8619
rect 10468 8588 10701 8616
rect 10468 8576 10474 8588
rect 10689 8585 10701 8588
rect 10735 8585 10747 8619
rect 10689 8579 10747 8585
rect 10965 8619 11023 8625
rect 10965 8585 10977 8619
rect 11011 8616 11023 8619
rect 13262 8616 13268 8628
rect 11011 8588 13268 8616
rect 11011 8585 11023 8588
rect 10965 8579 11023 8585
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 17402 8616 17408 8628
rect 17363 8588 17408 8616
rect 17402 8576 17408 8588
rect 17460 8576 17466 8628
rect 17862 8616 17868 8628
rect 17823 8588 17868 8616
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 19334 8616 19340 8628
rect 19295 8588 19340 8616
rect 19334 8576 19340 8588
rect 19392 8576 19398 8628
rect 21361 8619 21419 8625
rect 21361 8585 21373 8619
rect 21407 8616 21419 8619
rect 21450 8616 21456 8628
rect 21407 8588 21456 8616
rect 21407 8585 21419 8588
rect 21361 8579 21419 8585
rect 21450 8576 21456 8588
rect 21508 8616 21514 8628
rect 21637 8619 21695 8625
rect 21637 8616 21649 8619
rect 21508 8588 21649 8616
rect 21508 8576 21514 8588
rect 21637 8585 21649 8588
rect 21683 8585 21695 8619
rect 24670 8616 24676 8628
rect 24631 8588 24676 8616
rect 21637 8579 21695 8585
rect 24670 8576 24676 8588
rect 24728 8576 24734 8628
rect 24854 8576 24860 8628
rect 24912 8616 24918 8628
rect 24949 8619 25007 8625
rect 24949 8616 24961 8619
rect 24912 8588 24961 8616
rect 24912 8576 24918 8588
rect 24949 8585 24961 8588
rect 24995 8585 25007 8619
rect 26602 8616 26608 8628
rect 26563 8588 26608 8616
rect 24949 8579 25007 8585
rect 26602 8576 26608 8588
rect 26660 8576 26666 8628
rect 1578 8548 1584 8560
rect 1539 8520 1584 8548
rect 1578 8508 1584 8520
rect 1636 8508 1642 8560
rect 3053 8551 3111 8557
rect 3053 8517 3065 8551
rect 3099 8548 3111 8551
rect 3970 8548 3976 8560
rect 3099 8520 3976 8548
rect 3099 8517 3111 8520
rect 3053 8511 3111 8517
rect 2041 8483 2099 8489
rect 2041 8480 2053 8483
rect 1412 8452 2053 8480
rect 1412 8421 1440 8452
rect 2041 8449 2053 8452
rect 2087 8480 2099 8483
rect 2866 8480 2872 8492
rect 2087 8452 2872 8480
rect 2087 8449 2099 8452
rect 2041 8443 2099 8449
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 3620 8489 3648 8520
rect 3970 8508 3976 8520
rect 4028 8508 4034 8560
rect 4338 8508 4344 8560
rect 4396 8548 4402 8560
rect 4801 8551 4859 8557
rect 4801 8548 4813 8551
rect 4396 8520 4813 8548
rect 4396 8508 4402 8520
rect 4801 8517 4813 8520
rect 4847 8517 4859 8551
rect 4801 8511 4859 8517
rect 3605 8483 3663 8489
rect 3605 8449 3617 8483
rect 3651 8480 3663 8483
rect 3786 8480 3792 8492
rect 3651 8452 3685 8480
rect 3747 8452 3792 8480
rect 3651 8449 3663 8452
rect 3605 8443 3663 8449
rect 3786 8440 3792 8452
rect 3844 8440 3850 8492
rect 5353 8483 5411 8489
rect 5353 8480 5365 8483
rect 4632 8452 5365 8480
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8381 1455 8415
rect 3510 8412 3516 8424
rect 3423 8384 3516 8412
rect 1397 8375 1455 8381
rect 3510 8372 3516 8384
rect 3568 8412 3574 8424
rect 4062 8412 4068 8424
rect 3568 8384 4068 8412
rect 3568 8372 3574 8384
rect 4062 8372 4068 8384
rect 4120 8412 4126 8424
rect 4522 8412 4528 8424
rect 4120 8384 4528 8412
rect 4120 8372 4126 8384
rect 4522 8372 4528 8384
rect 4580 8372 4586 8424
rect 4632 8356 4660 8452
rect 5353 8449 5365 8452
rect 5399 8480 5411 8483
rect 5442 8480 5448 8492
rect 5399 8452 5448 8480
rect 5399 8449 5411 8452
rect 5353 8443 5411 8449
rect 5442 8440 5448 8452
rect 5500 8440 5506 8492
rect 6914 8480 6920 8492
rect 6875 8452 6920 8480
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 16482 8440 16488 8492
rect 16540 8480 16546 8492
rect 16850 8480 16856 8492
rect 16540 8452 16856 8480
rect 16540 8440 16546 8452
rect 16850 8440 16856 8452
rect 16908 8440 16914 8492
rect 17037 8483 17095 8489
rect 17037 8449 17049 8483
rect 17083 8480 17095 8483
rect 18506 8480 18512 8492
rect 17083 8452 18512 8480
rect 17083 8449 17095 8452
rect 17037 8443 17095 8449
rect 4890 8372 4896 8424
rect 4948 8412 4954 8424
rect 5169 8415 5227 8421
rect 5169 8412 5181 8415
rect 4948 8384 5181 8412
rect 4948 8372 4954 8384
rect 5169 8381 5181 8384
rect 5215 8381 5227 8415
rect 9030 8412 9036 8424
rect 8991 8384 9036 8412
rect 5169 8375 5227 8381
rect 9030 8372 9036 8384
rect 9088 8372 9094 8424
rect 10778 8372 10784 8424
rect 10836 8412 10842 8424
rect 14918 8412 14924 8424
rect 10836 8384 14924 8412
rect 10836 8372 10842 8384
rect 14918 8372 14924 8384
rect 14976 8372 14982 8424
rect 16574 8372 16580 8424
rect 16632 8412 16638 8424
rect 17052 8412 17080 8443
rect 18506 8440 18512 8452
rect 18564 8440 18570 8492
rect 22738 8440 22744 8492
rect 22796 8480 22802 8492
rect 22833 8483 22891 8489
rect 22833 8480 22845 8483
rect 22796 8452 22845 8480
rect 22796 8440 22802 8452
rect 22833 8449 22845 8452
rect 22879 8449 22891 8483
rect 22833 8443 22891 8449
rect 16632 8384 17080 8412
rect 16632 8372 16638 8384
rect 19702 8372 19708 8424
rect 19760 8412 19766 8424
rect 19981 8415 20039 8421
rect 19981 8412 19993 8415
rect 19760 8384 19993 8412
rect 19760 8372 19766 8384
rect 19981 8381 19993 8384
rect 20027 8381 20039 8415
rect 26418 8412 26424 8424
rect 26379 8384 26424 8412
rect 19981 8375 20039 8381
rect 26418 8372 26424 8384
rect 26476 8412 26482 8424
rect 26973 8415 27031 8421
rect 26973 8412 26985 8415
rect 26476 8384 26985 8412
rect 26476 8372 26482 8384
rect 26973 8381 26985 8384
rect 27019 8381 27031 8415
rect 26973 8375 27031 8381
rect 4614 8344 4620 8356
rect 4575 8316 4620 8344
rect 4614 8304 4620 8316
rect 4672 8304 4678 8356
rect 6454 8304 6460 8356
rect 6512 8344 6518 8356
rect 6549 8347 6607 8353
rect 6549 8344 6561 8347
rect 6512 8316 6561 8344
rect 6512 8304 6518 8316
rect 6549 8313 6561 8316
rect 6595 8313 6607 8347
rect 6549 8307 6607 8313
rect 8941 8347 8999 8353
rect 8941 8313 8953 8347
rect 8987 8344 8999 8347
rect 9278 8347 9336 8353
rect 9278 8344 9290 8347
rect 8987 8316 9290 8344
rect 8987 8313 8999 8316
rect 8941 8307 8999 8313
rect 9278 8313 9290 8316
rect 9324 8344 9336 8347
rect 9582 8344 9588 8356
rect 9324 8316 9588 8344
rect 9324 8313 9336 8316
rect 9278 8307 9336 8313
rect 9582 8304 9588 8316
rect 9640 8304 9646 8356
rect 15194 8304 15200 8356
rect 15252 8344 15258 8356
rect 16298 8344 16304 8356
rect 15252 8316 16304 8344
rect 15252 8304 15258 8316
rect 16298 8304 16304 8316
rect 16356 8344 16362 8356
rect 16761 8347 16819 8353
rect 16761 8344 16773 8347
rect 16356 8316 16773 8344
rect 16356 8304 16362 8316
rect 16761 8313 16773 8316
rect 16807 8313 16819 8347
rect 16761 8307 16819 8313
rect 19889 8347 19947 8353
rect 19889 8313 19901 8347
rect 19935 8344 19947 8347
rect 20226 8347 20284 8353
rect 20226 8344 20238 8347
rect 19935 8316 20238 8344
rect 19935 8313 19947 8316
rect 19889 8307 19947 8313
rect 20226 8313 20238 8316
rect 20272 8344 20284 8347
rect 20272 8316 22048 8344
rect 20272 8313 20284 8316
rect 20226 8307 20284 8313
rect 4246 8276 4252 8288
rect 4207 8248 4252 8276
rect 4246 8236 4252 8248
rect 4304 8236 4310 8288
rect 5258 8236 5264 8288
rect 5316 8276 5322 8288
rect 7466 8276 7472 8288
rect 5316 8248 5361 8276
rect 7379 8248 7472 8276
rect 5316 8236 5322 8248
rect 7466 8236 7472 8248
rect 7524 8276 7530 8288
rect 7926 8276 7932 8288
rect 7524 8248 7932 8276
rect 7524 8236 7530 8248
rect 7926 8236 7932 8248
rect 7984 8236 7990 8288
rect 10778 8236 10784 8288
rect 10836 8276 10842 8288
rect 10965 8279 11023 8285
rect 10965 8276 10977 8279
rect 10836 8248 10977 8276
rect 10836 8236 10842 8248
rect 10965 8245 10977 8248
rect 11011 8276 11023 8279
rect 11057 8279 11115 8285
rect 11057 8276 11069 8279
rect 11011 8248 11069 8276
rect 11011 8245 11023 8248
rect 10965 8239 11023 8245
rect 11057 8245 11069 8248
rect 11103 8245 11115 8279
rect 16390 8276 16396 8288
rect 16351 8248 16396 8276
rect 11057 8239 11115 8245
rect 16390 8236 16396 8248
rect 16448 8236 16454 8288
rect 22020 8276 22048 8316
rect 22094 8304 22100 8356
rect 22152 8344 22158 8356
rect 22830 8344 22836 8356
rect 22152 8316 22836 8344
rect 22152 8304 22158 8316
rect 22830 8304 22836 8316
rect 22888 8344 22894 8356
rect 23201 8347 23259 8353
rect 23201 8344 23213 8347
rect 22888 8316 23213 8344
rect 22888 8304 22894 8316
rect 23201 8313 23213 8316
rect 23247 8313 23259 8347
rect 23201 8307 23259 8313
rect 22465 8279 22523 8285
rect 22465 8276 22477 8279
rect 22020 8248 22477 8276
rect 22465 8245 22477 8248
rect 22511 8276 22523 8279
rect 23014 8276 23020 8288
rect 22511 8248 23020 8276
rect 22511 8245 22523 8248
rect 22465 8239 22523 8245
rect 23014 8236 23020 8248
rect 23072 8276 23078 8288
rect 24213 8279 24271 8285
rect 24213 8276 24225 8279
rect 23072 8248 24225 8276
rect 23072 8236 23078 8248
rect 24213 8245 24225 8248
rect 24259 8245 24271 8279
rect 24213 8239 24271 8245
rect 1104 8186 28888 8208
rect 1104 8134 10982 8186
rect 11034 8134 11046 8186
rect 11098 8134 11110 8186
rect 11162 8134 11174 8186
rect 11226 8134 20982 8186
rect 21034 8134 21046 8186
rect 21098 8134 21110 8186
rect 21162 8134 21174 8186
rect 21226 8134 28888 8186
rect 1104 8112 28888 8134
rect 3510 8072 3516 8084
rect 3471 8044 3516 8072
rect 3510 8032 3516 8044
rect 3568 8032 3574 8084
rect 4893 8075 4951 8081
rect 4893 8041 4905 8075
rect 4939 8072 4951 8075
rect 5258 8072 5264 8084
rect 4939 8044 5264 8072
rect 4939 8041 4951 8044
rect 4893 8035 4951 8041
rect 5258 8032 5264 8044
rect 5316 8032 5322 8084
rect 5534 8032 5540 8084
rect 5592 8072 5598 8084
rect 6549 8075 6607 8081
rect 6549 8072 6561 8075
rect 5592 8044 6561 8072
rect 5592 8032 5598 8044
rect 6549 8041 6561 8044
rect 6595 8041 6607 8075
rect 6549 8035 6607 8041
rect 6917 8075 6975 8081
rect 6917 8041 6929 8075
rect 6963 8072 6975 8075
rect 7374 8072 7380 8084
rect 6963 8044 7380 8072
rect 6963 8041 6975 8044
rect 6917 8035 6975 8041
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 16482 8072 16488 8084
rect 16443 8044 16488 8072
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 16850 8032 16856 8084
rect 16908 8072 16914 8084
rect 16945 8075 17003 8081
rect 16945 8072 16957 8075
rect 16908 8044 16957 8072
rect 16908 8032 16914 8044
rect 16945 8041 16957 8044
rect 16991 8041 17003 8075
rect 18506 8072 18512 8084
rect 18467 8044 18512 8072
rect 16945 8035 17003 8041
rect 18506 8032 18512 8044
rect 18564 8032 18570 8084
rect 20530 8072 20536 8084
rect 20491 8044 20536 8072
rect 20530 8032 20536 8044
rect 20588 8032 20594 8084
rect 21177 8075 21235 8081
rect 21177 8041 21189 8075
rect 21223 8072 21235 8075
rect 21358 8072 21364 8084
rect 21223 8044 21364 8072
rect 21223 8041 21235 8044
rect 21177 8035 21235 8041
rect 21358 8032 21364 8044
rect 21416 8032 21422 8084
rect 21542 8072 21548 8084
rect 21503 8044 21548 8072
rect 21542 8032 21548 8044
rect 21600 8032 21606 8084
rect 22002 8072 22008 8084
rect 21963 8044 22008 8072
rect 22002 8032 22008 8044
rect 22060 8032 22066 8084
rect 22465 8075 22523 8081
rect 22465 8041 22477 8075
rect 22511 8072 22523 8075
rect 22830 8072 22836 8084
rect 22511 8044 22836 8072
rect 22511 8041 22523 8044
rect 22465 8035 22523 8041
rect 22830 8032 22836 8044
rect 22888 8072 22894 8084
rect 23569 8075 23627 8081
rect 23569 8072 23581 8075
rect 22888 8044 23581 8072
rect 22888 8032 22894 8044
rect 23569 8041 23581 8044
rect 23615 8041 23627 8075
rect 26694 8072 26700 8084
rect 26655 8044 26700 8072
rect 23569 8035 23627 8041
rect 26694 8032 26700 8044
rect 26752 8032 26758 8084
rect 2774 7964 2780 8016
rect 2832 8004 2838 8016
rect 2832 7976 2877 8004
rect 2832 7964 2838 7976
rect 11330 7964 11336 8016
rect 11388 8013 11394 8016
rect 11388 8007 11452 8013
rect 11388 7973 11406 8007
rect 11440 7973 11452 8007
rect 17405 8007 17463 8013
rect 17405 8004 17417 8007
rect 11388 7967 11452 7973
rect 16960 7976 17417 8004
rect 11388 7964 11394 7967
rect 16960 7948 16988 7976
rect 17405 7973 17417 7976
rect 17451 8004 17463 8007
rect 18046 8004 18052 8016
rect 17451 7976 18052 8004
rect 17451 7973 17463 7976
rect 17405 7967 17463 7973
rect 18046 7964 18052 7976
rect 18104 7964 18110 8016
rect 2869 7939 2927 7945
rect 2869 7905 2881 7939
rect 2915 7936 2927 7939
rect 3418 7936 3424 7948
rect 2915 7908 3424 7936
rect 2915 7905 2927 7908
rect 2869 7899 2927 7905
rect 3418 7896 3424 7908
rect 3476 7896 3482 7948
rect 5166 7936 5172 7948
rect 5127 7908 5172 7936
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 5436 7939 5494 7945
rect 5436 7905 5448 7939
rect 5482 7936 5494 7939
rect 5810 7936 5816 7948
rect 5482 7908 5816 7936
rect 5482 7905 5494 7908
rect 5436 7899 5494 7905
rect 5810 7896 5816 7908
rect 5868 7896 5874 7948
rect 16942 7896 16948 7948
rect 17000 7896 17006 7948
rect 17310 7936 17316 7948
rect 17271 7908 17316 7936
rect 17310 7896 17316 7908
rect 17368 7896 17374 7948
rect 20714 7896 20720 7948
rect 20772 7936 20778 7948
rect 21818 7936 21824 7948
rect 20772 7908 21824 7936
rect 20772 7896 20778 7908
rect 21818 7896 21824 7908
rect 21876 7936 21882 7948
rect 22370 7936 22376 7948
rect 21876 7908 22376 7936
rect 21876 7896 21882 7908
rect 22370 7896 22376 7908
rect 22428 7896 22434 7948
rect 23842 7896 23848 7948
rect 23900 7936 23906 7948
rect 23937 7939 23995 7945
rect 23937 7936 23949 7939
rect 23900 7908 23949 7936
rect 23900 7896 23906 7908
rect 23937 7905 23949 7908
rect 23983 7936 23995 7939
rect 25222 7936 25228 7948
rect 23983 7908 25228 7936
rect 23983 7905 23995 7908
rect 23937 7899 23995 7905
rect 25222 7896 25228 7908
rect 25280 7896 25286 7948
rect 26510 7936 26516 7948
rect 26471 7908 26516 7936
rect 26510 7896 26516 7908
rect 26568 7896 26574 7948
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 4246 7868 4252 7880
rect 3099 7840 4252 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 2317 7803 2375 7809
rect 2317 7769 2329 7803
rect 2363 7800 2375 7803
rect 3068 7800 3096 7831
rect 4246 7828 4252 7840
rect 4304 7828 4310 7880
rect 10778 7828 10784 7880
rect 10836 7868 10842 7880
rect 11149 7871 11207 7877
rect 11149 7868 11161 7871
rect 10836 7840 11161 7868
rect 10836 7828 10842 7840
rect 11149 7837 11161 7840
rect 11195 7837 11207 7871
rect 13354 7868 13360 7880
rect 13315 7840 13360 7868
rect 11149 7831 11207 7837
rect 13354 7828 13360 7840
rect 13412 7828 13418 7880
rect 17494 7868 17500 7880
rect 17455 7840 17500 7868
rect 17494 7828 17500 7840
rect 17552 7828 17558 7880
rect 22646 7868 22652 7880
rect 22607 7840 22652 7868
rect 22646 7828 22652 7840
rect 22704 7868 22710 7880
rect 23382 7868 23388 7880
rect 22704 7840 23388 7868
rect 22704 7828 22710 7840
rect 23382 7828 23388 7840
rect 23440 7828 23446 7880
rect 24026 7868 24032 7880
rect 23987 7840 24032 7868
rect 24026 7828 24032 7840
rect 24084 7828 24090 7880
rect 24213 7871 24271 7877
rect 24213 7837 24225 7871
rect 24259 7868 24271 7871
rect 24302 7868 24308 7880
rect 24259 7840 24308 7868
rect 24259 7837 24271 7840
rect 24213 7831 24271 7837
rect 2363 7772 3096 7800
rect 23477 7803 23535 7809
rect 2363 7769 2375 7772
rect 2317 7763 2375 7769
rect 23477 7769 23489 7803
rect 23523 7800 23535 7803
rect 24228 7800 24256 7831
rect 24302 7828 24308 7840
rect 24360 7828 24366 7880
rect 23523 7772 24256 7800
rect 23523 7769 23535 7772
rect 23477 7763 23535 7769
rect 1673 7735 1731 7741
rect 1673 7701 1685 7735
rect 1719 7732 1731 7735
rect 1854 7732 1860 7744
rect 1719 7704 1860 7732
rect 1719 7701 1731 7704
rect 1673 7695 1731 7701
rect 1854 7692 1860 7704
rect 1912 7692 1918 7744
rect 2406 7732 2412 7744
rect 2367 7704 2412 7732
rect 2406 7692 2412 7704
rect 2464 7692 2470 7744
rect 3881 7735 3939 7741
rect 3881 7701 3893 7735
rect 3927 7732 3939 7735
rect 3970 7732 3976 7744
rect 3927 7704 3976 7732
rect 3927 7701 3939 7704
rect 3881 7695 3939 7701
rect 3970 7692 3976 7704
rect 4028 7692 4034 7744
rect 8294 7692 8300 7744
rect 8352 7732 8358 7744
rect 9030 7732 9036 7744
rect 8352 7704 9036 7732
rect 8352 7692 8358 7704
rect 9030 7692 9036 7704
rect 9088 7692 9094 7744
rect 12342 7692 12348 7744
rect 12400 7732 12406 7744
rect 12529 7735 12587 7741
rect 12529 7732 12541 7735
rect 12400 7704 12541 7732
rect 12400 7692 12406 7704
rect 12529 7701 12541 7704
rect 12575 7701 12587 7735
rect 18046 7732 18052 7744
rect 18007 7704 18052 7732
rect 12529 7695 12587 7701
rect 18046 7692 18052 7704
rect 18104 7692 18110 7744
rect 19702 7692 19708 7744
rect 19760 7732 19766 7744
rect 19981 7735 20039 7741
rect 19981 7732 19993 7735
rect 19760 7704 19993 7732
rect 19760 7692 19766 7704
rect 19981 7701 19993 7704
rect 20027 7701 20039 7735
rect 25314 7732 25320 7744
rect 25275 7704 25320 7732
rect 19981 7695 20039 7701
rect 25314 7692 25320 7704
rect 25372 7692 25378 7744
rect 1104 7642 28888 7664
rect 1104 7590 5982 7642
rect 6034 7590 6046 7642
rect 6098 7590 6110 7642
rect 6162 7590 6174 7642
rect 6226 7590 15982 7642
rect 16034 7590 16046 7642
rect 16098 7590 16110 7642
rect 16162 7590 16174 7642
rect 16226 7590 25982 7642
rect 26034 7590 26046 7642
rect 26098 7590 26110 7642
rect 26162 7590 26174 7642
rect 26226 7590 28888 7642
rect 1104 7568 28888 7590
rect 2774 7488 2780 7540
rect 2832 7528 2838 7540
rect 3053 7531 3111 7537
rect 3053 7528 3065 7531
rect 2832 7500 3065 7528
rect 2832 7488 2838 7500
rect 3053 7497 3065 7500
rect 3099 7497 3111 7531
rect 4982 7528 4988 7540
rect 4943 7500 4988 7528
rect 3053 7491 3111 7497
rect 4982 7488 4988 7500
rect 5040 7488 5046 7540
rect 5169 7531 5227 7537
rect 5169 7497 5181 7531
rect 5215 7528 5227 7531
rect 5258 7528 5264 7540
rect 5215 7500 5264 7528
rect 5215 7497 5227 7500
rect 5169 7491 5227 7497
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 15010 7528 15016 7540
rect 14660 7500 15016 7528
rect 14660 7404 14688 7500
rect 15010 7488 15016 7500
rect 15068 7488 15074 7540
rect 16669 7531 16727 7537
rect 16669 7497 16681 7531
rect 16715 7528 16727 7531
rect 17494 7528 17500 7540
rect 16715 7500 17500 7528
rect 16715 7497 16727 7500
rect 16669 7491 16727 7497
rect 17494 7488 17500 7500
rect 17552 7488 17558 7540
rect 21818 7528 21824 7540
rect 21779 7500 21824 7528
rect 21818 7488 21824 7500
rect 21876 7488 21882 7540
rect 22005 7531 22063 7537
rect 22005 7497 22017 7531
rect 22051 7528 22063 7531
rect 22738 7528 22744 7540
rect 22051 7500 22744 7528
rect 22051 7497 22063 7500
rect 22005 7491 22063 7497
rect 22738 7488 22744 7500
rect 22796 7488 22802 7540
rect 23106 7528 23112 7540
rect 23019 7500 23112 7528
rect 23106 7488 23112 7500
rect 23164 7528 23170 7540
rect 24026 7528 24032 7540
rect 23164 7500 24032 7528
rect 23164 7488 23170 7500
rect 24026 7488 24032 7500
rect 24084 7488 24090 7540
rect 24762 7528 24768 7540
rect 24723 7500 24768 7528
rect 24762 7488 24768 7500
rect 24820 7488 24826 7540
rect 25133 7531 25191 7537
rect 25133 7497 25145 7531
rect 25179 7528 25191 7531
rect 25222 7528 25228 7540
rect 25179 7500 25228 7528
rect 25179 7497 25191 7500
rect 25133 7491 25191 7497
rect 25222 7488 25228 7500
rect 25280 7488 25286 7540
rect 26510 7488 26516 7540
rect 26568 7528 26574 7540
rect 26973 7531 27031 7537
rect 26973 7528 26985 7531
rect 26568 7500 26985 7528
rect 26568 7488 26574 7500
rect 26973 7497 26985 7500
rect 27019 7497 27031 7531
rect 26973 7491 27031 7497
rect 23661 7463 23719 7469
rect 23661 7460 23673 7463
rect 22480 7432 23673 7460
rect 22480 7404 22508 7432
rect 23661 7429 23673 7432
rect 23707 7429 23719 7463
rect 23661 7423 23719 7429
rect 26326 7420 26332 7472
rect 26384 7460 26390 7472
rect 26697 7463 26755 7469
rect 26697 7460 26709 7463
rect 26384 7432 26709 7460
rect 26384 7420 26390 7432
rect 26697 7429 26709 7432
rect 26743 7429 26755 7463
rect 26697 7423 26755 7429
rect 2866 7352 2872 7404
rect 2924 7392 2930 7404
rect 4157 7395 4215 7401
rect 4157 7392 4169 7395
rect 2924 7364 4169 7392
rect 2924 7352 2930 7364
rect 4157 7361 4169 7364
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 4246 7352 4252 7404
rect 4304 7392 4310 7404
rect 4709 7395 4767 7401
rect 4709 7392 4721 7395
rect 4304 7364 4721 7392
rect 4304 7352 4310 7364
rect 4709 7361 4721 7364
rect 4755 7392 4767 7395
rect 5810 7392 5816 7404
rect 4755 7364 5816 7392
rect 4755 7361 4767 7364
rect 4709 7355 4767 7361
rect 5810 7352 5816 7364
rect 5868 7392 5874 7404
rect 6270 7392 6276 7404
rect 5868 7364 6276 7392
rect 5868 7352 5874 7364
rect 6270 7352 6276 7364
rect 6328 7352 6334 7404
rect 12158 7392 12164 7404
rect 12119 7364 12164 7392
rect 12158 7352 12164 7364
rect 12216 7352 12222 7404
rect 13078 7392 13084 7404
rect 13039 7364 13084 7392
rect 13078 7352 13084 7364
rect 13136 7352 13142 7404
rect 14642 7392 14648 7404
rect 14555 7364 14648 7392
rect 14642 7352 14648 7364
rect 14700 7352 14706 7404
rect 18598 7392 18604 7404
rect 18559 7364 18604 7392
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 21177 7395 21235 7401
rect 21177 7361 21189 7395
rect 21223 7392 21235 7395
rect 22278 7392 22284 7404
rect 21223 7364 22284 7392
rect 21223 7361 21235 7364
rect 21177 7355 21235 7361
rect 22278 7352 22284 7364
rect 22336 7352 22342 7404
rect 22462 7392 22468 7404
rect 22375 7364 22468 7392
rect 22462 7352 22468 7364
rect 22520 7352 22526 7404
rect 22557 7395 22615 7401
rect 22557 7361 22569 7395
rect 22603 7392 22615 7395
rect 22646 7392 22652 7404
rect 22603 7364 22652 7392
rect 22603 7361 22615 7364
rect 22557 7355 22615 7361
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7324 1455 7327
rect 3973 7327 4031 7333
rect 1443 7296 1900 7324
rect 1443 7293 1455 7296
rect 1397 7287 1455 7293
rect 1872 7268 1900 7296
rect 3973 7293 3985 7327
rect 4019 7324 4031 7327
rect 4062 7324 4068 7336
rect 4019 7296 4068 7324
rect 4019 7293 4031 7296
rect 3973 7287 4031 7293
rect 4062 7284 4068 7296
rect 4120 7284 4126 7336
rect 5166 7284 5172 7336
rect 5224 7324 5230 7336
rect 6549 7327 6607 7333
rect 6549 7324 6561 7327
rect 5224 7296 6561 7324
rect 5224 7284 5230 7296
rect 6549 7293 6561 7296
rect 6595 7293 6607 7327
rect 8294 7324 8300 7336
rect 8255 7296 8300 7324
rect 6549 7287 6607 7293
rect 8294 7284 8300 7296
rect 8352 7284 8358 7336
rect 14912 7327 14970 7333
rect 14912 7324 14924 7327
rect 14844 7296 14924 7324
rect 1670 7265 1676 7268
rect 1664 7219 1676 7265
rect 1728 7256 1734 7268
rect 1728 7228 1764 7256
rect 1670 7216 1676 7219
rect 1728 7216 1734 7228
rect 1854 7216 1860 7268
rect 1912 7216 1918 7268
rect 5626 7256 5632 7268
rect 5587 7228 5632 7256
rect 5626 7216 5632 7228
rect 5684 7216 5690 7268
rect 8205 7259 8263 7265
rect 8205 7225 8217 7259
rect 8251 7256 8263 7259
rect 8542 7259 8600 7265
rect 8542 7256 8554 7259
rect 8251 7228 8554 7256
rect 8251 7225 8263 7228
rect 8205 7219 8263 7225
rect 8542 7225 8554 7228
rect 8588 7256 8600 7259
rect 9858 7256 9864 7268
rect 8588 7228 9864 7256
rect 8588 7225 8600 7228
rect 8542 7219 8600 7225
rect 9858 7216 9864 7228
rect 9916 7216 9922 7268
rect 12894 7256 12900 7268
rect 11808 7228 12900 7256
rect 2777 7191 2835 7197
rect 2777 7157 2789 7191
rect 2823 7188 2835 7191
rect 2866 7188 2872 7200
rect 2823 7160 2872 7188
rect 2823 7157 2835 7160
rect 2777 7151 2835 7157
rect 2866 7148 2872 7160
rect 2924 7148 2930 7200
rect 3418 7188 3424 7200
rect 3379 7160 3424 7188
rect 3418 7148 3424 7160
rect 3476 7148 3482 7200
rect 3510 7148 3516 7200
rect 3568 7188 3574 7200
rect 3605 7191 3663 7197
rect 3605 7188 3617 7191
rect 3568 7160 3617 7188
rect 3568 7148 3574 7160
rect 3605 7157 3617 7160
rect 3651 7157 3663 7191
rect 4062 7188 4068 7200
rect 4023 7160 4068 7188
rect 3605 7151 3663 7157
rect 4062 7148 4068 7160
rect 4120 7148 4126 7200
rect 4982 7148 4988 7200
rect 5040 7188 5046 7200
rect 5537 7191 5595 7197
rect 5537 7188 5549 7191
rect 5040 7160 5549 7188
rect 5040 7148 5046 7160
rect 5537 7157 5549 7160
rect 5583 7157 5595 7191
rect 6270 7188 6276 7200
rect 6231 7160 6276 7188
rect 5537 7151 5595 7157
rect 6270 7148 6276 7160
rect 6328 7148 6334 7200
rect 6822 7188 6828 7200
rect 6783 7160 6828 7188
rect 6822 7148 6828 7160
rect 6880 7148 6886 7200
rect 9674 7188 9680 7200
rect 9635 7160 9680 7188
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 10778 7188 10784 7200
rect 10739 7160 10784 7188
rect 10778 7148 10784 7160
rect 10836 7148 10842 7200
rect 11241 7191 11299 7197
rect 11241 7157 11253 7191
rect 11287 7188 11299 7191
rect 11330 7188 11336 7200
rect 11287 7160 11336 7188
rect 11287 7157 11299 7160
rect 11241 7151 11299 7157
rect 11330 7148 11336 7160
rect 11388 7148 11394 7200
rect 11698 7148 11704 7200
rect 11756 7188 11762 7200
rect 11808 7197 11836 7228
rect 12894 7216 12900 7228
rect 12952 7216 12958 7268
rect 14553 7259 14611 7265
rect 14553 7225 14565 7259
rect 14599 7256 14611 7259
rect 14844 7256 14872 7296
rect 14912 7293 14924 7296
rect 14958 7324 14970 7327
rect 16482 7324 16488 7336
rect 14958 7296 16488 7324
rect 14958 7293 14970 7296
rect 14912 7287 14970 7293
rect 16482 7284 16488 7296
rect 16540 7284 16546 7336
rect 17773 7327 17831 7333
rect 17773 7324 17785 7327
rect 16592 7296 17785 7324
rect 16592 7256 16620 7296
rect 17773 7293 17785 7296
rect 17819 7324 17831 7327
rect 18414 7324 18420 7336
rect 17819 7296 18420 7324
rect 17819 7293 17831 7296
rect 17773 7287 17831 7293
rect 18414 7284 18420 7296
rect 18472 7284 18478 7336
rect 21545 7327 21603 7333
rect 21545 7293 21557 7327
rect 21591 7324 21603 7327
rect 22002 7324 22008 7336
rect 21591 7296 22008 7324
rect 21591 7293 21603 7296
rect 21545 7287 21603 7293
rect 22002 7284 22008 7296
rect 22060 7324 22066 7336
rect 22572 7324 22600 7355
rect 22646 7352 22652 7364
rect 22704 7352 22710 7404
rect 23474 7392 23480 7404
rect 23435 7364 23480 7392
rect 23474 7352 23480 7364
rect 23532 7392 23538 7404
rect 24118 7392 24124 7404
rect 23532 7364 24124 7392
rect 23532 7352 23538 7364
rect 24118 7352 24124 7364
rect 24176 7352 24182 7404
rect 24302 7392 24308 7404
rect 24263 7364 24308 7392
rect 24302 7352 24308 7364
rect 24360 7392 24366 7404
rect 24360 7364 25452 7392
rect 24360 7352 24366 7364
rect 22060 7296 22600 7324
rect 24029 7327 24087 7333
rect 22060 7284 22066 7296
rect 24029 7293 24041 7327
rect 24075 7324 24087 7327
rect 24762 7324 24768 7336
rect 24075 7296 24768 7324
rect 24075 7293 24087 7296
rect 24029 7287 24087 7293
rect 24762 7284 24768 7296
rect 24820 7284 24826 7336
rect 25314 7324 25320 7336
rect 25275 7296 25320 7324
rect 25314 7284 25320 7296
rect 25372 7284 25378 7336
rect 25424 7324 25452 7364
rect 25573 7327 25631 7333
rect 25573 7324 25585 7327
rect 25424 7296 25585 7324
rect 25573 7293 25585 7296
rect 25619 7293 25631 7327
rect 25573 7287 25631 7293
rect 14599 7228 14872 7256
rect 15028 7228 16620 7256
rect 14599 7225 14611 7228
rect 14553 7219 14611 7225
rect 11793 7191 11851 7197
rect 11793 7188 11805 7191
rect 11756 7160 11805 7188
rect 11756 7148 11762 7160
rect 11793 7157 11805 7160
rect 11839 7157 11851 7191
rect 11793 7151 11851 7157
rect 12250 7148 12256 7200
rect 12308 7188 12314 7200
rect 12437 7191 12495 7197
rect 12437 7188 12449 7191
rect 12308 7160 12449 7188
rect 12308 7148 12314 7160
rect 12437 7157 12449 7160
rect 12483 7157 12495 7191
rect 12802 7188 12808 7200
rect 12763 7160 12808 7188
rect 12437 7151 12495 7157
rect 12802 7148 12808 7160
rect 12860 7188 12866 7200
rect 15028 7188 15056 7228
rect 16666 7216 16672 7268
rect 16724 7256 16730 7268
rect 17310 7256 17316 7268
rect 16724 7228 17316 7256
rect 16724 7216 16730 7228
rect 17310 7216 17316 7228
rect 17368 7216 17374 7268
rect 18138 7216 18144 7268
rect 18196 7256 18202 7268
rect 18509 7259 18567 7265
rect 18509 7256 18521 7259
rect 18196 7228 18521 7256
rect 18196 7216 18202 7228
rect 18509 7225 18521 7228
rect 18555 7225 18567 7259
rect 18509 7219 18567 7225
rect 22278 7216 22284 7268
rect 22336 7256 22342 7268
rect 22373 7259 22431 7265
rect 22373 7256 22385 7259
rect 22336 7228 22385 7256
rect 22336 7216 22342 7228
rect 22373 7225 22385 7228
rect 22419 7225 22431 7259
rect 22373 7219 22431 7225
rect 12860 7160 15056 7188
rect 12860 7148 12866 7160
rect 15838 7148 15844 7200
rect 15896 7188 15902 7200
rect 16025 7191 16083 7197
rect 16025 7188 16037 7191
rect 15896 7160 16037 7188
rect 15896 7148 15902 7160
rect 16025 7157 16037 7160
rect 16071 7157 16083 7191
rect 16942 7188 16948 7200
rect 16903 7160 16948 7188
rect 16025 7151 16083 7157
rect 16942 7148 16948 7160
rect 17000 7148 17006 7200
rect 17862 7148 17868 7200
rect 17920 7188 17926 7200
rect 18049 7191 18107 7197
rect 18049 7188 18061 7191
rect 17920 7160 18061 7188
rect 17920 7148 17926 7160
rect 18049 7157 18061 7160
rect 18095 7157 18107 7191
rect 18049 7151 18107 7157
rect 1104 7098 28888 7120
rect 1104 7046 10982 7098
rect 11034 7046 11046 7098
rect 11098 7046 11110 7098
rect 11162 7046 11174 7098
rect 11226 7046 20982 7098
rect 21034 7046 21046 7098
rect 21098 7046 21110 7098
rect 21162 7046 21174 7098
rect 21226 7046 28888 7098
rect 1104 7024 28888 7046
rect 1670 6984 1676 6996
rect 1631 6956 1676 6984
rect 1670 6944 1676 6956
rect 1728 6944 1734 6996
rect 2317 6987 2375 6993
rect 2317 6953 2329 6987
rect 2363 6953 2375 6987
rect 2317 6947 2375 6953
rect 2332 6916 2360 6947
rect 2406 6944 2412 6996
rect 2464 6984 2470 6996
rect 2685 6987 2743 6993
rect 2685 6984 2697 6987
rect 2464 6956 2697 6984
rect 2464 6944 2470 6956
rect 2685 6953 2697 6956
rect 2731 6984 2743 6987
rect 2774 6984 2780 6996
rect 2731 6956 2780 6984
rect 2731 6953 2743 6956
rect 2685 6947 2743 6953
rect 2774 6944 2780 6956
rect 2832 6944 2838 6996
rect 5721 6987 5779 6993
rect 5721 6953 5733 6987
rect 5767 6984 5779 6987
rect 5810 6984 5816 6996
rect 5767 6956 5816 6984
rect 5767 6953 5779 6956
rect 5721 6947 5779 6953
rect 5810 6944 5816 6956
rect 5868 6984 5874 6996
rect 6822 6984 6828 6996
rect 5868 6956 6828 6984
rect 5868 6944 5874 6956
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 11330 6944 11336 6996
rect 11388 6984 11394 6996
rect 13078 6984 13084 6996
rect 11388 6956 13084 6984
rect 11388 6944 11394 6956
rect 13078 6944 13084 6956
rect 13136 6944 13142 6996
rect 13354 6944 13360 6996
rect 13412 6984 13418 6996
rect 13725 6987 13783 6993
rect 13725 6984 13737 6987
rect 13412 6956 13737 6984
rect 13412 6944 13418 6956
rect 13725 6953 13737 6956
rect 13771 6984 13783 6987
rect 13814 6984 13820 6996
rect 13771 6956 13820 6984
rect 13771 6953 13783 6956
rect 13725 6947 13783 6953
rect 13814 6944 13820 6956
rect 13872 6944 13878 6996
rect 14642 6984 14648 6996
rect 14603 6956 14648 6984
rect 14642 6944 14648 6956
rect 14700 6944 14706 6996
rect 22002 6984 22008 6996
rect 21963 6956 22008 6984
rect 22002 6944 22008 6956
rect 22060 6944 22066 6996
rect 22462 6984 22468 6996
rect 22423 6956 22468 6984
rect 22462 6944 22468 6956
rect 22520 6944 22526 6996
rect 23845 6987 23903 6993
rect 23845 6953 23857 6987
rect 23891 6984 23903 6987
rect 24578 6984 24584 6996
rect 23891 6956 24584 6984
rect 23891 6953 23903 6956
rect 23845 6947 23903 6953
rect 24578 6944 24584 6956
rect 24636 6944 24642 6996
rect 4062 6916 4068 6928
rect 2332 6888 4068 6916
rect 4062 6876 4068 6888
rect 4120 6876 4126 6928
rect 5626 6916 5632 6928
rect 5368 6888 5632 6916
rect 4338 6848 4344 6860
rect 4299 6820 4344 6848
rect 4338 6808 4344 6820
rect 4396 6808 4402 6860
rect 5261 6851 5319 6857
rect 5261 6817 5273 6851
rect 5307 6848 5319 6851
rect 5368 6848 5396 6888
rect 5626 6876 5632 6888
rect 5684 6876 5690 6928
rect 8294 6876 8300 6928
rect 8352 6916 8358 6928
rect 8389 6919 8447 6925
rect 8389 6916 8401 6919
rect 8352 6888 8401 6916
rect 8352 6876 8358 6888
rect 8389 6885 8401 6888
rect 8435 6916 8447 6919
rect 9674 6916 9680 6928
rect 8435 6888 9680 6916
rect 8435 6885 8447 6888
rect 8389 6879 8447 6885
rect 9674 6876 9680 6888
rect 9732 6916 9738 6928
rect 10778 6916 10784 6928
rect 9732 6888 10784 6916
rect 9732 6876 9738 6888
rect 10778 6876 10784 6888
rect 10836 6876 10842 6928
rect 12250 6876 12256 6928
rect 12308 6916 12314 6928
rect 21266 6916 21272 6928
rect 12308 6888 12353 6916
rect 21227 6888 21272 6916
rect 12308 6876 12314 6888
rect 21266 6876 21272 6888
rect 21324 6876 21330 6928
rect 22830 6916 22836 6928
rect 22791 6888 22836 6916
rect 22830 6876 22836 6888
rect 22888 6876 22894 6928
rect 5307 6820 5396 6848
rect 5307 6817 5319 6820
rect 5261 6811 5319 6817
rect 5442 6808 5448 6860
rect 5500 6848 5506 6860
rect 5813 6851 5871 6857
rect 5813 6848 5825 6851
rect 5500 6820 5825 6848
rect 5500 6808 5506 6820
rect 5813 6817 5825 6820
rect 5859 6848 5871 6851
rect 5994 6848 6000 6860
rect 5859 6820 6000 6848
rect 5859 6817 5871 6820
rect 5813 6811 5871 6817
rect 5994 6808 6000 6820
rect 6052 6808 6058 6860
rect 12161 6851 12219 6857
rect 12161 6817 12173 6851
rect 12207 6817 12219 6851
rect 12161 6811 12219 6817
rect 2777 6783 2835 6789
rect 2777 6749 2789 6783
rect 2823 6749 2835 6783
rect 2958 6780 2964 6792
rect 2919 6752 2964 6780
rect 2777 6743 2835 6749
rect 2590 6604 2596 6656
rect 2648 6644 2654 6656
rect 2792 6644 2820 6743
rect 2958 6740 2964 6752
rect 3016 6740 3022 6792
rect 5905 6783 5963 6789
rect 5905 6749 5917 6783
rect 5951 6780 5963 6783
rect 6270 6780 6276 6792
rect 5951 6752 6276 6780
rect 5951 6749 5963 6752
rect 5905 6743 5963 6749
rect 6270 6740 6276 6752
rect 6328 6740 6334 6792
rect 6917 6783 6975 6789
rect 6917 6749 6929 6783
rect 6963 6780 6975 6783
rect 7190 6780 7196 6792
rect 6963 6752 7196 6780
rect 6963 6749 6975 6752
rect 6917 6743 6975 6749
rect 7190 6740 7196 6752
rect 7248 6740 7254 6792
rect 4890 6672 4896 6724
rect 4948 6712 4954 6724
rect 5353 6715 5411 6721
rect 5353 6712 5365 6715
rect 4948 6684 5365 6712
rect 4948 6672 4954 6684
rect 5353 6681 5365 6684
rect 5399 6681 5411 6715
rect 5353 6675 5411 6681
rect 8849 6715 8907 6721
rect 8849 6681 8861 6715
rect 8895 6712 8907 6715
rect 9122 6712 9128 6724
rect 8895 6684 9128 6712
rect 8895 6681 8907 6684
rect 8849 6675 8907 6681
rect 9122 6672 9128 6684
rect 9180 6712 9186 6724
rect 11793 6715 11851 6721
rect 11793 6712 11805 6715
rect 9180 6684 11805 6712
rect 9180 6672 9186 6684
rect 11793 6681 11805 6684
rect 11839 6681 11851 6715
rect 11793 6675 11851 6681
rect 2648 6616 2820 6644
rect 2648 6604 2654 6616
rect 2866 6604 2872 6656
rect 2924 6644 2930 6656
rect 3605 6647 3663 6653
rect 3605 6644 3617 6647
rect 2924 6616 3617 6644
rect 2924 6604 2930 6616
rect 3605 6613 3617 6616
rect 3651 6613 3663 6647
rect 10410 6644 10416 6656
rect 10371 6616 10416 6644
rect 3605 6607 3663 6613
rect 10410 6604 10416 6616
rect 10468 6604 10474 6656
rect 12176 6644 12204 6811
rect 13722 6808 13728 6860
rect 13780 6848 13786 6860
rect 13817 6851 13875 6857
rect 13817 6848 13829 6851
rect 13780 6820 13829 6848
rect 13780 6808 13786 6820
rect 13817 6817 13829 6820
rect 13863 6817 13875 6851
rect 13817 6811 13875 6817
rect 16209 6851 16267 6857
rect 16209 6817 16221 6851
rect 16255 6848 16267 6851
rect 16390 6848 16396 6860
rect 16255 6820 16396 6848
rect 16255 6817 16267 6820
rect 16209 6811 16267 6817
rect 16390 6808 16396 6820
rect 16448 6808 16454 6860
rect 16853 6851 16911 6857
rect 16853 6817 16865 6851
rect 16899 6817 16911 6851
rect 16853 6811 16911 6817
rect 12342 6780 12348 6792
rect 12303 6752 12348 6780
rect 12342 6740 12348 6752
rect 12400 6740 12406 6792
rect 13998 6780 14004 6792
rect 13959 6752 14004 6780
rect 13998 6740 14004 6752
rect 14056 6740 14062 6792
rect 12897 6715 12955 6721
rect 12897 6681 12909 6715
rect 12943 6712 12955 6715
rect 13078 6712 13084 6724
rect 12943 6684 13084 6712
rect 12943 6681 12955 6684
rect 12897 6675 12955 6681
rect 13078 6672 13084 6684
rect 13136 6712 13142 6724
rect 14016 6712 14044 6740
rect 16868 6724 16896 6811
rect 16942 6808 16948 6860
rect 17000 6848 17006 6860
rect 17862 6848 17868 6860
rect 17000 6820 17868 6848
rect 17000 6808 17006 6820
rect 17862 6808 17868 6820
rect 17920 6808 17926 6860
rect 18414 6848 18420 6860
rect 18375 6820 18420 6848
rect 18414 6808 18420 6820
rect 18472 6808 18478 6860
rect 18506 6808 18512 6860
rect 18564 6848 18570 6860
rect 21358 6848 21364 6860
rect 18564 6820 18609 6848
rect 21319 6820 21364 6848
rect 18564 6808 18570 6820
rect 21358 6808 21364 6820
rect 21416 6808 21422 6860
rect 26513 6851 26571 6857
rect 26513 6817 26525 6851
rect 26559 6848 26571 6851
rect 26970 6848 26976 6860
rect 26559 6820 26976 6848
rect 26559 6817 26571 6820
rect 26513 6811 26571 6817
rect 26970 6808 26976 6820
rect 27028 6808 27034 6860
rect 17126 6780 17132 6792
rect 17087 6752 17132 6780
rect 17126 6740 17132 6752
rect 17184 6740 17190 6792
rect 18598 6780 18604 6792
rect 18559 6752 18604 6780
rect 18598 6740 18604 6752
rect 18656 6740 18662 6792
rect 21545 6783 21603 6789
rect 21545 6749 21557 6783
rect 21591 6780 21603 6783
rect 21818 6780 21824 6792
rect 21591 6752 21824 6780
rect 21591 6749 21603 6752
rect 21545 6743 21603 6749
rect 21818 6740 21824 6752
rect 21876 6740 21882 6792
rect 21910 6740 21916 6792
rect 21968 6780 21974 6792
rect 23934 6780 23940 6792
rect 21968 6752 23940 6780
rect 21968 6740 21974 6752
rect 23934 6740 23940 6752
rect 23992 6740 23998 6792
rect 24121 6783 24179 6789
rect 24121 6749 24133 6783
rect 24167 6780 24179 6783
rect 24302 6780 24308 6792
rect 24167 6752 24308 6780
rect 24167 6749 24179 6752
rect 24121 6743 24179 6749
rect 24302 6740 24308 6752
rect 24360 6780 24366 6792
rect 24360 6752 24624 6780
rect 24360 6740 24366 6752
rect 16850 6712 16856 6724
rect 13136 6684 14044 6712
rect 16763 6684 16856 6712
rect 13136 6672 13142 6684
rect 16850 6672 16856 6684
rect 16908 6712 16914 6724
rect 18049 6715 18107 6721
rect 18049 6712 18061 6715
rect 16908 6684 18061 6712
rect 16908 6672 16914 6684
rect 18049 6681 18061 6684
rect 18095 6681 18107 6715
rect 18049 6675 18107 6681
rect 22278 6672 22284 6724
rect 22336 6712 22342 6724
rect 23477 6715 23535 6721
rect 23477 6712 23489 6715
rect 22336 6684 23489 6712
rect 22336 6672 22342 6684
rect 23477 6681 23489 6684
rect 23523 6681 23535 6715
rect 23477 6675 23535 6681
rect 13354 6644 13360 6656
rect 12176 6616 13360 6644
rect 13354 6604 13360 6616
rect 13412 6604 13418 6656
rect 16485 6647 16543 6653
rect 16485 6613 16497 6647
rect 16531 6644 16543 6647
rect 16574 6644 16580 6656
rect 16531 6616 16580 6644
rect 16531 6613 16543 6616
rect 16485 6607 16543 6613
rect 16574 6604 16580 6616
rect 16632 6604 16638 6656
rect 20714 6604 20720 6656
rect 20772 6644 20778 6656
rect 24596 6653 24624 6752
rect 26694 6712 26700 6724
rect 26655 6684 26700 6712
rect 26694 6672 26700 6684
rect 26752 6672 26758 6724
rect 20901 6647 20959 6653
rect 20901 6644 20913 6647
rect 20772 6616 20913 6644
rect 20772 6604 20778 6616
rect 20901 6613 20913 6616
rect 20947 6613 20959 6647
rect 20901 6607 20959 6613
rect 24581 6647 24639 6653
rect 24581 6613 24593 6647
rect 24627 6644 24639 6647
rect 25038 6644 25044 6656
rect 24627 6616 25044 6644
rect 24627 6613 24639 6616
rect 24581 6607 24639 6613
rect 25038 6604 25044 6616
rect 25096 6644 25102 6656
rect 25317 6647 25375 6653
rect 25317 6644 25329 6647
rect 25096 6616 25329 6644
rect 25096 6604 25102 6616
rect 25317 6613 25329 6616
rect 25363 6613 25375 6647
rect 25317 6607 25375 6613
rect 1104 6554 28888 6576
rect 1104 6502 5982 6554
rect 6034 6502 6046 6554
rect 6098 6502 6110 6554
rect 6162 6502 6174 6554
rect 6226 6502 15982 6554
rect 16034 6502 16046 6554
rect 16098 6502 16110 6554
rect 16162 6502 16174 6554
rect 16226 6502 25982 6554
rect 26034 6502 26046 6554
rect 26098 6502 26110 6554
rect 26162 6502 26174 6554
rect 26226 6502 28888 6554
rect 1104 6480 28888 6502
rect 1486 6400 1492 6452
rect 1544 6440 1550 6452
rect 1581 6443 1639 6449
rect 1581 6440 1593 6443
rect 1544 6412 1593 6440
rect 1544 6400 1550 6412
rect 1581 6409 1593 6412
rect 1627 6409 1639 6443
rect 2038 6440 2044 6452
rect 1999 6412 2044 6440
rect 1581 6403 1639 6409
rect 2038 6400 2044 6412
rect 2096 6400 2102 6452
rect 2590 6400 2596 6452
rect 2648 6440 2654 6452
rect 2685 6443 2743 6449
rect 2685 6440 2697 6443
rect 2648 6412 2697 6440
rect 2648 6400 2654 6412
rect 2685 6409 2697 6412
rect 2731 6409 2743 6443
rect 2685 6403 2743 6409
rect 2774 6400 2780 6452
rect 2832 6440 2838 6452
rect 3053 6443 3111 6449
rect 3053 6440 3065 6443
rect 2832 6412 3065 6440
rect 2832 6400 2838 6412
rect 3053 6409 3065 6412
rect 3099 6409 3111 6443
rect 5442 6440 5448 6452
rect 5403 6412 5448 6440
rect 3053 6403 3111 6409
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 5810 6440 5816 6452
rect 5771 6412 5816 6440
rect 5810 6400 5816 6412
rect 5868 6400 5874 6452
rect 6181 6443 6239 6449
rect 6181 6409 6193 6443
rect 6227 6440 6239 6443
rect 6270 6440 6276 6452
rect 6227 6412 6276 6440
rect 6227 6409 6239 6412
rect 6181 6403 6239 6409
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 6546 6440 6552 6452
rect 6507 6412 6552 6440
rect 6546 6400 6552 6412
rect 6604 6440 6610 6452
rect 6604 6412 7328 6440
rect 6604 6400 6610 6412
rect 1670 6332 1676 6384
rect 1728 6372 1734 6384
rect 2317 6375 2375 6381
rect 2317 6372 2329 6375
rect 1728 6344 2329 6372
rect 1728 6332 1734 6344
rect 2317 6341 2329 6344
rect 2363 6372 2375 6375
rect 2958 6372 2964 6384
rect 2363 6344 2964 6372
rect 2363 6341 2375 6344
rect 2317 6335 2375 6341
rect 2958 6332 2964 6344
rect 3016 6332 3022 6384
rect 6546 6264 6552 6316
rect 6604 6304 6610 6316
rect 6730 6304 6736 6316
rect 6604 6276 6736 6304
rect 6604 6264 6610 6276
rect 6730 6264 6736 6276
rect 6788 6264 6794 6316
rect 7300 6313 7328 6412
rect 9858 6400 9864 6452
rect 9916 6440 9922 6452
rect 10137 6443 10195 6449
rect 10137 6440 10149 6443
rect 9916 6412 10149 6440
rect 9916 6400 9922 6412
rect 10137 6409 10149 6412
rect 10183 6440 10195 6443
rect 12250 6440 12256 6452
rect 10183 6412 10824 6440
rect 12211 6412 12256 6440
rect 10183 6409 10195 6412
rect 10137 6403 10195 6409
rect 8294 6332 8300 6384
rect 8352 6372 8358 6384
rect 8757 6375 8815 6381
rect 8757 6372 8769 6375
rect 8352 6344 8769 6372
rect 8352 6332 8358 6344
rect 8757 6341 8769 6344
rect 8803 6341 8815 6375
rect 10321 6375 10379 6381
rect 10321 6372 10333 6375
rect 8757 6335 8815 6341
rect 9232 6344 10333 6372
rect 7285 6307 7343 6313
rect 7285 6273 7297 6307
rect 7331 6273 7343 6307
rect 7285 6267 7343 6273
rect 7469 6307 7527 6313
rect 7469 6273 7481 6307
rect 7515 6304 7527 6307
rect 7558 6304 7564 6316
rect 7515 6276 7564 6304
rect 7515 6273 7527 6276
rect 7469 6267 7527 6273
rect 7558 6264 7564 6276
rect 7616 6304 7622 6316
rect 7837 6307 7895 6313
rect 7837 6304 7849 6307
rect 7616 6276 7849 6304
rect 7616 6264 7622 6276
rect 7837 6273 7849 6276
rect 7883 6273 7895 6307
rect 7837 6267 7895 6273
rect 8846 6264 8852 6316
rect 8904 6304 8910 6316
rect 9232 6313 9260 6344
rect 10321 6341 10333 6344
rect 10367 6341 10379 6375
rect 10796 6372 10824 6412
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 12713 6443 12771 6449
rect 12713 6409 12725 6443
rect 12759 6440 12771 6443
rect 13354 6440 13360 6452
rect 12759 6412 13360 6440
rect 12759 6409 12771 6412
rect 12713 6403 12771 6409
rect 13354 6400 13360 6412
rect 13412 6400 13418 6452
rect 13814 6440 13820 6452
rect 13775 6412 13820 6440
rect 13814 6400 13820 6412
rect 13872 6400 13878 6452
rect 18506 6440 18512 6452
rect 18467 6412 18512 6440
rect 18506 6400 18512 6412
rect 18564 6400 18570 6452
rect 21266 6400 21272 6452
rect 21324 6440 21330 6452
rect 21729 6443 21787 6449
rect 21729 6440 21741 6443
rect 21324 6412 21741 6440
rect 21324 6400 21330 6412
rect 21729 6409 21741 6412
rect 21775 6409 21787 6443
rect 21729 6403 21787 6409
rect 11793 6375 11851 6381
rect 11793 6372 11805 6375
rect 10796 6344 11805 6372
rect 10321 6335 10379 6341
rect 9217 6307 9275 6313
rect 9217 6304 9229 6307
rect 8904 6276 9229 6304
rect 8904 6264 8910 6276
rect 9217 6273 9229 6276
rect 9263 6273 9275 6307
rect 9217 6267 9275 6273
rect 9309 6307 9367 6313
rect 9309 6273 9321 6307
rect 9355 6304 9367 6307
rect 9582 6304 9588 6316
rect 9355 6276 9588 6304
rect 9355 6273 9367 6276
rect 9309 6267 9367 6273
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 2038 6236 2044 6248
rect 1443 6208 2044 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 2038 6196 2044 6208
rect 2096 6196 2102 6248
rect 7190 6236 7196 6248
rect 7151 6208 7196 6236
rect 7190 6196 7196 6208
rect 7248 6196 7254 6248
rect 8665 6239 8723 6245
rect 8665 6205 8677 6239
rect 8711 6236 8723 6239
rect 9324 6236 9352 6267
rect 9582 6264 9588 6276
rect 9640 6264 9646 6316
rect 10410 6264 10416 6316
rect 10468 6304 10474 6316
rect 10686 6304 10692 6316
rect 10468 6276 10692 6304
rect 10468 6264 10474 6276
rect 10686 6264 10692 6276
rect 10744 6304 10750 6316
rect 10888 6313 10916 6344
rect 11793 6341 11805 6344
rect 11839 6372 11851 6375
rect 12342 6372 12348 6384
rect 11839 6344 12348 6372
rect 11839 6341 11851 6344
rect 11793 6335 11851 6341
rect 12342 6332 12348 6344
rect 12400 6332 12406 6384
rect 13449 6375 13507 6381
rect 13449 6341 13461 6375
rect 13495 6372 13507 6375
rect 13722 6372 13728 6384
rect 13495 6344 13728 6372
rect 13495 6341 13507 6344
rect 13449 6335 13507 6341
rect 13722 6332 13728 6344
rect 13780 6332 13786 6384
rect 17586 6332 17592 6384
rect 17644 6372 17650 6384
rect 17865 6375 17923 6381
rect 17865 6372 17877 6375
rect 17644 6344 17877 6372
rect 17644 6332 17650 6344
rect 17865 6341 17877 6344
rect 17911 6372 17923 6375
rect 18598 6372 18604 6384
rect 17911 6344 18604 6372
rect 17911 6341 17923 6344
rect 17865 6335 17923 6341
rect 18598 6332 18604 6344
rect 18656 6332 18662 6384
rect 21358 6372 21364 6384
rect 21319 6344 21364 6372
rect 21358 6332 21364 6344
rect 21416 6332 21422 6384
rect 10781 6307 10839 6313
rect 10781 6304 10793 6307
rect 10744 6276 10793 6304
rect 10744 6264 10750 6276
rect 10781 6273 10793 6276
rect 10827 6273 10839 6307
rect 10781 6267 10839 6273
rect 10873 6307 10931 6313
rect 10873 6273 10885 6307
rect 10919 6273 10931 6307
rect 10873 6267 10931 6273
rect 16390 6264 16396 6316
rect 16448 6304 16454 6316
rect 16577 6307 16635 6313
rect 16577 6304 16589 6307
rect 16448 6276 16589 6304
rect 16448 6264 16454 6276
rect 16577 6273 16589 6276
rect 16623 6273 16635 6307
rect 16577 6267 16635 6273
rect 16669 6307 16727 6313
rect 16669 6273 16681 6307
rect 16715 6273 16727 6307
rect 16669 6267 16727 6273
rect 18049 6307 18107 6313
rect 18049 6273 18061 6307
rect 18095 6304 18107 6307
rect 18414 6304 18420 6316
rect 18095 6276 18420 6304
rect 18095 6273 18107 6276
rect 18049 6267 18107 6273
rect 15838 6236 15844 6248
rect 8711 6208 9352 6236
rect 15751 6208 15844 6236
rect 8711 6205 8723 6208
rect 8665 6199 8723 6205
rect 15838 6196 15844 6208
rect 15896 6236 15902 6248
rect 16684 6236 16712 6267
rect 18414 6264 18420 6276
rect 18472 6304 18478 6316
rect 18877 6307 18935 6313
rect 18877 6304 18889 6307
rect 18472 6276 18889 6304
rect 18472 6264 18478 6276
rect 18877 6273 18889 6276
rect 18923 6273 18935 6307
rect 21744 6304 21772 6403
rect 21818 6400 21824 6452
rect 21876 6440 21882 6452
rect 22373 6443 22431 6449
rect 22373 6440 22385 6443
rect 21876 6412 22385 6440
rect 21876 6400 21882 6412
rect 22373 6409 22385 6412
rect 22419 6409 22431 6443
rect 22373 6403 22431 6409
rect 23477 6443 23535 6449
rect 23477 6409 23489 6443
rect 23523 6440 23535 6443
rect 24302 6440 24308 6452
rect 23523 6412 24308 6440
rect 23523 6409 23535 6412
rect 23477 6403 23535 6409
rect 24302 6400 24308 6412
rect 24360 6400 24366 6452
rect 26970 6440 26976 6452
rect 26931 6412 26976 6440
rect 26970 6400 26976 6412
rect 27028 6400 27034 6452
rect 23934 6372 23940 6384
rect 23895 6344 23940 6372
rect 23934 6332 23940 6344
rect 23992 6332 23998 6384
rect 21913 6307 21971 6313
rect 21913 6304 21925 6307
rect 21744 6276 21925 6304
rect 18877 6267 18935 6273
rect 21913 6273 21925 6276
rect 21959 6273 21971 6307
rect 21913 6267 21971 6273
rect 23566 6264 23572 6316
rect 23624 6304 23630 6316
rect 24305 6307 24363 6313
rect 24305 6304 24317 6307
rect 23624 6276 24317 6304
rect 23624 6264 23630 6276
rect 24305 6273 24317 6276
rect 24351 6304 24363 6307
rect 24578 6304 24584 6316
rect 24351 6276 24584 6304
rect 24351 6273 24363 6276
rect 24305 6267 24363 6273
rect 24578 6264 24584 6276
rect 24636 6264 24642 6316
rect 17126 6236 17132 6248
rect 15896 6208 17132 6236
rect 15896 6196 15902 6208
rect 17126 6196 17132 6208
rect 17184 6196 17190 6248
rect 19702 6236 19708 6248
rect 19663 6208 19708 6236
rect 19702 6196 19708 6208
rect 19760 6196 19766 6248
rect 26421 6239 26479 6245
rect 26421 6205 26433 6239
rect 26467 6205 26479 6239
rect 26421 6199 26479 6205
rect 9122 6168 9128 6180
rect 9083 6140 9128 6168
rect 9122 6128 9128 6140
rect 9180 6128 9186 6180
rect 9861 6171 9919 6177
rect 9861 6137 9873 6171
rect 9907 6168 9919 6171
rect 10410 6168 10416 6180
rect 9907 6140 10416 6168
rect 9907 6137 9919 6140
rect 9861 6131 9919 6137
rect 10410 6128 10416 6140
rect 10468 6168 10474 6180
rect 10689 6171 10747 6177
rect 10689 6168 10701 6171
rect 10468 6140 10701 6168
rect 10468 6128 10474 6140
rect 10689 6137 10701 6140
rect 10735 6137 10747 6171
rect 10689 6131 10747 6137
rect 15657 6171 15715 6177
rect 15657 6137 15669 6171
rect 15703 6168 15715 6171
rect 16485 6171 16543 6177
rect 16485 6168 16497 6171
rect 15703 6140 16497 6168
rect 15703 6137 15715 6140
rect 15657 6131 15715 6137
rect 16485 6137 16497 6140
rect 16531 6168 16543 6171
rect 17034 6168 17040 6180
rect 16531 6140 17040 6168
rect 16531 6137 16543 6140
rect 16485 6131 16543 6137
rect 17034 6128 17040 6140
rect 17092 6128 17098 6180
rect 19613 6171 19671 6177
rect 19613 6137 19625 6171
rect 19659 6168 19671 6171
rect 19972 6171 20030 6177
rect 19972 6168 19984 6171
rect 19659 6140 19984 6168
rect 19659 6137 19671 6140
rect 19613 6131 19671 6137
rect 19972 6137 19984 6140
rect 20018 6168 20030 6171
rect 21818 6168 21824 6180
rect 20018 6140 21824 6168
rect 20018 6137 20030 6140
rect 19972 6131 20030 6137
rect 21818 6128 21824 6140
rect 21876 6128 21882 6180
rect 26234 6168 26240 6180
rect 26195 6140 26240 6168
rect 26234 6128 26240 6140
rect 26292 6168 26298 6180
rect 26436 6168 26464 6199
rect 26292 6140 26464 6168
rect 26292 6128 26298 6140
rect 6822 6100 6828 6112
rect 6783 6072 6828 6100
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 13998 6060 14004 6112
rect 14056 6100 14062 6112
rect 14093 6103 14151 6109
rect 14093 6100 14105 6103
rect 14056 6072 14105 6100
rect 14056 6060 14062 6072
rect 14093 6069 14105 6072
rect 14139 6069 14151 6103
rect 14093 6063 14151 6069
rect 15194 6060 15200 6112
rect 15252 6100 15258 6112
rect 15841 6103 15899 6109
rect 15841 6100 15853 6103
rect 15252 6072 15853 6100
rect 15252 6060 15258 6072
rect 15841 6069 15853 6072
rect 15887 6100 15899 6103
rect 15933 6103 15991 6109
rect 15933 6100 15945 6103
rect 15887 6072 15945 6100
rect 15887 6069 15899 6072
rect 15841 6063 15899 6069
rect 15933 6069 15945 6072
rect 15979 6069 15991 6103
rect 16114 6100 16120 6112
rect 16075 6072 16120 6100
rect 15933 6063 15991 6069
rect 16114 6060 16120 6072
rect 16172 6060 16178 6112
rect 21085 6103 21143 6109
rect 21085 6069 21097 6103
rect 21131 6100 21143 6103
rect 21266 6100 21272 6112
rect 21131 6072 21272 6100
rect 21131 6069 21143 6072
rect 21085 6063 21143 6069
rect 21266 6060 21272 6072
rect 21324 6060 21330 6112
rect 26602 6100 26608 6112
rect 26563 6072 26608 6100
rect 26602 6060 26608 6072
rect 26660 6060 26666 6112
rect 1104 6010 28888 6032
rect 1104 5958 10982 6010
rect 11034 5958 11046 6010
rect 11098 5958 11110 6010
rect 11162 5958 11174 6010
rect 11226 5958 20982 6010
rect 21034 5958 21046 6010
rect 21098 5958 21110 6010
rect 21162 5958 21174 6010
rect 21226 5958 28888 6010
rect 1104 5936 28888 5958
rect 6917 5899 6975 5905
rect 6917 5865 6929 5899
rect 6963 5896 6975 5899
rect 7190 5896 7196 5908
rect 6963 5868 7196 5896
rect 6963 5865 6975 5868
rect 6917 5859 6975 5865
rect 7190 5856 7196 5868
rect 7248 5856 7254 5908
rect 8846 5896 8852 5908
rect 8807 5868 8852 5896
rect 8846 5856 8852 5868
rect 8904 5856 8910 5908
rect 10410 5896 10416 5908
rect 10371 5868 10416 5896
rect 10410 5856 10416 5868
rect 10468 5856 10474 5908
rect 10502 5856 10508 5908
rect 10560 5896 10566 5908
rect 10873 5899 10931 5905
rect 10873 5896 10885 5899
rect 10560 5868 10885 5896
rect 10560 5856 10566 5868
rect 10873 5865 10885 5868
rect 10919 5896 10931 5899
rect 11977 5899 12035 5905
rect 11977 5896 11989 5899
rect 10919 5868 11989 5896
rect 10919 5865 10931 5868
rect 10873 5859 10931 5865
rect 11977 5865 11989 5868
rect 12023 5865 12035 5899
rect 11977 5859 12035 5865
rect 15838 5856 15844 5908
rect 15896 5896 15902 5908
rect 15933 5899 15991 5905
rect 15933 5896 15945 5899
rect 15896 5868 15945 5896
rect 15896 5856 15902 5868
rect 15933 5865 15945 5868
rect 15979 5896 15991 5899
rect 16114 5896 16120 5908
rect 15979 5868 16120 5896
rect 15979 5865 15991 5868
rect 15933 5859 15991 5865
rect 16114 5856 16120 5868
rect 16172 5856 16178 5908
rect 16850 5896 16856 5908
rect 16811 5868 16856 5896
rect 16850 5856 16856 5868
rect 16908 5856 16914 5908
rect 17034 5896 17040 5908
rect 16995 5868 17040 5896
rect 17034 5856 17040 5868
rect 17092 5856 17098 5908
rect 17402 5896 17408 5908
rect 17363 5868 17408 5896
rect 17402 5856 17408 5868
rect 17460 5856 17466 5908
rect 2032 5831 2090 5837
rect 2032 5797 2044 5831
rect 2078 5828 2090 5831
rect 2314 5828 2320 5840
rect 2078 5800 2320 5828
rect 2078 5797 2090 5800
rect 2032 5791 2090 5797
rect 2314 5788 2320 5800
rect 2372 5828 2378 5840
rect 2866 5828 2872 5840
rect 2372 5800 2872 5828
rect 2372 5788 2378 5800
rect 2866 5788 2872 5800
rect 2924 5788 2930 5840
rect 4798 5788 4804 5840
rect 4856 5828 4862 5840
rect 5046 5831 5104 5837
rect 5046 5828 5058 5831
rect 4856 5800 5058 5828
rect 4856 5788 4862 5800
rect 5046 5797 5058 5800
rect 5092 5797 5104 5831
rect 5046 5791 5104 5797
rect 5166 5788 5172 5840
rect 5224 5788 5230 5840
rect 7377 5831 7435 5837
rect 7377 5797 7389 5831
rect 7423 5828 7435 5831
rect 7926 5828 7932 5840
rect 7423 5800 7932 5828
rect 7423 5797 7435 5800
rect 7377 5791 7435 5797
rect 7926 5788 7932 5800
rect 7984 5788 7990 5840
rect 10226 5788 10232 5840
rect 10284 5828 10290 5840
rect 10781 5831 10839 5837
rect 10781 5828 10793 5831
rect 10284 5800 10793 5828
rect 10284 5788 10290 5800
rect 10781 5797 10793 5800
rect 10827 5797 10839 5831
rect 10781 5791 10839 5797
rect 16577 5831 16635 5837
rect 16577 5797 16589 5831
rect 16623 5828 16635 5831
rect 16942 5828 16948 5840
rect 16623 5800 16948 5828
rect 16623 5797 16635 5800
rect 16577 5791 16635 5797
rect 16942 5788 16948 5800
rect 17000 5788 17006 5840
rect 19702 5788 19708 5840
rect 19760 5828 19766 5840
rect 19797 5831 19855 5837
rect 19797 5828 19809 5831
rect 19760 5800 19809 5828
rect 19760 5788 19766 5800
rect 19797 5797 19809 5800
rect 19843 5828 19855 5831
rect 22186 5828 22192 5840
rect 19843 5800 22192 5828
rect 19843 5797 19855 5800
rect 19797 5791 19855 5797
rect 22186 5788 22192 5800
rect 22244 5788 22250 5840
rect 5184 5760 5212 5788
rect 4816 5732 5212 5760
rect 7469 5763 7527 5769
rect 1762 5692 1768 5704
rect 1723 5664 1768 5692
rect 1762 5652 1768 5664
rect 1820 5652 1826 5704
rect 4816 5701 4844 5732
rect 7469 5729 7481 5763
rect 7515 5760 7527 5763
rect 7650 5760 7656 5772
rect 7515 5732 7656 5760
rect 7515 5729 7527 5732
rect 7469 5723 7527 5729
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 11974 5720 11980 5772
rect 12032 5760 12038 5772
rect 12342 5760 12348 5772
rect 12032 5732 12348 5760
rect 12032 5720 12038 5732
rect 12342 5720 12348 5732
rect 12400 5720 12406 5772
rect 15841 5763 15899 5769
rect 15841 5729 15853 5763
rect 15887 5760 15899 5763
rect 16482 5760 16488 5772
rect 15887 5732 16488 5760
rect 15887 5729 15899 5732
rect 15841 5723 15899 5729
rect 16482 5720 16488 5732
rect 16540 5720 16546 5772
rect 21174 5720 21180 5772
rect 21232 5760 21238 5772
rect 21269 5763 21327 5769
rect 21269 5760 21281 5763
rect 21232 5732 21281 5760
rect 21232 5720 21238 5732
rect 21269 5729 21281 5732
rect 21315 5729 21327 5763
rect 26510 5760 26516 5772
rect 26423 5732 26516 5760
rect 21269 5723 21327 5729
rect 26510 5720 26516 5732
rect 26568 5760 26574 5772
rect 26970 5760 26976 5772
rect 26568 5732 26976 5760
rect 26568 5720 26574 5732
rect 26970 5720 26976 5732
rect 27028 5720 27034 5772
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5661 4859 5695
rect 7558 5692 7564 5704
rect 7519 5664 7564 5692
rect 4801 5655 4859 5661
rect 7558 5652 7564 5664
rect 7616 5652 7622 5704
rect 10965 5695 11023 5701
rect 10965 5661 10977 5695
rect 11011 5692 11023 5695
rect 11330 5692 11336 5704
rect 11011 5664 11336 5692
rect 11011 5661 11023 5664
rect 10965 5655 11023 5661
rect 11330 5652 11336 5664
rect 11388 5652 11394 5704
rect 12066 5652 12072 5704
rect 12124 5692 12130 5704
rect 12437 5695 12495 5701
rect 12437 5692 12449 5695
rect 12124 5664 12449 5692
rect 12124 5652 12130 5664
rect 12437 5661 12449 5664
rect 12483 5661 12495 5695
rect 12437 5655 12495 5661
rect 12621 5695 12679 5701
rect 12621 5661 12633 5695
rect 12667 5692 12679 5695
rect 16117 5695 16175 5701
rect 12667 5664 12940 5692
rect 12667 5661 12679 5664
rect 12621 5655 12679 5661
rect 12912 5568 12940 5664
rect 16117 5661 16129 5695
rect 16163 5692 16175 5695
rect 16298 5692 16304 5704
rect 16163 5664 16304 5692
rect 16163 5661 16175 5664
rect 16117 5655 16175 5661
rect 16298 5652 16304 5664
rect 16356 5652 16362 5704
rect 17494 5692 17500 5704
rect 17455 5664 17500 5692
rect 17494 5652 17500 5664
rect 17552 5652 17558 5704
rect 17586 5652 17592 5704
rect 17644 5692 17650 5704
rect 17644 5664 17689 5692
rect 17644 5652 17650 5664
rect 20254 5652 20260 5704
rect 20312 5692 20318 5704
rect 21361 5695 21419 5701
rect 21361 5692 21373 5695
rect 20312 5664 21373 5692
rect 20312 5652 20318 5664
rect 21361 5661 21373 5664
rect 21407 5661 21419 5695
rect 21361 5655 21419 5661
rect 21545 5695 21603 5701
rect 21545 5661 21557 5695
rect 21591 5692 21603 5695
rect 21818 5692 21824 5704
rect 21591 5664 21824 5692
rect 21591 5661 21603 5664
rect 21545 5655 21603 5661
rect 21818 5652 21824 5664
rect 21876 5652 21882 5704
rect 3142 5556 3148 5568
rect 3103 5528 3148 5556
rect 3142 5516 3148 5528
rect 3200 5516 3206 5568
rect 6181 5559 6239 5565
rect 6181 5525 6193 5559
rect 6227 5556 6239 5559
rect 6270 5556 6276 5568
rect 6227 5528 6276 5556
rect 6227 5525 6239 5528
rect 6181 5519 6239 5525
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 7006 5556 7012 5568
rect 6967 5528 7012 5556
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 11422 5556 11428 5568
rect 11383 5528 11428 5556
rect 11422 5516 11428 5528
rect 11480 5516 11486 5568
rect 12894 5516 12900 5568
rect 12952 5556 12958 5568
rect 12989 5559 13047 5565
rect 12989 5556 13001 5559
rect 12952 5528 13001 5556
rect 12952 5516 12958 5528
rect 12989 5525 13001 5528
rect 13035 5525 13047 5559
rect 13354 5556 13360 5568
rect 13315 5528 13360 5556
rect 12989 5519 13047 5525
rect 13354 5516 13360 5528
rect 13412 5516 13418 5568
rect 15470 5556 15476 5568
rect 15431 5528 15476 5556
rect 15470 5516 15476 5528
rect 15528 5516 15534 5568
rect 20533 5559 20591 5565
rect 20533 5525 20545 5559
rect 20579 5556 20591 5559
rect 20898 5556 20904 5568
rect 20579 5528 20904 5556
rect 20579 5525 20591 5528
rect 20533 5519 20591 5525
rect 20898 5516 20904 5528
rect 20956 5516 20962 5568
rect 23658 5556 23664 5568
rect 23619 5528 23664 5556
rect 23658 5516 23664 5528
rect 23716 5516 23722 5568
rect 26697 5559 26755 5565
rect 26697 5525 26709 5559
rect 26743 5556 26755 5559
rect 26786 5556 26792 5568
rect 26743 5528 26792 5556
rect 26743 5525 26755 5528
rect 26697 5519 26755 5525
rect 26786 5516 26792 5528
rect 26844 5516 26850 5568
rect 1104 5466 28888 5488
rect 1104 5414 5982 5466
rect 6034 5414 6046 5466
rect 6098 5414 6110 5466
rect 6162 5414 6174 5466
rect 6226 5414 15982 5466
rect 16034 5414 16046 5466
rect 16098 5414 16110 5466
rect 16162 5414 16174 5466
rect 16226 5414 25982 5466
rect 26034 5414 26046 5466
rect 26098 5414 26110 5466
rect 26162 5414 26174 5466
rect 26226 5414 28888 5466
rect 1104 5392 28888 5414
rect 1578 5352 1584 5364
rect 1539 5324 1584 5352
rect 1578 5312 1584 5324
rect 1636 5312 1642 5364
rect 2314 5352 2320 5364
rect 2275 5324 2320 5352
rect 2314 5312 2320 5324
rect 2372 5312 2378 5364
rect 2869 5355 2927 5361
rect 2869 5321 2881 5355
rect 2915 5352 2927 5355
rect 3142 5352 3148 5364
rect 2915 5324 3148 5352
rect 2915 5321 2927 5324
rect 2869 5315 2927 5321
rect 3142 5312 3148 5324
rect 3200 5312 3206 5364
rect 5166 5352 5172 5364
rect 5127 5324 5172 5352
rect 5166 5312 5172 5324
rect 5224 5312 5230 5364
rect 6270 5352 6276 5364
rect 6231 5324 6276 5352
rect 6270 5312 6276 5324
rect 6328 5312 6334 5364
rect 7926 5352 7932 5364
rect 7887 5324 7932 5352
rect 7926 5312 7932 5324
rect 7984 5312 7990 5364
rect 9769 5355 9827 5361
rect 9769 5321 9781 5355
rect 9815 5352 9827 5355
rect 10502 5352 10508 5364
rect 9815 5324 10508 5352
rect 9815 5321 9827 5324
rect 9769 5315 9827 5321
rect 10502 5312 10508 5324
rect 10560 5312 10566 5364
rect 10686 5352 10692 5364
rect 10647 5324 10692 5352
rect 10686 5312 10692 5324
rect 10744 5312 10750 5364
rect 12066 5352 12072 5364
rect 12027 5324 12072 5352
rect 12066 5312 12072 5324
rect 12124 5312 12130 5364
rect 13998 5352 14004 5364
rect 13959 5324 14004 5352
rect 13998 5312 14004 5324
rect 14056 5312 14062 5364
rect 16209 5355 16267 5361
rect 16209 5321 16221 5355
rect 16255 5352 16267 5355
rect 16298 5352 16304 5364
rect 16255 5324 16304 5352
rect 16255 5321 16267 5324
rect 16209 5315 16267 5321
rect 16298 5312 16304 5324
rect 16356 5312 16362 5364
rect 16574 5352 16580 5364
rect 16535 5324 16580 5352
rect 16574 5312 16580 5324
rect 16632 5312 16638 5364
rect 17494 5352 17500 5364
rect 17455 5324 17500 5352
rect 17494 5312 17500 5324
rect 17552 5312 17558 5364
rect 17586 5312 17592 5364
rect 17644 5352 17650 5364
rect 17773 5355 17831 5361
rect 17773 5352 17785 5355
rect 17644 5324 17785 5352
rect 17644 5312 17650 5324
rect 17773 5321 17785 5324
rect 17819 5321 17831 5355
rect 17773 5315 17831 5321
rect 21174 5312 21180 5364
rect 21232 5352 21238 5364
rect 21453 5355 21511 5361
rect 21453 5352 21465 5355
rect 21232 5324 21465 5352
rect 21232 5312 21238 5324
rect 21453 5321 21465 5324
rect 21499 5321 21511 5355
rect 25038 5352 25044 5364
rect 24999 5324 25044 5352
rect 21453 5315 21511 5321
rect 25038 5312 25044 5324
rect 25096 5312 25102 5364
rect 26970 5352 26976 5364
rect 26931 5324 26976 5352
rect 26970 5312 26976 5324
rect 27028 5312 27034 5364
rect 6288 5284 6316 5312
rect 6288 5256 7420 5284
rect 2038 5216 2044 5228
rect 1412 5188 2044 5216
rect 1412 5157 1440 5188
rect 2038 5176 2044 5188
rect 2096 5176 2102 5228
rect 6638 5216 6644 5228
rect 6599 5188 6644 5216
rect 6638 5176 6644 5188
rect 6696 5176 6702 5228
rect 7006 5176 7012 5228
rect 7064 5216 7070 5228
rect 7392 5225 7420 5256
rect 10226 5244 10232 5296
rect 10284 5284 10290 5296
rect 10413 5287 10471 5293
rect 10413 5284 10425 5287
rect 10284 5256 10425 5284
rect 10284 5244 10290 5256
rect 10413 5253 10425 5256
rect 10459 5253 10471 5287
rect 10413 5247 10471 5253
rect 17129 5287 17187 5293
rect 17129 5253 17141 5287
rect 17175 5284 17187 5287
rect 17402 5284 17408 5296
rect 17175 5256 17408 5284
rect 17175 5253 17187 5256
rect 17129 5247 17187 5253
rect 17402 5244 17408 5256
rect 17460 5244 17466 5296
rect 20254 5284 20260 5296
rect 20215 5256 20260 5284
rect 20254 5244 20260 5256
rect 20312 5244 20318 5296
rect 20622 5244 20628 5296
rect 20680 5284 20686 5296
rect 21358 5284 21364 5296
rect 20680 5256 21364 5284
rect 20680 5244 20686 5256
rect 21358 5244 21364 5256
rect 21416 5244 21422 5296
rect 7285 5219 7343 5225
rect 7285 5216 7297 5219
rect 7064 5188 7297 5216
rect 7064 5176 7070 5188
rect 7285 5185 7297 5188
rect 7331 5185 7343 5219
rect 7285 5179 7343 5185
rect 7377 5219 7435 5225
rect 7377 5185 7389 5219
rect 7423 5216 7435 5219
rect 7466 5216 7472 5228
rect 7423 5188 7472 5216
rect 7423 5185 7435 5188
rect 7377 5179 7435 5185
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 10137 5219 10195 5225
rect 10137 5185 10149 5219
rect 10183 5216 10195 5219
rect 10778 5216 10784 5228
rect 10183 5188 10784 5216
rect 10183 5185 10195 5188
rect 10137 5179 10195 5185
rect 10778 5176 10784 5188
rect 10836 5216 10842 5228
rect 11330 5216 11336 5228
rect 10836 5188 11336 5216
rect 10836 5176 10842 5188
rect 11330 5176 11336 5188
rect 11388 5176 11394 5228
rect 14642 5176 14648 5228
rect 14700 5216 14706 5228
rect 14829 5219 14887 5225
rect 14829 5216 14841 5219
rect 14700 5188 14841 5216
rect 14700 5176 14706 5188
rect 14829 5185 14841 5188
rect 14875 5185 14887 5219
rect 20898 5216 20904 5228
rect 20859 5188 20904 5216
rect 14829 5179 14887 5185
rect 20898 5176 20904 5188
rect 20956 5176 20962 5228
rect 21085 5219 21143 5225
rect 21085 5185 21097 5219
rect 21131 5216 21143 5219
rect 21266 5216 21272 5228
rect 21131 5188 21272 5216
rect 21131 5185 21143 5188
rect 21085 5179 21143 5185
rect 21266 5176 21272 5188
rect 21324 5176 21330 5228
rect 22186 5176 22192 5228
rect 22244 5216 22250 5228
rect 23658 5216 23664 5228
rect 22244 5188 23664 5216
rect 22244 5176 22250 5188
rect 23658 5176 23664 5188
rect 23716 5176 23722 5228
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5117 1455 5151
rect 1397 5111 1455 5117
rect 2961 5151 3019 5157
rect 2961 5117 2973 5151
rect 3007 5148 3019 5151
rect 3602 5148 3608 5160
rect 3007 5120 3608 5148
rect 3007 5117 3019 5120
rect 2961 5111 3019 5117
rect 3602 5108 3608 5120
rect 3660 5108 3666 5160
rect 6914 5108 6920 5160
rect 6972 5148 6978 5160
rect 7193 5151 7251 5157
rect 7193 5148 7205 5151
rect 6972 5120 7205 5148
rect 6972 5108 6978 5120
rect 7193 5117 7205 5120
rect 7239 5148 7251 5151
rect 8205 5151 8263 5157
rect 8205 5148 8217 5151
rect 7239 5120 8217 5148
rect 7239 5117 7251 5120
rect 7193 5111 7251 5117
rect 8205 5117 8217 5120
rect 8251 5117 8263 5151
rect 8205 5111 8263 5117
rect 12621 5151 12679 5157
rect 12621 5117 12633 5151
rect 12667 5148 12679 5151
rect 13354 5148 13360 5160
rect 12667 5120 13360 5148
rect 12667 5117 12679 5120
rect 12621 5111 12679 5117
rect 13354 5108 13360 5120
rect 13412 5108 13418 5160
rect 19981 5151 20039 5157
rect 19981 5117 19993 5151
rect 20027 5148 20039 5151
rect 20714 5148 20720 5160
rect 20027 5120 20720 5148
rect 20027 5117 20039 5120
rect 19981 5111 20039 5117
rect 20714 5108 20720 5120
rect 20772 5148 20778 5160
rect 20809 5151 20867 5157
rect 20809 5148 20821 5151
rect 20772 5120 20821 5148
rect 20772 5108 20778 5120
rect 20809 5117 20821 5120
rect 20855 5117 20867 5151
rect 21284 5148 21312 5176
rect 22370 5148 22376 5160
rect 21284 5120 22376 5148
rect 20809 5111 20867 5117
rect 22370 5108 22376 5120
rect 22428 5108 22434 5160
rect 26421 5151 26479 5157
rect 26421 5117 26433 5151
rect 26467 5117 26479 5151
rect 26421 5111 26479 5117
rect 3142 5040 3148 5092
rect 3200 5089 3206 5092
rect 3200 5083 3264 5089
rect 3200 5049 3218 5083
rect 3252 5049 3264 5083
rect 3200 5043 3264 5049
rect 11057 5083 11115 5089
rect 11057 5049 11069 5083
rect 11103 5080 11115 5083
rect 11422 5080 11428 5092
rect 11103 5052 11428 5080
rect 11103 5049 11115 5052
rect 11057 5043 11115 5049
rect 3200 5040 3206 5043
rect 11422 5040 11428 5052
rect 11480 5040 11486 5092
rect 12894 5089 12900 5092
rect 12888 5080 12900 5089
rect 12855 5052 12900 5080
rect 12888 5043 12900 5052
rect 12894 5040 12900 5043
rect 12952 5040 12958 5092
rect 15102 5089 15108 5092
rect 14737 5083 14795 5089
rect 14737 5049 14749 5083
rect 14783 5080 14795 5083
rect 15074 5083 15108 5089
rect 15074 5080 15086 5083
rect 14783 5052 15086 5080
rect 14783 5049 14795 5052
rect 14737 5043 14795 5049
rect 15074 5049 15086 5052
rect 15160 5080 15166 5092
rect 23906 5083 23964 5089
rect 23906 5080 23918 5083
rect 15160 5052 15222 5080
rect 23584 5052 23918 5080
rect 15074 5043 15108 5049
rect 15102 5040 15108 5043
rect 15160 5040 15166 5052
rect 23584 5024 23612 5052
rect 23906 5049 23918 5052
rect 23952 5049 23964 5083
rect 26234 5080 26240 5092
rect 26195 5052 26240 5080
rect 23906 5043 23964 5049
rect 26234 5040 26240 5052
rect 26292 5080 26298 5092
rect 26436 5080 26464 5111
rect 26292 5052 26464 5080
rect 26292 5040 26298 5052
rect 3694 4972 3700 5024
rect 3752 5012 3758 5024
rect 4341 5015 4399 5021
rect 4341 5012 4353 5015
rect 3752 4984 4353 5012
rect 3752 4972 3758 4984
rect 4341 4981 4353 4984
rect 4387 5012 4399 5015
rect 4798 5012 4804 5024
rect 4387 4984 4804 5012
rect 4387 4981 4399 4984
rect 4341 4975 4399 4981
rect 4798 4972 4804 4984
rect 4856 4972 4862 5024
rect 6822 5012 6828 5024
rect 6783 4984 6828 5012
rect 6822 4972 6828 4984
rect 6880 4972 6886 5024
rect 11149 5015 11207 5021
rect 11149 4981 11161 5015
rect 11195 5012 11207 5015
rect 11330 5012 11336 5024
rect 11195 4984 11336 5012
rect 11195 4981 11207 4984
rect 11149 4975 11207 4981
rect 11330 4972 11336 4984
rect 11388 4972 11394 5024
rect 11606 4972 11612 5024
rect 11664 5012 11670 5024
rect 16666 5012 16672 5024
rect 11664 4984 16672 5012
rect 11664 4972 11670 4984
rect 16666 4972 16672 4984
rect 16724 4972 16730 5024
rect 20438 5012 20444 5024
rect 20399 4984 20444 5012
rect 20438 4972 20444 4984
rect 20496 4972 20502 5024
rect 23477 5015 23535 5021
rect 23477 4981 23489 5015
rect 23523 5012 23535 5015
rect 23566 5012 23572 5024
rect 23523 4984 23572 5012
rect 23523 4981 23535 4984
rect 23477 4975 23535 4981
rect 23566 4972 23572 4984
rect 23624 4972 23630 5024
rect 26602 5012 26608 5024
rect 26563 4984 26608 5012
rect 26602 4972 26608 4984
rect 26660 4972 26666 5024
rect 1104 4922 28888 4944
rect 1104 4870 10982 4922
rect 11034 4870 11046 4922
rect 11098 4870 11110 4922
rect 11162 4870 11174 4922
rect 11226 4870 20982 4922
rect 21034 4870 21046 4922
rect 21098 4870 21110 4922
rect 21162 4870 21174 4922
rect 21226 4870 28888 4922
rect 1104 4848 28888 4870
rect 1578 4808 1584 4820
rect 1539 4780 1584 4808
rect 1578 4768 1584 4780
rect 1636 4768 1642 4820
rect 3142 4808 3148 4820
rect 3103 4780 3148 4808
rect 3142 4768 3148 4780
rect 3200 4768 3206 4820
rect 3513 4811 3571 4817
rect 3513 4777 3525 4811
rect 3559 4808 3571 4811
rect 3602 4808 3608 4820
rect 3559 4780 3608 4808
rect 3559 4777 3571 4780
rect 3513 4771 3571 4777
rect 1762 4700 1768 4752
rect 1820 4740 1826 4752
rect 2409 4743 2467 4749
rect 2409 4740 2421 4743
rect 1820 4712 2421 4740
rect 1820 4700 1826 4712
rect 2409 4709 2421 4712
rect 2455 4740 2467 4743
rect 3528 4740 3556 4771
rect 3602 4768 3608 4780
rect 3660 4808 3666 4820
rect 5166 4808 5172 4820
rect 3660 4780 5172 4808
rect 3660 4768 3666 4780
rect 5166 4768 5172 4780
rect 5224 4768 5230 4820
rect 6362 4808 6368 4820
rect 6323 4780 6368 4808
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 7006 4768 7012 4820
rect 7064 4808 7070 4820
rect 7377 4811 7435 4817
rect 7377 4808 7389 4811
rect 7064 4780 7389 4808
rect 7064 4768 7070 4780
rect 7377 4777 7389 4780
rect 7423 4777 7435 4811
rect 10778 4808 10784 4820
rect 10739 4780 10784 4808
rect 7377 4771 7435 4777
rect 10778 4768 10784 4780
rect 10836 4768 10842 4820
rect 11149 4811 11207 4817
rect 11149 4777 11161 4811
rect 11195 4808 11207 4811
rect 11330 4808 11336 4820
rect 11195 4780 11336 4808
rect 11195 4777 11207 4780
rect 11149 4771 11207 4777
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 11422 4768 11428 4820
rect 11480 4808 11486 4820
rect 12897 4811 12955 4817
rect 12897 4808 12909 4811
rect 11480 4780 12909 4808
rect 11480 4768 11486 4780
rect 12897 4777 12909 4780
rect 12943 4777 12955 4811
rect 13262 4808 13268 4820
rect 13223 4780 13268 4808
rect 12897 4771 12955 4777
rect 13262 4768 13268 4780
rect 13320 4768 13326 4820
rect 13357 4811 13415 4817
rect 13357 4777 13369 4811
rect 13403 4808 13415 4811
rect 13446 4808 13452 4820
rect 13403 4780 13452 4808
rect 13403 4777 13415 4780
rect 13357 4771 13415 4777
rect 13446 4768 13452 4780
rect 13504 4768 13510 4820
rect 14642 4768 14648 4820
rect 14700 4808 14706 4820
rect 14829 4811 14887 4817
rect 14829 4808 14841 4811
rect 14700 4780 14841 4808
rect 14700 4768 14706 4780
rect 14829 4777 14841 4780
rect 14875 4777 14887 4811
rect 15838 4808 15844 4820
rect 15799 4780 15844 4808
rect 14829 4771 14887 4777
rect 2455 4712 3556 4740
rect 2455 4709 2467 4712
rect 2409 4703 2467 4709
rect 5718 4700 5724 4752
rect 5776 4740 5782 4752
rect 8110 4740 8116 4752
rect 5776 4712 8116 4740
rect 5776 4700 5782 4712
rect 8110 4700 8116 4712
rect 8168 4700 8174 4752
rect 11790 4740 11796 4752
rect 11751 4712 11796 4740
rect 11790 4700 11796 4712
rect 11848 4700 11854 4752
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4672 1455 4675
rect 2038 4672 2044 4684
rect 1443 4644 2044 4672
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 2038 4632 2044 4644
rect 2096 4632 2102 4684
rect 2498 4672 2504 4684
rect 2459 4644 2504 4672
rect 2498 4632 2504 4644
rect 2556 4632 2562 4684
rect 4062 4672 4068 4684
rect 4023 4644 4068 4672
rect 4062 4632 4068 4644
rect 4120 4632 4126 4684
rect 11606 4632 11612 4684
rect 11664 4672 11670 4684
rect 11701 4675 11759 4681
rect 11701 4672 11713 4675
rect 11664 4644 11713 4672
rect 11664 4632 11670 4644
rect 11701 4641 11713 4644
rect 11747 4641 11759 4675
rect 14844 4672 14872 4771
rect 15838 4768 15844 4780
rect 15896 4768 15902 4820
rect 19613 4811 19671 4817
rect 19613 4777 19625 4811
rect 19659 4808 19671 4811
rect 19702 4808 19708 4820
rect 19659 4780 19708 4808
rect 19659 4777 19671 4780
rect 19613 4771 19671 4777
rect 19702 4768 19708 4780
rect 19760 4808 19766 4820
rect 20438 4808 20444 4820
rect 19760 4780 20444 4808
rect 19760 4768 19766 4780
rect 20438 4768 20444 4780
rect 20496 4768 20502 4820
rect 20533 4811 20591 4817
rect 20533 4777 20545 4811
rect 20579 4808 20591 4811
rect 21266 4808 21272 4820
rect 20579 4780 21272 4808
rect 20579 4777 20591 4780
rect 20533 4771 20591 4777
rect 21266 4768 21272 4780
rect 21324 4768 21330 4820
rect 21358 4768 21364 4820
rect 21416 4808 21422 4820
rect 21913 4811 21971 4817
rect 21913 4808 21925 4811
rect 21416 4780 21925 4808
rect 21416 4768 21422 4780
rect 21913 4777 21925 4780
rect 21959 4808 21971 4811
rect 22094 4808 22100 4820
rect 21959 4780 22100 4808
rect 21959 4777 21971 4780
rect 21913 4771 21971 4777
rect 22094 4768 22100 4780
rect 22152 4768 22158 4820
rect 27338 4768 27344 4820
rect 27396 4808 27402 4820
rect 27798 4808 27804 4820
rect 27396 4780 27804 4808
rect 27396 4768 27402 4780
rect 27798 4768 27804 4780
rect 27856 4768 27862 4820
rect 16298 4749 16304 4752
rect 15565 4743 15623 4749
rect 15565 4709 15577 4743
rect 15611 4740 15623 4743
rect 16292 4740 16304 4749
rect 15611 4712 16304 4740
rect 15611 4709 15623 4712
rect 15565 4703 15623 4709
rect 16292 4703 16304 4712
rect 16298 4700 16304 4703
rect 16356 4700 16362 4752
rect 16390 4700 16396 4752
rect 16448 4700 16454 4752
rect 22370 4700 22376 4752
rect 22428 4749 22434 4752
rect 22428 4743 22492 4749
rect 22428 4709 22446 4743
rect 22480 4709 22492 4743
rect 22428 4703 22492 4709
rect 22428 4700 22434 4703
rect 16025 4675 16083 4681
rect 16025 4672 16037 4675
rect 14844 4644 16037 4672
rect 11701 4635 11759 4641
rect 16025 4641 16037 4644
rect 16071 4672 16083 4675
rect 16408 4672 16436 4700
rect 18046 4672 18052 4684
rect 16071 4644 18052 4672
rect 16071 4641 16083 4644
rect 16025 4635 16083 4641
rect 18046 4632 18052 4644
rect 18104 4632 18110 4684
rect 21177 4675 21235 4681
rect 21177 4641 21189 4675
rect 21223 4672 21235 4675
rect 21358 4672 21364 4684
rect 21223 4644 21364 4672
rect 21223 4641 21235 4644
rect 21177 4635 21235 4641
rect 21358 4632 21364 4644
rect 21416 4672 21422 4684
rect 21818 4672 21824 4684
rect 21416 4644 21824 4672
rect 21416 4632 21422 4644
rect 21818 4632 21824 4644
rect 21876 4632 21882 4684
rect 26510 4672 26516 4684
rect 26471 4644 26516 4672
rect 26510 4632 26516 4644
rect 26568 4632 26574 4684
rect 6454 4604 6460 4616
rect 6415 4576 6460 4604
rect 6454 4564 6460 4576
rect 6512 4564 6518 4616
rect 6546 4564 6552 4616
rect 6604 4604 6610 4616
rect 7009 4607 7067 4613
rect 7009 4604 7021 4607
rect 6604 4576 7021 4604
rect 6604 4564 6610 4576
rect 7009 4573 7021 4576
rect 7055 4604 7067 4607
rect 7558 4604 7564 4616
rect 7055 4576 7564 4604
rect 7055 4573 7067 4576
rect 7009 4567 7067 4573
rect 7558 4564 7564 4576
rect 7616 4564 7622 4616
rect 11974 4604 11980 4616
rect 11887 4576 11980 4604
rect 11974 4564 11980 4576
rect 12032 4604 12038 4616
rect 12805 4607 12863 4613
rect 12805 4604 12817 4607
rect 12032 4576 12817 4604
rect 12032 4564 12038 4576
rect 12805 4573 12817 4576
rect 12851 4604 12863 4607
rect 12894 4604 12900 4616
rect 12851 4576 12900 4604
rect 12851 4573 12863 4576
rect 12805 4567 12863 4573
rect 12894 4564 12900 4576
rect 12952 4604 12958 4616
rect 13538 4604 13544 4616
rect 12952 4576 13544 4604
rect 12952 4564 12958 4576
rect 13538 4564 13544 4576
rect 13596 4564 13602 4616
rect 19610 4564 19616 4616
rect 19668 4604 19674 4616
rect 19705 4607 19763 4613
rect 19705 4604 19717 4607
rect 19668 4576 19717 4604
rect 19668 4564 19674 4576
rect 19705 4573 19717 4576
rect 19751 4573 19763 4607
rect 19886 4604 19892 4616
rect 19847 4576 19892 4604
rect 19705 4567 19763 4573
rect 19886 4564 19892 4576
rect 19944 4564 19950 4616
rect 22186 4604 22192 4616
rect 22147 4576 22192 4604
rect 22186 4564 22192 4576
rect 22244 4564 22250 4616
rect 23566 4536 23572 4548
rect 23527 4508 23572 4536
rect 23566 4496 23572 4508
rect 23624 4496 23630 4548
rect 2682 4468 2688 4480
rect 2643 4440 2688 4468
rect 2682 4428 2688 4440
rect 2740 4428 2746 4480
rect 4154 4428 4160 4480
rect 4212 4468 4218 4480
rect 4249 4471 4307 4477
rect 4249 4468 4261 4471
rect 4212 4440 4261 4468
rect 4212 4428 4218 4440
rect 4249 4437 4261 4440
rect 4295 4437 4307 4471
rect 4249 4431 4307 4437
rect 5997 4471 6055 4477
rect 5997 4437 6009 4471
rect 6043 4468 6055 4471
rect 6270 4468 6276 4480
rect 6043 4440 6276 4468
rect 6043 4437 6055 4440
rect 5997 4431 6055 4437
rect 6270 4428 6276 4440
rect 6328 4428 6334 4480
rect 12434 4428 12440 4480
rect 12492 4468 12498 4480
rect 17405 4471 17463 4477
rect 12492 4440 12537 4468
rect 12492 4428 12498 4440
rect 17405 4437 17417 4471
rect 17451 4468 17463 4471
rect 17770 4468 17776 4480
rect 17451 4440 17776 4468
rect 17451 4437 17463 4440
rect 17405 4431 17463 4437
rect 17770 4428 17776 4440
rect 17828 4428 17834 4480
rect 19242 4468 19248 4480
rect 19203 4440 19248 4468
rect 19242 4428 19248 4440
rect 19300 4428 19306 4480
rect 26697 4471 26755 4477
rect 26697 4437 26709 4471
rect 26743 4468 26755 4471
rect 26878 4468 26884 4480
rect 26743 4440 26884 4468
rect 26743 4437 26755 4440
rect 26697 4431 26755 4437
rect 26878 4428 26884 4440
rect 26936 4428 26942 4480
rect 1104 4378 28888 4400
rect 1104 4326 5982 4378
rect 6034 4326 6046 4378
rect 6098 4326 6110 4378
rect 6162 4326 6174 4378
rect 6226 4326 15982 4378
rect 16034 4326 16046 4378
rect 16098 4326 16110 4378
rect 16162 4326 16174 4378
rect 16226 4326 25982 4378
rect 26034 4326 26046 4378
rect 26098 4326 26110 4378
rect 26162 4326 26174 4378
rect 26226 4326 28888 4378
rect 1104 4304 28888 4326
rect 2317 4267 2375 4273
rect 2317 4233 2329 4267
rect 2363 4264 2375 4267
rect 2498 4264 2504 4276
rect 2363 4236 2504 4264
rect 2363 4233 2375 4236
rect 2317 4227 2375 4233
rect 2498 4224 2504 4236
rect 2556 4224 2562 4276
rect 4798 4224 4804 4276
rect 4856 4264 4862 4276
rect 5629 4267 5687 4273
rect 5629 4264 5641 4267
rect 4856 4236 5641 4264
rect 4856 4224 4862 4236
rect 5629 4233 5641 4236
rect 5675 4264 5687 4267
rect 6546 4264 6552 4276
rect 5675 4236 6552 4264
rect 5675 4233 5687 4236
rect 5629 4227 5687 4233
rect 6546 4224 6552 4236
rect 6604 4224 6610 4276
rect 7466 4264 7472 4276
rect 7427 4236 7472 4264
rect 7466 4224 7472 4236
rect 7524 4224 7530 4276
rect 11241 4267 11299 4273
rect 11241 4233 11253 4267
rect 11287 4264 11299 4267
rect 11422 4264 11428 4276
rect 11287 4236 11428 4264
rect 11287 4233 11299 4236
rect 11241 4227 11299 4233
rect 11422 4224 11428 4236
rect 11480 4264 11486 4276
rect 11974 4264 11980 4276
rect 11480 4236 11980 4264
rect 11480 4224 11486 4236
rect 11974 4224 11980 4236
rect 12032 4224 12038 4276
rect 13262 4264 13268 4276
rect 13223 4236 13268 4264
rect 13262 4224 13268 4236
rect 13320 4224 13326 4276
rect 13538 4224 13544 4276
rect 13596 4264 13602 4276
rect 13633 4267 13691 4273
rect 13633 4264 13645 4267
rect 13596 4236 13645 4264
rect 13596 4224 13602 4236
rect 13633 4233 13645 4236
rect 13679 4233 13691 4267
rect 16390 4264 16396 4276
rect 16351 4236 16396 4264
rect 13633 4227 13691 4233
rect 16390 4224 16396 4236
rect 16448 4224 16454 4276
rect 17770 4264 17776 4276
rect 17731 4236 17776 4264
rect 17770 4224 17776 4236
rect 17828 4224 17834 4276
rect 19797 4267 19855 4273
rect 19797 4233 19809 4267
rect 19843 4264 19855 4267
rect 19886 4264 19892 4276
rect 19843 4236 19892 4264
rect 19843 4233 19855 4236
rect 19797 4227 19855 4233
rect 19886 4224 19892 4236
rect 19944 4224 19950 4276
rect 21634 4264 21640 4276
rect 21595 4236 21640 4264
rect 21634 4224 21640 4236
rect 21692 4224 21698 4276
rect 22370 4224 22376 4276
rect 22428 4264 22434 4276
rect 22833 4267 22891 4273
rect 22833 4264 22845 4267
rect 22428 4236 22845 4264
rect 22428 4224 22434 4236
rect 22833 4233 22845 4236
rect 22879 4233 22891 4267
rect 22833 4227 22891 4233
rect 26510 4224 26516 4276
rect 26568 4264 26574 4276
rect 27341 4267 27399 4273
rect 27341 4264 27353 4267
rect 26568 4236 27353 4264
rect 26568 4224 26574 4236
rect 27341 4233 27353 4236
rect 27387 4233 27399 4267
rect 27341 4227 27399 4233
rect 3142 4156 3148 4208
rect 3200 4196 3206 4208
rect 6089 4199 6147 4205
rect 3200 4168 3372 4196
rect 3200 4156 3206 4168
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4128 2743 4131
rect 3234 4128 3240 4140
rect 2731 4100 3240 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 3234 4088 3240 4100
rect 3292 4088 3298 4140
rect 3344 4137 3372 4168
rect 6089 4165 6101 4199
rect 6135 4196 6147 4199
rect 6362 4196 6368 4208
rect 6135 4168 6368 4196
rect 6135 4165 6147 4168
rect 6089 4159 6147 4165
rect 6362 4156 6368 4168
rect 6420 4156 6426 4208
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4097 3387 4131
rect 4985 4131 5043 4137
rect 4985 4128 4997 4131
rect 3329 4091 3387 4097
rect 4356 4100 4997 4128
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4060 1455 4063
rect 1854 4060 1860 4072
rect 1443 4032 1860 4060
rect 1443 4029 1455 4032
rect 1397 4023 1455 4029
rect 1854 4020 1860 4032
rect 1912 4020 1918 4072
rect 4356 4069 4384 4100
rect 4985 4097 4997 4100
rect 5031 4128 5043 4131
rect 5442 4128 5448 4140
rect 5031 4100 5448 4128
rect 5031 4097 5043 4100
rect 4985 4091 5043 4097
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 7484 4128 7512 4224
rect 11609 4199 11667 4205
rect 11609 4165 11621 4199
rect 11655 4196 11667 4199
rect 11790 4196 11796 4208
rect 11655 4168 11796 4196
rect 11655 4165 11667 4168
rect 11609 4159 11667 4165
rect 11790 4156 11796 4168
rect 11848 4156 11854 4208
rect 12989 4199 13047 4205
rect 12989 4165 13001 4199
rect 13035 4196 13047 4199
rect 13446 4196 13452 4208
rect 13035 4168 13452 4196
rect 13035 4165 13047 4168
rect 12989 4159 13047 4165
rect 13446 4156 13452 4168
rect 13504 4156 13510 4208
rect 16117 4199 16175 4205
rect 16117 4165 16129 4199
rect 16163 4196 16175 4199
rect 16298 4196 16304 4208
rect 16163 4168 16304 4196
rect 16163 4165 16175 4168
rect 16117 4159 16175 4165
rect 16298 4156 16304 4168
rect 16356 4156 16362 4208
rect 17788 4128 17816 4224
rect 19429 4199 19487 4205
rect 19429 4165 19441 4199
rect 19475 4196 19487 4199
rect 20346 4196 20352 4208
rect 19475 4168 20352 4196
rect 19475 4165 19487 4168
rect 19429 4159 19487 4165
rect 20346 4156 20352 4168
rect 20404 4196 20410 4208
rect 21358 4196 21364 4208
rect 20404 4168 21364 4196
rect 20404 4156 20410 4168
rect 20162 4128 20168 4140
rect 7484 4100 7788 4128
rect 17788 4100 18184 4128
rect 20123 4100 20168 4128
rect 4341 4063 4399 4069
rect 4341 4029 4353 4063
rect 4387 4029 4399 4063
rect 4341 4023 4399 4029
rect 7193 4063 7251 4069
rect 7193 4029 7205 4063
rect 7239 4060 7251 4063
rect 7653 4063 7711 4069
rect 7653 4060 7665 4063
rect 7239 4032 7665 4060
rect 7239 4029 7251 4032
rect 7193 4023 7251 4029
rect 7653 4029 7665 4032
rect 7699 4029 7711 4063
rect 7760 4060 7788 4100
rect 7909 4063 7967 4069
rect 7909 4060 7921 4063
rect 7760 4032 7921 4060
rect 7653 4023 7711 4029
rect 7909 4029 7921 4032
rect 7955 4029 7967 4063
rect 9674 4060 9680 4072
rect 7909 4023 7967 4029
rect 8128 4032 9680 4060
rect 7668 3992 7696 4023
rect 8128 3992 8156 4032
rect 9674 4020 9680 4032
rect 9732 4060 9738 4072
rect 9858 4060 9864 4072
rect 9732 4032 9864 4060
rect 9732 4020 9738 4032
rect 9858 4020 9864 4032
rect 9916 4020 9922 4072
rect 11606 4020 11612 4072
rect 11664 4060 11670 4072
rect 11885 4063 11943 4069
rect 11885 4060 11897 4063
rect 11664 4032 11897 4060
rect 11664 4020 11670 4032
rect 11885 4029 11897 4032
rect 11931 4029 11943 4063
rect 18046 4060 18052 4072
rect 18007 4032 18052 4060
rect 11885 4023 11943 4029
rect 18046 4020 18052 4032
rect 18104 4020 18110 4072
rect 18156 4060 18184 4100
rect 20162 4088 20168 4100
rect 20220 4128 20226 4140
rect 20916 4137 20944 4168
rect 21358 4156 21364 4168
rect 21416 4196 21422 4208
rect 21416 4168 22416 4196
rect 21416 4156 21422 4168
rect 20901 4131 20959 4137
rect 20220 4100 20668 4128
rect 20220 4088 20226 4100
rect 20640 4072 20668 4100
rect 20901 4097 20913 4131
rect 20947 4097 20959 4131
rect 20901 4091 20959 4097
rect 22094 4088 22100 4140
rect 22152 4128 22158 4140
rect 22388 4137 22416 4168
rect 22281 4131 22339 4137
rect 22281 4128 22293 4131
rect 22152 4100 22293 4128
rect 22152 4088 22158 4100
rect 22281 4097 22293 4100
rect 22327 4097 22339 4131
rect 22281 4091 22339 4097
rect 22373 4131 22431 4137
rect 22373 4097 22385 4131
rect 22419 4097 22431 4131
rect 22373 4091 22431 4097
rect 18322 4069 18328 4072
rect 18305 4063 18328 4069
rect 18305 4060 18317 4063
rect 18156 4032 18317 4060
rect 18305 4029 18317 4032
rect 18380 4060 18386 4072
rect 20622 4060 20628 4072
rect 18380 4032 18453 4060
rect 20535 4032 20628 4060
rect 18305 4023 18328 4029
rect 18322 4020 18328 4023
rect 18380 4020 18386 4032
rect 20622 4020 20628 4032
rect 20680 4020 20686 4072
rect 21634 4020 21640 4072
rect 21692 4060 21698 4072
rect 22189 4063 22247 4069
rect 22189 4060 22201 4063
rect 21692 4032 22201 4060
rect 21692 4020 21698 4032
rect 22189 4029 22201 4032
rect 22235 4029 22247 4063
rect 26418 4060 26424 4072
rect 26379 4032 26424 4060
rect 22189 4023 22247 4029
rect 10106 3995 10164 4001
rect 10106 3992 10118 3995
rect 7668 3964 8156 3992
rect 9692 3964 10118 3992
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 2774 3884 2780 3936
rect 2832 3924 2838 3936
rect 3142 3924 3148 3936
rect 2832 3896 2877 3924
rect 3055 3896 3148 3924
rect 2832 3884 2838 3896
rect 3142 3884 3148 3896
rect 3200 3924 3206 3936
rect 4062 3924 4068 3936
rect 3200 3896 4068 3924
rect 3200 3884 3206 3896
rect 4062 3884 4068 3896
rect 4120 3924 4126 3936
rect 4157 3927 4215 3933
rect 4157 3924 4169 3927
rect 4120 3896 4169 3924
rect 4120 3884 4126 3896
rect 4157 3893 4169 3896
rect 4203 3924 4215 3927
rect 4246 3924 4252 3936
rect 4203 3896 4252 3924
rect 4203 3893 4215 3896
rect 4157 3887 4215 3893
rect 4246 3884 4252 3896
rect 4304 3884 4310 3936
rect 4522 3924 4528 3936
rect 4483 3896 4528 3924
rect 4522 3884 4528 3896
rect 4580 3884 4586 3936
rect 6454 3924 6460 3936
rect 6415 3896 6460 3924
rect 6454 3884 6460 3896
rect 6512 3884 6518 3936
rect 9030 3924 9036 3936
rect 8991 3896 9036 3924
rect 9030 3884 9036 3896
rect 9088 3924 9094 3936
rect 9692 3933 9720 3964
rect 10106 3961 10118 3964
rect 10152 3961 10164 3995
rect 22204 3992 22232 4023
rect 26418 4020 26424 4032
rect 26476 4060 26482 4072
rect 26973 4063 27031 4069
rect 26973 4060 26985 4063
rect 26476 4032 26985 4060
rect 26476 4020 26482 4032
rect 26973 4029 26985 4032
rect 27019 4029 27031 4063
rect 26973 4023 27031 4029
rect 27525 4063 27583 4069
rect 27525 4029 27537 4063
rect 27571 4060 27583 4063
rect 28077 4063 28135 4069
rect 28077 4060 28089 4063
rect 27571 4032 28089 4060
rect 27571 4029 27583 4032
rect 27525 4023 27583 4029
rect 28077 4029 28089 4032
rect 28123 4029 28135 4063
rect 28077 4023 28135 4029
rect 27540 3992 27568 4023
rect 22204 3964 27568 3992
rect 10106 3955 10164 3961
rect 9677 3927 9735 3933
rect 9677 3924 9689 3927
rect 9088 3896 9689 3924
rect 9088 3884 9094 3896
rect 9677 3893 9689 3896
rect 9723 3893 9735 3927
rect 20254 3924 20260 3936
rect 20215 3896 20260 3924
rect 9677 3887 9735 3893
rect 20254 3884 20260 3896
rect 20312 3884 20318 3936
rect 20714 3884 20720 3936
rect 20772 3924 20778 3936
rect 21818 3924 21824 3936
rect 20772 3896 20817 3924
rect 21779 3896 21824 3924
rect 20772 3884 20778 3896
rect 21818 3884 21824 3896
rect 21876 3884 21882 3936
rect 26605 3927 26663 3933
rect 26605 3893 26617 3927
rect 26651 3924 26663 3927
rect 26694 3924 26700 3936
rect 26651 3896 26700 3924
rect 26651 3893 26663 3896
rect 26605 3887 26663 3893
rect 26694 3884 26700 3896
rect 26752 3884 26758 3936
rect 27706 3924 27712 3936
rect 27667 3896 27712 3924
rect 27706 3884 27712 3896
rect 27764 3884 27770 3936
rect 1104 3834 28888 3856
rect 1104 3782 10982 3834
rect 11034 3782 11046 3834
rect 11098 3782 11110 3834
rect 11162 3782 11174 3834
rect 11226 3782 20982 3834
rect 21034 3782 21046 3834
rect 21098 3782 21110 3834
rect 21162 3782 21174 3834
rect 21226 3782 28888 3834
rect 1104 3760 28888 3782
rect 1673 3723 1731 3729
rect 1673 3689 1685 3723
rect 1719 3720 1731 3723
rect 1854 3720 1860 3732
rect 1719 3692 1860 3720
rect 1719 3689 1731 3692
rect 1673 3683 1731 3689
rect 1854 3680 1860 3692
rect 1912 3680 1918 3732
rect 2774 3680 2780 3732
rect 2832 3720 2838 3732
rect 3329 3723 3387 3729
rect 3329 3720 3341 3723
rect 2832 3692 3341 3720
rect 2832 3680 2838 3692
rect 3329 3689 3341 3692
rect 3375 3720 3387 3723
rect 3786 3720 3792 3732
rect 3375 3692 3792 3720
rect 3375 3689 3387 3692
rect 3329 3683 3387 3689
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 5442 3680 5448 3732
rect 5500 3720 5506 3732
rect 5813 3723 5871 3729
rect 5813 3720 5825 3723
rect 5500 3692 5825 3720
rect 5500 3680 5506 3692
rect 5813 3689 5825 3692
rect 5859 3720 5871 3723
rect 6917 3723 6975 3729
rect 6917 3720 6929 3723
rect 5859 3692 6929 3720
rect 5859 3689 5871 3692
rect 5813 3683 5871 3689
rect 6917 3689 6929 3692
rect 6963 3689 6975 3723
rect 9858 3720 9864 3732
rect 9819 3692 9864 3720
rect 6917 3683 6975 3689
rect 9858 3680 9864 3692
rect 9916 3680 9922 3732
rect 11422 3720 11428 3732
rect 11383 3692 11428 3720
rect 11422 3680 11428 3692
rect 11480 3680 11486 3732
rect 19702 3720 19708 3732
rect 19663 3692 19708 3720
rect 19702 3680 19708 3692
rect 19760 3680 19766 3732
rect 20346 3720 20352 3732
rect 20307 3692 20352 3720
rect 20346 3680 20352 3692
rect 20404 3680 20410 3732
rect 21269 3723 21327 3729
rect 21269 3689 21281 3723
rect 21315 3720 21327 3723
rect 21818 3720 21824 3732
rect 21315 3692 21824 3720
rect 21315 3689 21327 3692
rect 21269 3683 21327 3689
rect 21818 3680 21824 3692
rect 21876 3680 21882 3732
rect 22278 3720 22284 3732
rect 22239 3692 22284 3720
rect 22278 3680 22284 3692
rect 22336 3680 22342 3732
rect 2869 3655 2927 3661
rect 2869 3621 2881 3655
rect 2915 3652 2927 3655
rect 3142 3652 3148 3664
rect 2915 3624 3148 3652
rect 2915 3621 2927 3624
rect 2869 3615 2927 3621
rect 3142 3612 3148 3624
rect 3200 3612 3206 3664
rect 6270 3612 6276 3664
rect 6328 3652 6334 3664
rect 7285 3655 7343 3661
rect 7285 3652 7297 3655
rect 6328 3624 7297 3652
rect 6328 3612 6334 3624
rect 7285 3621 7297 3624
rect 7331 3621 7343 3655
rect 7285 3615 7343 3621
rect 20254 3612 20260 3664
rect 20312 3652 20318 3664
rect 21358 3652 21364 3664
rect 20312 3624 21364 3652
rect 20312 3612 20318 3624
rect 21358 3612 21364 3624
rect 21416 3612 21422 3664
rect 1946 3584 1952 3596
rect 1907 3556 1952 3584
rect 1946 3544 1952 3556
rect 2004 3544 2010 3596
rect 4062 3584 4068 3596
rect 4023 3556 4068 3584
rect 4062 3544 4068 3556
rect 4120 3544 4126 3596
rect 4798 3544 4804 3596
rect 4856 3584 4862 3596
rect 5721 3587 5779 3593
rect 5721 3584 5733 3587
rect 4856 3556 5733 3584
rect 4856 3544 4862 3556
rect 5721 3553 5733 3556
rect 5767 3584 5779 3587
rect 6822 3584 6828 3596
rect 5767 3556 6828 3584
rect 5767 3553 5779 3556
rect 5721 3547 5779 3553
rect 6822 3544 6828 3556
rect 6880 3544 6886 3596
rect 15654 3584 15660 3596
rect 15615 3556 15660 3584
rect 15654 3544 15660 3556
rect 15712 3544 15718 3596
rect 17310 3544 17316 3596
rect 17368 3584 17374 3596
rect 18049 3587 18107 3593
rect 18049 3584 18061 3587
rect 17368 3556 18061 3584
rect 17368 3544 17374 3556
rect 18049 3553 18061 3556
rect 18095 3553 18107 3587
rect 18049 3547 18107 3553
rect 23934 3544 23940 3596
rect 23992 3584 23998 3596
rect 26513 3587 26571 3593
rect 26513 3584 26525 3587
rect 23992 3556 26525 3584
rect 23992 3544 23998 3556
rect 26513 3553 26525 3556
rect 26559 3584 26571 3587
rect 27338 3584 27344 3596
rect 26559 3556 27344 3584
rect 26559 3553 26571 3556
rect 26513 3547 26571 3553
rect 27338 3544 27344 3556
rect 27396 3544 27402 3596
rect 5810 3476 5816 3528
rect 5868 3516 5874 3528
rect 5905 3519 5963 3525
rect 5905 3516 5917 3519
rect 5868 3488 5917 3516
rect 5868 3476 5874 3488
rect 5905 3485 5917 3488
rect 5951 3485 5963 3519
rect 5905 3479 5963 3485
rect 6546 3476 6552 3528
rect 6604 3516 6610 3528
rect 7377 3519 7435 3525
rect 7377 3516 7389 3519
rect 6604 3488 7389 3516
rect 6604 3476 6610 3488
rect 7377 3485 7389 3488
rect 7423 3485 7435 3519
rect 7377 3479 7435 3485
rect 7466 3476 7472 3528
rect 7524 3516 7530 3528
rect 15933 3519 15991 3525
rect 7524 3488 7569 3516
rect 7524 3476 7530 3488
rect 15933 3485 15945 3519
rect 15979 3516 15991 3519
rect 16298 3516 16304 3528
rect 15979 3488 16304 3516
rect 15979 3485 15991 3488
rect 15933 3479 15991 3485
rect 16298 3476 16304 3488
rect 16356 3476 16362 3528
rect 17862 3476 17868 3528
rect 17920 3516 17926 3528
rect 18141 3519 18199 3525
rect 18141 3516 18153 3519
rect 17920 3488 18153 3516
rect 17920 3476 17926 3488
rect 18141 3485 18153 3488
rect 18187 3485 18199 3519
rect 18322 3516 18328 3528
rect 18283 3488 18328 3516
rect 18141 3479 18199 3485
rect 18322 3476 18328 3488
rect 18380 3476 18386 3528
rect 19337 3519 19395 3525
rect 19337 3485 19349 3519
rect 19383 3516 19395 3519
rect 19610 3516 19616 3528
rect 19383 3488 19616 3516
rect 19383 3485 19395 3488
rect 19337 3479 19395 3485
rect 19610 3476 19616 3488
rect 19668 3516 19674 3528
rect 19668 3488 20944 3516
rect 19668 3476 19674 3488
rect 17681 3451 17739 3457
rect 17681 3417 17693 3451
rect 17727 3448 17739 3451
rect 20625 3451 20683 3457
rect 20625 3448 20637 3451
rect 17727 3420 20637 3448
rect 17727 3417 17739 3420
rect 17681 3411 17739 3417
rect 20625 3417 20637 3420
rect 20671 3448 20683 3451
rect 20714 3448 20720 3460
rect 20671 3420 20720 3448
rect 20671 3417 20683 3420
rect 20625 3411 20683 3417
rect 20714 3408 20720 3420
rect 20772 3408 20778 3460
rect 20916 3457 20944 3488
rect 21266 3476 21272 3528
rect 21324 3516 21330 3528
rect 21453 3519 21511 3525
rect 21453 3516 21465 3519
rect 21324 3488 21465 3516
rect 21324 3476 21330 3488
rect 21453 3485 21465 3488
rect 21499 3485 21511 3519
rect 21453 3479 21511 3485
rect 20901 3451 20959 3457
rect 20901 3417 20913 3451
rect 20947 3417 20959 3451
rect 20901 3411 20959 3417
rect 2130 3380 2136 3392
rect 2091 3352 2136 3380
rect 2130 3340 2136 3352
rect 2188 3340 2194 3392
rect 4062 3340 4068 3392
rect 4120 3380 4126 3392
rect 4249 3383 4307 3389
rect 4249 3380 4261 3383
rect 4120 3352 4261 3380
rect 4120 3340 4126 3352
rect 4249 3349 4261 3352
rect 4295 3349 4307 3383
rect 5350 3380 5356 3392
rect 5311 3352 5356 3380
rect 4249 3343 4307 3349
rect 5350 3340 5356 3352
rect 5408 3340 5414 3392
rect 26697 3383 26755 3389
rect 26697 3349 26709 3383
rect 26743 3380 26755 3383
rect 26786 3380 26792 3392
rect 26743 3352 26792 3380
rect 26743 3349 26755 3352
rect 26697 3343 26755 3349
rect 26786 3340 26792 3352
rect 26844 3340 26850 3392
rect 1104 3290 28888 3312
rect 1104 3238 5982 3290
rect 6034 3238 6046 3290
rect 6098 3238 6110 3290
rect 6162 3238 6174 3290
rect 6226 3238 15982 3290
rect 16034 3238 16046 3290
rect 16098 3238 16110 3290
rect 16162 3238 16174 3290
rect 16226 3238 25982 3290
rect 26034 3238 26046 3290
rect 26098 3238 26110 3290
rect 26162 3238 26174 3290
rect 26226 3238 28888 3290
rect 1104 3216 28888 3238
rect 1946 3136 1952 3188
rect 2004 3176 2010 3188
rect 2133 3179 2191 3185
rect 2133 3176 2145 3179
rect 2004 3148 2145 3176
rect 2004 3136 2010 3148
rect 2133 3145 2145 3148
rect 2179 3145 2191 3179
rect 4430 3176 4436 3188
rect 4391 3148 4436 3176
rect 2133 3139 2191 3145
rect 4430 3136 4436 3148
rect 4488 3136 4494 3188
rect 4798 3176 4804 3188
rect 4759 3148 4804 3176
rect 4798 3136 4804 3148
rect 4856 3136 4862 3188
rect 5810 3176 5816 3188
rect 5771 3148 5816 3176
rect 5810 3136 5816 3148
rect 5868 3136 5874 3188
rect 6270 3176 6276 3188
rect 6231 3148 6276 3176
rect 6270 3136 6276 3148
rect 6328 3136 6334 3188
rect 7466 3136 7472 3188
rect 7524 3176 7530 3188
rect 7561 3179 7619 3185
rect 7561 3176 7573 3179
rect 7524 3148 7573 3176
rect 7524 3136 7530 3148
rect 7561 3145 7573 3148
rect 7607 3145 7619 3179
rect 13630 3176 13636 3188
rect 13591 3148 13636 3176
rect 7561 3139 7619 3145
rect 13630 3136 13636 3148
rect 13688 3136 13694 3188
rect 15289 3179 15347 3185
rect 15289 3145 15301 3179
rect 15335 3176 15347 3179
rect 15470 3176 15476 3188
rect 15335 3148 15476 3176
rect 15335 3145 15347 3148
rect 15289 3139 15347 3145
rect 3326 3108 3332 3120
rect 3287 3080 3332 3108
rect 3326 3068 3332 3080
rect 3384 3068 3390 3120
rect 3970 3068 3976 3120
rect 4028 3108 4034 3120
rect 5077 3111 5135 3117
rect 5077 3108 5089 3111
rect 4028 3080 5089 3108
rect 4028 3068 4034 3080
rect 5077 3077 5089 3080
rect 5123 3077 5135 3111
rect 5077 3071 5135 3077
rect 3786 3040 3792 3052
rect 3747 3012 3792 3040
rect 3786 3000 3792 3012
rect 3844 3000 3850 3052
rect 3881 3043 3939 3049
rect 3881 3009 3893 3043
rect 3927 3009 3939 3043
rect 6546 3040 6552 3052
rect 6507 3012 6552 3040
rect 3881 3003 3939 3009
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2972 1455 2975
rect 1946 2972 1952 2984
rect 1443 2944 1952 2972
rect 1443 2941 1455 2944
rect 1397 2935 1455 2941
rect 1946 2932 1952 2944
rect 2004 2932 2010 2984
rect 3694 2932 3700 2984
rect 3752 2972 3758 2984
rect 3896 2972 3924 3003
rect 6546 3000 6552 3012
rect 6604 3000 6610 3052
rect 3752 2944 3924 2972
rect 3752 2932 3758 2944
rect 1673 2907 1731 2913
rect 1673 2873 1685 2907
rect 1719 2904 1731 2907
rect 2038 2904 2044 2916
rect 1719 2876 2044 2904
rect 1719 2873 1731 2876
rect 1673 2867 1731 2873
rect 2038 2864 2044 2876
rect 2096 2864 2102 2916
rect 3896 2848 3924 2944
rect 4614 2932 4620 2984
rect 4672 2972 4678 2984
rect 4893 2975 4951 2981
rect 4893 2972 4905 2975
rect 4672 2944 4905 2972
rect 4672 2932 4678 2944
rect 4893 2941 4905 2944
rect 4939 2972 4951 2975
rect 5445 2975 5503 2981
rect 5445 2972 5457 2975
rect 4939 2944 5457 2972
rect 4939 2941 4951 2944
rect 4893 2935 4951 2941
rect 5445 2941 5457 2944
rect 5491 2941 5503 2975
rect 5445 2935 5503 2941
rect 6730 2932 6736 2984
rect 6788 2972 6794 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6788 2944 6837 2972
rect 6788 2932 6794 2944
rect 6825 2941 6837 2944
rect 6871 2972 6883 2975
rect 7929 2975 7987 2981
rect 7929 2972 7941 2975
rect 6871 2944 7941 2972
rect 6871 2941 6883 2944
rect 6825 2935 6883 2941
rect 7929 2941 7941 2944
rect 7975 2941 7987 2975
rect 7929 2935 7987 2941
rect 12897 2975 12955 2981
rect 12897 2941 12909 2975
rect 12943 2972 12955 2975
rect 13630 2972 13636 2984
rect 12943 2944 13636 2972
rect 12943 2941 12955 2944
rect 12897 2935 12955 2941
rect 13630 2932 13636 2944
rect 13688 2932 13694 2984
rect 14461 2975 14519 2981
rect 14461 2941 14473 2975
rect 14507 2972 14519 2975
rect 15304 2972 15332 3139
rect 15470 3136 15476 3148
rect 15528 3136 15534 3188
rect 15654 3176 15660 3188
rect 15615 3148 15660 3176
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 17310 3176 17316 3188
rect 17271 3148 17316 3176
rect 17310 3136 17316 3148
rect 17368 3136 17374 3188
rect 21358 3176 21364 3188
rect 21319 3148 21364 3176
rect 21358 3136 21364 3148
rect 21416 3136 21422 3188
rect 21729 3179 21787 3185
rect 21729 3145 21741 3179
rect 21775 3176 21787 3179
rect 21818 3176 21824 3188
rect 21775 3148 21824 3176
rect 21775 3145 21787 3148
rect 21729 3139 21787 3145
rect 21818 3136 21824 3148
rect 21876 3136 21882 3188
rect 27338 3176 27344 3188
rect 27299 3148 27344 3176
rect 27338 3136 27344 3148
rect 27396 3136 27402 3188
rect 17773 3111 17831 3117
rect 17773 3077 17785 3111
rect 17819 3108 17831 3111
rect 17862 3108 17868 3120
rect 17819 3080 17868 3108
rect 17819 3077 17831 3080
rect 17773 3071 17831 3077
rect 17862 3068 17868 3080
rect 17920 3068 17926 3120
rect 20993 3111 21051 3117
rect 20993 3077 21005 3111
rect 21039 3108 21051 3111
rect 21266 3108 21272 3120
rect 21039 3080 21272 3108
rect 21039 3077 21051 3080
rect 20993 3071 21051 3077
rect 21266 3068 21272 3080
rect 21324 3068 21330 3120
rect 24949 3111 25007 3117
rect 24949 3077 24961 3111
rect 24995 3108 25007 3111
rect 26326 3108 26332 3120
rect 24995 3080 26332 3108
rect 24995 3077 25007 3080
rect 24949 3071 25007 3077
rect 26326 3068 26332 3080
rect 26384 3068 26390 3120
rect 14507 2944 15332 2972
rect 14507 2941 14519 2944
rect 14461 2935 14519 2941
rect 17954 2932 17960 2984
rect 18012 2972 18018 2984
rect 18049 2975 18107 2981
rect 18049 2972 18061 2975
rect 18012 2944 18061 2972
rect 18012 2932 18018 2944
rect 18049 2941 18061 2944
rect 18095 2972 18107 2975
rect 18785 2975 18843 2981
rect 18785 2972 18797 2975
rect 18095 2944 18797 2972
rect 18095 2941 18107 2944
rect 18049 2935 18107 2941
rect 18785 2941 18797 2944
rect 18831 2941 18843 2975
rect 18785 2935 18843 2941
rect 23661 2975 23719 2981
rect 23661 2941 23673 2975
rect 23707 2972 23719 2975
rect 24305 2975 24363 2981
rect 24305 2972 24317 2975
rect 23707 2944 24317 2972
rect 23707 2941 23719 2944
rect 23661 2935 23719 2941
rect 24305 2941 24317 2944
rect 24351 2972 24363 2975
rect 24765 2975 24823 2981
rect 24765 2972 24777 2975
rect 24351 2944 24777 2972
rect 24351 2941 24363 2944
rect 24305 2935 24363 2941
rect 24765 2941 24777 2944
rect 24811 2972 24823 2975
rect 24946 2972 24952 2984
rect 24811 2944 24952 2972
rect 24811 2941 24823 2944
rect 24765 2935 24823 2941
rect 24946 2932 24952 2944
rect 25004 2972 25010 2984
rect 25317 2975 25375 2981
rect 25317 2972 25329 2975
rect 25004 2944 25329 2972
rect 25004 2932 25010 2944
rect 25317 2941 25329 2944
rect 25363 2941 25375 2975
rect 26418 2972 26424 2984
rect 26379 2944 26424 2972
rect 25317 2935 25375 2941
rect 26418 2932 26424 2944
rect 26476 2972 26482 2984
rect 26973 2975 27031 2981
rect 26973 2972 26985 2975
rect 26476 2944 26985 2972
rect 26476 2932 26482 2944
rect 26973 2941 26985 2944
rect 27019 2941 27031 2975
rect 27522 2972 27528 2984
rect 27483 2944 27528 2972
rect 26973 2935 27031 2941
rect 27522 2932 27528 2944
rect 27580 2972 27586 2984
rect 28077 2975 28135 2981
rect 28077 2972 28089 2975
rect 27580 2944 28089 2972
rect 27580 2932 27586 2944
rect 28077 2941 28089 2944
rect 28123 2941 28135 2975
rect 28077 2935 28135 2941
rect 7101 2907 7159 2913
rect 7101 2873 7113 2907
rect 7147 2904 7159 2907
rect 7742 2904 7748 2916
rect 7147 2876 7748 2904
rect 7147 2873 7159 2876
rect 7101 2867 7159 2873
rect 7742 2864 7748 2876
rect 7800 2864 7806 2916
rect 13173 2907 13231 2913
rect 13173 2873 13185 2907
rect 13219 2904 13231 2907
rect 13446 2904 13452 2916
rect 13219 2876 13452 2904
rect 13219 2873 13231 2876
rect 13173 2867 13231 2873
rect 13446 2864 13452 2876
rect 13504 2864 13510 2916
rect 14737 2907 14795 2913
rect 14737 2873 14749 2907
rect 14783 2904 14795 2907
rect 14918 2904 14924 2916
rect 14783 2876 14924 2904
rect 14783 2873 14795 2876
rect 14737 2867 14795 2873
rect 14918 2864 14924 2876
rect 14976 2864 14982 2916
rect 18325 2907 18383 2913
rect 18325 2873 18337 2907
rect 18371 2904 18383 2907
rect 19150 2904 19156 2916
rect 18371 2876 19156 2904
rect 18371 2873 18383 2876
rect 18325 2867 18383 2873
rect 19150 2864 19156 2876
rect 19208 2864 19214 2916
rect 21726 2864 21732 2916
rect 21784 2904 21790 2916
rect 24026 2904 24032 2916
rect 21784 2876 24032 2904
rect 21784 2864 21790 2876
rect 24026 2864 24032 2876
rect 24084 2864 24090 2916
rect 3237 2839 3295 2845
rect 3237 2805 3249 2839
rect 3283 2836 3295 2839
rect 3697 2839 3755 2845
rect 3697 2836 3709 2839
rect 3283 2808 3709 2836
rect 3283 2805 3295 2808
rect 3237 2799 3295 2805
rect 3697 2805 3709 2808
rect 3743 2836 3755 2839
rect 3786 2836 3792 2848
rect 3743 2808 3792 2836
rect 3743 2805 3755 2808
rect 3697 2799 3755 2805
rect 3786 2796 3792 2808
rect 3844 2796 3850 2848
rect 3878 2796 3884 2848
rect 3936 2796 3942 2848
rect 23842 2836 23848 2848
rect 23803 2808 23848 2836
rect 23842 2796 23848 2808
rect 23900 2796 23906 2848
rect 26602 2836 26608 2848
rect 26563 2808 26608 2836
rect 26602 2796 26608 2808
rect 26660 2796 26666 2848
rect 27706 2836 27712 2848
rect 27667 2808 27712 2836
rect 27706 2796 27712 2808
rect 27764 2796 27770 2848
rect 1104 2746 28888 2768
rect 1104 2694 10982 2746
rect 11034 2694 11046 2746
rect 11098 2694 11110 2746
rect 11162 2694 11174 2746
rect 11226 2694 20982 2746
rect 21034 2694 21046 2746
rect 21098 2694 21110 2746
rect 21162 2694 21174 2746
rect 21226 2694 28888 2746
rect 1104 2672 28888 2694
rect 1673 2635 1731 2641
rect 1673 2601 1685 2635
rect 1719 2632 1731 2635
rect 1946 2632 1952 2644
rect 1719 2604 1952 2632
rect 1719 2601 1731 2604
rect 1673 2595 1731 2601
rect 1946 2592 1952 2604
rect 2004 2592 2010 2644
rect 2961 2635 3019 2641
rect 2961 2601 2973 2635
rect 3007 2632 3019 2635
rect 3510 2632 3516 2644
rect 3007 2604 3516 2632
rect 3007 2601 3019 2604
rect 2961 2595 3019 2601
rect 2133 2499 2191 2505
rect 2133 2465 2145 2499
rect 2179 2496 2191 2499
rect 2976 2496 3004 2595
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 3878 2592 3884 2644
rect 3936 2592 3942 2644
rect 5442 2632 5448 2644
rect 5403 2604 5448 2632
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 6273 2635 6331 2641
rect 6273 2601 6285 2635
rect 6319 2632 6331 2635
rect 6454 2632 6460 2644
rect 6319 2604 6460 2632
rect 6319 2601 6331 2604
rect 6273 2595 6331 2601
rect 3421 2567 3479 2573
rect 3421 2533 3433 2567
rect 3467 2564 3479 2567
rect 3896 2564 3924 2592
rect 3467 2536 3924 2564
rect 3467 2533 3479 2536
rect 3421 2527 3479 2533
rect 2179 2468 3004 2496
rect 3881 2499 3939 2505
rect 2179 2465 2191 2468
rect 2133 2459 2191 2465
rect 3881 2465 3893 2499
rect 3927 2496 3939 2499
rect 4341 2499 4399 2505
rect 4341 2496 4353 2499
rect 3927 2468 4353 2496
rect 3927 2465 3939 2468
rect 3881 2459 3939 2465
rect 4341 2465 4353 2468
rect 4387 2496 4399 2499
rect 5350 2496 5356 2508
rect 4387 2468 5356 2496
rect 4387 2465 4399 2468
rect 4341 2459 4399 2465
rect 5350 2456 5356 2468
rect 5408 2456 5414 2508
rect 5629 2499 5687 2505
rect 5629 2465 5641 2499
rect 5675 2496 5687 2499
rect 6288 2496 6316 2595
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 7745 2635 7803 2641
rect 7745 2601 7757 2635
rect 7791 2632 7803 2635
rect 8202 2632 8208 2644
rect 7791 2604 8208 2632
rect 7791 2601 7803 2604
rect 7745 2595 7803 2601
rect 5675 2468 6316 2496
rect 6917 2499 6975 2505
rect 5675 2465 5687 2468
rect 5629 2459 5687 2465
rect 6917 2465 6929 2499
rect 6963 2496 6975 2499
rect 7760 2496 7788 2595
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 16850 2632 16856 2644
rect 16811 2604 16856 2632
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 17770 2632 17776 2644
rect 17731 2604 17776 2632
rect 17770 2592 17776 2604
rect 17828 2592 17834 2644
rect 22554 2632 22560 2644
rect 22515 2604 22560 2632
rect 22554 2592 22560 2604
rect 22612 2592 22618 2644
rect 6963 2468 7788 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 8110 2456 8116 2508
rect 8168 2496 8174 2508
rect 8205 2499 8263 2505
rect 8205 2496 8217 2499
rect 8168 2468 8217 2496
rect 8168 2456 8174 2468
rect 8205 2465 8217 2468
rect 8251 2496 8263 2499
rect 8941 2499 8999 2505
rect 8941 2496 8953 2499
rect 8251 2468 8953 2496
rect 8251 2465 8263 2468
rect 8205 2459 8263 2465
rect 8941 2465 8953 2468
rect 8987 2465 8999 2499
rect 9766 2496 9772 2508
rect 9727 2468 9772 2496
rect 8941 2459 8999 2465
rect 9766 2456 9772 2468
rect 9824 2496 9830 2508
rect 10505 2499 10563 2505
rect 10505 2496 10517 2499
rect 9824 2468 10517 2496
rect 9824 2456 9830 2468
rect 10505 2465 10517 2468
rect 10551 2465 10563 2499
rect 10505 2459 10563 2465
rect 12621 2499 12679 2505
rect 12621 2465 12633 2499
rect 12667 2496 12679 2499
rect 12710 2496 12716 2508
rect 12667 2468 12716 2496
rect 12667 2465 12679 2468
rect 12621 2459 12679 2465
rect 12710 2456 12716 2468
rect 12768 2496 12774 2508
rect 13357 2499 13415 2505
rect 13357 2496 13369 2499
rect 12768 2468 13369 2496
rect 12768 2456 12774 2468
rect 13357 2465 13369 2468
rect 13403 2465 13415 2499
rect 16868 2496 16896 2592
rect 16945 2499 17003 2505
rect 16945 2496 16957 2499
rect 16868 2468 16957 2496
rect 13357 2459 13415 2465
rect 16945 2465 16957 2468
rect 16991 2465 17003 2499
rect 16945 2459 17003 2465
rect 18230 2456 18236 2508
rect 18288 2496 18294 2508
rect 19153 2499 19211 2505
rect 19153 2496 19165 2499
rect 18288 2468 19165 2496
rect 18288 2456 18294 2468
rect 19153 2465 19165 2468
rect 19199 2496 19211 2499
rect 19889 2499 19947 2505
rect 19889 2496 19901 2499
rect 19199 2468 19901 2496
rect 19199 2465 19211 2468
rect 19153 2459 19211 2465
rect 19889 2465 19901 2468
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 21821 2499 21879 2505
rect 21821 2465 21833 2499
rect 21867 2496 21879 2499
rect 22572 2496 22600 2592
rect 24026 2496 24032 2508
rect 21867 2468 22600 2496
rect 23987 2468 24032 2496
rect 21867 2465 21879 2468
rect 21821 2459 21879 2465
rect 24026 2456 24032 2468
rect 24084 2496 24090 2508
rect 24765 2499 24823 2505
rect 24765 2496 24777 2499
rect 24084 2468 24777 2496
rect 24084 2456 24090 2468
rect 24765 2465 24777 2468
rect 24811 2465 24823 2499
rect 25682 2496 25688 2508
rect 25643 2468 25688 2496
rect 24765 2459 24823 2465
rect 25682 2456 25688 2468
rect 25740 2496 25746 2508
rect 26237 2499 26295 2505
rect 26237 2496 26249 2499
rect 25740 2468 26249 2496
rect 25740 2456 25746 2468
rect 26237 2465 26249 2468
rect 26283 2465 26295 2499
rect 26237 2459 26295 2465
rect 2409 2431 2467 2437
rect 2409 2397 2421 2431
rect 2455 2428 2467 2431
rect 3510 2428 3516 2440
rect 2455 2400 3516 2428
rect 2455 2397 2467 2400
rect 2409 2391 2467 2397
rect 3510 2388 3516 2400
rect 3568 2388 3574 2440
rect 4617 2431 4675 2437
rect 4617 2397 4629 2431
rect 4663 2428 4675 2431
rect 4890 2428 4896 2440
rect 4663 2400 4896 2428
rect 4663 2397 4675 2400
rect 4617 2391 4675 2397
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 6362 2388 6368 2440
rect 6420 2428 6426 2440
rect 7101 2431 7159 2437
rect 7101 2428 7113 2431
rect 6420 2400 7113 2428
rect 6420 2388 6426 2400
rect 7101 2397 7113 2400
rect 7147 2397 7159 2431
rect 7101 2391 7159 2397
rect 8481 2431 8539 2437
rect 8481 2397 8493 2431
rect 8527 2428 8539 2431
rect 9214 2428 9220 2440
rect 8527 2400 9220 2428
rect 8527 2397 8539 2400
rect 8481 2391 8539 2397
rect 9214 2388 9220 2400
rect 9272 2388 9278 2440
rect 10045 2431 10103 2437
rect 10045 2397 10057 2431
rect 10091 2428 10103 2431
rect 10594 2428 10600 2440
rect 10091 2400 10600 2428
rect 10091 2397 10103 2400
rect 10045 2391 10103 2397
rect 10594 2388 10600 2400
rect 10652 2388 10658 2440
rect 12066 2388 12072 2440
rect 12124 2428 12130 2440
rect 12805 2431 12863 2437
rect 12805 2428 12817 2431
rect 12124 2400 12817 2428
rect 12124 2388 12130 2400
rect 12805 2397 12817 2400
rect 12851 2397 12863 2431
rect 12805 2391 12863 2397
rect 17221 2431 17279 2437
rect 17221 2397 17233 2431
rect 17267 2428 17279 2431
rect 17770 2428 17776 2440
rect 17267 2400 17776 2428
rect 17267 2397 17279 2400
rect 17221 2391 17279 2397
rect 17770 2388 17776 2400
rect 17828 2388 17834 2440
rect 19429 2431 19487 2437
rect 19429 2397 19441 2431
rect 19475 2428 19487 2431
rect 20622 2428 20628 2440
rect 19475 2400 20628 2428
rect 19475 2397 19487 2400
rect 19429 2391 19487 2397
rect 20622 2388 20628 2400
rect 20680 2388 20686 2440
rect 22002 2388 22008 2440
rect 22060 2428 22066 2440
rect 22097 2431 22155 2437
rect 22097 2428 22109 2431
rect 22060 2400 22109 2428
rect 22060 2388 22066 2400
rect 22097 2397 22109 2400
rect 22143 2397 22155 2431
rect 22097 2391 22155 2397
rect 23474 2388 23480 2440
rect 23532 2428 23538 2440
rect 24213 2431 24271 2437
rect 24213 2428 24225 2431
rect 23532 2400 24225 2428
rect 23532 2388 23538 2400
rect 24213 2397 24225 2400
rect 24259 2397 24271 2431
rect 24213 2391 24271 2397
rect 5810 2292 5816 2304
rect 5771 2264 5816 2292
rect 5810 2252 5816 2264
rect 5868 2252 5874 2304
rect 25866 2292 25872 2304
rect 25827 2264 25872 2292
rect 25866 2252 25872 2264
rect 25924 2252 25930 2304
rect 27065 2295 27123 2301
rect 27065 2261 27077 2295
rect 27111 2292 27123 2295
rect 29178 2292 29184 2304
rect 27111 2264 29184 2292
rect 27111 2261 27123 2264
rect 27065 2255 27123 2261
rect 29178 2252 29184 2264
rect 29236 2252 29242 2304
rect 1104 2202 28888 2224
rect 1104 2150 5982 2202
rect 6034 2150 6046 2202
rect 6098 2150 6110 2202
rect 6162 2150 6174 2202
rect 6226 2150 15982 2202
rect 16034 2150 16046 2202
rect 16098 2150 16110 2202
rect 16162 2150 16174 2202
rect 16226 2150 25982 2202
rect 26034 2150 26046 2202
rect 26098 2150 26110 2202
rect 26162 2150 26174 2202
rect 26226 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 3976 22176 4028 22228
rect 12532 22176 12584 22228
rect 21456 22108 21508 22160
rect 25780 22108 25832 22160
rect 5982 21734 6034 21786
rect 6046 21734 6098 21786
rect 6110 21734 6162 21786
rect 6174 21734 6226 21786
rect 15982 21734 16034 21786
rect 16046 21734 16098 21786
rect 16110 21734 16162 21786
rect 16174 21734 16226 21786
rect 25982 21734 26034 21786
rect 26046 21734 26098 21786
rect 26110 21734 26162 21786
rect 26174 21734 26226 21786
rect 10982 21190 11034 21242
rect 11046 21190 11098 21242
rect 11110 21190 11162 21242
rect 11174 21190 11226 21242
rect 20982 21190 21034 21242
rect 21046 21190 21098 21242
rect 21110 21190 21162 21242
rect 21174 21190 21226 21242
rect 10508 20952 10560 21004
rect 22376 20952 22428 21004
rect 10140 20927 10192 20936
rect 10140 20893 10149 20927
rect 10149 20893 10183 20927
rect 10183 20893 10192 20927
rect 10140 20884 10192 20893
rect 10232 20927 10284 20936
rect 10232 20893 10241 20927
rect 10241 20893 10275 20927
rect 10275 20893 10284 20927
rect 10232 20884 10284 20893
rect 19708 20884 19760 20936
rect 22284 20927 22336 20936
rect 22284 20893 22293 20927
rect 22293 20893 22327 20927
rect 22327 20893 22336 20927
rect 22284 20884 22336 20893
rect 4068 20816 4120 20868
rect 9956 20816 10008 20868
rect 8760 20791 8812 20800
rect 8760 20757 8769 20791
rect 8769 20757 8803 20791
rect 8803 20757 8812 20791
rect 8760 20748 8812 20757
rect 8852 20748 8904 20800
rect 22652 20748 22704 20800
rect 5982 20646 6034 20698
rect 6046 20646 6098 20698
rect 6110 20646 6162 20698
rect 6174 20646 6226 20698
rect 15982 20646 16034 20698
rect 16046 20646 16098 20698
rect 16110 20646 16162 20698
rect 16174 20646 16226 20698
rect 25982 20646 26034 20698
rect 26046 20646 26098 20698
rect 26110 20646 26162 20698
rect 26174 20646 26226 20698
rect 8208 20544 8260 20596
rect 10140 20544 10192 20596
rect 22376 20587 22428 20596
rect 22376 20553 22385 20587
rect 22385 20553 22419 20587
rect 22419 20553 22428 20587
rect 22376 20544 22428 20553
rect 28264 20544 28316 20596
rect 11612 20476 11664 20528
rect 8760 20451 8812 20460
rect 8760 20417 8769 20451
rect 8769 20417 8803 20451
rect 8803 20417 8812 20451
rect 8760 20408 8812 20417
rect 10784 20340 10836 20392
rect 9312 20272 9364 20324
rect 10508 20272 10560 20324
rect 22284 20476 22336 20528
rect 12440 20451 12492 20460
rect 12440 20417 12449 20451
rect 12449 20417 12483 20451
rect 12483 20417 12492 20451
rect 16120 20451 16172 20460
rect 12440 20408 12492 20417
rect 16120 20417 16129 20451
rect 16129 20417 16163 20451
rect 16163 20417 16172 20451
rect 16120 20408 16172 20417
rect 19708 20451 19760 20460
rect 19708 20417 19717 20451
rect 19717 20417 19751 20451
rect 19751 20417 19760 20451
rect 19708 20408 19760 20417
rect 15844 20383 15896 20392
rect 15844 20349 15853 20383
rect 15853 20349 15887 20383
rect 15887 20349 15896 20383
rect 15844 20340 15896 20349
rect 20720 20272 20772 20324
rect 9680 20204 9732 20256
rect 10232 20204 10284 20256
rect 13820 20247 13872 20256
rect 13820 20213 13829 20247
rect 13829 20213 13863 20247
rect 13863 20213 13872 20247
rect 13820 20204 13872 20213
rect 20812 20204 20864 20256
rect 26056 20247 26108 20256
rect 26056 20213 26065 20247
rect 26065 20213 26099 20247
rect 26099 20213 26108 20247
rect 26056 20204 26108 20213
rect 27252 20204 27304 20256
rect 27436 20204 27488 20256
rect 10982 20102 11034 20154
rect 11046 20102 11098 20154
rect 11110 20102 11162 20154
rect 11174 20102 11226 20154
rect 20982 20102 21034 20154
rect 21046 20102 21098 20154
rect 21110 20102 21162 20154
rect 21174 20102 21226 20154
rect 8024 20043 8076 20052
rect 8024 20009 8033 20043
rect 8033 20009 8067 20043
rect 8067 20009 8076 20043
rect 8024 20000 8076 20009
rect 8484 20000 8536 20052
rect 8852 20000 8904 20052
rect 10508 20043 10560 20052
rect 10508 20009 10517 20043
rect 10517 20009 10551 20043
rect 10551 20009 10560 20043
rect 10508 20000 10560 20009
rect 12440 20043 12492 20052
rect 12440 20009 12449 20043
rect 12449 20009 12483 20043
rect 12483 20009 12492 20043
rect 12440 20000 12492 20009
rect 21640 20000 21692 20052
rect 5724 19864 5776 19916
rect 8852 19864 8904 19916
rect 10784 19864 10836 19916
rect 12440 19864 12492 19916
rect 13820 19864 13872 19916
rect 20812 19864 20864 19916
rect 22284 19864 22336 19916
rect 22836 19907 22888 19916
rect 22836 19873 22845 19907
rect 22845 19873 22879 19907
rect 22879 19873 22888 19907
rect 22836 19864 22888 19873
rect 23112 19907 23164 19916
rect 23112 19873 23146 19907
rect 23146 19873 23164 19907
rect 23112 19864 23164 19873
rect 1676 19796 1728 19848
rect 2688 19796 2740 19848
rect 5632 19839 5684 19848
rect 5632 19805 5641 19839
rect 5641 19805 5675 19839
rect 5675 19805 5684 19839
rect 5632 19796 5684 19805
rect 8576 19839 8628 19848
rect 8576 19805 8585 19839
rect 8585 19805 8619 19839
rect 8619 19805 8628 19839
rect 8576 19796 8628 19805
rect 10968 19839 11020 19848
rect 10968 19805 10977 19839
rect 10977 19805 11011 19839
rect 11011 19805 11020 19839
rect 10968 19796 11020 19805
rect 10876 19728 10928 19780
rect 12624 19796 12676 19848
rect 14188 19771 14240 19780
rect 14188 19737 14197 19771
rect 14197 19737 14231 19771
rect 14231 19737 14240 19771
rect 14188 19728 14240 19737
rect 7104 19660 7156 19712
rect 10600 19660 10652 19712
rect 16488 19660 16540 19712
rect 19616 19703 19668 19712
rect 19616 19669 19625 19703
rect 19625 19669 19659 19703
rect 19659 19669 19668 19703
rect 19616 19660 19668 19669
rect 22100 19703 22152 19712
rect 22100 19669 22109 19703
rect 22109 19669 22143 19703
rect 22143 19669 22152 19703
rect 24216 19703 24268 19712
rect 22100 19660 22152 19669
rect 24216 19669 24225 19703
rect 24225 19669 24259 19703
rect 24259 19669 24268 19703
rect 24216 19660 24268 19669
rect 25412 19660 25464 19712
rect 5982 19558 6034 19610
rect 6046 19558 6098 19610
rect 6110 19558 6162 19610
rect 6174 19558 6226 19610
rect 15982 19558 16034 19610
rect 16046 19558 16098 19610
rect 16110 19558 16162 19610
rect 16174 19558 16226 19610
rect 25982 19558 26034 19610
rect 26046 19558 26098 19610
rect 26110 19558 26162 19610
rect 26174 19558 26226 19610
rect 5724 19499 5776 19508
rect 5724 19465 5733 19499
rect 5733 19465 5767 19499
rect 5767 19465 5776 19499
rect 5724 19456 5776 19465
rect 10140 19499 10192 19508
rect 10140 19465 10149 19499
rect 10149 19465 10183 19499
rect 10183 19465 10192 19499
rect 10140 19456 10192 19465
rect 20812 19456 20864 19508
rect 22376 19456 22428 19508
rect 23572 19456 23624 19508
rect 24216 19456 24268 19508
rect 10048 19388 10100 19440
rect 10968 19388 11020 19440
rect 9312 19363 9364 19372
rect 6828 19295 6880 19304
rect 6828 19261 6837 19295
rect 6837 19261 6871 19295
rect 6871 19261 6880 19295
rect 6828 19252 6880 19261
rect 9312 19329 9321 19363
rect 9321 19329 9355 19363
rect 9355 19329 9364 19363
rect 9312 19320 9364 19329
rect 10876 19320 10928 19372
rect 9956 19295 10008 19304
rect 5724 19184 5776 19236
rect 9956 19261 9965 19295
rect 9965 19261 9999 19295
rect 9999 19261 10008 19295
rect 10508 19295 10560 19304
rect 9956 19252 10008 19261
rect 10508 19261 10517 19295
rect 10517 19261 10551 19295
rect 10551 19261 10560 19295
rect 10508 19252 10560 19261
rect 5632 19116 5684 19168
rect 6920 19116 6972 19168
rect 8024 19184 8076 19236
rect 12624 19184 12676 19236
rect 8576 19116 8628 19168
rect 8852 19159 8904 19168
rect 8852 19125 8861 19159
rect 8861 19125 8895 19159
rect 8895 19125 8904 19159
rect 8852 19116 8904 19125
rect 10600 19159 10652 19168
rect 10600 19125 10609 19159
rect 10609 19125 10643 19159
rect 10643 19125 10652 19159
rect 10600 19116 10652 19125
rect 12440 19116 12492 19168
rect 15200 19116 15252 19168
rect 19616 19363 19668 19372
rect 19616 19329 19625 19363
rect 19625 19329 19659 19363
rect 19659 19329 19668 19363
rect 19616 19320 19668 19329
rect 22652 19363 22704 19372
rect 20720 19252 20772 19304
rect 22652 19329 22661 19363
rect 22661 19329 22695 19363
rect 22695 19329 22704 19363
rect 22652 19320 22704 19329
rect 25504 19431 25556 19440
rect 25504 19397 25513 19431
rect 25513 19397 25547 19431
rect 25547 19397 25556 19431
rect 25504 19388 25556 19397
rect 24952 19320 25004 19372
rect 25228 19320 25280 19372
rect 25412 19320 25464 19372
rect 22100 19252 22152 19304
rect 15844 19184 15896 19236
rect 15752 19116 15804 19168
rect 19984 19184 20036 19236
rect 24584 19252 24636 19304
rect 27528 19295 27580 19304
rect 16488 19116 16540 19168
rect 16856 19116 16908 19168
rect 21272 19116 21324 19168
rect 21732 19116 21784 19168
rect 22468 19159 22520 19168
rect 22468 19125 22477 19159
rect 22477 19125 22511 19159
rect 22511 19125 22520 19159
rect 22468 19116 22520 19125
rect 23112 19159 23164 19168
rect 23112 19125 23121 19159
rect 23121 19125 23155 19159
rect 23155 19125 23164 19159
rect 23112 19116 23164 19125
rect 24124 19184 24176 19236
rect 25504 19184 25556 19236
rect 25688 19184 25740 19236
rect 25320 19159 25372 19168
rect 25320 19125 25329 19159
rect 25329 19125 25363 19159
rect 25363 19125 25372 19159
rect 25320 19116 25372 19125
rect 26424 19116 26476 19168
rect 27528 19261 27537 19295
rect 27537 19261 27571 19295
rect 27571 19261 27580 19295
rect 27528 19252 27580 19261
rect 26976 19227 27028 19236
rect 26976 19193 26985 19227
rect 26985 19193 27019 19227
rect 27019 19193 27028 19227
rect 26976 19184 27028 19193
rect 27160 19116 27212 19168
rect 10982 19014 11034 19066
rect 11046 19014 11098 19066
rect 11110 19014 11162 19066
rect 11174 19014 11226 19066
rect 20982 19014 21034 19066
rect 21046 19014 21098 19066
rect 21110 19014 21162 19066
rect 21174 19014 21226 19066
rect 8484 18955 8536 18964
rect 8484 18921 8493 18955
rect 8493 18921 8527 18955
rect 8527 18921 8536 18955
rect 8484 18912 8536 18921
rect 10784 18955 10836 18964
rect 10784 18921 10793 18955
rect 10793 18921 10827 18955
rect 10827 18921 10836 18955
rect 10784 18912 10836 18921
rect 22468 18912 22520 18964
rect 24124 18955 24176 18964
rect 24124 18921 24133 18955
rect 24133 18921 24167 18955
rect 24167 18921 24176 18955
rect 24124 18912 24176 18921
rect 24584 18912 24636 18964
rect 27160 18955 27212 18964
rect 27160 18921 27169 18955
rect 27169 18921 27203 18955
rect 27203 18921 27212 18955
rect 27160 18912 27212 18921
rect 22836 18887 22888 18896
rect 22836 18853 22845 18887
rect 22845 18853 22879 18887
rect 22879 18853 22888 18887
rect 22836 18844 22888 18853
rect 4252 18776 4304 18828
rect 9772 18776 9824 18828
rect 15200 18776 15252 18828
rect 23296 18776 23348 18828
rect 23480 18819 23532 18828
rect 23480 18785 23489 18819
rect 23489 18785 23523 18819
rect 23523 18785 23532 18819
rect 23480 18776 23532 18785
rect 4528 18751 4580 18760
rect 4528 18717 4537 18751
rect 4537 18717 4571 18751
rect 4571 18717 4580 18751
rect 4528 18708 4580 18717
rect 4804 18708 4856 18760
rect 10140 18751 10192 18760
rect 10140 18717 10149 18751
rect 10149 18717 10183 18751
rect 10183 18717 10192 18751
rect 10140 18708 10192 18717
rect 10876 18708 10928 18760
rect 15292 18751 15344 18760
rect 15292 18717 15301 18751
rect 15301 18717 15335 18751
rect 15335 18717 15344 18751
rect 15292 18708 15344 18717
rect 20444 18708 20496 18760
rect 23572 18751 23624 18760
rect 23572 18717 23581 18751
rect 23581 18717 23615 18751
rect 23615 18717 23624 18751
rect 23572 18708 23624 18717
rect 8392 18640 8444 18692
rect 4160 18572 4212 18624
rect 5080 18615 5132 18624
rect 5080 18581 5089 18615
rect 5089 18581 5123 18615
rect 5123 18581 5132 18615
rect 5080 18572 5132 18581
rect 6920 18615 6972 18624
rect 6920 18581 6929 18615
rect 6929 18581 6963 18615
rect 6963 18581 6972 18615
rect 6920 18572 6972 18581
rect 7196 18572 7248 18624
rect 12624 18572 12676 18624
rect 16672 18615 16724 18624
rect 16672 18581 16681 18615
rect 16681 18581 16715 18615
rect 16715 18581 16724 18615
rect 16672 18572 16724 18581
rect 25688 18572 25740 18624
rect 5982 18470 6034 18522
rect 6046 18470 6098 18522
rect 6110 18470 6162 18522
rect 6174 18470 6226 18522
rect 15982 18470 16034 18522
rect 16046 18470 16098 18522
rect 16110 18470 16162 18522
rect 16174 18470 16226 18522
rect 25982 18470 26034 18522
rect 26046 18470 26098 18522
rect 26110 18470 26162 18522
rect 26174 18470 26226 18522
rect 4528 18368 4580 18420
rect 5356 18411 5408 18420
rect 5356 18377 5365 18411
rect 5365 18377 5399 18411
rect 5399 18377 5408 18411
rect 5356 18368 5408 18377
rect 8852 18368 8904 18420
rect 3976 18232 4028 18284
rect 4804 18232 4856 18284
rect 8208 18232 8260 18284
rect 2228 18164 2280 18216
rect 4068 18164 4120 18216
rect 5080 18164 5132 18216
rect 8392 18164 8444 18216
rect 2780 18096 2832 18148
rect 4252 18096 4304 18148
rect 8024 18139 8076 18148
rect 8024 18105 8033 18139
rect 8033 18105 8067 18139
rect 8067 18105 8076 18139
rect 9588 18232 9640 18284
rect 10876 18368 10928 18420
rect 18880 18411 18932 18420
rect 18880 18377 18889 18411
rect 18889 18377 18923 18411
rect 18923 18377 18932 18411
rect 20444 18411 20496 18420
rect 18880 18368 18932 18377
rect 15844 18275 15896 18284
rect 15844 18241 15853 18275
rect 15853 18241 15887 18275
rect 15887 18241 15896 18275
rect 15844 18232 15896 18241
rect 10324 18164 10376 18216
rect 12624 18164 12676 18216
rect 8024 18096 8076 18105
rect 10232 18096 10284 18148
rect 14464 18164 14516 18216
rect 16672 18232 16724 18284
rect 20444 18377 20453 18411
rect 20453 18377 20487 18411
rect 20487 18377 20496 18411
rect 20444 18368 20496 18377
rect 23572 18368 23624 18420
rect 20720 18300 20772 18352
rect 19984 18275 20036 18284
rect 19984 18241 19993 18275
rect 19993 18241 20027 18275
rect 20027 18241 20036 18275
rect 19984 18232 20036 18241
rect 20812 18232 20864 18284
rect 19340 18207 19392 18216
rect 19340 18173 19349 18207
rect 19349 18173 19383 18207
rect 19383 18173 19392 18207
rect 19340 18164 19392 18173
rect 18604 18139 18656 18148
rect 18604 18105 18613 18139
rect 18613 18105 18647 18139
rect 18647 18105 18656 18139
rect 20444 18164 20496 18216
rect 18604 18096 18656 18105
rect 23296 18096 23348 18148
rect 3516 18071 3568 18080
rect 3516 18037 3525 18071
rect 3525 18037 3559 18071
rect 3559 18037 3568 18071
rect 3516 18028 3568 18037
rect 4436 18028 4488 18080
rect 5172 18028 5224 18080
rect 9680 18028 9732 18080
rect 13820 18028 13872 18080
rect 15200 18071 15252 18080
rect 15200 18037 15209 18071
rect 15209 18037 15243 18071
rect 15243 18037 15252 18071
rect 15200 18028 15252 18037
rect 15384 18071 15436 18080
rect 15384 18037 15393 18071
rect 15393 18037 15427 18071
rect 15427 18037 15436 18071
rect 15384 18028 15436 18037
rect 16212 18028 16264 18080
rect 16948 18071 17000 18080
rect 16948 18037 16957 18071
rect 16957 18037 16991 18071
rect 16991 18037 17000 18071
rect 16948 18028 17000 18037
rect 19708 18028 19760 18080
rect 21364 18028 21416 18080
rect 23480 18071 23532 18080
rect 23480 18037 23489 18071
rect 23489 18037 23523 18071
rect 23523 18037 23532 18071
rect 23480 18028 23532 18037
rect 24768 18028 24820 18080
rect 10982 17926 11034 17978
rect 11046 17926 11098 17978
rect 11110 17926 11162 17978
rect 11174 17926 11226 17978
rect 20982 17926 21034 17978
rect 21046 17926 21098 17978
rect 21110 17926 21162 17978
rect 21174 17926 21226 17978
rect 4068 17824 4120 17876
rect 4160 17824 4212 17876
rect 4620 17824 4672 17876
rect 8208 17867 8260 17876
rect 8208 17833 8217 17867
rect 8217 17833 8251 17867
rect 8251 17833 8260 17867
rect 8208 17824 8260 17833
rect 10232 17867 10284 17876
rect 10232 17833 10241 17867
rect 10241 17833 10275 17867
rect 10275 17833 10284 17867
rect 10232 17824 10284 17833
rect 13268 17867 13320 17876
rect 13268 17833 13277 17867
rect 13277 17833 13311 17867
rect 13311 17833 13320 17867
rect 13268 17824 13320 17833
rect 16212 17867 16264 17876
rect 16212 17833 16221 17867
rect 16221 17833 16255 17867
rect 16255 17833 16264 17867
rect 16212 17824 16264 17833
rect 19708 17867 19760 17876
rect 19708 17833 19717 17867
rect 19717 17833 19751 17867
rect 19751 17833 19760 17867
rect 19708 17824 19760 17833
rect 20812 17824 20864 17876
rect 23296 17824 23348 17876
rect 24860 17867 24912 17876
rect 24860 17833 24869 17867
rect 24869 17833 24903 17867
rect 24903 17833 24912 17867
rect 24860 17824 24912 17833
rect 2780 17756 2832 17808
rect 3976 17756 4028 17808
rect 16672 17799 16724 17808
rect 16672 17765 16681 17799
rect 16681 17765 16715 17799
rect 16715 17765 16724 17799
rect 16672 17756 16724 17765
rect 24676 17756 24728 17808
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 4436 17731 4488 17740
rect 4436 17697 4445 17731
rect 4445 17697 4479 17731
rect 4479 17697 4488 17731
rect 4436 17688 4488 17697
rect 6368 17731 6420 17740
rect 3516 17620 3568 17672
rect 4344 17620 4396 17672
rect 6368 17697 6402 17731
rect 6402 17697 6420 17731
rect 6368 17688 6420 17697
rect 10140 17688 10192 17740
rect 10600 17731 10652 17740
rect 10600 17697 10609 17731
rect 10609 17697 10643 17731
rect 10643 17697 10652 17731
rect 10600 17688 10652 17697
rect 10784 17688 10836 17740
rect 16948 17688 17000 17740
rect 20628 17688 20680 17740
rect 23204 17688 23256 17740
rect 24860 17688 24912 17740
rect 5172 17663 5224 17672
rect 5172 17629 5181 17663
rect 5181 17629 5215 17663
rect 5215 17629 5224 17663
rect 5172 17620 5224 17629
rect 5724 17620 5776 17672
rect 10876 17663 10928 17672
rect 10876 17629 10885 17663
rect 10885 17629 10919 17663
rect 10919 17629 10928 17663
rect 10876 17620 10928 17629
rect 13360 17663 13412 17672
rect 13360 17629 13369 17663
rect 13369 17629 13403 17663
rect 13403 17629 13412 17663
rect 13360 17620 13412 17629
rect 13728 17620 13780 17672
rect 16764 17663 16816 17672
rect 16764 17629 16773 17663
rect 16773 17629 16807 17663
rect 16807 17629 16816 17663
rect 16764 17620 16816 17629
rect 19800 17620 19852 17672
rect 21272 17620 21324 17672
rect 23480 17663 23532 17672
rect 23480 17629 23489 17663
rect 23489 17629 23523 17663
rect 23523 17629 23532 17663
rect 23480 17620 23532 17629
rect 25412 17663 25464 17672
rect 16396 17552 16448 17604
rect 23112 17552 23164 17604
rect 25412 17629 25421 17663
rect 25421 17629 25455 17663
rect 25455 17629 25464 17663
rect 25412 17620 25464 17629
rect 1400 17484 1452 17536
rect 2320 17484 2372 17536
rect 4068 17527 4120 17536
rect 4068 17493 4077 17527
rect 4077 17493 4111 17527
rect 4111 17493 4120 17527
rect 4068 17484 4120 17493
rect 7472 17527 7524 17536
rect 7472 17493 7481 17527
rect 7481 17493 7515 17527
rect 7515 17493 7524 17527
rect 7472 17484 7524 17493
rect 10416 17484 10468 17536
rect 12716 17484 12768 17536
rect 13820 17484 13872 17536
rect 15292 17484 15344 17536
rect 16304 17484 16356 17536
rect 19524 17484 19576 17536
rect 25780 17484 25832 17536
rect 5982 17382 6034 17434
rect 6046 17382 6098 17434
rect 6110 17382 6162 17434
rect 6174 17382 6226 17434
rect 15982 17382 16034 17434
rect 16046 17382 16098 17434
rect 16110 17382 16162 17434
rect 16174 17382 16226 17434
rect 25982 17382 26034 17434
rect 26046 17382 26098 17434
rect 26110 17382 26162 17434
rect 26174 17382 26226 17434
rect 2044 17323 2096 17332
rect 2044 17289 2053 17323
rect 2053 17289 2087 17323
rect 2087 17289 2096 17323
rect 2044 17280 2096 17289
rect 4344 17323 4396 17332
rect 4344 17289 4353 17323
rect 4353 17289 4387 17323
rect 4387 17289 4396 17323
rect 4344 17280 4396 17289
rect 4436 17280 4488 17332
rect 6368 17280 6420 17332
rect 10140 17280 10192 17332
rect 13360 17323 13412 17332
rect 13360 17289 13369 17323
rect 13369 17289 13403 17323
rect 13403 17289 13412 17323
rect 13360 17280 13412 17289
rect 14464 17323 14516 17332
rect 14464 17289 14473 17323
rect 14473 17289 14507 17323
rect 14507 17289 14516 17323
rect 14464 17280 14516 17289
rect 16672 17323 16724 17332
rect 16672 17289 16681 17323
rect 16681 17289 16715 17323
rect 16715 17289 16724 17323
rect 16672 17280 16724 17289
rect 16948 17323 17000 17332
rect 16948 17289 16957 17323
rect 16957 17289 16991 17323
rect 16991 17289 17000 17323
rect 16948 17280 17000 17289
rect 19708 17280 19760 17332
rect 22744 17323 22796 17332
rect 3792 17212 3844 17264
rect 4620 17255 4672 17264
rect 4620 17221 4629 17255
rect 4629 17221 4663 17255
rect 4663 17221 4672 17255
rect 4620 17212 4672 17221
rect 9588 17255 9640 17264
rect 9588 17221 9597 17255
rect 9597 17221 9631 17255
rect 9631 17221 9640 17255
rect 9588 17212 9640 17221
rect 10600 17212 10652 17264
rect 10876 17212 10928 17264
rect 12348 17212 12400 17264
rect 13728 17212 13780 17264
rect 13268 17144 13320 17196
rect 16764 17212 16816 17264
rect 17500 17212 17552 17264
rect 18236 17212 18288 17264
rect 16396 17144 16448 17196
rect 22744 17289 22753 17323
rect 22753 17289 22787 17323
rect 22787 17289 22796 17323
rect 22744 17280 22796 17289
rect 23480 17280 23532 17332
rect 25412 17280 25464 17332
rect 20628 17255 20680 17264
rect 20628 17221 20637 17255
rect 20637 17221 20671 17255
rect 20671 17221 20680 17255
rect 20628 17212 20680 17221
rect 21272 17255 21324 17264
rect 21272 17221 21281 17255
rect 21281 17221 21315 17255
rect 21315 17221 21324 17255
rect 21272 17212 21324 17221
rect 23112 17212 23164 17264
rect 24216 17187 24268 17196
rect 2044 17076 2096 17128
rect 7196 17119 7248 17128
rect 4068 17008 4120 17060
rect 3240 16983 3292 16992
rect 3240 16949 3249 16983
rect 3249 16949 3283 16983
rect 3283 16949 3292 16983
rect 3240 16940 3292 16949
rect 3700 16983 3752 16992
rect 3700 16949 3709 16983
rect 3709 16949 3743 16983
rect 3743 16949 3752 16983
rect 3700 16940 3752 16949
rect 5724 16940 5776 16992
rect 7196 17085 7205 17119
rect 7205 17085 7239 17119
rect 7239 17085 7248 17119
rect 7196 17076 7248 17085
rect 19524 17119 19576 17128
rect 19524 17085 19533 17119
rect 19533 17085 19567 17119
rect 19567 17085 19576 17119
rect 19524 17076 19576 17085
rect 21364 17119 21416 17128
rect 21364 17085 21373 17119
rect 21373 17085 21407 17119
rect 21407 17085 21416 17119
rect 21364 17076 21416 17085
rect 24216 17153 24225 17187
rect 24225 17153 24259 17187
rect 24259 17153 24268 17187
rect 24216 17144 24268 17153
rect 25412 17144 25464 17196
rect 24768 17076 24820 17128
rect 7472 17051 7524 17060
rect 7472 17017 7484 17051
rect 7484 17017 7524 17051
rect 7472 17008 7524 17017
rect 11612 17008 11664 17060
rect 13452 17008 13504 17060
rect 19800 17008 19852 17060
rect 23480 17051 23532 17060
rect 23480 17017 23489 17051
rect 23489 17017 23523 17051
rect 23523 17017 23532 17051
rect 23480 17008 23532 17017
rect 25780 17008 25832 17060
rect 7012 16983 7064 16992
rect 7012 16949 7021 16983
rect 7021 16949 7055 16983
rect 7055 16949 7064 16983
rect 7012 16940 7064 16949
rect 8576 16983 8628 16992
rect 8576 16949 8585 16983
rect 8585 16949 8619 16983
rect 8619 16949 8628 16983
rect 8576 16940 8628 16949
rect 9864 16983 9916 16992
rect 9864 16949 9873 16983
rect 9873 16949 9907 16983
rect 9907 16949 9916 16983
rect 9864 16940 9916 16949
rect 10416 16983 10468 16992
rect 10416 16949 10425 16983
rect 10425 16949 10459 16983
rect 10459 16949 10468 16983
rect 10416 16940 10468 16949
rect 10784 16940 10836 16992
rect 13820 16983 13872 16992
rect 13820 16949 13829 16983
rect 13829 16949 13863 16983
rect 13863 16949 13872 16983
rect 13820 16940 13872 16949
rect 15384 16983 15436 16992
rect 15384 16949 15393 16983
rect 15393 16949 15427 16983
rect 15427 16949 15436 16983
rect 15384 16940 15436 16949
rect 15476 16940 15528 16992
rect 15844 16940 15896 16992
rect 18328 16983 18380 16992
rect 18328 16949 18337 16983
rect 18337 16949 18371 16983
rect 18371 16949 18380 16983
rect 18328 16940 18380 16949
rect 19616 16983 19668 16992
rect 19616 16949 19625 16983
rect 19625 16949 19659 16983
rect 19659 16949 19668 16983
rect 19616 16940 19668 16949
rect 23204 16940 23256 16992
rect 23664 16940 23716 16992
rect 10982 16838 11034 16890
rect 11046 16838 11098 16890
rect 11110 16838 11162 16890
rect 11174 16838 11226 16890
rect 20982 16838 21034 16890
rect 21046 16838 21098 16890
rect 21110 16838 21162 16890
rect 21174 16838 21226 16890
rect 1492 16736 1544 16788
rect 3700 16736 3752 16788
rect 4068 16779 4120 16788
rect 4068 16745 4077 16779
rect 4077 16745 4111 16779
rect 4111 16745 4120 16779
rect 4068 16736 4120 16745
rect 4712 16736 4764 16788
rect 6828 16779 6880 16788
rect 6828 16745 6837 16779
rect 6837 16745 6871 16779
rect 6871 16745 6880 16779
rect 6828 16736 6880 16745
rect 7196 16736 7248 16788
rect 10324 16736 10376 16788
rect 13452 16779 13504 16788
rect 13452 16745 13461 16779
rect 13461 16745 13495 16779
rect 13495 16745 13504 16779
rect 13452 16736 13504 16745
rect 17500 16779 17552 16788
rect 17500 16745 17509 16779
rect 17509 16745 17543 16779
rect 17543 16745 17552 16779
rect 17500 16736 17552 16745
rect 18328 16736 18380 16788
rect 19616 16736 19668 16788
rect 21364 16779 21416 16788
rect 21364 16745 21373 16779
rect 21373 16745 21407 16779
rect 21407 16745 21416 16779
rect 21364 16736 21416 16745
rect 23112 16779 23164 16788
rect 23112 16745 23121 16779
rect 23121 16745 23155 16779
rect 23155 16745 23164 16779
rect 23112 16736 23164 16745
rect 24216 16736 24268 16788
rect 24860 16779 24912 16788
rect 24860 16745 24869 16779
rect 24869 16745 24903 16779
rect 24903 16745 24912 16779
rect 24860 16736 24912 16745
rect 25780 16736 25832 16788
rect 5816 16668 5868 16720
rect 13360 16668 13412 16720
rect 13636 16668 13688 16720
rect 13912 16668 13964 16720
rect 14464 16668 14516 16720
rect 5080 16600 5132 16652
rect 7012 16600 7064 16652
rect 10508 16643 10560 16652
rect 10508 16609 10517 16643
rect 10517 16609 10551 16643
rect 10551 16609 10560 16643
rect 10508 16600 10560 16609
rect 15844 16600 15896 16652
rect 16212 16600 16264 16652
rect 16396 16643 16448 16652
rect 16396 16609 16430 16643
rect 16430 16609 16448 16643
rect 16396 16600 16448 16609
rect 19432 16600 19484 16652
rect 23664 16643 23716 16652
rect 10600 16575 10652 16584
rect 3976 16464 4028 16516
rect 6460 16464 6512 16516
rect 10600 16541 10609 16575
rect 10609 16541 10643 16575
rect 10643 16541 10652 16575
rect 10600 16532 10652 16541
rect 10876 16532 10928 16584
rect 13360 16532 13412 16584
rect 14004 16575 14056 16584
rect 14004 16541 14013 16575
rect 14013 16541 14047 16575
rect 14047 16541 14056 16575
rect 19800 16575 19852 16584
rect 14004 16532 14056 16541
rect 19800 16541 19809 16575
rect 19809 16541 19843 16575
rect 19843 16541 19852 16575
rect 19800 16532 19852 16541
rect 23664 16609 23673 16643
rect 23673 16609 23707 16643
rect 23707 16609 23716 16643
rect 23664 16600 23716 16609
rect 24400 16600 24452 16652
rect 26516 16643 26568 16652
rect 26516 16609 26525 16643
rect 26525 16609 26559 16643
rect 26559 16609 26568 16643
rect 26516 16600 26568 16609
rect 20996 16532 21048 16584
rect 25320 16532 25372 16584
rect 25412 16464 25464 16516
rect 2320 16396 2372 16448
rect 3700 16439 3752 16448
rect 3700 16405 3709 16439
rect 3709 16405 3743 16439
rect 3743 16405 3752 16439
rect 3700 16396 3752 16405
rect 6368 16439 6420 16448
rect 6368 16405 6377 16439
rect 6377 16405 6411 16439
rect 6411 16405 6420 16439
rect 6368 16396 6420 16405
rect 15384 16396 15436 16448
rect 15844 16396 15896 16448
rect 18788 16396 18840 16448
rect 24676 16439 24728 16448
rect 24676 16405 24685 16439
rect 24685 16405 24719 16439
rect 24719 16405 24728 16439
rect 24676 16396 24728 16405
rect 5982 16294 6034 16346
rect 6046 16294 6098 16346
rect 6110 16294 6162 16346
rect 6174 16294 6226 16346
rect 15982 16294 16034 16346
rect 16046 16294 16098 16346
rect 16110 16294 16162 16346
rect 16174 16294 16226 16346
rect 25982 16294 26034 16346
rect 26046 16294 26098 16346
rect 26110 16294 26162 16346
rect 26174 16294 26226 16346
rect 3608 16235 3660 16244
rect 3608 16201 3617 16235
rect 3617 16201 3651 16235
rect 3651 16201 3660 16235
rect 3608 16192 3660 16201
rect 4712 16235 4764 16244
rect 4712 16201 4721 16235
rect 4721 16201 4755 16235
rect 4755 16201 4764 16235
rect 4712 16192 4764 16201
rect 5080 16235 5132 16244
rect 5080 16201 5089 16235
rect 5089 16201 5123 16235
rect 5123 16201 5132 16235
rect 5080 16192 5132 16201
rect 5816 16192 5868 16244
rect 6460 16235 6512 16244
rect 6460 16201 6469 16235
rect 6469 16201 6503 16235
rect 6503 16201 6512 16235
rect 6460 16192 6512 16201
rect 6920 16192 6972 16244
rect 10508 16235 10560 16244
rect 10508 16201 10517 16235
rect 10517 16201 10551 16235
rect 10551 16201 10560 16235
rect 10508 16192 10560 16201
rect 10876 16235 10928 16244
rect 10876 16201 10885 16235
rect 10885 16201 10919 16235
rect 10919 16201 10928 16235
rect 10876 16192 10928 16201
rect 13636 16192 13688 16244
rect 13820 16192 13872 16244
rect 18604 16235 18656 16244
rect 18604 16201 18613 16235
rect 18613 16201 18647 16235
rect 18647 16201 18656 16235
rect 18604 16192 18656 16201
rect 3976 16124 4028 16176
rect 3700 16056 3752 16108
rect 4068 16099 4120 16108
rect 4068 16065 4077 16099
rect 4077 16065 4111 16099
rect 4111 16065 4120 16099
rect 4068 16056 4120 16065
rect 10600 16124 10652 16176
rect 16120 16167 16172 16176
rect 13268 16056 13320 16108
rect 16120 16133 16129 16167
rect 16129 16133 16163 16167
rect 16163 16133 16172 16167
rect 16120 16124 16172 16133
rect 16396 16124 16448 16176
rect 19340 16167 19392 16176
rect 19340 16133 19349 16167
rect 19349 16133 19383 16167
rect 19383 16133 19392 16167
rect 19340 16124 19392 16133
rect 15476 16099 15528 16108
rect 15476 16065 15485 16099
rect 15485 16065 15519 16099
rect 15519 16065 15528 16099
rect 15476 16056 15528 16065
rect 8208 15988 8260 16040
rect 14004 15988 14056 16040
rect 15384 16031 15436 16040
rect 1676 15963 1728 15972
rect 1676 15929 1710 15963
rect 1710 15929 1728 15963
rect 1676 15920 1728 15929
rect 2320 15920 2372 15972
rect 2688 15920 2740 15972
rect 8760 15920 8812 15972
rect 15384 15997 15393 16031
rect 15393 15997 15427 16031
rect 15427 15997 15436 16031
rect 15384 15988 15436 15997
rect 20996 16235 21048 16244
rect 20996 16201 21005 16235
rect 21005 16201 21039 16235
rect 21039 16201 21048 16235
rect 20996 16192 21048 16201
rect 22652 16192 22704 16244
rect 22836 16192 22888 16244
rect 20720 16056 20772 16108
rect 24768 16192 24820 16244
rect 25412 16192 25464 16244
rect 25688 16235 25740 16244
rect 25688 16201 25697 16235
rect 25697 16201 25731 16235
rect 25731 16201 25740 16235
rect 25688 16192 25740 16201
rect 24676 16124 24728 16176
rect 26516 16192 26568 16244
rect 15200 15920 15252 15972
rect 25320 16031 25372 16040
rect 19892 15963 19944 15972
rect 19892 15929 19901 15963
rect 19901 15929 19935 15963
rect 19935 15929 19944 15963
rect 19892 15920 19944 15929
rect 3608 15852 3660 15904
rect 8392 15852 8444 15904
rect 9680 15852 9732 15904
rect 12808 15895 12860 15904
rect 12808 15861 12817 15895
rect 12817 15861 12851 15895
rect 12851 15861 12860 15895
rect 12808 15852 12860 15861
rect 13360 15895 13412 15904
rect 13360 15861 13369 15895
rect 13369 15861 13403 15895
rect 13403 15861 13412 15895
rect 13360 15852 13412 15861
rect 13636 15852 13688 15904
rect 16304 15852 16356 15904
rect 17776 15852 17828 15904
rect 18880 15895 18932 15904
rect 18880 15861 18889 15895
rect 18889 15861 18923 15895
rect 18923 15861 18932 15895
rect 18880 15852 18932 15861
rect 19432 15895 19484 15904
rect 19432 15861 19441 15895
rect 19441 15861 19475 15895
rect 19475 15861 19484 15895
rect 19432 15852 19484 15861
rect 19616 15852 19668 15904
rect 25320 15997 25329 16031
rect 25329 15997 25363 16031
rect 25363 15997 25372 16031
rect 25320 15988 25372 15997
rect 25412 15988 25464 16040
rect 21456 15895 21508 15904
rect 21456 15861 21465 15895
rect 21465 15861 21499 15895
rect 21499 15861 21508 15895
rect 21456 15852 21508 15861
rect 23756 15852 23808 15904
rect 26240 15895 26292 15904
rect 26240 15861 26249 15895
rect 26249 15861 26283 15895
rect 26283 15861 26292 15895
rect 26240 15852 26292 15861
rect 10982 15750 11034 15802
rect 11046 15750 11098 15802
rect 11110 15750 11162 15802
rect 11174 15750 11226 15802
rect 20982 15750 21034 15802
rect 21046 15750 21098 15802
rect 21110 15750 21162 15802
rect 21174 15750 21226 15802
rect 4068 15691 4120 15700
rect 4068 15657 4077 15691
rect 4077 15657 4111 15691
rect 4111 15657 4120 15691
rect 4068 15648 4120 15657
rect 4436 15691 4488 15700
rect 4436 15657 4445 15691
rect 4445 15657 4479 15691
rect 4479 15657 4488 15691
rect 4436 15648 4488 15657
rect 4528 15691 4580 15700
rect 4528 15657 4537 15691
rect 4537 15657 4571 15691
rect 4571 15657 4580 15691
rect 13268 15691 13320 15700
rect 4528 15648 4580 15657
rect 13268 15657 13277 15691
rect 13277 15657 13311 15691
rect 13311 15657 13320 15691
rect 13268 15648 13320 15657
rect 13360 15648 13412 15700
rect 15384 15648 15436 15700
rect 15752 15648 15804 15700
rect 16028 15691 16080 15700
rect 16028 15657 16037 15691
rect 16037 15657 16071 15691
rect 16071 15657 16080 15691
rect 16028 15648 16080 15657
rect 19432 15648 19484 15700
rect 19524 15648 19576 15700
rect 21364 15648 21416 15700
rect 21916 15648 21968 15700
rect 25136 15648 25188 15700
rect 25412 15648 25464 15700
rect 3976 15580 4028 15632
rect 11888 15580 11940 15632
rect 14004 15623 14056 15632
rect 14004 15589 14013 15623
rect 14013 15589 14047 15623
rect 14047 15589 14056 15623
rect 14004 15580 14056 15589
rect 15476 15580 15528 15632
rect 19800 15580 19852 15632
rect 22744 15580 22796 15632
rect 5816 15512 5868 15564
rect 6552 15512 6604 15564
rect 9680 15555 9732 15564
rect 9680 15521 9689 15555
rect 9689 15521 9723 15555
rect 9723 15521 9732 15555
rect 9680 15512 9732 15521
rect 9956 15555 10008 15564
rect 9956 15521 9990 15555
rect 9990 15521 10008 15555
rect 9956 15512 10008 15521
rect 13176 15512 13228 15564
rect 13636 15555 13688 15564
rect 13636 15521 13645 15555
rect 13645 15521 13679 15555
rect 13679 15521 13688 15555
rect 13636 15512 13688 15521
rect 17960 15512 18012 15564
rect 19248 15512 19300 15564
rect 19616 15555 19668 15564
rect 1860 15487 1912 15496
rect 1860 15453 1869 15487
rect 1869 15453 1903 15487
rect 1903 15453 1912 15487
rect 1860 15444 1912 15453
rect 1676 15419 1728 15428
rect 1676 15385 1685 15419
rect 1685 15385 1719 15419
rect 1719 15385 1728 15419
rect 5724 15444 5776 15496
rect 10692 15444 10744 15496
rect 11796 15444 11848 15496
rect 16120 15487 16172 15496
rect 16120 15453 16129 15487
rect 16129 15453 16163 15487
rect 16163 15453 16172 15487
rect 16120 15444 16172 15453
rect 16304 15444 16356 15496
rect 18880 15444 18932 15496
rect 19616 15521 19625 15555
rect 19625 15521 19659 15555
rect 19659 15521 19668 15555
rect 19616 15512 19668 15521
rect 21824 15555 21876 15564
rect 21824 15521 21833 15555
rect 21833 15521 21867 15555
rect 21867 15521 21876 15555
rect 21824 15512 21876 15521
rect 22652 15555 22704 15564
rect 22652 15521 22661 15555
rect 22661 15521 22695 15555
rect 22695 15521 22704 15555
rect 22652 15512 22704 15521
rect 26332 15512 26384 15564
rect 27344 15512 27396 15564
rect 19800 15487 19852 15496
rect 19800 15453 19809 15487
rect 19809 15453 19843 15487
rect 19843 15453 19852 15487
rect 19800 15444 19852 15453
rect 1676 15376 1728 15385
rect 4896 15376 4948 15428
rect 2320 15308 2372 15360
rect 5724 15351 5776 15360
rect 5724 15317 5733 15351
rect 5733 15317 5767 15351
rect 5767 15317 5776 15351
rect 5724 15308 5776 15317
rect 21456 15376 21508 15428
rect 24400 15376 24452 15428
rect 8392 15351 8444 15360
rect 8392 15317 8401 15351
rect 8401 15317 8435 15351
rect 8435 15317 8444 15351
rect 8392 15308 8444 15317
rect 11060 15351 11112 15360
rect 11060 15317 11069 15351
rect 11069 15317 11103 15351
rect 11103 15317 11112 15351
rect 11060 15308 11112 15317
rect 17776 15308 17828 15360
rect 21364 15308 21416 15360
rect 22652 15308 22704 15360
rect 24768 15308 24820 15360
rect 25412 15308 25464 15360
rect 26332 15308 26384 15360
rect 26792 15308 26844 15360
rect 5982 15206 6034 15258
rect 6046 15206 6098 15258
rect 6110 15206 6162 15258
rect 6174 15206 6226 15258
rect 15982 15206 16034 15258
rect 16046 15206 16098 15258
rect 16110 15206 16162 15258
rect 16174 15206 16226 15258
rect 25982 15206 26034 15258
rect 26046 15206 26098 15258
rect 26110 15206 26162 15258
rect 26174 15206 26226 15258
rect 4160 15104 4212 15156
rect 4436 15147 4488 15156
rect 4436 15113 4445 15147
rect 4445 15113 4479 15147
rect 4479 15113 4488 15147
rect 4436 15104 4488 15113
rect 4896 15147 4948 15156
rect 4896 15113 4905 15147
rect 4905 15113 4939 15147
rect 4939 15113 4948 15147
rect 4896 15104 4948 15113
rect 5724 15147 5776 15156
rect 5724 15113 5733 15147
rect 5733 15113 5767 15147
rect 5767 15113 5776 15147
rect 5724 15104 5776 15113
rect 5816 15104 5868 15156
rect 8208 15104 8260 15156
rect 8576 15104 8628 15156
rect 9680 15104 9732 15156
rect 10600 15104 10652 15156
rect 11796 15104 11848 15156
rect 12624 15147 12676 15156
rect 12624 15113 12633 15147
rect 12633 15113 12667 15147
rect 12667 15113 12676 15147
rect 12624 15104 12676 15113
rect 13820 15104 13872 15156
rect 15752 15104 15804 15156
rect 16304 15147 16356 15156
rect 16304 15113 16313 15147
rect 16313 15113 16347 15147
rect 16347 15113 16356 15147
rect 16304 15104 16356 15113
rect 17868 15147 17920 15156
rect 17868 15113 17877 15147
rect 17877 15113 17911 15147
rect 17911 15113 17920 15147
rect 17868 15104 17920 15113
rect 18880 15147 18932 15156
rect 18880 15113 18889 15147
rect 18889 15113 18923 15147
rect 18923 15113 18932 15147
rect 18880 15104 18932 15113
rect 19156 15147 19208 15156
rect 19156 15113 19165 15147
rect 19165 15113 19199 15147
rect 19199 15113 19208 15147
rect 19156 15104 19208 15113
rect 15292 15036 15344 15088
rect 15844 15036 15896 15088
rect 17960 15036 18012 15088
rect 2320 15011 2372 15020
rect 2320 14977 2329 15011
rect 2329 14977 2363 15011
rect 2363 14977 2372 15011
rect 2320 14968 2372 14977
rect 4344 14968 4396 15020
rect 4528 14968 4580 15020
rect 8392 15011 8444 15020
rect 8392 14977 8401 15011
rect 8401 14977 8435 15011
rect 8435 14977 8444 15011
rect 8392 14968 8444 14977
rect 17776 14968 17828 15020
rect 18880 14968 18932 15020
rect 19708 15104 19760 15156
rect 20720 15147 20772 15156
rect 20720 15113 20729 15147
rect 20729 15113 20763 15147
rect 20763 15113 20772 15147
rect 20720 15104 20772 15113
rect 21824 15104 21876 15156
rect 22744 15147 22796 15156
rect 22744 15113 22753 15147
rect 22753 15113 22787 15147
rect 22787 15113 22796 15147
rect 22744 15104 22796 15113
rect 24492 15104 24544 15156
rect 25872 15104 25924 15156
rect 27344 15147 27396 15156
rect 27344 15113 27353 15147
rect 27353 15113 27387 15147
rect 27387 15113 27396 15147
rect 27344 15104 27396 15113
rect 22652 15036 22704 15088
rect 25412 14968 25464 15020
rect 13820 14943 13872 14952
rect 13820 14909 13854 14943
rect 13854 14909 13872 14943
rect 2504 14832 2556 14884
rect 6552 14832 6604 14884
rect 8576 14832 8628 14884
rect 13820 14900 13872 14909
rect 13728 14832 13780 14884
rect 19800 14832 19852 14884
rect 25504 14832 25556 14884
rect 1676 14807 1728 14816
rect 1676 14773 1685 14807
rect 1685 14773 1719 14807
rect 1719 14773 1728 14807
rect 1676 14764 1728 14773
rect 1768 14764 1820 14816
rect 3700 14807 3752 14816
rect 3700 14773 3709 14807
rect 3709 14773 3743 14807
rect 3743 14773 3752 14807
rect 3700 14764 3752 14773
rect 9220 14764 9272 14816
rect 9956 14764 10008 14816
rect 11888 14807 11940 14816
rect 11888 14773 11897 14807
rect 11897 14773 11931 14807
rect 11931 14773 11940 14807
rect 11888 14764 11940 14773
rect 14924 14807 14976 14816
rect 14924 14773 14933 14807
rect 14933 14773 14967 14807
rect 14967 14773 14976 14807
rect 14924 14764 14976 14773
rect 24584 14764 24636 14816
rect 10982 14662 11034 14714
rect 11046 14662 11098 14714
rect 11110 14662 11162 14714
rect 11174 14662 11226 14714
rect 20982 14662 21034 14714
rect 21046 14662 21098 14714
rect 21110 14662 21162 14714
rect 21174 14662 21226 14714
rect 1768 14560 1820 14612
rect 1860 14560 1912 14612
rect 2964 14560 3016 14612
rect 8208 14560 8260 14612
rect 19800 14603 19852 14612
rect 19800 14569 19809 14603
rect 19809 14569 19843 14603
rect 19843 14569 19852 14603
rect 19800 14560 19852 14569
rect 25412 14560 25464 14612
rect 2596 14492 2648 14544
rect 3240 14492 3292 14544
rect 5816 14535 5868 14544
rect 5816 14501 5850 14535
rect 5850 14501 5868 14535
rect 5816 14492 5868 14501
rect 6828 14492 6880 14544
rect 10784 14492 10836 14544
rect 15200 14492 15252 14544
rect 5632 14424 5684 14476
rect 8300 14467 8352 14476
rect 8300 14433 8309 14467
rect 8309 14433 8343 14467
rect 8343 14433 8352 14467
rect 8300 14424 8352 14433
rect 10600 14467 10652 14476
rect 10600 14433 10609 14467
rect 10609 14433 10643 14467
rect 10643 14433 10652 14467
rect 10600 14424 10652 14433
rect 16304 14424 16356 14476
rect 18144 14424 18196 14476
rect 22652 14492 22704 14544
rect 22376 14424 22428 14476
rect 24584 14424 24636 14476
rect 2504 14399 2556 14408
rect 2504 14365 2513 14399
rect 2513 14365 2547 14399
rect 2547 14365 2556 14399
rect 2504 14356 2556 14365
rect 15844 14399 15896 14408
rect 15844 14365 15853 14399
rect 15853 14365 15887 14399
rect 15887 14365 15896 14399
rect 15844 14356 15896 14365
rect 1952 14220 2004 14272
rect 5080 14263 5132 14272
rect 5080 14229 5089 14263
rect 5089 14229 5123 14263
rect 5123 14229 5132 14263
rect 5080 14220 5132 14229
rect 6920 14263 6972 14272
rect 6920 14229 6929 14263
rect 6929 14229 6963 14263
rect 6963 14229 6972 14263
rect 6920 14220 6972 14229
rect 9220 14220 9272 14272
rect 10876 14220 10928 14272
rect 11888 14220 11940 14272
rect 13728 14220 13780 14272
rect 15108 14220 15160 14272
rect 18788 14220 18840 14272
rect 23756 14220 23808 14272
rect 5982 14118 6034 14170
rect 6046 14118 6098 14170
rect 6110 14118 6162 14170
rect 6174 14118 6226 14170
rect 15982 14118 16034 14170
rect 16046 14118 16098 14170
rect 16110 14118 16162 14170
rect 16174 14118 16226 14170
rect 25982 14118 26034 14170
rect 26046 14118 26098 14170
rect 26110 14118 26162 14170
rect 26174 14118 26226 14170
rect 2596 14059 2648 14068
rect 2596 14025 2605 14059
rect 2605 14025 2639 14059
rect 2639 14025 2648 14059
rect 2596 14016 2648 14025
rect 2964 14059 3016 14068
rect 2964 14025 2973 14059
rect 2973 14025 3007 14059
rect 3007 14025 3016 14059
rect 2964 14016 3016 14025
rect 5816 14016 5868 14068
rect 10600 14016 10652 14068
rect 16304 14016 16356 14068
rect 18880 14059 18932 14068
rect 18880 14025 18889 14059
rect 18889 14025 18923 14059
rect 18923 14025 18932 14059
rect 18880 14016 18932 14025
rect 19248 14016 19300 14068
rect 21824 14016 21876 14068
rect 22376 14059 22428 14068
rect 22376 14025 22385 14059
rect 22385 14025 22419 14059
rect 22419 14025 22428 14059
rect 22376 14016 22428 14025
rect 22652 14059 22704 14068
rect 22652 14025 22661 14059
rect 22661 14025 22695 14059
rect 22695 14025 22704 14059
rect 22652 14016 22704 14025
rect 24860 14016 24912 14068
rect 1768 13948 1820 14000
rect 1676 13880 1728 13932
rect 4068 13948 4120 14000
rect 5724 13948 5776 14000
rect 16580 13948 16632 14000
rect 5080 13880 5132 13932
rect 5356 13880 5408 13932
rect 2504 13812 2556 13864
rect 4988 13812 5040 13864
rect 6920 13880 6972 13932
rect 8300 13880 8352 13932
rect 9220 13923 9272 13932
rect 9220 13889 9229 13923
rect 9229 13889 9263 13923
rect 9263 13889 9272 13923
rect 9220 13880 9272 13889
rect 24860 13880 24912 13932
rect 25228 13880 25280 13932
rect 8024 13812 8076 13864
rect 10784 13812 10836 13864
rect 15200 13855 15252 13864
rect 15200 13821 15209 13855
rect 15209 13821 15243 13855
rect 15243 13821 15252 13855
rect 15200 13812 15252 13821
rect 15384 13812 15436 13864
rect 19708 13855 19760 13864
rect 19708 13821 19717 13855
rect 19717 13821 19751 13855
rect 19751 13821 19760 13855
rect 19708 13812 19760 13821
rect 25412 13812 25464 13864
rect 25780 13855 25832 13864
rect 25780 13821 25803 13855
rect 25803 13821 25832 13855
rect 25780 13812 25832 13821
rect 5172 13744 5224 13796
rect 1584 13719 1636 13728
rect 1584 13685 1593 13719
rect 1593 13685 1627 13719
rect 1627 13685 1636 13719
rect 1584 13676 1636 13685
rect 1952 13719 2004 13728
rect 1952 13685 1961 13719
rect 1961 13685 1995 13719
rect 1995 13685 2004 13719
rect 1952 13676 2004 13685
rect 4804 13676 4856 13728
rect 9404 13744 9456 13796
rect 5724 13676 5776 13728
rect 6368 13676 6420 13728
rect 8576 13719 8628 13728
rect 8576 13685 8585 13719
rect 8585 13685 8619 13719
rect 8619 13685 8628 13719
rect 8576 13676 8628 13685
rect 14188 13676 14240 13728
rect 14924 13744 14976 13796
rect 15844 13744 15896 13796
rect 18144 13676 18196 13728
rect 26516 13676 26568 13728
rect 10982 13574 11034 13626
rect 11046 13574 11098 13626
rect 11110 13574 11162 13626
rect 11174 13574 11226 13626
rect 20982 13574 21034 13626
rect 21046 13574 21098 13626
rect 21110 13574 21162 13626
rect 21174 13574 21226 13626
rect 1676 13472 1728 13524
rect 1952 13472 2004 13524
rect 4068 13472 4120 13524
rect 6644 13472 6696 13524
rect 8024 13515 8076 13524
rect 8024 13481 8033 13515
rect 8033 13481 8067 13515
rect 8067 13481 8076 13515
rect 8024 13472 8076 13481
rect 15016 13515 15068 13524
rect 15016 13481 15025 13515
rect 15025 13481 15059 13515
rect 15059 13481 15068 13515
rect 15016 13472 15068 13481
rect 18144 13472 18196 13524
rect 4896 13447 4948 13456
rect 4896 13413 4905 13447
rect 4905 13413 4939 13447
rect 4939 13413 4948 13447
rect 4896 13404 4948 13413
rect 5816 13404 5868 13456
rect 2228 13379 2280 13388
rect 2228 13345 2237 13379
rect 2237 13345 2271 13379
rect 2271 13345 2280 13379
rect 2228 13336 2280 13345
rect 2872 13336 2924 13388
rect 11336 13404 11388 13456
rect 15752 13447 15804 13456
rect 15752 13413 15761 13447
rect 15761 13413 15795 13447
rect 15795 13413 15804 13447
rect 15752 13404 15804 13413
rect 22928 13404 22980 13456
rect 23664 13447 23716 13456
rect 23664 13413 23673 13447
rect 23673 13413 23707 13447
rect 23707 13413 23716 13447
rect 23664 13404 23716 13413
rect 8392 13379 8444 13388
rect 2504 13311 2556 13320
rect 2504 13277 2513 13311
rect 2513 13277 2547 13311
rect 2547 13277 2556 13311
rect 2504 13268 2556 13277
rect 4988 13268 5040 13320
rect 5540 13268 5592 13320
rect 6368 13268 6420 13320
rect 8392 13345 8401 13379
rect 8401 13345 8435 13379
rect 8435 13345 8444 13379
rect 8392 13336 8444 13345
rect 10784 13336 10836 13388
rect 11152 13336 11204 13388
rect 7012 13268 7064 13320
rect 8024 13268 8076 13320
rect 8668 13311 8720 13320
rect 8668 13277 8677 13311
rect 8677 13277 8711 13311
rect 8711 13277 8720 13311
rect 8668 13268 8720 13277
rect 13912 13336 13964 13388
rect 14096 13379 14148 13388
rect 14096 13345 14105 13379
rect 14105 13345 14139 13379
rect 14139 13345 14148 13379
rect 14096 13336 14148 13345
rect 16396 13336 16448 13388
rect 17776 13379 17828 13388
rect 17776 13345 17785 13379
rect 17785 13345 17819 13379
rect 17819 13345 17828 13379
rect 17776 13336 17828 13345
rect 18052 13379 18104 13388
rect 18052 13345 18086 13379
rect 18086 13345 18104 13379
rect 18052 13336 18104 13345
rect 21272 13379 21324 13388
rect 21272 13345 21281 13379
rect 21281 13345 21315 13379
rect 21315 13345 21324 13379
rect 21272 13336 21324 13345
rect 23572 13379 23624 13388
rect 23572 13345 23581 13379
rect 23581 13345 23615 13379
rect 23615 13345 23624 13379
rect 23572 13336 23624 13345
rect 25136 13336 25188 13388
rect 9496 13200 9548 13252
rect 12348 13268 12400 13320
rect 14188 13311 14240 13320
rect 14188 13277 14197 13311
rect 14197 13277 14231 13311
rect 14231 13277 14240 13311
rect 14188 13268 14240 13277
rect 15844 13311 15896 13320
rect 15844 13277 15853 13311
rect 15853 13277 15887 13311
rect 15887 13277 15896 13311
rect 15844 13268 15896 13277
rect 21364 13311 21416 13320
rect 21364 13277 21373 13311
rect 21373 13277 21407 13311
rect 21407 13277 21416 13311
rect 21364 13268 21416 13277
rect 21456 13311 21508 13320
rect 21456 13277 21465 13311
rect 21465 13277 21499 13311
rect 21499 13277 21508 13311
rect 23756 13311 23808 13320
rect 21456 13268 21508 13277
rect 23756 13277 23765 13311
rect 23765 13277 23799 13311
rect 23799 13277 23808 13311
rect 23756 13268 23808 13277
rect 25320 13311 25372 13320
rect 25320 13277 25329 13311
rect 25329 13277 25363 13311
rect 25363 13277 25372 13311
rect 25320 13268 25372 13277
rect 25504 13311 25556 13320
rect 25504 13277 25513 13311
rect 25513 13277 25547 13311
rect 25547 13277 25556 13311
rect 25504 13268 25556 13277
rect 26516 13268 26568 13320
rect 11520 13200 11572 13252
rect 4528 13175 4580 13184
rect 4528 13141 4537 13175
rect 4537 13141 4571 13175
rect 4571 13141 4580 13175
rect 4528 13132 4580 13141
rect 9128 13175 9180 13184
rect 9128 13141 9137 13175
rect 9137 13141 9171 13175
rect 9171 13141 9180 13175
rect 9128 13132 9180 13141
rect 10048 13132 10100 13184
rect 10508 13132 10560 13184
rect 13820 13132 13872 13184
rect 15660 13132 15712 13184
rect 20904 13175 20956 13184
rect 20904 13141 20913 13175
rect 20913 13141 20947 13175
rect 20947 13141 20956 13175
rect 20904 13132 20956 13141
rect 22560 13132 22612 13184
rect 24308 13175 24360 13184
rect 24308 13141 24317 13175
rect 24317 13141 24351 13175
rect 24351 13141 24360 13175
rect 24308 13132 24360 13141
rect 24860 13175 24912 13184
rect 24860 13141 24869 13175
rect 24869 13141 24903 13175
rect 24903 13141 24912 13175
rect 24860 13132 24912 13141
rect 25044 13132 25096 13184
rect 25504 13132 25556 13184
rect 5982 13030 6034 13082
rect 6046 13030 6098 13082
rect 6110 13030 6162 13082
rect 6174 13030 6226 13082
rect 15982 13030 16034 13082
rect 16046 13030 16098 13082
rect 16110 13030 16162 13082
rect 16174 13030 16226 13082
rect 25982 13030 26034 13082
rect 26046 13030 26098 13082
rect 26110 13030 26162 13082
rect 26174 13030 26226 13082
rect 4896 12928 4948 12980
rect 5172 12971 5224 12980
rect 5172 12937 5181 12971
rect 5181 12937 5215 12971
rect 5215 12937 5224 12971
rect 5172 12928 5224 12937
rect 6368 12928 6420 12980
rect 7012 12971 7064 12980
rect 7012 12937 7021 12971
rect 7021 12937 7055 12971
rect 7055 12937 7064 12971
rect 7012 12928 7064 12937
rect 10048 12928 10100 12980
rect 11520 12971 11572 12980
rect 2044 12792 2096 12844
rect 4804 12860 4856 12912
rect 3056 12792 3108 12844
rect 3700 12792 3752 12844
rect 8668 12860 8720 12912
rect 8760 12860 8812 12912
rect 9772 12860 9824 12912
rect 5816 12835 5868 12844
rect 5816 12801 5825 12835
rect 5825 12801 5859 12835
rect 5859 12801 5868 12835
rect 5816 12792 5868 12801
rect 8576 12792 8628 12844
rect 8852 12792 8904 12844
rect 1584 12724 1636 12776
rect 2596 12724 2648 12776
rect 3884 12724 3936 12776
rect 4528 12724 4580 12776
rect 8668 12724 8720 12776
rect 9588 12792 9640 12844
rect 11520 12937 11529 12971
rect 11529 12937 11563 12971
rect 11563 12937 11572 12971
rect 11520 12928 11572 12937
rect 12440 12928 12492 12980
rect 14832 12971 14884 12980
rect 14832 12937 14841 12971
rect 14841 12937 14875 12971
rect 14875 12937 14884 12971
rect 14832 12928 14884 12937
rect 15568 12928 15620 12980
rect 15752 12928 15804 12980
rect 15844 12928 15896 12980
rect 21272 12928 21324 12980
rect 22928 12971 22980 12980
rect 22928 12937 22937 12971
rect 22937 12937 22971 12971
rect 22971 12937 22980 12971
rect 22928 12928 22980 12937
rect 23572 12928 23624 12980
rect 25320 12928 25372 12980
rect 26516 12971 26568 12980
rect 26516 12937 26525 12971
rect 26525 12937 26559 12971
rect 26559 12937 26568 12971
rect 26516 12928 26568 12937
rect 27344 12928 27396 12980
rect 10784 12860 10836 12912
rect 9496 12724 9548 12776
rect 10508 12767 10560 12776
rect 10508 12733 10517 12767
rect 10517 12733 10551 12767
rect 10551 12733 10560 12767
rect 10508 12724 10560 12733
rect 10876 12792 10928 12844
rect 11152 12767 11204 12776
rect 2228 12656 2280 12708
rect 2964 12656 3016 12708
rect 9128 12656 9180 12708
rect 9588 12656 9640 12708
rect 11152 12733 11161 12767
rect 11161 12733 11195 12767
rect 11195 12733 11204 12767
rect 11152 12724 11204 12733
rect 15660 12724 15712 12776
rect 16396 12860 16448 12912
rect 21364 12860 21416 12912
rect 23756 12860 23808 12912
rect 18052 12792 18104 12844
rect 18788 12835 18840 12844
rect 18788 12801 18797 12835
rect 18797 12801 18831 12835
rect 18831 12801 18840 12835
rect 18788 12792 18840 12801
rect 20352 12835 20404 12844
rect 20352 12801 20361 12835
rect 20361 12801 20395 12835
rect 20395 12801 20404 12835
rect 20352 12792 20404 12801
rect 20444 12724 20496 12776
rect 24584 12835 24636 12844
rect 24584 12801 24593 12835
rect 24593 12801 24627 12835
rect 24627 12801 24636 12835
rect 24584 12792 24636 12801
rect 24400 12724 24452 12776
rect 24768 12724 24820 12776
rect 10784 12656 10836 12708
rect 14280 12656 14332 12708
rect 18512 12699 18564 12708
rect 18512 12665 18521 12699
rect 18521 12665 18555 12699
rect 18555 12665 18564 12699
rect 18512 12656 18564 12665
rect 19616 12656 19668 12708
rect 22100 12656 22152 12708
rect 1952 12588 2004 12640
rect 2872 12631 2924 12640
rect 2872 12597 2881 12631
rect 2881 12597 2915 12631
rect 2915 12597 2924 12631
rect 2872 12588 2924 12597
rect 4068 12588 4120 12640
rect 5264 12588 5316 12640
rect 6644 12631 6696 12640
rect 6644 12597 6653 12631
rect 6653 12597 6687 12631
rect 6687 12597 6696 12631
rect 6644 12588 6696 12597
rect 8024 12631 8076 12640
rect 8024 12597 8033 12631
rect 8033 12597 8067 12631
rect 8067 12597 8076 12631
rect 8024 12588 8076 12597
rect 8392 12588 8444 12640
rect 9496 12588 9548 12640
rect 10600 12588 10652 12640
rect 11428 12588 11480 12640
rect 13452 12631 13504 12640
rect 13452 12597 13461 12631
rect 13461 12597 13495 12631
rect 13495 12597 13504 12631
rect 13452 12588 13504 12597
rect 17408 12588 17460 12640
rect 18604 12631 18656 12640
rect 18604 12597 18613 12631
rect 18613 12597 18647 12631
rect 18647 12597 18656 12631
rect 18604 12588 18656 12597
rect 20812 12588 20864 12640
rect 21456 12588 21508 12640
rect 24308 12588 24360 12640
rect 25044 12656 25096 12708
rect 25228 12656 25280 12708
rect 25136 12588 25188 12640
rect 26148 12860 26200 12912
rect 25780 12792 25832 12844
rect 25412 12724 25464 12776
rect 25964 12724 26016 12776
rect 27528 12767 27580 12776
rect 27528 12733 27537 12767
rect 27537 12733 27571 12767
rect 27571 12733 27580 12767
rect 27528 12724 27580 12733
rect 25596 12656 25648 12708
rect 26424 12656 26476 12708
rect 26884 12631 26936 12640
rect 26884 12597 26893 12631
rect 26893 12597 26927 12631
rect 26927 12597 26936 12631
rect 26884 12588 26936 12597
rect 10982 12486 11034 12538
rect 11046 12486 11098 12538
rect 11110 12486 11162 12538
rect 11174 12486 11226 12538
rect 20982 12486 21034 12538
rect 21046 12486 21098 12538
rect 21110 12486 21162 12538
rect 21174 12486 21226 12538
rect 3884 12427 3936 12436
rect 3884 12393 3893 12427
rect 3893 12393 3927 12427
rect 3927 12393 3936 12427
rect 3884 12384 3936 12393
rect 4988 12384 5040 12436
rect 5540 12384 5592 12436
rect 8668 12427 8720 12436
rect 8668 12393 8677 12427
rect 8677 12393 8711 12427
rect 8711 12393 8720 12427
rect 8668 12384 8720 12393
rect 8852 12384 8904 12436
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 10784 12427 10836 12436
rect 10784 12393 10793 12427
rect 10793 12393 10827 12427
rect 10827 12393 10836 12427
rect 10784 12384 10836 12393
rect 11336 12384 11388 12436
rect 11888 12384 11940 12436
rect 12348 12384 12400 12436
rect 12440 12427 12492 12436
rect 12440 12393 12449 12427
rect 12449 12393 12483 12427
rect 12483 12393 12492 12427
rect 12440 12384 12492 12393
rect 14188 12384 14240 12436
rect 17408 12427 17460 12436
rect 17408 12393 17417 12427
rect 17417 12393 17451 12427
rect 17451 12393 17460 12427
rect 17408 12384 17460 12393
rect 17776 12384 17828 12436
rect 18512 12427 18564 12436
rect 18512 12393 18521 12427
rect 18521 12393 18555 12427
rect 18555 12393 18564 12427
rect 18512 12384 18564 12393
rect 20352 12427 20404 12436
rect 20352 12393 20361 12427
rect 20361 12393 20395 12427
rect 20395 12393 20404 12427
rect 20352 12384 20404 12393
rect 20812 12384 20864 12436
rect 21364 12384 21416 12436
rect 21640 12384 21692 12436
rect 21824 12384 21876 12436
rect 23572 12427 23624 12436
rect 23572 12393 23581 12427
rect 23581 12393 23615 12427
rect 23615 12393 23624 12427
rect 23572 12384 23624 12393
rect 23664 12384 23716 12436
rect 1768 12316 1820 12368
rect 3700 12316 3752 12368
rect 8024 12316 8076 12368
rect 15844 12316 15896 12368
rect 18420 12316 18472 12368
rect 24124 12316 24176 12368
rect 2228 12248 2280 12300
rect 5632 12248 5684 12300
rect 6000 12291 6052 12300
rect 6000 12257 6009 12291
rect 6009 12257 6043 12291
rect 6043 12257 6052 12291
rect 6000 12248 6052 12257
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 10048 12248 10100 12257
rect 12532 12248 12584 12300
rect 12808 12291 12860 12300
rect 12808 12257 12817 12291
rect 12817 12257 12851 12291
rect 12851 12257 12860 12291
rect 12808 12248 12860 12257
rect 13636 12291 13688 12300
rect 13636 12257 13645 12291
rect 13645 12257 13679 12291
rect 13679 12257 13688 12291
rect 13636 12248 13688 12257
rect 13820 12248 13872 12300
rect 14096 12248 14148 12300
rect 5816 12180 5868 12232
rect 6368 12180 6420 12232
rect 9680 12180 9732 12232
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 11428 12180 11480 12232
rect 12900 12223 12952 12232
rect 12900 12189 12909 12223
rect 12909 12189 12943 12223
rect 12943 12189 12952 12223
rect 12900 12180 12952 12189
rect 12440 12112 12492 12164
rect 14556 12180 14608 12232
rect 15108 12248 15160 12300
rect 15752 12291 15804 12300
rect 15752 12257 15761 12291
rect 15761 12257 15795 12291
rect 15795 12257 15804 12291
rect 15752 12248 15804 12257
rect 17040 12248 17092 12300
rect 17316 12291 17368 12300
rect 17316 12257 17325 12291
rect 17325 12257 17359 12291
rect 17359 12257 17368 12291
rect 17316 12248 17368 12257
rect 21640 12248 21692 12300
rect 14924 12223 14976 12232
rect 14924 12189 14933 12223
rect 14933 12189 14967 12223
rect 14967 12189 14976 12223
rect 14924 12180 14976 12189
rect 16580 12180 16632 12232
rect 17132 12180 17184 12232
rect 18144 12180 18196 12232
rect 18972 12223 19024 12232
rect 18972 12189 18981 12223
rect 18981 12189 19015 12223
rect 19015 12189 19024 12223
rect 18972 12180 19024 12189
rect 19156 12223 19208 12232
rect 19156 12189 19165 12223
rect 19165 12189 19199 12223
rect 19199 12189 19208 12223
rect 19156 12180 19208 12189
rect 22100 12223 22152 12232
rect 22100 12189 22109 12223
rect 22109 12189 22143 12223
rect 22143 12189 22152 12223
rect 22100 12180 22152 12189
rect 23020 12223 23072 12232
rect 23020 12189 23029 12223
rect 23029 12189 23063 12223
rect 23063 12189 23072 12223
rect 23020 12180 23072 12189
rect 24584 12316 24636 12368
rect 24584 12180 24636 12232
rect 24768 12384 24820 12436
rect 25780 12384 25832 12436
rect 27528 12384 27580 12436
rect 3056 12044 3108 12096
rect 5264 12087 5316 12096
rect 5264 12053 5273 12087
rect 5273 12053 5307 12087
rect 5307 12053 5316 12087
rect 5264 12044 5316 12053
rect 5448 12044 5500 12096
rect 14280 12087 14332 12096
rect 14280 12053 14289 12087
rect 14289 12053 14323 12087
rect 14323 12053 14332 12087
rect 14280 12044 14332 12053
rect 14372 12044 14424 12096
rect 16396 12087 16448 12096
rect 16396 12053 16405 12087
rect 16405 12053 16439 12087
rect 16439 12053 16448 12087
rect 16396 12044 16448 12053
rect 17684 12044 17736 12096
rect 24308 12087 24360 12096
rect 24308 12053 24317 12087
rect 24317 12053 24351 12087
rect 24351 12053 24360 12087
rect 24308 12044 24360 12053
rect 24952 12044 25004 12096
rect 26148 12316 26200 12368
rect 26884 12248 26936 12300
rect 25412 12044 25464 12096
rect 25780 12044 25832 12096
rect 5982 11942 6034 11994
rect 6046 11942 6098 11994
rect 6110 11942 6162 11994
rect 6174 11942 6226 11994
rect 15982 11942 16034 11994
rect 16046 11942 16098 11994
rect 16110 11942 16162 11994
rect 16174 11942 16226 11994
rect 25982 11942 26034 11994
rect 26046 11942 26098 11994
rect 26110 11942 26162 11994
rect 26174 11942 26226 11994
rect 1768 11840 1820 11892
rect 2596 11840 2648 11892
rect 3240 11840 3292 11892
rect 5632 11883 5684 11892
rect 5632 11849 5641 11883
rect 5641 11849 5675 11883
rect 5675 11849 5684 11883
rect 5632 11840 5684 11849
rect 6368 11883 6420 11892
rect 6368 11849 6377 11883
rect 6377 11849 6411 11883
rect 6411 11849 6420 11883
rect 6368 11840 6420 11849
rect 10048 11840 10100 11892
rect 11888 11883 11940 11892
rect 11888 11849 11897 11883
rect 11897 11849 11931 11883
rect 11931 11849 11940 11883
rect 11888 11840 11940 11849
rect 12900 11840 12952 11892
rect 15384 11883 15436 11892
rect 15384 11849 15393 11883
rect 15393 11849 15427 11883
rect 15427 11849 15436 11883
rect 15384 11840 15436 11849
rect 15844 11840 15896 11892
rect 17132 11840 17184 11892
rect 17408 11883 17460 11892
rect 17408 11849 17417 11883
rect 17417 11849 17451 11883
rect 17451 11849 17460 11883
rect 17408 11840 17460 11849
rect 18604 11840 18656 11892
rect 20536 11840 20588 11892
rect 2504 11772 2556 11824
rect 6276 11772 6328 11824
rect 12808 11772 12860 11824
rect 16672 11815 16724 11824
rect 10416 11704 10468 11756
rect 14188 11704 14240 11756
rect 10784 11636 10836 11688
rect 13820 11636 13872 11688
rect 14280 11636 14332 11688
rect 16672 11781 16681 11815
rect 16681 11781 16715 11815
rect 16715 11781 16724 11815
rect 16672 11772 16724 11781
rect 19616 11815 19668 11824
rect 19616 11781 19625 11815
rect 19625 11781 19659 11815
rect 19659 11781 19668 11815
rect 19616 11772 19668 11781
rect 16120 11747 16172 11756
rect 16120 11713 16129 11747
rect 16129 11713 16163 11747
rect 16163 11713 16172 11747
rect 16120 11704 16172 11713
rect 19156 11747 19208 11756
rect 19156 11713 19165 11747
rect 19165 11713 19199 11747
rect 19199 11713 19208 11747
rect 21272 11840 21324 11892
rect 24124 11883 24176 11892
rect 24124 11849 24133 11883
rect 24133 11849 24167 11883
rect 24167 11849 24176 11883
rect 24124 11840 24176 11849
rect 25044 11840 25096 11892
rect 26884 11840 26936 11892
rect 25228 11772 25280 11824
rect 19156 11704 19208 11713
rect 22100 11747 22152 11756
rect 22100 11713 22109 11747
rect 22109 11713 22143 11747
rect 22143 11713 22152 11747
rect 22100 11704 22152 11713
rect 25136 11747 25188 11756
rect 25136 11713 25145 11747
rect 25145 11713 25179 11747
rect 25179 11713 25188 11747
rect 25136 11704 25188 11713
rect 27436 11747 27488 11756
rect 25688 11679 25740 11688
rect 25688 11645 25697 11679
rect 25697 11645 25731 11679
rect 25731 11645 25740 11679
rect 25688 11636 25740 11645
rect 9312 11568 9364 11620
rect 1584 11543 1636 11552
rect 1584 11509 1593 11543
rect 1593 11509 1627 11543
rect 1627 11509 1636 11543
rect 1584 11500 1636 11509
rect 10140 11543 10192 11552
rect 10140 11509 10149 11543
rect 10149 11509 10183 11543
rect 10183 11509 10192 11543
rect 10140 11500 10192 11509
rect 13912 11568 13964 11620
rect 14372 11611 14424 11620
rect 14372 11577 14381 11611
rect 14381 11577 14415 11611
rect 14415 11577 14424 11611
rect 14372 11568 14424 11577
rect 15292 11568 15344 11620
rect 16396 11568 16448 11620
rect 19064 11568 19116 11620
rect 23020 11568 23072 11620
rect 27436 11713 27445 11747
rect 27445 11713 27479 11747
rect 27479 11713 27488 11747
rect 27436 11704 27488 11713
rect 27068 11636 27120 11688
rect 10784 11500 10836 11552
rect 11428 11543 11480 11552
rect 11428 11509 11437 11543
rect 11437 11509 11471 11543
rect 11471 11509 11480 11543
rect 11428 11500 11480 11509
rect 12440 11500 12492 11552
rect 13544 11543 13596 11552
rect 13544 11509 13553 11543
rect 13553 11509 13587 11543
rect 13587 11509 13596 11543
rect 13544 11500 13596 11509
rect 13820 11543 13872 11552
rect 13820 11509 13829 11543
rect 13829 11509 13863 11543
rect 13863 11509 13872 11543
rect 13820 11500 13872 11509
rect 14004 11543 14056 11552
rect 14004 11509 14013 11543
rect 14013 11509 14047 11543
rect 14047 11509 14056 11543
rect 14004 11500 14056 11509
rect 15384 11500 15436 11552
rect 18420 11543 18472 11552
rect 18420 11509 18429 11543
rect 18429 11509 18463 11543
rect 18463 11509 18472 11543
rect 18420 11500 18472 11509
rect 18512 11500 18564 11552
rect 20812 11500 20864 11552
rect 21640 11500 21692 11552
rect 22928 11543 22980 11552
rect 22928 11509 22937 11543
rect 22937 11509 22971 11543
rect 22971 11509 22980 11543
rect 22928 11500 22980 11509
rect 26240 11500 26292 11552
rect 27252 11543 27304 11552
rect 27252 11509 27261 11543
rect 27261 11509 27295 11543
rect 27295 11509 27304 11543
rect 27252 11500 27304 11509
rect 10982 11398 11034 11450
rect 11046 11398 11098 11450
rect 11110 11398 11162 11450
rect 11174 11398 11226 11450
rect 20982 11398 21034 11450
rect 21046 11398 21098 11450
rect 21110 11398 21162 11450
rect 21174 11398 21226 11450
rect 2044 11339 2096 11348
rect 2044 11305 2053 11339
rect 2053 11305 2087 11339
rect 2087 11305 2096 11339
rect 2044 11296 2096 11305
rect 2228 11296 2280 11348
rect 2688 11339 2740 11348
rect 2688 11305 2697 11339
rect 2697 11305 2731 11339
rect 2731 11305 2740 11339
rect 2688 11296 2740 11305
rect 6552 11339 6604 11348
rect 6552 11305 6561 11339
rect 6561 11305 6595 11339
rect 6595 11305 6604 11339
rect 6552 11296 6604 11305
rect 9220 11296 9272 11348
rect 10232 11296 10284 11348
rect 12440 11339 12492 11348
rect 12440 11305 12449 11339
rect 12449 11305 12483 11339
rect 12483 11305 12492 11339
rect 14556 11339 14608 11348
rect 12440 11296 12492 11305
rect 14556 11305 14565 11339
rect 14565 11305 14599 11339
rect 14599 11305 14608 11339
rect 14556 11296 14608 11305
rect 17040 11339 17092 11348
rect 17040 11305 17049 11339
rect 17049 11305 17083 11339
rect 17083 11305 17092 11339
rect 17040 11296 17092 11305
rect 18972 11339 19024 11348
rect 18972 11305 18981 11339
rect 18981 11305 19015 11339
rect 19015 11305 19024 11339
rect 18972 11296 19024 11305
rect 21824 11296 21876 11348
rect 22928 11296 22980 11348
rect 24584 11339 24636 11348
rect 24584 11305 24593 11339
rect 24593 11305 24627 11339
rect 24627 11305 24636 11339
rect 24584 11296 24636 11305
rect 24952 11339 25004 11348
rect 24952 11305 24961 11339
rect 24961 11305 24995 11339
rect 24995 11305 25004 11339
rect 24952 11296 25004 11305
rect 27252 11296 27304 11348
rect 27436 11339 27488 11348
rect 27436 11305 27445 11339
rect 27445 11305 27479 11339
rect 27479 11305 27488 11339
rect 27436 11296 27488 11305
rect 1492 11160 1544 11212
rect 2688 11160 2740 11212
rect 7380 11228 7432 11280
rect 9680 11228 9732 11280
rect 15936 11228 15988 11280
rect 22100 11228 22152 11280
rect 26424 11228 26476 11280
rect 27068 11271 27120 11280
rect 27068 11237 27077 11271
rect 27077 11237 27111 11271
rect 27111 11237 27120 11271
rect 27068 11228 27120 11237
rect 5264 11160 5316 11212
rect 10968 11160 11020 11212
rect 12900 11160 12952 11212
rect 13820 11160 13872 11212
rect 14924 11160 14976 11212
rect 15476 11160 15528 11212
rect 15752 11203 15804 11212
rect 15752 11169 15761 11203
rect 15761 11169 15795 11203
rect 15795 11169 15804 11203
rect 15752 11160 15804 11169
rect 20076 11160 20128 11212
rect 20260 11160 20312 11212
rect 25688 11160 25740 11212
rect 27252 11160 27304 11212
rect 5172 11135 5224 11144
rect 5172 11101 5181 11135
rect 5181 11101 5215 11135
rect 5215 11101 5224 11135
rect 5172 11092 5224 11101
rect 1768 11024 1820 11076
rect 7288 10956 7340 11008
rect 9864 11092 9916 11144
rect 10232 11092 10284 11144
rect 10508 11135 10560 11144
rect 10508 11101 10517 11135
rect 10517 11101 10551 11135
rect 10551 11101 10560 11135
rect 10508 11092 10560 11101
rect 10600 11135 10652 11144
rect 10600 11101 10609 11135
rect 10609 11101 10643 11135
rect 10643 11101 10652 11135
rect 12808 11135 12860 11144
rect 10600 11092 10652 11101
rect 12808 11101 12817 11135
rect 12817 11101 12851 11135
rect 12851 11101 12860 11135
rect 12808 11092 12860 11101
rect 16120 11092 16172 11144
rect 19524 11092 19576 11144
rect 21916 11135 21968 11144
rect 7748 10956 7800 11008
rect 8392 10956 8444 11008
rect 9588 10956 9640 11008
rect 14188 10999 14240 11008
rect 14188 10965 14197 10999
rect 14197 10965 14231 10999
rect 14231 10965 14240 10999
rect 14188 10956 14240 10965
rect 15108 10956 15160 11008
rect 18512 10999 18564 11008
rect 18512 10965 18521 10999
rect 18521 10965 18555 10999
rect 18555 10965 18564 10999
rect 18512 10956 18564 10965
rect 21916 11101 21925 11135
rect 21925 11101 21959 11135
rect 21959 11101 21968 11135
rect 21916 11092 21968 11101
rect 26700 11067 26752 11076
rect 26700 11033 26709 11067
rect 26709 11033 26743 11067
rect 26743 11033 26752 11067
rect 26700 11024 26752 11033
rect 19616 10956 19668 11008
rect 5982 10854 6034 10906
rect 6046 10854 6098 10906
rect 6110 10854 6162 10906
rect 6174 10854 6226 10906
rect 15982 10854 16034 10906
rect 16046 10854 16098 10906
rect 16110 10854 16162 10906
rect 16174 10854 16226 10906
rect 25982 10854 26034 10906
rect 26046 10854 26098 10906
rect 26110 10854 26162 10906
rect 26174 10854 26226 10906
rect 1492 10752 1544 10804
rect 2688 10752 2740 10804
rect 5264 10795 5316 10804
rect 5264 10761 5273 10795
rect 5273 10761 5307 10795
rect 5307 10761 5316 10795
rect 5264 10752 5316 10761
rect 6552 10795 6604 10804
rect 6552 10761 6561 10795
rect 6561 10761 6595 10795
rect 6595 10761 6604 10795
rect 6552 10752 6604 10761
rect 5172 10684 5224 10736
rect 5816 10684 5868 10736
rect 7748 10752 7800 10804
rect 10508 10752 10560 10804
rect 12900 10795 12952 10804
rect 12900 10761 12909 10795
rect 12909 10761 12943 10795
rect 12943 10761 12952 10795
rect 12900 10752 12952 10761
rect 13728 10795 13780 10804
rect 13728 10761 13737 10795
rect 13737 10761 13771 10795
rect 13771 10761 13780 10795
rect 13728 10752 13780 10761
rect 14096 10795 14148 10804
rect 14096 10761 14105 10795
rect 14105 10761 14139 10795
rect 14139 10761 14148 10795
rect 14096 10752 14148 10761
rect 15752 10752 15804 10804
rect 9864 10727 9916 10736
rect 9864 10693 9873 10727
rect 9873 10693 9907 10727
rect 9907 10693 9916 10727
rect 9864 10684 9916 10693
rect 10324 10684 10376 10736
rect 2228 10616 2280 10668
rect 5632 10616 5684 10668
rect 6644 10616 6696 10668
rect 7288 10659 7340 10668
rect 7288 10625 7297 10659
rect 7297 10625 7331 10659
rect 7331 10625 7340 10659
rect 7288 10616 7340 10625
rect 6552 10548 6604 10600
rect 8392 10616 8444 10668
rect 9496 10616 9548 10668
rect 10140 10616 10192 10668
rect 15844 10684 15896 10736
rect 10600 10659 10652 10668
rect 10600 10625 10609 10659
rect 10609 10625 10643 10659
rect 10643 10625 10652 10659
rect 10600 10616 10652 10625
rect 11060 10616 11112 10668
rect 13728 10616 13780 10668
rect 14188 10616 14240 10668
rect 19064 10752 19116 10804
rect 22008 10795 22060 10804
rect 22008 10761 22017 10795
rect 22017 10761 22051 10795
rect 22051 10761 22060 10795
rect 22008 10752 22060 10761
rect 27252 10752 27304 10804
rect 19616 10659 19668 10668
rect 19616 10625 19625 10659
rect 19625 10625 19659 10659
rect 19659 10625 19668 10659
rect 19616 10616 19668 10625
rect 8576 10548 8628 10600
rect 9588 10548 9640 10600
rect 9864 10548 9916 10600
rect 10048 10548 10100 10600
rect 11336 10548 11388 10600
rect 14740 10548 14792 10600
rect 15384 10548 15436 10600
rect 19340 10591 19392 10600
rect 19340 10557 19349 10591
rect 19349 10557 19383 10591
rect 19383 10557 19392 10591
rect 19340 10548 19392 10557
rect 26424 10591 26476 10600
rect 26424 10557 26433 10591
rect 26433 10557 26467 10591
rect 26467 10557 26476 10591
rect 26424 10548 26476 10557
rect 27528 10591 27580 10600
rect 27528 10557 27537 10591
rect 27537 10557 27571 10591
rect 27571 10557 27580 10591
rect 27528 10548 27580 10557
rect 3056 10480 3108 10532
rect 3884 10480 3936 10532
rect 4804 10480 4856 10532
rect 6368 10480 6420 10532
rect 8852 10523 8904 10532
rect 3792 10455 3844 10464
rect 3792 10421 3801 10455
rect 3801 10421 3835 10455
rect 3835 10421 3844 10455
rect 3792 10412 3844 10421
rect 6644 10412 6696 10464
rect 7380 10412 7432 10464
rect 8392 10455 8444 10464
rect 8392 10421 8401 10455
rect 8401 10421 8435 10455
rect 8435 10421 8444 10455
rect 8392 10412 8444 10421
rect 8852 10489 8861 10523
rect 8861 10489 8895 10523
rect 8895 10489 8904 10523
rect 8852 10480 8904 10489
rect 9496 10455 9548 10464
rect 9496 10421 9505 10455
rect 9505 10421 9539 10455
rect 9539 10421 9548 10455
rect 9496 10412 9548 10421
rect 10324 10480 10376 10532
rect 15108 10480 15160 10532
rect 18420 10523 18472 10532
rect 18420 10489 18429 10523
rect 18429 10489 18463 10523
rect 18463 10489 18472 10523
rect 18420 10480 18472 10489
rect 13820 10412 13872 10464
rect 14188 10412 14240 10464
rect 14556 10455 14608 10464
rect 14556 10421 14565 10455
rect 14565 10421 14599 10455
rect 14599 10421 14608 10455
rect 14556 10412 14608 10421
rect 18880 10455 18932 10464
rect 18880 10421 18889 10455
rect 18889 10421 18923 10455
rect 18923 10421 18932 10455
rect 20444 10480 20496 10532
rect 21916 10480 21968 10532
rect 22100 10480 22152 10532
rect 18880 10412 18932 10421
rect 20260 10412 20312 10464
rect 25228 10455 25280 10464
rect 25228 10421 25237 10455
rect 25237 10421 25271 10455
rect 25271 10421 25280 10455
rect 25228 10412 25280 10421
rect 26608 10455 26660 10464
rect 26608 10421 26617 10455
rect 26617 10421 26651 10455
rect 26651 10421 26660 10455
rect 26608 10412 26660 10421
rect 27712 10455 27764 10464
rect 27712 10421 27721 10455
rect 27721 10421 27755 10455
rect 27755 10421 27764 10455
rect 27712 10412 27764 10421
rect 10982 10310 11034 10362
rect 11046 10310 11098 10362
rect 11110 10310 11162 10362
rect 11174 10310 11226 10362
rect 20982 10310 21034 10362
rect 21046 10310 21098 10362
rect 21110 10310 21162 10362
rect 21174 10310 21226 10362
rect 3056 10251 3108 10260
rect 3056 10217 3065 10251
rect 3065 10217 3099 10251
rect 3099 10217 3108 10251
rect 3056 10208 3108 10217
rect 6368 10251 6420 10260
rect 6368 10217 6377 10251
rect 6377 10217 6411 10251
rect 6411 10217 6420 10251
rect 6368 10208 6420 10217
rect 7748 10251 7800 10260
rect 7748 10217 7757 10251
rect 7757 10217 7791 10251
rect 7791 10217 7800 10251
rect 7748 10208 7800 10217
rect 8576 10251 8628 10260
rect 8576 10217 8585 10251
rect 8585 10217 8619 10251
rect 8619 10217 8628 10251
rect 8576 10208 8628 10217
rect 8852 10251 8904 10260
rect 8852 10217 8861 10251
rect 8861 10217 8895 10251
rect 8895 10217 8904 10251
rect 8852 10208 8904 10217
rect 9496 10208 9548 10260
rect 10048 10251 10100 10260
rect 10048 10217 10057 10251
rect 10057 10217 10091 10251
rect 10091 10217 10100 10251
rect 10048 10208 10100 10217
rect 10416 10251 10468 10260
rect 10416 10217 10425 10251
rect 10425 10217 10459 10251
rect 10459 10217 10468 10251
rect 10416 10208 10468 10217
rect 10508 10208 10560 10260
rect 10692 10208 10744 10260
rect 14096 10208 14148 10260
rect 14556 10208 14608 10260
rect 14740 10251 14792 10260
rect 14740 10217 14749 10251
rect 14749 10217 14783 10251
rect 14783 10217 14792 10251
rect 14740 10208 14792 10217
rect 15108 10251 15160 10260
rect 15108 10217 15117 10251
rect 15117 10217 15151 10251
rect 15151 10217 15160 10251
rect 15108 10208 15160 10217
rect 15476 10251 15528 10260
rect 15476 10217 15485 10251
rect 15485 10217 15519 10251
rect 15519 10217 15528 10251
rect 15476 10208 15528 10217
rect 18512 10208 18564 10260
rect 25504 10208 25556 10260
rect 2228 10140 2280 10192
rect 3516 10183 3568 10192
rect 3516 10149 3525 10183
rect 3525 10149 3559 10183
rect 3559 10149 3568 10183
rect 3516 10140 3568 10149
rect 9864 10140 9916 10192
rect 11520 10140 11572 10192
rect 1676 10072 1728 10124
rect 2504 10115 2556 10124
rect 2504 10081 2513 10115
rect 2513 10081 2547 10115
rect 2547 10081 2556 10115
rect 2504 10072 2556 10081
rect 6736 10115 6788 10124
rect 6736 10081 6745 10115
rect 6745 10081 6779 10115
rect 6779 10081 6788 10115
rect 6736 10072 6788 10081
rect 8208 10072 8260 10124
rect 13728 10072 13780 10124
rect 14004 10072 14056 10124
rect 18696 10072 18748 10124
rect 19340 10115 19392 10124
rect 19340 10081 19349 10115
rect 19349 10081 19383 10115
rect 19383 10081 19392 10115
rect 19340 10072 19392 10081
rect 19708 10072 19760 10124
rect 25228 10115 25280 10124
rect 25228 10081 25237 10115
rect 25237 10081 25271 10115
rect 25271 10081 25280 10115
rect 25228 10072 25280 10081
rect 26516 10115 26568 10124
rect 26516 10081 26525 10115
rect 26525 10081 26559 10115
rect 26559 10081 26568 10115
rect 26516 10072 26568 10081
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 5264 9936 5316 9988
rect 6460 9936 6512 9988
rect 10416 10004 10468 10056
rect 14188 10047 14240 10056
rect 14188 10013 14197 10047
rect 14197 10013 14231 10047
rect 14231 10013 14240 10047
rect 14188 10004 14240 10013
rect 19432 10047 19484 10056
rect 19432 10013 19441 10047
rect 19441 10013 19475 10047
rect 19475 10013 19484 10047
rect 19432 10004 19484 10013
rect 19616 10047 19668 10056
rect 19616 10013 19625 10047
rect 19625 10013 19659 10047
rect 19659 10013 19668 10047
rect 19616 10004 19668 10013
rect 10968 9936 11020 9988
rect 20168 9936 20220 9988
rect 25872 10047 25924 10056
rect 25872 10013 25881 10047
rect 25881 10013 25915 10047
rect 25915 10013 25924 10047
rect 25872 10004 25924 10013
rect 1584 9911 1636 9920
rect 1584 9877 1593 9911
rect 1593 9877 1627 9911
rect 1627 9877 1636 9911
rect 1584 9868 1636 9877
rect 2688 9911 2740 9920
rect 2688 9877 2697 9911
rect 2697 9877 2731 9911
rect 2731 9877 2740 9911
rect 2688 9868 2740 9877
rect 7380 9911 7432 9920
rect 7380 9877 7389 9911
rect 7389 9877 7423 9911
rect 7423 9877 7432 9911
rect 7380 9868 7432 9877
rect 8116 9868 8168 9920
rect 12808 9911 12860 9920
rect 12808 9877 12817 9911
rect 12817 9877 12851 9911
rect 12851 9877 12860 9911
rect 12808 9868 12860 9877
rect 13636 9911 13688 9920
rect 13636 9877 13645 9911
rect 13645 9877 13679 9911
rect 13679 9877 13688 9911
rect 13636 9868 13688 9877
rect 19248 9868 19300 9920
rect 24676 9911 24728 9920
rect 24676 9877 24685 9911
rect 24685 9877 24719 9911
rect 24719 9877 24728 9911
rect 24676 9868 24728 9877
rect 24860 9911 24912 9920
rect 24860 9877 24869 9911
rect 24869 9877 24903 9911
rect 24903 9877 24912 9911
rect 24860 9868 24912 9877
rect 26700 9911 26752 9920
rect 26700 9877 26709 9911
rect 26709 9877 26743 9911
rect 26743 9877 26752 9911
rect 26700 9868 26752 9877
rect 5982 9766 6034 9818
rect 6046 9766 6098 9818
rect 6110 9766 6162 9818
rect 6174 9766 6226 9818
rect 15982 9766 16034 9818
rect 16046 9766 16098 9818
rect 16110 9766 16162 9818
rect 16174 9766 16226 9818
rect 25982 9766 26034 9818
rect 26046 9766 26098 9818
rect 26110 9766 26162 9818
rect 26174 9766 26226 9818
rect 2504 9707 2556 9716
rect 2504 9673 2513 9707
rect 2513 9673 2547 9707
rect 2547 9673 2556 9707
rect 2504 9664 2556 9673
rect 5816 9664 5868 9716
rect 6736 9596 6788 9648
rect 2044 9571 2096 9580
rect 2044 9537 2053 9571
rect 2053 9537 2087 9571
rect 2087 9537 2096 9571
rect 2044 9528 2096 9537
rect 3516 9571 3568 9580
rect 3516 9537 3525 9571
rect 3525 9537 3559 9571
rect 3559 9537 3568 9571
rect 3516 9528 3568 9537
rect 8024 9664 8076 9716
rect 8208 9707 8260 9716
rect 8208 9673 8217 9707
rect 8217 9673 8251 9707
rect 8251 9673 8260 9707
rect 8208 9664 8260 9673
rect 9864 9664 9916 9716
rect 10692 9664 10744 9716
rect 13176 9664 13228 9716
rect 13452 9664 13504 9716
rect 14188 9707 14240 9716
rect 14188 9673 14197 9707
rect 14197 9673 14231 9707
rect 14231 9673 14240 9707
rect 14188 9664 14240 9673
rect 7288 9596 7340 9648
rect 7472 9596 7524 9648
rect 10876 9596 10928 9648
rect 7380 9571 7432 9580
rect 3792 9503 3844 9512
rect 3792 9469 3826 9503
rect 3826 9469 3844 9503
rect 3792 9460 3844 9469
rect 6092 9460 6144 9512
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 10968 9528 11020 9580
rect 6552 9460 6604 9512
rect 7748 9460 7800 9512
rect 9680 9460 9732 9512
rect 12808 9503 12860 9512
rect 6828 9392 6880 9444
rect 6920 9392 6972 9444
rect 1400 9324 1452 9376
rect 4252 9324 4304 9376
rect 5540 9324 5592 9376
rect 6736 9324 6788 9376
rect 12808 9469 12817 9503
rect 12817 9469 12851 9503
rect 12851 9469 12860 9503
rect 12808 9460 12860 9469
rect 12900 9460 12952 9512
rect 13452 9460 13504 9512
rect 15016 9503 15068 9512
rect 15016 9469 15025 9503
rect 15025 9469 15059 9503
rect 15059 9469 15068 9503
rect 15016 9460 15068 9469
rect 16304 9528 16356 9580
rect 16856 9664 16908 9716
rect 18696 9707 18748 9716
rect 18696 9673 18705 9707
rect 18705 9673 18739 9707
rect 18739 9673 18748 9707
rect 18696 9664 18748 9673
rect 19616 9664 19668 9716
rect 22008 9664 22060 9716
rect 25504 9664 25556 9716
rect 26516 9664 26568 9716
rect 19340 9528 19392 9580
rect 20628 9528 20680 9580
rect 25872 9528 25924 9580
rect 26332 9528 26384 9580
rect 13544 9392 13596 9444
rect 19432 9392 19484 9444
rect 22100 9460 22152 9512
rect 23664 9503 23716 9512
rect 23664 9469 23673 9503
rect 23673 9469 23707 9503
rect 23707 9469 23716 9503
rect 23664 9460 23716 9469
rect 26516 9460 26568 9512
rect 21456 9392 21508 9444
rect 24676 9392 24728 9444
rect 25964 9392 26016 9444
rect 16396 9367 16448 9376
rect 16396 9333 16405 9367
rect 16405 9333 16439 9367
rect 16439 9333 16448 9367
rect 16396 9324 16448 9333
rect 20444 9367 20496 9376
rect 20444 9333 20453 9367
rect 20453 9333 20487 9367
rect 20487 9333 20496 9367
rect 20444 9324 20496 9333
rect 23480 9367 23532 9376
rect 23480 9333 23489 9367
rect 23489 9333 23523 9367
rect 23523 9333 23532 9367
rect 23480 9324 23532 9333
rect 25044 9367 25096 9376
rect 25044 9333 25053 9367
rect 25053 9333 25087 9367
rect 25087 9333 25096 9367
rect 25044 9324 25096 9333
rect 25872 9367 25924 9376
rect 25872 9333 25881 9367
rect 25881 9333 25915 9367
rect 25915 9333 25924 9367
rect 25872 9324 25924 9333
rect 10982 9222 11034 9274
rect 11046 9222 11098 9274
rect 11110 9222 11162 9274
rect 11174 9222 11226 9274
rect 20982 9222 21034 9274
rect 21046 9222 21098 9274
rect 21110 9222 21162 9274
rect 21174 9222 21226 9274
rect 1676 9163 1728 9172
rect 1676 9129 1685 9163
rect 1685 9129 1719 9163
rect 1719 9129 1728 9163
rect 1676 9120 1728 9129
rect 3792 9120 3844 9172
rect 6092 9163 6144 9172
rect 6092 9129 6101 9163
rect 6101 9129 6135 9163
rect 6135 9129 6144 9163
rect 6092 9120 6144 9129
rect 6460 9163 6512 9172
rect 6460 9129 6469 9163
rect 6469 9129 6503 9163
rect 6503 9129 6512 9163
rect 6460 9120 6512 9129
rect 6828 9163 6880 9172
rect 6828 9129 6837 9163
rect 6837 9129 6871 9163
rect 6871 9129 6880 9163
rect 6828 9120 6880 9129
rect 11336 9120 11388 9172
rect 13728 9163 13780 9172
rect 13728 9129 13737 9163
rect 13737 9129 13771 9163
rect 13771 9129 13780 9163
rect 13728 9120 13780 9129
rect 14096 9163 14148 9172
rect 14096 9129 14105 9163
rect 14105 9129 14139 9163
rect 14139 9129 14148 9163
rect 14096 9120 14148 9129
rect 21364 9120 21416 9172
rect 22744 9120 22796 9172
rect 2504 9052 2556 9104
rect 3608 9052 3660 9104
rect 7288 9095 7340 9104
rect 7288 9061 7297 9095
rect 7297 9061 7331 9095
rect 7331 9061 7340 9095
rect 7288 9052 7340 9061
rect 10416 9052 10468 9104
rect 16396 9052 16448 9104
rect 17408 9095 17460 9104
rect 17408 9061 17420 9095
rect 17420 9061 17460 9095
rect 17408 9052 17460 9061
rect 21548 9052 21600 9104
rect 24860 9120 24912 9172
rect 25228 9163 25280 9172
rect 25228 9129 25237 9163
rect 25237 9129 25271 9163
rect 25271 9129 25280 9163
rect 25228 9120 25280 9129
rect 24676 9095 24728 9104
rect 24676 9061 24685 9095
rect 24685 9061 24719 9095
rect 24719 9061 24728 9095
rect 24676 9052 24728 9061
rect 25872 9052 25924 9104
rect 6460 8984 6512 9036
rect 7472 8984 7524 9036
rect 8116 8984 8168 9036
rect 8576 8984 8628 9036
rect 15016 8984 15068 9036
rect 17868 8984 17920 9036
rect 19340 8984 19392 9036
rect 20536 8984 20588 9036
rect 22836 9027 22888 9036
rect 22836 8993 22845 9027
rect 22845 8993 22879 9027
rect 22879 8993 22888 9027
rect 22836 8984 22888 8993
rect 2872 8959 2924 8968
rect 2872 8925 2881 8959
rect 2881 8925 2915 8959
rect 2915 8925 2924 8959
rect 2872 8916 2924 8925
rect 4252 8916 4304 8968
rect 7380 8959 7432 8968
rect 7380 8925 7389 8959
rect 7389 8925 7423 8959
rect 7423 8925 7432 8959
rect 7380 8916 7432 8925
rect 21364 8959 21416 8968
rect 21364 8925 21373 8959
rect 21373 8925 21407 8959
rect 21407 8925 21416 8959
rect 21364 8916 21416 8925
rect 21456 8959 21508 8968
rect 21456 8925 21465 8959
rect 21465 8925 21499 8959
rect 21499 8925 21508 8959
rect 23020 8959 23072 8968
rect 21456 8916 21508 8925
rect 23020 8925 23029 8959
rect 23029 8925 23063 8959
rect 23063 8925 23072 8959
rect 23020 8916 23072 8925
rect 25044 8916 25096 8968
rect 25872 8959 25924 8968
rect 25872 8925 25881 8959
rect 25881 8925 25915 8959
rect 25915 8925 25924 8959
rect 25872 8916 25924 8925
rect 2596 8780 2648 8832
rect 4896 8823 4948 8832
rect 4896 8789 4905 8823
rect 4905 8789 4939 8823
rect 4939 8789 4948 8823
rect 4896 8780 4948 8789
rect 9036 8780 9088 8832
rect 12808 8780 12860 8832
rect 13268 8780 13320 8832
rect 16488 8823 16540 8832
rect 16488 8789 16497 8823
rect 16497 8789 16531 8823
rect 16531 8789 16540 8823
rect 16488 8780 16540 8789
rect 18512 8823 18564 8832
rect 18512 8789 18521 8823
rect 18521 8789 18555 8823
rect 18555 8789 18564 8823
rect 18512 8780 18564 8789
rect 19432 8780 19484 8832
rect 19708 8780 19760 8832
rect 20444 8780 20496 8832
rect 20812 8780 20864 8832
rect 23664 8823 23716 8832
rect 23664 8789 23673 8823
rect 23673 8789 23707 8823
rect 23707 8789 23716 8823
rect 23664 8780 23716 8789
rect 5982 8678 6034 8730
rect 6046 8678 6098 8730
rect 6110 8678 6162 8730
rect 6174 8678 6226 8730
rect 15982 8678 16034 8730
rect 16046 8678 16098 8730
rect 16110 8678 16162 8730
rect 16174 8678 16226 8730
rect 25982 8678 26034 8730
rect 26046 8678 26098 8730
rect 26110 8678 26162 8730
rect 26174 8678 26226 8730
rect 2504 8619 2556 8628
rect 2504 8585 2513 8619
rect 2513 8585 2547 8619
rect 2547 8585 2556 8619
rect 2504 8576 2556 8585
rect 2872 8576 2924 8628
rect 8576 8619 8628 8628
rect 8576 8585 8585 8619
rect 8585 8585 8619 8619
rect 8619 8585 8628 8619
rect 8576 8576 8628 8585
rect 10416 8619 10468 8628
rect 10416 8585 10425 8619
rect 10425 8585 10459 8619
rect 10459 8585 10468 8619
rect 10416 8576 10468 8585
rect 13268 8576 13320 8628
rect 17408 8619 17460 8628
rect 17408 8585 17417 8619
rect 17417 8585 17451 8619
rect 17451 8585 17460 8619
rect 17408 8576 17460 8585
rect 17868 8619 17920 8628
rect 17868 8585 17877 8619
rect 17877 8585 17911 8619
rect 17911 8585 17920 8619
rect 17868 8576 17920 8585
rect 19340 8619 19392 8628
rect 19340 8585 19349 8619
rect 19349 8585 19383 8619
rect 19383 8585 19392 8619
rect 19340 8576 19392 8585
rect 21456 8576 21508 8628
rect 24676 8619 24728 8628
rect 24676 8585 24685 8619
rect 24685 8585 24719 8619
rect 24719 8585 24728 8619
rect 24676 8576 24728 8585
rect 24860 8576 24912 8628
rect 26608 8619 26660 8628
rect 26608 8585 26617 8619
rect 26617 8585 26651 8619
rect 26651 8585 26660 8619
rect 26608 8576 26660 8585
rect 1584 8551 1636 8560
rect 1584 8517 1593 8551
rect 1593 8517 1627 8551
rect 1627 8517 1636 8551
rect 1584 8508 1636 8517
rect 2872 8440 2924 8492
rect 3976 8508 4028 8560
rect 4344 8508 4396 8560
rect 3792 8483 3844 8492
rect 3792 8449 3801 8483
rect 3801 8449 3835 8483
rect 3835 8449 3844 8483
rect 3792 8440 3844 8449
rect 3516 8415 3568 8424
rect 3516 8381 3525 8415
rect 3525 8381 3559 8415
rect 3559 8381 3568 8415
rect 3516 8372 3568 8381
rect 4068 8372 4120 8424
rect 4528 8372 4580 8424
rect 5448 8440 5500 8492
rect 6920 8483 6972 8492
rect 6920 8449 6929 8483
rect 6929 8449 6963 8483
rect 6963 8449 6972 8483
rect 6920 8440 6972 8449
rect 16488 8440 16540 8492
rect 16856 8483 16908 8492
rect 16856 8449 16865 8483
rect 16865 8449 16899 8483
rect 16899 8449 16908 8483
rect 16856 8440 16908 8449
rect 4896 8372 4948 8424
rect 9036 8415 9088 8424
rect 9036 8381 9045 8415
rect 9045 8381 9079 8415
rect 9079 8381 9088 8415
rect 9036 8372 9088 8381
rect 10784 8372 10836 8424
rect 14924 8372 14976 8424
rect 16580 8372 16632 8424
rect 18512 8440 18564 8492
rect 22744 8440 22796 8492
rect 19708 8372 19760 8424
rect 26424 8415 26476 8424
rect 26424 8381 26433 8415
rect 26433 8381 26467 8415
rect 26467 8381 26476 8415
rect 26424 8372 26476 8381
rect 4620 8347 4672 8356
rect 4620 8313 4629 8347
rect 4629 8313 4663 8347
rect 4663 8313 4672 8347
rect 4620 8304 4672 8313
rect 6460 8304 6512 8356
rect 9588 8304 9640 8356
rect 15200 8304 15252 8356
rect 16304 8347 16356 8356
rect 16304 8313 16313 8347
rect 16313 8313 16347 8347
rect 16347 8313 16356 8347
rect 16304 8304 16356 8313
rect 4252 8279 4304 8288
rect 4252 8245 4261 8279
rect 4261 8245 4295 8279
rect 4295 8245 4304 8279
rect 4252 8236 4304 8245
rect 5264 8279 5316 8288
rect 5264 8245 5273 8279
rect 5273 8245 5307 8279
rect 5307 8245 5316 8279
rect 7472 8279 7524 8288
rect 5264 8236 5316 8245
rect 7472 8245 7481 8279
rect 7481 8245 7515 8279
rect 7515 8245 7524 8279
rect 7472 8236 7524 8245
rect 7932 8236 7984 8288
rect 10784 8236 10836 8288
rect 16396 8279 16448 8288
rect 16396 8245 16405 8279
rect 16405 8245 16439 8279
rect 16439 8245 16448 8279
rect 16396 8236 16448 8245
rect 22100 8304 22152 8356
rect 22836 8304 22888 8356
rect 23020 8236 23072 8288
rect 10982 8134 11034 8186
rect 11046 8134 11098 8186
rect 11110 8134 11162 8186
rect 11174 8134 11226 8186
rect 20982 8134 21034 8186
rect 21046 8134 21098 8186
rect 21110 8134 21162 8186
rect 21174 8134 21226 8186
rect 3516 8075 3568 8084
rect 3516 8041 3525 8075
rect 3525 8041 3559 8075
rect 3559 8041 3568 8075
rect 3516 8032 3568 8041
rect 5264 8032 5316 8084
rect 5540 8032 5592 8084
rect 7380 8032 7432 8084
rect 16488 8075 16540 8084
rect 16488 8041 16497 8075
rect 16497 8041 16531 8075
rect 16531 8041 16540 8075
rect 16488 8032 16540 8041
rect 16856 8032 16908 8084
rect 18512 8075 18564 8084
rect 18512 8041 18521 8075
rect 18521 8041 18555 8075
rect 18555 8041 18564 8075
rect 18512 8032 18564 8041
rect 20536 8075 20588 8084
rect 20536 8041 20545 8075
rect 20545 8041 20579 8075
rect 20579 8041 20588 8075
rect 20536 8032 20588 8041
rect 21364 8032 21416 8084
rect 21548 8075 21600 8084
rect 21548 8041 21557 8075
rect 21557 8041 21591 8075
rect 21591 8041 21600 8075
rect 21548 8032 21600 8041
rect 22008 8075 22060 8084
rect 22008 8041 22017 8075
rect 22017 8041 22051 8075
rect 22051 8041 22060 8075
rect 22008 8032 22060 8041
rect 22836 8032 22888 8084
rect 26700 8075 26752 8084
rect 26700 8041 26709 8075
rect 26709 8041 26743 8075
rect 26743 8041 26752 8075
rect 26700 8032 26752 8041
rect 2780 8007 2832 8016
rect 2780 7973 2789 8007
rect 2789 7973 2823 8007
rect 2823 7973 2832 8007
rect 2780 7964 2832 7973
rect 11336 7964 11388 8016
rect 18052 7964 18104 8016
rect 3424 7896 3476 7948
rect 5172 7939 5224 7948
rect 5172 7905 5181 7939
rect 5181 7905 5215 7939
rect 5215 7905 5224 7939
rect 5172 7896 5224 7905
rect 5816 7896 5868 7948
rect 16948 7896 17000 7948
rect 17316 7939 17368 7948
rect 17316 7905 17325 7939
rect 17325 7905 17359 7939
rect 17359 7905 17368 7939
rect 17316 7896 17368 7905
rect 20720 7896 20772 7948
rect 21824 7896 21876 7948
rect 22376 7939 22428 7948
rect 22376 7905 22385 7939
rect 22385 7905 22419 7939
rect 22419 7905 22428 7939
rect 22376 7896 22428 7905
rect 23848 7896 23900 7948
rect 25228 7896 25280 7948
rect 26516 7939 26568 7948
rect 26516 7905 26525 7939
rect 26525 7905 26559 7939
rect 26559 7905 26568 7939
rect 26516 7896 26568 7905
rect 4252 7828 4304 7880
rect 10784 7828 10836 7880
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 17500 7871 17552 7880
rect 17500 7837 17509 7871
rect 17509 7837 17543 7871
rect 17543 7837 17552 7871
rect 17500 7828 17552 7837
rect 22652 7871 22704 7880
rect 22652 7837 22661 7871
rect 22661 7837 22695 7871
rect 22695 7837 22704 7871
rect 22652 7828 22704 7837
rect 23388 7828 23440 7880
rect 24032 7871 24084 7880
rect 24032 7837 24041 7871
rect 24041 7837 24075 7871
rect 24075 7837 24084 7871
rect 24032 7828 24084 7837
rect 24308 7828 24360 7880
rect 1860 7692 1912 7744
rect 2412 7735 2464 7744
rect 2412 7701 2421 7735
rect 2421 7701 2455 7735
rect 2455 7701 2464 7735
rect 2412 7692 2464 7701
rect 3976 7692 4028 7744
rect 8300 7692 8352 7744
rect 9036 7735 9088 7744
rect 9036 7701 9045 7735
rect 9045 7701 9079 7735
rect 9079 7701 9088 7735
rect 9036 7692 9088 7701
rect 12348 7692 12400 7744
rect 18052 7735 18104 7744
rect 18052 7701 18061 7735
rect 18061 7701 18095 7735
rect 18095 7701 18104 7735
rect 18052 7692 18104 7701
rect 19708 7692 19760 7744
rect 25320 7735 25372 7744
rect 25320 7701 25329 7735
rect 25329 7701 25363 7735
rect 25363 7701 25372 7735
rect 25320 7692 25372 7701
rect 5982 7590 6034 7642
rect 6046 7590 6098 7642
rect 6110 7590 6162 7642
rect 6174 7590 6226 7642
rect 15982 7590 16034 7642
rect 16046 7590 16098 7642
rect 16110 7590 16162 7642
rect 16174 7590 16226 7642
rect 25982 7590 26034 7642
rect 26046 7590 26098 7642
rect 26110 7590 26162 7642
rect 26174 7590 26226 7642
rect 2780 7488 2832 7540
rect 4988 7531 5040 7540
rect 4988 7497 4997 7531
rect 4997 7497 5031 7531
rect 5031 7497 5040 7531
rect 4988 7488 5040 7497
rect 5264 7488 5316 7540
rect 15016 7488 15068 7540
rect 17500 7488 17552 7540
rect 21824 7531 21876 7540
rect 21824 7497 21833 7531
rect 21833 7497 21867 7531
rect 21867 7497 21876 7531
rect 21824 7488 21876 7497
rect 22744 7488 22796 7540
rect 23112 7531 23164 7540
rect 23112 7497 23121 7531
rect 23121 7497 23155 7531
rect 23155 7497 23164 7531
rect 23112 7488 23164 7497
rect 24032 7488 24084 7540
rect 24768 7531 24820 7540
rect 24768 7497 24777 7531
rect 24777 7497 24811 7531
rect 24811 7497 24820 7531
rect 24768 7488 24820 7497
rect 25228 7488 25280 7540
rect 26516 7488 26568 7540
rect 26332 7420 26384 7472
rect 2872 7352 2924 7404
rect 4252 7352 4304 7404
rect 5816 7395 5868 7404
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 6276 7352 6328 7404
rect 12164 7395 12216 7404
rect 12164 7361 12173 7395
rect 12173 7361 12207 7395
rect 12207 7361 12216 7395
rect 12164 7352 12216 7361
rect 13084 7395 13136 7404
rect 13084 7361 13093 7395
rect 13093 7361 13127 7395
rect 13127 7361 13136 7395
rect 13084 7352 13136 7361
rect 14648 7395 14700 7404
rect 14648 7361 14657 7395
rect 14657 7361 14691 7395
rect 14691 7361 14700 7395
rect 14648 7352 14700 7361
rect 18604 7395 18656 7404
rect 18604 7361 18613 7395
rect 18613 7361 18647 7395
rect 18647 7361 18656 7395
rect 18604 7352 18656 7361
rect 22284 7352 22336 7404
rect 22468 7395 22520 7404
rect 22468 7361 22477 7395
rect 22477 7361 22511 7395
rect 22511 7361 22520 7395
rect 22468 7352 22520 7361
rect 4068 7284 4120 7336
rect 5172 7284 5224 7336
rect 8300 7327 8352 7336
rect 8300 7293 8309 7327
rect 8309 7293 8343 7327
rect 8343 7293 8352 7327
rect 8300 7284 8352 7293
rect 1676 7259 1728 7268
rect 1676 7225 1710 7259
rect 1710 7225 1728 7259
rect 1676 7216 1728 7225
rect 1860 7216 1912 7268
rect 5632 7259 5684 7268
rect 5632 7225 5641 7259
rect 5641 7225 5675 7259
rect 5675 7225 5684 7259
rect 5632 7216 5684 7225
rect 9864 7216 9916 7268
rect 12900 7259 12952 7268
rect 2872 7148 2924 7200
rect 3424 7191 3476 7200
rect 3424 7157 3433 7191
rect 3433 7157 3467 7191
rect 3467 7157 3476 7191
rect 3424 7148 3476 7157
rect 3516 7148 3568 7200
rect 4068 7191 4120 7200
rect 4068 7157 4077 7191
rect 4077 7157 4111 7191
rect 4111 7157 4120 7191
rect 4068 7148 4120 7157
rect 4988 7148 5040 7200
rect 6276 7191 6328 7200
rect 6276 7157 6285 7191
rect 6285 7157 6319 7191
rect 6319 7157 6328 7191
rect 6276 7148 6328 7157
rect 6828 7191 6880 7200
rect 6828 7157 6837 7191
rect 6837 7157 6871 7191
rect 6871 7157 6880 7191
rect 6828 7148 6880 7157
rect 9680 7191 9732 7200
rect 9680 7157 9689 7191
rect 9689 7157 9723 7191
rect 9723 7157 9732 7191
rect 9680 7148 9732 7157
rect 10784 7191 10836 7200
rect 10784 7157 10793 7191
rect 10793 7157 10827 7191
rect 10827 7157 10836 7191
rect 10784 7148 10836 7157
rect 11336 7148 11388 7200
rect 11704 7148 11756 7200
rect 12900 7225 12909 7259
rect 12909 7225 12943 7259
rect 12943 7225 12952 7259
rect 12900 7216 12952 7225
rect 16488 7284 16540 7336
rect 18420 7327 18472 7336
rect 18420 7293 18429 7327
rect 18429 7293 18463 7327
rect 18463 7293 18472 7327
rect 18420 7284 18472 7293
rect 22008 7284 22060 7336
rect 22652 7352 22704 7404
rect 23480 7395 23532 7404
rect 23480 7361 23489 7395
rect 23489 7361 23523 7395
rect 23523 7361 23532 7395
rect 24124 7395 24176 7404
rect 23480 7352 23532 7361
rect 24124 7361 24133 7395
rect 24133 7361 24167 7395
rect 24167 7361 24176 7395
rect 24124 7352 24176 7361
rect 24308 7395 24360 7404
rect 24308 7361 24317 7395
rect 24317 7361 24351 7395
rect 24351 7361 24360 7395
rect 24308 7352 24360 7361
rect 24768 7284 24820 7336
rect 25320 7327 25372 7336
rect 25320 7293 25329 7327
rect 25329 7293 25363 7327
rect 25363 7293 25372 7327
rect 25320 7284 25372 7293
rect 12256 7148 12308 7200
rect 12808 7191 12860 7200
rect 12808 7157 12817 7191
rect 12817 7157 12851 7191
rect 12851 7157 12860 7191
rect 16672 7216 16724 7268
rect 17316 7259 17368 7268
rect 17316 7225 17325 7259
rect 17325 7225 17359 7259
rect 17359 7225 17368 7259
rect 17316 7216 17368 7225
rect 18144 7216 18196 7268
rect 22284 7216 22336 7268
rect 12808 7148 12860 7157
rect 15844 7148 15896 7200
rect 16948 7191 17000 7200
rect 16948 7157 16957 7191
rect 16957 7157 16991 7191
rect 16991 7157 17000 7191
rect 16948 7148 17000 7157
rect 17868 7148 17920 7200
rect 10982 7046 11034 7098
rect 11046 7046 11098 7098
rect 11110 7046 11162 7098
rect 11174 7046 11226 7098
rect 20982 7046 21034 7098
rect 21046 7046 21098 7098
rect 21110 7046 21162 7098
rect 21174 7046 21226 7098
rect 1676 6987 1728 6996
rect 1676 6953 1685 6987
rect 1685 6953 1719 6987
rect 1719 6953 1728 6987
rect 1676 6944 1728 6953
rect 2412 6944 2464 6996
rect 2780 6944 2832 6996
rect 5816 6944 5868 6996
rect 6828 6944 6880 6996
rect 11336 6944 11388 6996
rect 13084 6944 13136 6996
rect 13360 6944 13412 6996
rect 13820 6944 13872 6996
rect 14648 6987 14700 6996
rect 14648 6953 14657 6987
rect 14657 6953 14691 6987
rect 14691 6953 14700 6987
rect 14648 6944 14700 6953
rect 22008 6987 22060 6996
rect 22008 6953 22017 6987
rect 22017 6953 22051 6987
rect 22051 6953 22060 6987
rect 22008 6944 22060 6953
rect 22468 6987 22520 6996
rect 22468 6953 22477 6987
rect 22477 6953 22511 6987
rect 22511 6953 22520 6987
rect 22468 6944 22520 6953
rect 24584 6944 24636 6996
rect 4068 6876 4120 6928
rect 4344 6851 4396 6860
rect 4344 6817 4353 6851
rect 4353 6817 4387 6851
rect 4387 6817 4396 6851
rect 4344 6808 4396 6817
rect 5632 6876 5684 6928
rect 8300 6876 8352 6928
rect 9680 6876 9732 6928
rect 10784 6876 10836 6928
rect 12256 6919 12308 6928
rect 12256 6885 12265 6919
rect 12265 6885 12299 6919
rect 12299 6885 12308 6919
rect 21272 6919 21324 6928
rect 12256 6876 12308 6885
rect 21272 6885 21281 6919
rect 21281 6885 21315 6919
rect 21315 6885 21324 6919
rect 21272 6876 21324 6885
rect 22836 6919 22888 6928
rect 22836 6885 22845 6919
rect 22845 6885 22879 6919
rect 22879 6885 22888 6919
rect 22836 6876 22888 6885
rect 5448 6808 5500 6860
rect 6000 6808 6052 6860
rect 2964 6783 3016 6792
rect 2596 6604 2648 6656
rect 2964 6749 2973 6783
rect 2973 6749 3007 6783
rect 3007 6749 3016 6783
rect 2964 6740 3016 6749
rect 6276 6740 6328 6792
rect 7196 6740 7248 6792
rect 4896 6672 4948 6724
rect 9128 6672 9180 6724
rect 2872 6604 2924 6656
rect 10416 6647 10468 6656
rect 10416 6613 10425 6647
rect 10425 6613 10459 6647
rect 10459 6613 10468 6647
rect 10416 6604 10468 6613
rect 13728 6808 13780 6860
rect 16396 6808 16448 6860
rect 12348 6783 12400 6792
rect 12348 6749 12357 6783
rect 12357 6749 12391 6783
rect 12391 6749 12400 6783
rect 12348 6740 12400 6749
rect 14004 6783 14056 6792
rect 14004 6749 14013 6783
rect 14013 6749 14047 6783
rect 14047 6749 14056 6783
rect 14004 6740 14056 6749
rect 13084 6672 13136 6724
rect 16948 6851 17000 6860
rect 16948 6817 16957 6851
rect 16957 6817 16991 6851
rect 16991 6817 17000 6851
rect 16948 6808 17000 6817
rect 17868 6808 17920 6860
rect 18420 6851 18472 6860
rect 18420 6817 18429 6851
rect 18429 6817 18463 6851
rect 18463 6817 18472 6851
rect 18420 6808 18472 6817
rect 18512 6851 18564 6860
rect 18512 6817 18521 6851
rect 18521 6817 18555 6851
rect 18555 6817 18564 6851
rect 21364 6851 21416 6860
rect 18512 6808 18564 6817
rect 21364 6817 21373 6851
rect 21373 6817 21407 6851
rect 21407 6817 21416 6851
rect 21364 6808 21416 6817
rect 26976 6808 27028 6860
rect 17132 6783 17184 6792
rect 17132 6749 17141 6783
rect 17141 6749 17175 6783
rect 17175 6749 17184 6783
rect 17132 6740 17184 6749
rect 18604 6783 18656 6792
rect 18604 6749 18613 6783
rect 18613 6749 18647 6783
rect 18647 6749 18656 6783
rect 18604 6740 18656 6749
rect 21824 6740 21876 6792
rect 21916 6740 21968 6792
rect 23940 6783 23992 6792
rect 23940 6749 23949 6783
rect 23949 6749 23983 6783
rect 23983 6749 23992 6783
rect 23940 6740 23992 6749
rect 24308 6740 24360 6792
rect 16856 6672 16908 6724
rect 22284 6672 22336 6724
rect 13360 6647 13412 6656
rect 13360 6613 13369 6647
rect 13369 6613 13403 6647
rect 13403 6613 13412 6647
rect 13360 6604 13412 6613
rect 16580 6604 16632 6656
rect 20720 6604 20772 6656
rect 26700 6715 26752 6724
rect 26700 6681 26709 6715
rect 26709 6681 26743 6715
rect 26743 6681 26752 6715
rect 26700 6672 26752 6681
rect 25044 6604 25096 6656
rect 5982 6502 6034 6554
rect 6046 6502 6098 6554
rect 6110 6502 6162 6554
rect 6174 6502 6226 6554
rect 15982 6502 16034 6554
rect 16046 6502 16098 6554
rect 16110 6502 16162 6554
rect 16174 6502 16226 6554
rect 25982 6502 26034 6554
rect 26046 6502 26098 6554
rect 26110 6502 26162 6554
rect 26174 6502 26226 6554
rect 1492 6400 1544 6452
rect 2044 6443 2096 6452
rect 2044 6409 2053 6443
rect 2053 6409 2087 6443
rect 2087 6409 2096 6443
rect 2044 6400 2096 6409
rect 2596 6400 2648 6452
rect 2780 6400 2832 6452
rect 5448 6443 5500 6452
rect 5448 6409 5457 6443
rect 5457 6409 5491 6443
rect 5491 6409 5500 6443
rect 5448 6400 5500 6409
rect 5816 6443 5868 6452
rect 5816 6409 5825 6443
rect 5825 6409 5859 6443
rect 5859 6409 5868 6443
rect 5816 6400 5868 6409
rect 6276 6400 6328 6452
rect 6552 6443 6604 6452
rect 6552 6409 6561 6443
rect 6561 6409 6595 6443
rect 6595 6409 6604 6443
rect 6552 6400 6604 6409
rect 1676 6332 1728 6384
rect 2964 6332 3016 6384
rect 6552 6264 6604 6316
rect 6736 6264 6788 6316
rect 9864 6400 9916 6452
rect 12256 6443 12308 6452
rect 8300 6332 8352 6384
rect 7564 6264 7616 6316
rect 8852 6264 8904 6316
rect 12256 6409 12265 6443
rect 12265 6409 12299 6443
rect 12299 6409 12308 6443
rect 12256 6400 12308 6409
rect 13360 6400 13412 6452
rect 13820 6443 13872 6452
rect 13820 6409 13829 6443
rect 13829 6409 13863 6443
rect 13863 6409 13872 6443
rect 13820 6400 13872 6409
rect 18512 6443 18564 6452
rect 18512 6409 18521 6443
rect 18521 6409 18555 6443
rect 18555 6409 18564 6443
rect 18512 6400 18564 6409
rect 21272 6400 21324 6452
rect 2044 6196 2096 6248
rect 7196 6239 7248 6248
rect 7196 6205 7205 6239
rect 7205 6205 7239 6239
rect 7239 6205 7248 6239
rect 7196 6196 7248 6205
rect 9588 6264 9640 6316
rect 10416 6264 10468 6316
rect 10692 6264 10744 6316
rect 12348 6332 12400 6384
rect 13728 6332 13780 6384
rect 17592 6332 17644 6384
rect 18604 6332 18656 6384
rect 21364 6375 21416 6384
rect 21364 6341 21373 6375
rect 21373 6341 21407 6375
rect 21407 6341 21416 6375
rect 21364 6332 21416 6341
rect 16396 6264 16448 6316
rect 15844 6239 15896 6248
rect 15844 6205 15853 6239
rect 15853 6205 15887 6239
rect 15887 6205 15896 6239
rect 18420 6264 18472 6316
rect 21824 6400 21876 6452
rect 24308 6400 24360 6452
rect 26976 6443 27028 6452
rect 26976 6409 26985 6443
rect 26985 6409 27019 6443
rect 27019 6409 27028 6443
rect 26976 6400 27028 6409
rect 23940 6375 23992 6384
rect 23940 6341 23949 6375
rect 23949 6341 23983 6375
rect 23983 6341 23992 6375
rect 23940 6332 23992 6341
rect 23572 6264 23624 6316
rect 24584 6264 24636 6316
rect 17132 6239 17184 6248
rect 15844 6196 15896 6205
rect 17132 6205 17141 6239
rect 17141 6205 17175 6239
rect 17175 6205 17184 6239
rect 17132 6196 17184 6205
rect 19708 6239 19760 6248
rect 19708 6205 19717 6239
rect 19717 6205 19751 6239
rect 19751 6205 19760 6239
rect 19708 6196 19760 6205
rect 9128 6171 9180 6180
rect 9128 6137 9137 6171
rect 9137 6137 9171 6171
rect 9171 6137 9180 6171
rect 9128 6128 9180 6137
rect 10416 6128 10468 6180
rect 17040 6128 17092 6180
rect 21824 6128 21876 6180
rect 26240 6171 26292 6180
rect 26240 6137 26249 6171
rect 26249 6137 26283 6171
rect 26283 6137 26292 6171
rect 26240 6128 26292 6137
rect 6828 6103 6880 6112
rect 6828 6069 6837 6103
rect 6837 6069 6871 6103
rect 6871 6069 6880 6103
rect 6828 6060 6880 6069
rect 14004 6060 14056 6112
rect 15200 6060 15252 6112
rect 16120 6103 16172 6112
rect 16120 6069 16129 6103
rect 16129 6069 16163 6103
rect 16163 6069 16172 6103
rect 16120 6060 16172 6069
rect 21272 6060 21324 6112
rect 26608 6103 26660 6112
rect 26608 6069 26617 6103
rect 26617 6069 26651 6103
rect 26651 6069 26660 6103
rect 26608 6060 26660 6069
rect 10982 5958 11034 6010
rect 11046 5958 11098 6010
rect 11110 5958 11162 6010
rect 11174 5958 11226 6010
rect 20982 5958 21034 6010
rect 21046 5958 21098 6010
rect 21110 5958 21162 6010
rect 21174 5958 21226 6010
rect 7196 5856 7248 5908
rect 8852 5899 8904 5908
rect 8852 5865 8861 5899
rect 8861 5865 8895 5899
rect 8895 5865 8904 5899
rect 8852 5856 8904 5865
rect 10416 5899 10468 5908
rect 10416 5865 10425 5899
rect 10425 5865 10459 5899
rect 10459 5865 10468 5899
rect 10416 5856 10468 5865
rect 10508 5856 10560 5908
rect 15844 5856 15896 5908
rect 16120 5856 16172 5908
rect 16856 5899 16908 5908
rect 16856 5865 16865 5899
rect 16865 5865 16899 5899
rect 16899 5865 16908 5899
rect 16856 5856 16908 5865
rect 17040 5899 17092 5908
rect 17040 5865 17049 5899
rect 17049 5865 17083 5899
rect 17083 5865 17092 5899
rect 17040 5856 17092 5865
rect 17408 5899 17460 5908
rect 17408 5865 17417 5899
rect 17417 5865 17451 5899
rect 17451 5865 17460 5899
rect 17408 5856 17460 5865
rect 2320 5788 2372 5840
rect 2872 5788 2924 5840
rect 4804 5788 4856 5840
rect 5172 5788 5224 5840
rect 7932 5788 7984 5840
rect 10232 5788 10284 5840
rect 16948 5788 17000 5840
rect 19708 5788 19760 5840
rect 22192 5788 22244 5840
rect 1768 5695 1820 5704
rect 1768 5661 1777 5695
rect 1777 5661 1811 5695
rect 1811 5661 1820 5695
rect 1768 5652 1820 5661
rect 7656 5720 7708 5772
rect 11980 5720 12032 5772
rect 12348 5763 12400 5772
rect 12348 5729 12357 5763
rect 12357 5729 12391 5763
rect 12391 5729 12400 5763
rect 12348 5720 12400 5729
rect 16488 5720 16540 5772
rect 21180 5720 21232 5772
rect 26516 5763 26568 5772
rect 26516 5729 26525 5763
rect 26525 5729 26559 5763
rect 26559 5729 26568 5763
rect 26516 5720 26568 5729
rect 26976 5720 27028 5772
rect 7564 5695 7616 5704
rect 7564 5661 7573 5695
rect 7573 5661 7607 5695
rect 7607 5661 7616 5695
rect 7564 5652 7616 5661
rect 11336 5652 11388 5704
rect 12072 5652 12124 5704
rect 16304 5652 16356 5704
rect 17500 5695 17552 5704
rect 17500 5661 17509 5695
rect 17509 5661 17543 5695
rect 17543 5661 17552 5695
rect 17500 5652 17552 5661
rect 17592 5695 17644 5704
rect 17592 5661 17601 5695
rect 17601 5661 17635 5695
rect 17635 5661 17644 5695
rect 17592 5652 17644 5661
rect 20260 5652 20312 5704
rect 21824 5652 21876 5704
rect 3148 5559 3200 5568
rect 3148 5525 3157 5559
rect 3157 5525 3191 5559
rect 3191 5525 3200 5559
rect 3148 5516 3200 5525
rect 6276 5516 6328 5568
rect 7012 5559 7064 5568
rect 7012 5525 7021 5559
rect 7021 5525 7055 5559
rect 7055 5525 7064 5559
rect 7012 5516 7064 5525
rect 11428 5559 11480 5568
rect 11428 5525 11437 5559
rect 11437 5525 11471 5559
rect 11471 5525 11480 5559
rect 11428 5516 11480 5525
rect 12900 5516 12952 5568
rect 13360 5559 13412 5568
rect 13360 5525 13369 5559
rect 13369 5525 13403 5559
rect 13403 5525 13412 5559
rect 13360 5516 13412 5525
rect 15476 5559 15528 5568
rect 15476 5525 15485 5559
rect 15485 5525 15519 5559
rect 15519 5525 15528 5559
rect 15476 5516 15528 5525
rect 20904 5559 20956 5568
rect 20904 5525 20913 5559
rect 20913 5525 20947 5559
rect 20947 5525 20956 5559
rect 20904 5516 20956 5525
rect 23664 5559 23716 5568
rect 23664 5525 23673 5559
rect 23673 5525 23707 5559
rect 23707 5525 23716 5559
rect 23664 5516 23716 5525
rect 26792 5516 26844 5568
rect 5982 5414 6034 5466
rect 6046 5414 6098 5466
rect 6110 5414 6162 5466
rect 6174 5414 6226 5466
rect 15982 5414 16034 5466
rect 16046 5414 16098 5466
rect 16110 5414 16162 5466
rect 16174 5414 16226 5466
rect 25982 5414 26034 5466
rect 26046 5414 26098 5466
rect 26110 5414 26162 5466
rect 26174 5414 26226 5466
rect 1584 5355 1636 5364
rect 1584 5321 1593 5355
rect 1593 5321 1627 5355
rect 1627 5321 1636 5355
rect 1584 5312 1636 5321
rect 2320 5355 2372 5364
rect 2320 5321 2329 5355
rect 2329 5321 2363 5355
rect 2363 5321 2372 5355
rect 2320 5312 2372 5321
rect 3148 5312 3200 5364
rect 5172 5355 5224 5364
rect 5172 5321 5181 5355
rect 5181 5321 5215 5355
rect 5215 5321 5224 5355
rect 5172 5312 5224 5321
rect 6276 5355 6328 5364
rect 6276 5321 6285 5355
rect 6285 5321 6319 5355
rect 6319 5321 6328 5355
rect 6276 5312 6328 5321
rect 7932 5355 7984 5364
rect 7932 5321 7941 5355
rect 7941 5321 7975 5355
rect 7975 5321 7984 5355
rect 7932 5312 7984 5321
rect 10508 5312 10560 5364
rect 10692 5355 10744 5364
rect 10692 5321 10701 5355
rect 10701 5321 10735 5355
rect 10735 5321 10744 5355
rect 10692 5312 10744 5321
rect 12072 5355 12124 5364
rect 12072 5321 12081 5355
rect 12081 5321 12115 5355
rect 12115 5321 12124 5355
rect 12072 5312 12124 5321
rect 14004 5355 14056 5364
rect 14004 5321 14013 5355
rect 14013 5321 14047 5355
rect 14047 5321 14056 5355
rect 14004 5312 14056 5321
rect 16304 5312 16356 5364
rect 16580 5355 16632 5364
rect 16580 5321 16589 5355
rect 16589 5321 16623 5355
rect 16623 5321 16632 5355
rect 16580 5312 16632 5321
rect 17500 5355 17552 5364
rect 17500 5321 17509 5355
rect 17509 5321 17543 5355
rect 17543 5321 17552 5355
rect 17500 5312 17552 5321
rect 17592 5312 17644 5364
rect 21180 5312 21232 5364
rect 25044 5355 25096 5364
rect 25044 5321 25053 5355
rect 25053 5321 25087 5355
rect 25087 5321 25096 5355
rect 25044 5312 25096 5321
rect 26976 5355 27028 5364
rect 26976 5321 26985 5355
rect 26985 5321 27019 5355
rect 27019 5321 27028 5355
rect 26976 5312 27028 5321
rect 2044 5219 2096 5228
rect 2044 5185 2053 5219
rect 2053 5185 2087 5219
rect 2087 5185 2096 5219
rect 2044 5176 2096 5185
rect 6644 5219 6696 5228
rect 6644 5185 6653 5219
rect 6653 5185 6687 5219
rect 6687 5185 6696 5219
rect 6644 5176 6696 5185
rect 7012 5176 7064 5228
rect 10232 5244 10284 5296
rect 17408 5244 17460 5296
rect 20260 5287 20312 5296
rect 20260 5253 20269 5287
rect 20269 5253 20303 5287
rect 20303 5253 20312 5287
rect 20260 5244 20312 5253
rect 20628 5244 20680 5296
rect 21364 5244 21416 5296
rect 7472 5176 7524 5228
rect 10784 5176 10836 5228
rect 11336 5219 11388 5228
rect 11336 5185 11345 5219
rect 11345 5185 11379 5219
rect 11379 5185 11388 5219
rect 11336 5176 11388 5185
rect 14648 5176 14700 5228
rect 20904 5219 20956 5228
rect 20904 5185 20913 5219
rect 20913 5185 20947 5219
rect 20947 5185 20956 5219
rect 20904 5176 20956 5185
rect 21272 5176 21324 5228
rect 22192 5176 22244 5228
rect 23664 5219 23716 5228
rect 23664 5185 23673 5219
rect 23673 5185 23707 5219
rect 23707 5185 23716 5219
rect 23664 5176 23716 5185
rect 3608 5108 3660 5160
rect 6920 5108 6972 5160
rect 13360 5108 13412 5160
rect 20720 5108 20772 5160
rect 22376 5108 22428 5160
rect 3148 5040 3200 5092
rect 11428 5040 11480 5092
rect 12900 5083 12952 5092
rect 12900 5049 12934 5083
rect 12934 5049 12952 5083
rect 12900 5040 12952 5049
rect 15108 5083 15160 5092
rect 15108 5049 15120 5083
rect 15120 5049 15160 5083
rect 15108 5040 15160 5049
rect 26240 5083 26292 5092
rect 26240 5049 26249 5083
rect 26249 5049 26283 5083
rect 26283 5049 26292 5083
rect 26240 5040 26292 5049
rect 3700 4972 3752 5024
rect 4804 5015 4856 5024
rect 4804 4981 4813 5015
rect 4813 4981 4847 5015
rect 4847 4981 4856 5015
rect 4804 4972 4856 4981
rect 6828 5015 6880 5024
rect 6828 4981 6837 5015
rect 6837 4981 6871 5015
rect 6871 4981 6880 5015
rect 6828 4972 6880 4981
rect 11336 4972 11388 5024
rect 11612 4972 11664 5024
rect 16672 4972 16724 5024
rect 20444 5015 20496 5024
rect 20444 4981 20453 5015
rect 20453 4981 20487 5015
rect 20487 4981 20496 5015
rect 20444 4972 20496 4981
rect 23572 4972 23624 5024
rect 26608 5015 26660 5024
rect 26608 4981 26617 5015
rect 26617 4981 26651 5015
rect 26651 4981 26660 5015
rect 26608 4972 26660 4981
rect 10982 4870 11034 4922
rect 11046 4870 11098 4922
rect 11110 4870 11162 4922
rect 11174 4870 11226 4922
rect 20982 4870 21034 4922
rect 21046 4870 21098 4922
rect 21110 4870 21162 4922
rect 21174 4870 21226 4922
rect 1584 4811 1636 4820
rect 1584 4777 1593 4811
rect 1593 4777 1627 4811
rect 1627 4777 1636 4811
rect 1584 4768 1636 4777
rect 3148 4811 3200 4820
rect 3148 4777 3157 4811
rect 3157 4777 3191 4811
rect 3191 4777 3200 4811
rect 3148 4768 3200 4777
rect 1768 4700 1820 4752
rect 3608 4768 3660 4820
rect 5172 4768 5224 4820
rect 6368 4811 6420 4820
rect 6368 4777 6377 4811
rect 6377 4777 6411 4811
rect 6411 4777 6420 4811
rect 6368 4768 6420 4777
rect 7012 4768 7064 4820
rect 10784 4811 10836 4820
rect 10784 4777 10793 4811
rect 10793 4777 10827 4811
rect 10827 4777 10836 4811
rect 10784 4768 10836 4777
rect 11336 4811 11388 4820
rect 11336 4777 11345 4811
rect 11345 4777 11379 4811
rect 11379 4777 11388 4811
rect 11336 4768 11388 4777
rect 11428 4768 11480 4820
rect 13268 4811 13320 4820
rect 13268 4777 13277 4811
rect 13277 4777 13311 4811
rect 13311 4777 13320 4811
rect 13268 4768 13320 4777
rect 13452 4768 13504 4820
rect 14648 4768 14700 4820
rect 15844 4811 15896 4820
rect 5724 4700 5776 4752
rect 8116 4700 8168 4752
rect 11796 4743 11848 4752
rect 11796 4709 11805 4743
rect 11805 4709 11839 4743
rect 11839 4709 11848 4743
rect 11796 4700 11848 4709
rect 2044 4675 2096 4684
rect 2044 4641 2053 4675
rect 2053 4641 2087 4675
rect 2087 4641 2096 4675
rect 2044 4632 2096 4641
rect 2504 4675 2556 4684
rect 2504 4641 2513 4675
rect 2513 4641 2547 4675
rect 2547 4641 2556 4675
rect 2504 4632 2556 4641
rect 4068 4675 4120 4684
rect 4068 4641 4077 4675
rect 4077 4641 4111 4675
rect 4111 4641 4120 4675
rect 4068 4632 4120 4641
rect 11612 4632 11664 4684
rect 15844 4777 15853 4811
rect 15853 4777 15887 4811
rect 15887 4777 15896 4811
rect 15844 4768 15896 4777
rect 19708 4768 19760 4820
rect 20444 4768 20496 4820
rect 21272 4768 21324 4820
rect 21364 4768 21416 4820
rect 22100 4768 22152 4820
rect 27344 4768 27396 4820
rect 27804 4768 27856 4820
rect 16304 4743 16356 4752
rect 16304 4709 16338 4743
rect 16338 4709 16356 4743
rect 16304 4700 16356 4709
rect 16396 4700 16448 4752
rect 22376 4700 22428 4752
rect 18052 4675 18104 4684
rect 18052 4641 18061 4675
rect 18061 4641 18095 4675
rect 18095 4641 18104 4675
rect 18052 4632 18104 4641
rect 21364 4632 21416 4684
rect 21824 4632 21876 4684
rect 26516 4675 26568 4684
rect 26516 4641 26525 4675
rect 26525 4641 26559 4675
rect 26559 4641 26568 4675
rect 26516 4632 26568 4641
rect 6460 4607 6512 4616
rect 6460 4573 6469 4607
rect 6469 4573 6503 4607
rect 6503 4573 6512 4607
rect 6460 4564 6512 4573
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 7564 4564 7616 4616
rect 11980 4607 12032 4616
rect 11980 4573 11989 4607
rect 11989 4573 12023 4607
rect 12023 4573 12032 4607
rect 11980 4564 12032 4573
rect 12900 4564 12952 4616
rect 13544 4607 13596 4616
rect 13544 4573 13553 4607
rect 13553 4573 13587 4607
rect 13587 4573 13596 4607
rect 13544 4564 13596 4573
rect 19616 4564 19668 4616
rect 19892 4607 19944 4616
rect 19892 4573 19901 4607
rect 19901 4573 19935 4607
rect 19935 4573 19944 4607
rect 19892 4564 19944 4573
rect 22192 4607 22244 4616
rect 22192 4573 22201 4607
rect 22201 4573 22235 4607
rect 22235 4573 22244 4607
rect 22192 4564 22244 4573
rect 23572 4539 23624 4548
rect 23572 4505 23581 4539
rect 23581 4505 23615 4539
rect 23615 4505 23624 4539
rect 23572 4496 23624 4505
rect 2688 4471 2740 4480
rect 2688 4437 2697 4471
rect 2697 4437 2731 4471
rect 2731 4437 2740 4471
rect 2688 4428 2740 4437
rect 4160 4428 4212 4480
rect 6276 4428 6328 4480
rect 12440 4471 12492 4480
rect 12440 4437 12449 4471
rect 12449 4437 12483 4471
rect 12483 4437 12492 4471
rect 12440 4428 12492 4437
rect 17776 4428 17828 4480
rect 19248 4471 19300 4480
rect 19248 4437 19257 4471
rect 19257 4437 19291 4471
rect 19291 4437 19300 4471
rect 19248 4428 19300 4437
rect 26884 4428 26936 4480
rect 5982 4326 6034 4378
rect 6046 4326 6098 4378
rect 6110 4326 6162 4378
rect 6174 4326 6226 4378
rect 15982 4326 16034 4378
rect 16046 4326 16098 4378
rect 16110 4326 16162 4378
rect 16174 4326 16226 4378
rect 25982 4326 26034 4378
rect 26046 4326 26098 4378
rect 26110 4326 26162 4378
rect 26174 4326 26226 4378
rect 2504 4224 2556 4276
rect 4804 4224 4856 4276
rect 6552 4224 6604 4276
rect 7472 4267 7524 4276
rect 7472 4233 7481 4267
rect 7481 4233 7515 4267
rect 7515 4233 7524 4267
rect 7472 4224 7524 4233
rect 11428 4224 11480 4276
rect 11980 4224 12032 4276
rect 13268 4267 13320 4276
rect 13268 4233 13277 4267
rect 13277 4233 13311 4267
rect 13311 4233 13320 4267
rect 13268 4224 13320 4233
rect 13544 4224 13596 4276
rect 16396 4267 16448 4276
rect 16396 4233 16405 4267
rect 16405 4233 16439 4267
rect 16439 4233 16448 4267
rect 16396 4224 16448 4233
rect 17776 4267 17828 4276
rect 17776 4233 17785 4267
rect 17785 4233 17819 4267
rect 17819 4233 17828 4267
rect 17776 4224 17828 4233
rect 19892 4224 19944 4276
rect 21640 4267 21692 4276
rect 21640 4233 21649 4267
rect 21649 4233 21683 4267
rect 21683 4233 21692 4267
rect 21640 4224 21692 4233
rect 22376 4224 22428 4276
rect 26516 4224 26568 4276
rect 3148 4156 3200 4208
rect 3240 4131 3292 4140
rect 3240 4097 3249 4131
rect 3249 4097 3283 4131
rect 3283 4097 3292 4131
rect 3240 4088 3292 4097
rect 6368 4156 6420 4208
rect 1860 4020 1912 4072
rect 5448 4088 5500 4140
rect 11796 4156 11848 4208
rect 13452 4156 13504 4208
rect 16304 4156 16356 4208
rect 20352 4156 20404 4208
rect 21364 4199 21416 4208
rect 20168 4131 20220 4140
rect 9680 4020 9732 4072
rect 9864 4063 9916 4072
rect 9864 4029 9873 4063
rect 9873 4029 9907 4063
rect 9907 4029 9916 4063
rect 9864 4020 9916 4029
rect 11612 4020 11664 4072
rect 18052 4063 18104 4072
rect 18052 4029 18061 4063
rect 18061 4029 18095 4063
rect 18095 4029 18104 4063
rect 18052 4020 18104 4029
rect 20168 4097 20177 4131
rect 20177 4097 20211 4131
rect 20211 4097 20220 4131
rect 21364 4165 21373 4199
rect 21373 4165 21407 4199
rect 21407 4165 21416 4199
rect 21364 4156 21416 4165
rect 20168 4088 20220 4097
rect 22100 4088 22152 4140
rect 18328 4063 18380 4072
rect 18328 4029 18351 4063
rect 18351 4029 18380 4063
rect 20628 4063 20680 4072
rect 18328 4020 18380 4029
rect 20628 4029 20637 4063
rect 20637 4029 20671 4063
rect 20671 4029 20680 4063
rect 20628 4020 20680 4029
rect 21640 4020 21692 4072
rect 26424 4063 26476 4072
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 2780 3927 2832 3936
rect 2780 3893 2789 3927
rect 2789 3893 2823 3927
rect 2823 3893 2832 3927
rect 3148 3927 3200 3936
rect 2780 3884 2832 3893
rect 3148 3893 3157 3927
rect 3157 3893 3191 3927
rect 3191 3893 3200 3927
rect 3148 3884 3200 3893
rect 4068 3884 4120 3936
rect 4252 3884 4304 3936
rect 4528 3927 4580 3936
rect 4528 3893 4537 3927
rect 4537 3893 4571 3927
rect 4571 3893 4580 3927
rect 4528 3884 4580 3893
rect 6460 3927 6512 3936
rect 6460 3893 6469 3927
rect 6469 3893 6503 3927
rect 6503 3893 6512 3927
rect 6460 3884 6512 3893
rect 9036 3927 9088 3936
rect 9036 3893 9045 3927
rect 9045 3893 9079 3927
rect 9079 3893 9088 3927
rect 26424 4029 26433 4063
rect 26433 4029 26467 4063
rect 26467 4029 26476 4063
rect 26424 4020 26476 4029
rect 9036 3884 9088 3893
rect 20260 3927 20312 3936
rect 20260 3893 20269 3927
rect 20269 3893 20303 3927
rect 20303 3893 20312 3927
rect 20260 3884 20312 3893
rect 20720 3927 20772 3936
rect 20720 3893 20729 3927
rect 20729 3893 20763 3927
rect 20763 3893 20772 3927
rect 21824 3927 21876 3936
rect 20720 3884 20772 3893
rect 21824 3893 21833 3927
rect 21833 3893 21867 3927
rect 21867 3893 21876 3927
rect 21824 3884 21876 3893
rect 26700 3884 26752 3936
rect 27712 3927 27764 3936
rect 27712 3893 27721 3927
rect 27721 3893 27755 3927
rect 27755 3893 27764 3927
rect 27712 3884 27764 3893
rect 10982 3782 11034 3834
rect 11046 3782 11098 3834
rect 11110 3782 11162 3834
rect 11174 3782 11226 3834
rect 20982 3782 21034 3834
rect 21046 3782 21098 3834
rect 21110 3782 21162 3834
rect 21174 3782 21226 3834
rect 1860 3680 1912 3732
rect 2780 3680 2832 3732
rect 3792 3680 3844 3732
rect 5448 3680 5500 3732
rect 9864 3723 9916 3732
rect 9864 3689 9873 3723
rect 9873 3689 9907 3723
rect 9907 3689 9916 3723
rect 9864 3680 9916 3689
rect 11428 3723 11480 3732
rect 11428 3689 11437 3723
rect 11437 3689 11471 3723
rect 11471 3689 11480 3723
rect 11428 3680 11480 3689
rect 19708 3723 19760 3732
rect 19708 3689 19717 3723
rect 19717 3689 19751 3723
rect 19751 3689 19760 3723
rect 19708 3680 19760 3689
rect 20352 3723 20404 3732
rect 20352 3689 20361 3723
rect 20361 3689 20395 3723
rect 20395 3689 20404 3723
rect 20352 3680 20404 3689
rect 21824 3680 21876 3732
rect 22284 3723 22336 3732
rect 22284 3689 22293 3723
rect 22293 3689 22327 3723
rect 22327 3689 22336 3723
rect 22284 3680 22336 3689
rect 3148 3612 3200 3664
rect 6276 3612 6328 3664
rect 20260 3612 20312 3664
rect 21364 3655 21416 3664
rect 21364 3621 21373 3655
rect 21373 3621 21407 3655
rect 21407 3621 21416 3655
rect 21364 3612 21416 3621
rect 1952 3587 2004 3596
rect 1952 3553 1961 3587
rect 1961 3553 1995 3587
rect 1995 3553 2004 3587
rect 1952 3544 2004 3553
rect 4068 3587 4120 3596
rect 4068 3553 4077 3587
rect 4077 3553 4111 3587
rect 4111 3553 4120 3587
rect 4068 3544 4120 3553
rect 4804 3544 4856 3596
rect 6828 3544 6880 3596
rect 15660 3587 15712 3596
rect 15660 3553 15669 3587
rect 15669 3553 15703 3587
rect 15703 3553 15712 3587
rect 15660 3544 15712 3553
rect 17316 3544 17368 3596
rect 23940 3544 23992 3596
rect 27344 3544 27396 3596
rect 5816 3476 5868 3528
rect 6552 3476 6604 3528
rect 7472 3519 7524 3528
rect 7472 3485 7481 3519
rect 7481 3485 7515 3519
rect 7515 3485 7524 3519
rect 7472 3476 7524 3485
rect 16304 3476 16356 3528
rect 17868 3476 17920 3528
rect 18328 3519 18380 3528
rect 18328 3485 18337 3519
rect 18337 3485 18371 3519
rect 18371 3485 18380 3519
rect 18328 3476 18380 3485
rect 19616 3476 19668 3528
rect 20720 3408 20772 3460
rect 21272 3476 21324 3528
rect 2136 3383 2188 3392
rect 2136 3349 2145 3383
rect 2145 3349 2179 3383
rect 2179 3349 2188 3383
rect 2136 3340 2188 3349
rect 4068 3340 4120 3392
rect 5356 3383 5408 3392
rect 5356 3349 5365 3383
rect 5365 3349 5399 3383
rect 5399 3349 5408 3383
rect 5356 3340 5408 3349
rect 26792 3340 26844 3392
rect 5982 3238 6034 3290
rect 6046 3238 6098 3290
rect 6110 3238 6162 3290
rect 6174 3238 6226 3290
rect 15982 3238 16034 3290
rect 16046 3238 16098 3290
rect 16110 3238 16162 3290
rect 16174 3238 16226 3290
rect 25982 3238 26034 3290
rect 26046 3238 26098 3290
rect 26110 3238 26162 3290
rect 26174 3238 26226 3290
rect 1952 3136 2004 3188
rect 4436 3179 4488 3188
rect 4436 3145 4445 3179
rect 4445 3145 4479 3179
rect 4479 3145 4488 3179
rect 4436 3136 4488 3145
rect 4804 3179 4856 3188
rect 4804 3145 4813 3179
rect 4813 3145 4847 3179
rect 4847 3145 4856 3179
rect 4804 3136 4856 3145
rect 5816 3179 5868 3188
rect 5816 3145 5825 3179
rect 5825 3145 5859 3179
rect 5859 3145 5868 3179
rect 5816 3136 5868 3145
rect 6276 3179 6328 3188
rect 6276 3145 6285 3179
rect 6285 3145 6319 3179
rect 6319 3145 6328 3179
rect 6276 3136 6328 3145
rect 7472 3136 7524 3188
rect 13636 3179 13688 3188
rect 13636 3145 13645 3179
rect 13645 3145 13679 3179
rect 13679 3145 13688 3179
rect 13636 3136 13688 3145
rect 3332 3111 3384 3120
rect 3332 3077 3341 3111
rect 3341 3077 3375 3111
rect 3375 3077 3384 3111
rect 3332 3068 3384 3077
rect 3976 3068 4028 3120
rect 3792 3043 3844 3052
rect 3792 3009 3801 3043
rect 3801 3009 3835 3043
rect 3835 3009 3844 3043
rect 3792 3000 3844 3009
rect 6552 3043 6604 3052
rect 1952 2932 2004 2984
rect 3700 2932 3752 2984
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 2044 2864 2096 2916
rect 4620 2932 4672 2984
rect 6736 2932 6788 2984
rect 13636 2932 13688 2984
rect 15476 3136 15528 3188
rect 15660 3179 15712 3188
rect 15660 3145 15669 3179
rect 15669 3145 15703 3179
rect 15703 3145 15712 3179
rect 15660 3136 15712 3145
rect 17316 3179 17368 3188
rect 17316 3145 17325 3179
rect 17325 3145 17359 3179
rect 17359 3145 17368 3179
rect 17316 3136 17368 3145
rect 21364 3179 21416 3188
rect 21364 3145 21373 3179
rect 21373 3145 21407 3179
rect 21407 3145 21416 3179
rect 21364 3136 21416 3145
rect 21824 3136 21876 3188
rect 27344 3179 27396 3188
rect 27344 3145 27353 3179
rect 27353 3145 27387 3179
rect 27387 3145 27396 3179
rect 27344 3136 27396 3145
rect 17868 3068 17920 3120
rect 21272 3068 21324 3120
rect 26332 3068 26384 3120
rect 17960 2932 18012 2984
rect 24952 2932 25004 2984
rect 26424 2975 26476 2984
rect 26424 2941 26433 2975
rect 26433 2941 26467 2975
rect 26467 2941 26476 2975
rect 26424 2932 26476 2941
rect 27528 2975 27580 2984
rect 27528 2941 27537 2975
rect 27537 2941 27571 2975
rect 27571 2941 27580 2975
rect 27528 2932 27580 2941
rect 7748 2864 7800 2916
rect 13452 2864 13504 2916
rect 14924 2864 14976 2916
rect 19156 2864 19208 2916
rect 21732 2864 21784 2916
rect 24032 2864 24084 2916
rect 3792 2796 3844 2848
rect 3884 2796 3936 2848
rect 23848 2839 23900 2848
rect 23848 2805 23857 2839
rect 23857 2805 23891 2839
rect 23891 2805 23900 2839
rect 23848 2796 23900 2805
rect 26608 2839 26660 2848
rect 26608 2805 26617 2839
rect 26617 2805 26651 2839
rect 26651 2805 26660 2839
rect 26608 2796 26660 2805
rect 27712 2839 27764 2848
rect 27712 2805 27721 2839
rect 27721 2805 27755 2839
rect 27755 2805 27764 2839
rect 27712 2796 27764 2805
rect 10982 2694 11034 2746
rect 11046 2694 11098 2746
rect 11110 2694 11162 2746
rect 11174 2694 11226 2746
rect 20982 2694 21034 2746
rect 21046 2694 21098 2746
rect 21110 2694 21162 2746
rect 21174 2694 21226 2746
rect 1952 2592 2004 2644
rect 3516 2592 3568 2644
rect 3884 2592 3936 2644
rect 5448 2635 5500 2644
rect 5448 2601 5457 2635
rect 5457 2601 5491 2635
rect 5491 2601 5500 2635
rect 5448 2592 5500 2601
rect 5356 2456 5408 2508
rect 6460 2592 6512 2644
rect 8208 2592 8260 2644
rect 16856 2635 16908 2644
rect 16856 2601 16865 2635
rect 16865 2601 16899 2635
rect 16899 2601 16908 2635
rect 16856 2592 16908 2601
rect 17776 2635 17828 2644
rect 17776 2601 17785 2635
rect 17785 2601 17819 2635
rect 17819 2601 17828 2635
rect 17776 2592 17828 2601
rect 22560 2635 22612 2644
rect 22560 2601 22569 2635
rect 22569 2601 22603 2635
rect 22603 2601 22612 2635
rect 22560 2592 22612 2601
rect 8116 2456 8168 2508
rect 9772 2499 9824 2508
rect 9772 2465 9781 2499
rect 9781 2465 9815 2499
rect 9815 2465 9824 2499
rect 9772 2456 9824 2465
rect 12716 2456 12768 2508
rect 18236 2456 18288 2508
rect 24032 2499 24084 2508
rect 24032 2465 24041 2499
rect 24041 2465 24075 2499
rect 24075 2465 24084 2499
rect 24032 2456 24084 2465
rect 25688 2499 25740 2508
rect 25688 2465 25697 2499
rect 25697 2465 25731 2499
rect 25731 2465 25740 2499
rect 25688 2456 25740 2465
rect 3516 2388 3568 2440
rect 4896 2388 4948 2440
rect 6368 2388 6420 2440
rect 9220 2388 9272 2440
rect 10600 2388 10652 2440
rect 12072 2388 12124 2440
rect 17776 2388 17828 2440
rect 20628 2388 20680 2440
rect 22008 2388 22060 2440
rect 23480 2388 23532 2440
rect 5816 2295 5868 2304
rect 5816 2261 5825 2295
rect 5825 2261 5859 2295
rect 5859 2261 5868 2295
rect 5816 2252 5868 2261
rect 25872 2295 25924 2304
rect 25872 2261 25881 2295
rect 25881 2261 25915 2295
rect 25915 2261 25924 2295
rect 25872 2252 25924 2261
rect 29184 2252 29236 2304
rect 5982 2150 6034 2202
rect 6046 2150 6098 2202
rect 6110 2150 6162 2202
rect 6174 2150 6226 2202
rect 15982 2150 16034 2202
rect 16046 2150 16098 2202
rect 16110 2150 16162 2202
rect 16174 2150 16226 2202
rect 25982 2150 26034 2202
rect 26046 2150 26098 2202
rect 26110 2150 26162 2202
rect 26174 2150 26226 2202
<< metal2 >>
rect 1674 23520 1730 24000
rect 3974 23624 4030 23633
rect 3974 23559 4030 23568
rect 1688 19854 1716 23520
rect 2870 22400 2926 22409
rect 2870 22335 2926 22344
rect 1676 19848 1728 19854
rect 1676 19790 1728 19796
rect 2688 19848 2740 19854
rect 2688 19790 2740 19796
rect 2228 18216 2280 18222
rect 2280 18164 2360 18170
rect 2228 18158 2360 18164
rect 2240 18142 2360 18158
rect 2042 18048 2098 18057
rect 2042 17983 2098 17992
rect 1398 17776 1454 17785
rect 1398 17711 1400 17720
rect 1452 17711 1454 17720
rect 1400 17682 1452 17688
rect 1412 17626 1440 17682
rect 1412 17598 1532 17626
rect 1400 17536 1452 17542
rect 1400 17478 1452 17484
rect 1412 11121 1440 17478
rect 1504 16794 1532 17598
rect 2056 17338 2084 17983
rect 2332 17542 2360 18142
rect 2320 17536 2372 17542
rect 2320 17478 2372 17484
rect 2044 17332 2096 17338
rect 2044 17274 2096 17280
rect 2056 17134 2084 17274
rect 2044 17128 2096 17134
rect 2044 17070 2096 17076
rect 1492 16788 1544 16794
rect 1492 16730 1544 16736
rect 2332 16454 2360 17478
rect 2320 16448 2372 16454
rect 2320 16390 2372 16396
rect 2332 15978 2360 16390
rect 2700 15978 2728 19790
rect 2780 18148 2832 18154
rect 2780 18090 2832 18096
rect 2792 17814 2820 18090
rect 2780 17808 2832 17814
rect 2780 17750 2832 17756
rect 1676 15972 1728 15978
rect 1676 15914 1728 15920
rect 2320 15972 2372 15978
rect 2320 15914 2372 15920
rect 2688 15972 2740 15978
rect 2688 15914 2740 15920
rect 1688 15434 1716 15914
rect 1860 15496 1912 15502
rect 1860 15438 1912 15444
rect 1676 15428 1728 15434
rect 1676 15370 1728 15376
rect 1676 14816 1728 14822
rect 1676 14758 1728 14764
rect 1768 14816 1820 14822
rect 1768 14758 1820 14764
rect 1688 13938 1716 14758
rect 1780 14618 1808 14758
rect 1872 14618 1900 15438
rect 2332 15366 2360 15914
rect 2778 15872 2834 15881
rect 2778 15807 2834 15816
rect 2320 15360 2372 15366
rect 2320 15302 2372 15308
rect 2332 15026 2360 15302
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2504 14884 2556 14890
rect 2504 14826 2556 14832
rect 1768 14612 1820 14618
rect 1768 14554 1820 14560
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 1780 14006 1808 14554
rect 2516 14414 2544 14826
rect 2596 14544 2648 14550
rect 2596 14486 2648 14492
rect 2504 14408 2556 14414
rect 2504 14350 2556 14356
rect 1952 14272 2004 14278
rect 1952 14214 2004 14220
rect 1768 14000 1820 14006
rect 1768 13942 1820 13948
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1584 13728 1636 13734
rect 1584 13670 1636 13676
rect 1596 12782 1624 13670
rect 1688 13530 1716 13874
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1584 12776 1636 12782
rect 1584 12718 1636 12724
rect 1780 12374 1808 13942
rect 1964 13734 1992 14214
rect 2516 13870 2544 14350
rect 2608 14074 2636 14486
rect 2596 14068 2648 14074
rect 2596 14010 2648 14016
rect 2504 13864 2556 13870
rect 2504 13806 2556 13812
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1964 13530 1992 13670
rect 1952 13524 2004 13530
rect 1952 13466 2004 13472
rect 2228 13388 2280 13394
rect 2228 13330 2280 13336
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 1952 12640 2004 12646
rect 1952 12582 2004 12588
rect 1768 12368 1820 12374
rect 1768 12310 1820 12316
rect 1490 12200 1546 12209
rect 1490 12135 1546 12144
rect 1504 11218 1532 12135
rect 1780 11898 1808 12310
rect 1768 11892 1820 11898
rect 1768 11834 1820 11840
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1492 11212 1544 11218
rect 1492 11154 1544 11160
rect 1398 11112 1454 11121
rect 1398 11047 1454 11056
rect 1504 10810 1532 11154
rect 1492 10804 1544 10810
rect 1492 10746 1544 10752
rect 1596 10441 1624 11494
rect 1768 11076 1820 11082
rect 1768 11018 1820 11024
rect 1582 10432 1638 10441
rect 1582 10367 1638 10376
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1584 9920 1636 9926
rect 1584 9862 1636 9868
rect 1400 9376 1452 9382
rect 1596 9353 1624 9862
rect 1688 9489 1716 10066
rect 1674 9480 1730 9489
rect 1674 9415 1730 9424
rect 1400 9318 1452 9324
rect 1582 9344 1638 9353
rect 1412 8129 1440 9318
rect 1582 9279 1638 9288
rect 1688 9178 1716 9415
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 1490 8664 1546 8673
rect 1490 8599 1546 8608
rect 1398 8120 1454 8129
rect 1398 8055 1454 8064
rect 1504 6458 1532 8599
rect 1584 8560 1636 8566
rect 1584 8502 1636 8508
rect 1596 7449 1624 8502
rect 1582 7440 1638 7449
rect 1582 7375 1638 7384
rect 1676 7268 1728 7274
rect 1676 7210 1728 7216
rect 1688 7002 1716 7210
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1492 6452 1544 6458
rect 1492 6394 1544 6400
rect 1688 6390 1716 6938
rect 1780 6905 1808 11018
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1872 7274 1900 7686
rect 1860 7268 1912 7274
rect 1860 7210 1912 7216
rect 1766 6896 1822 6905
rect 1766 6831 1822 6840
rect 1676 6384 1728 6390
rect 1676 6326 1728 6332
rect 1768 5704 1820 5710
rect 1582 5672 1638 5681
rect 1872 5692 1900 7210
rect 1820 5664 1900 5692
rect 1768 5646 1820 5652
rect 1582 5607 1638 5616
rect 1596 5370 1624 5607
rect 1584 5364 1636 5370
rect 1584 5306 1636 5312
rect 1582 5128 1638 5137
rect 1582 5063 1638 5072
rect 1596 4826 1624 5063
rect 1584 4820 1636 4826
rect 1584 4762 1636 4768
rect 1780 4758 1808 5646
rect 1858 5128 1914 5137
rect 1858 5063 1914 5072
rect 1768 4752 1820 4758
rect 1768 4694 1820 4700
rect 1582 4448 1638 4457
rect 1582 4383 1638 4392
rect 1596 3942 1624 4383
rect 1872 4078 1900 5063
rect 1964 4434 1992 12582
rect 2056 11354 2084 12786
rect 2240 12714 2268 13330
rect 2516 13326 2544 13806
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2608 12968 2636 14010
rect 2516 12940 2636 12968
rect 2228 12708 2280 12714
rect 2228 12650 2280 12656
rect 2228 12300 2280 12306
rect 2228 12242 2280 12248
rect 2240 11354 2268 12242
rect 2516 11830 2544 12940
rect 2596 12776 2648 12782
rect 2792 12730 2820 15807
rect 2884 13954 2912 22335
rect 3988 22234 4016 23559
rect 4986 23520 5042 24000
rect 8298 23520 8354 24000
rect 11610 23520 11666 24000
rect 14922 23520 14978 24000
rect 18326 23520 18382 24000
rect 21638 23520 21694 24000
rect 24950 23520 25006 24000
rect 25870 23624 25926 23633
rect 25870 23559 25926 23568
rect 4250 23080 4306 23089
rect 4250 23015 4306 23024
rect 3976 22228 4028 22234
rect 3976 22170 4028 22176
rect 4066 21856 4122 21865
rect 4066 21791 4122 21800
rect 4080 20874 4108 21791
rect 4068 20868 4120 20874
rect 4068 20810 4120 20816
rect 3238 20632 3294 20641
rect 3238 20567 3294 20576
rect 3252 17252 3280 20567
rect 3330 20088 3386 20097
rect 3330 20023 3386 20032
rect 3344 17354 3372 20023
rect 4264 18834 4292 23015
rect 5000 20369 5028 23520
rect 5956 21788 6252 21808
rect 6012 21786 6036 21788
rect 6092 21786 6116 21788
rect 6172 21786 6196 21788
rect 6034 21734 6036 21786
rect 6098 21734 6110 21786
rect 6172 21734 6174 21786
rect 6012 21732 6036 21734
rect 6092 21732 6116 21734
rect 6172 21732 6196 21734
rect 5956 21712 6252 21732
rect 7286 21312 7342 21321
rect 7286 21247 7342 21256
rect 5956 20700 6252 20720
rect 6012 20698 6036 20700
rect 6092 20698 6116 20700
rect 6172 20698 6196 20700
rect 6034 20646 6036 20698
rect 6098 20646 6110 20698
rect 6172 20646 6174 20698
rect 6012 20644 6036 20646
rect 6092 20644 6116 20646
rect 6172 20644 6196 20646
rect 5956 20624 6252 20644
rect 4986 20360 5042 20369
rect 4986 20295 5042 20304
rect 5724 19916 5776 19922
rect 5724 19858 5776 19864
rect 5632 19848 5684 19854
rect 5632 19790 5684 19796
rect 5644 19174 5672 19790
rect 5736 19514 5764 19858
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 5956 19612 6252 19632
rect 6012 19610 6036 19612
rect 6092 19610 6116 19612
rect 6172 19610 6196 19612
rect 6034 19558 6036 19610
rect 6098 19558 6110 19610
rect 6172 19558 6174 19610
rect 6012 19556 6036 19558
rect 6092 19556 6116 19558
rect 6172 19556 6196 19558
rect 5956 19536 6252 19556
rect 5724 19508 5776 19514
rect 5724 19450 5776 19456
rect 5736 19242 5764 19450
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 5724 19236 5776 19242
rect 5724 19178 5776 19184
rect 5632 19168 5684 19174
rect 5354 19136 5410 19145
rect 6840 19156 6868 19246
rect 6920 19168 6972 19174
rect 6840 19128 6920 19156
rect 5632 19110 5684 19116
rect 6920 19110 6972 19116
rect 5354 19071 5410 19080
rect 4986 18864 5042 18873
rect 4252 18828 4304 18834
rect 4986 18799 5042 18808
rect 4252 18770 4304 18776
rect 4160 18624 4212 18630
rect 4160 18566 4212 18572
rect 3976 18284 4028 18290
rect 3976 18226 4028 18232
rect 3516 18080 3568 18086
rect 3516 18022 3568 18028
rect 3528 17678 3556 18022
rect 3988 17814 4016 18226
rect 4068 18216 4120 18222
rect 4068 18158 4120 18164
rect 4080 17882 4108 18158
rect 4172 17882 4200 18566
rect 4264 18193 4292 18770
rect 4528 18760 4580 18766
rect 4528 18702 4580 18708
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 4540 18426 4568 18702
rect 4528 18420 4580 18426
rect 4528 18362 4580 18368
rect 4250 18184 4306 18193
rect 4250 18119 4252 18128
rect 4304 18119 4306 18128
rect 4252 18090 4304 18096
rect 4436 18080 4488 18086
rect 4540 18057 4568 18362
rect 4710 18320 4766 18329
rect 4816 18290 4844 18702
rect 4710 18255 4766 18264
rect 4804 18284 4856 18290
rect 4724 18057 4752 18255
rect 4804 18226 4856 18232
rect 4436 18022 4488 18028
rect 4526 18048 4582 18057
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 4160 17876 4212 17882
rect 4160 17818 4212 17824
rect 3976 17808 4028 17814
rect 3976 17750 4028 17756
rect 3516 17672 3568 17678
rect 3422 17640 3478 17649
rect 3516 17614 3568 17620
rect 3422 17575 3478 17584
rect 3436 17524 3464 17575
rect 3436 17496 3556 17524
rect 3344 17326 3464 17354
rect 3252 17224 3372 17252
rect 3146 17096 3202 17105
rect 3146 17031 3202 17040
rect 3160 15473 3188 17031
rect 3240 16992 3292 16998
rect 3240 16934 3292 16940
rect 3252 16833 3280 16934
rect 3238 16824 3294 16833
rect 3238 16759 3294 16768
rect 3146 15464 3202 15473
rect 3146 15399 3202 15408
rect 3238 14920 3294 14929
rect 3238 14855 3294 14864
rect 2964 14612 3016 14618
rect 2964 14554 3016 14560
rect 2976 14074 3004 14554
rect 3252 14550 3280 14855
rect 3240 14544 3292 14550
rect 3240 14486 3292 14492
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 2884 13926 3004 13954
rect 2872 13388 2924 13394
rect 2872 13330 2924 13336
rect 2596 12718 2648 12724
rect 2608 11898 2636 12718
rect 2700 12702 2820 12730
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2504 11824 2556 11830
rect 2504 11766 2556 11772
rect 2700 11778 2728 12702
rect 2884 12646 2912 13330
rect 2976 12714 3004 13926
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 2964 12708 3016 12714
rect 2964 12650 3016 12656
rect 2872 12640 2924 12646
rect 2872 12582 2924 12588
rect 2884 12209 2912 12582
rect 2870 12200 2926 12209
rect 2870 12135 2926 12144
rect 2976 11801 3004 12650
rect 3068 12102 3096 12786
rect 3238 12608 3294 12617
rect 3238 12543 3294 12552
rect 3056 12096 3108 12102
rect 3056 12038 3108 12044
rect 2962 11792 3018 11801
rect 2700 11750 2820 11778
rect 2686 11656 2742 11665
rect 2686 11591 2742 11600
rect 2700 11354 2728 11591
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2240 10674 2268 11290
rect 2686 11248 2742 11257
rect 2686 11183 2688 11192
rect 2740 11183 2742 11192
rect 2688 11154 2740 11160
rect 2700 10810 2728 11154
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 2240 10198 2268 10610
rect 2502 10296 2558 10305
rect 2502 10231 2558 10240
rect 2228 10192 2280 10198
rect 2228 10134 2280 10140
rect 2516 10130 2544 10231
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2516 9722 2544 10066
rect 2688 9920 2740 9926
rect 2686 9888 2688 9897
rect 2740 9888 2742 9897
rect 2686 9823 2742 9832
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 2042 9616 2098 9625
rect 2042 9551 2044 9560
rect 2096 9551 2098 9560
rect 2044 9522 2096 9528
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2516 8634 2544 9046
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2424 7002 2452 7686
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2502 6896 2558 6905
rect 2502 6831 2558 6840
rect 2042 6488 2098 6497
rect 2042 6423 2044 6432
rect 2096 6423 2098 6432
rect 2044 6394 2096 6400
rect 2056 6254 2084 6394
rect 2044 6248 2096 6254
rect 2044 6190 2096 6196
rect 2320 5840 2372 5846
rect 2320 5782 2372 5788
rect 2332 5370 2360 5782
rect 2320 5364 2372 5370
rect 2320 5306 2372 5312
rect 2042 5264 2098 5273
rect 2042 5199 2044 5208
rect 2096 5199 2098 5208
rect 2044 5170 2096 5176
rect 2042 4720 2098 4729
rect 2516 4690 2544 6831
rect 2608 6662 2636 8774
rect 2792 8022 2820 11750
rect 2962 11727 3018 11736
rect 3068 10538 3096 12038
rect 3252 11898 3280 12543
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3056 10532 3108 10538
rect 3056 10474 3108 10480
rect 3068 10266 3096 10474
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2884 8634 2912 8910
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2870 8528 2926 8537
rect 2870 8463 2872 8472
rect 2924 8463 2926 8472
rect 2872 8434 2924 8440
rect 2780 8016 2832 8022
rect 2778 7984 2780 7993
rect 2832 7984 2834 7993
rect 2778 7919 2834 7928
rect 2792 7546 2820 7919
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2884 7206 2912 7346
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2780 6996 2832 7002
rect 2780 6938 2832 6944
rect 2596 6656 2648 6662
rect 2596 6598 2648 6604
rect 2608 6458 2636 6598
rect 2792 6458 2820 6938
rect 2884 6662 2912 7142
rect 2962 7032 3018 7041
rect 2962 6967 3018 6976
rect 2976 6798 3004 6967
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2884 5846 2912 6598
rect 2976 6390 3004 6734
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 2872 5840 2924 5846
rect 2872 5782 2924 5788
rect 3148 5568 3200 5574
rect 3148 5510 3200 5516
rect 3160 5370 3188 5510
rect 3148 5364 3200 5370
rect 3148 5306 3200 5312
rect 3160 5098 3188 5306
rect 3148 5092 3200 5098
rect 3148 5034 3200 5040
rect 3160 4826 3188 5034
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 2042 4655 2044 4664
rect 2096 4655 2098 4664
rect 2504 4684 2556 4690
rect 2044 4626 2096 4632
rect 2504 4626 2556 4632
rect 1964 4406 2084 4434
rect 1950 4176 2006 4185
rect 1950 4111 2006 4120
rect 1860 4072 1912 4078
rect 1860 4014 1912 4020
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1872 3738 1900 4014
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 1964 3602 1992 4111
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 1964 3194 1992 3538
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 2056 3074 2084 4406
rect 2516 4282 2544 4626
rect 2688 4480 2740 4486
rect 2688 4422 2740 4428
rect 2504 4276 2556 4282
rect 2504 4218 2556 4224
rect 2700 3913 2728 4422
rect 3160 4214 3188 4762
rect 3148 4208 3200 4214
rect 3148 4150 3200 4156
rect 3252 4146 3280 11834
rect 3344 7585 3372 17224
rect 3436 11665 3464 17326
rect 3422 11656 3478 11665
rect 3422 11591 3478 11600
rect 3528 10713 3556 17496
rect 3792 17264 3844 17270
rect 3792 17206 3844 17212
rect 3700 16992 3752 16998
rect 3700 16934 3752 16940
rect 3712 16794 3740 16934
rect 3700 16788 3752 16794
rect 3700 16730 3752 16736
rect 3712 16538 3740 16730
rect 3620 16510 3740 16538
rect 3620 16250 3648 16510
rect 3700 16448 3752 16454
rect 3700 16390 3752 16396
rect 3608 16244 3660 16250
rect 3608 16186 3660 16192
rect 3712 16114 3740 16390
rect 3700 16108 3752 16114
rect 3700 16050 3752 16056
rect 3606 16008 3662 16017
rect 3606 15943 3662 15952
rect 3620 15910 3648 15943
rect 3608 15904 3660 15910
rect 3608 15846 3660 15852
rect 3620 13433 3648 15846
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3606 13424 3662 13433
rect 3606 13359 3662 13368
rect 3514 10704 3570 10713
rect 3514 10639 3570 10648
rect 3516 10192 3568 10198
rect 3516 10134 3568 10140
rect 3528 9586 3556 10134
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3620 9110 3648 13359
rect 3712 12850 3740 14758
rect 3700 12844 3752 12850
rect 3700 12786 3752 12792
rect 3712 12374 3740 12786
rect 3700 12368 3752 12374
rect 3700 12310 3752 12316
rect 3804 12220 3832 17206
rect 3988 16522 4016 17750
rect 4448 17746 4476 18022
rect 4526 17983 4582 17992
rect 4710 18048 4766 18057
rect 4710 17983 4766 17992
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 4436 17740 4488 17746
rect 4436 17682 4488 17688
rect 4344 17672 4396 17678
rect 4344 17614 4396 17620
rect 4068 17536 4120 17542
rect 4068 17478 4120 17484
rect 4080 17241 4108 17478
rect 4356 17338 4384 17614
rect 4448 17338 4476 17682
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4436 17332 4488 17338
rect 4436 17274 4488 17280
rect 4632 17270 4660 17818
rect 4620 17264 4672 17270
rect 4066 17232 4122 17241
rect 4620 17206 4672 17212
rect 4066 17167 4122 17176
rect 4068 17060 4120 17066
rect 4068 17002 4120 17008
rect 4080 16794 4108 17002
rect 4724 16794 4752 17983
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4526 16552 4582 16561
rect 3976 16516 4028 16522
rect 4526 16487 4582 16496
rect 3976 16458 4028 16464
rect 3882 16416 3938 16425
rect 3882 16351 3938 16360
rect 3896 13705 3924 16351
rect 3988 16182 4016 16458
rect 3976 16176 4028 16182
rect 3976 16118 4028 16124
rect 3988 15638 4016 16118
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 4080 15706 4108 16050
rect 4434 15736 4490 15745
rect 4068 15700 4120 15706
rect 4540 15706 4568 16487
rect 4724 16250 4752 16730
rect 4712 16244 4764 16250
rect 4712 16186 4764 16192
rect 4434 15671 4436 15680
rect 4068 15642 4120 15648
rect 4488 15671 4490 15680
rect 4528 15700 4580 15706
rect 4436 15642 4488 15648
rect 4528 15642 4580 15648
rect 3976 15632 4028 15638
rect 3976 15574 4028 15580
rect 4448 15162 4476 15642
rect 4160 15156 4212 15162
rect 4160 15098 4212 15104
rect 4436 15156 4488 15162
rect 4436 15098 4488 15104
rect 4068 14000 4120 14006
rect 4068 13942 4120 13948
rect 3882 13696 3938 13705
rect 3882 13631 3938 13640
rect 4080 13530 4108 13942
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 3896 12442 3924 12718
rect 4080 12646 4108 13466
rect 4068 12640 4120 12646
rect 3974 12608 4030 12617
rect 4068 12582 4120 12588
rect 3974 12543 4030 12552
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 3988 12345 4016 12543
rect 3974 12336 4030 12345
rect 3974 12271 4030 12280
rect 3712 12192 3832 12220
rect 3608 9104 3660 9110
rect 3608 9046 3660 9052
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3528 8090 3556 8366
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 3330 7576 3386 7585
rect 3330 7511 3386 7520
rect 3436 7206 3464 7890
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3436 4185 3464 7142
rect 3422 4176 3478 4185
rect 3240 4140 3292 4146
rect 3422 4111 3478 4120
rect 3240 4082 3292 4088
rect 2780 3936 2832 3942
rect 2686 3904 2742 3913
rect 2780 3878 2832 3884
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 2686 3839 2742 3848
rect 2792 3738 2820 3878
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 3160 3670 3188 3878
rect 3148 3664 3200 3670
rect 3148 3606 3200 3612
rect 2136 3392 2188 3398
rect 2136 3334 2188 3340
rect 1964 3046 2084 3074
rect 1964 2990 1992 3046
rect 1952 2984 2004 2990
rect 662 2952 718 2961
rect 1952 2926 2004 2932
rect 662 2887 718 2896
rect 676 480 704 2887
rect 1964 2650 1992 2926
rect 2044 2916 2096 2922
rect 2044 2858 2096 2864
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 2056 480 2084 2858
rect 2148 1465 2176 3334
rect 3332 3120 3384 3126
rect 3330 3088 3332 3097
rect 3384 3088 3386 3097
rect 3330 3023 3386 3032
rect 3528 2650 3556 7142
rect 3712 6361 3740 12192
rect 3884 10532 3936 10538
rect 3884 10474 3936 10480
rect 3792 10464 3844 10470
rect 3792 10406 3844 10412
rect 3804 9518 3832 10406
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3804 9178 3832 9454
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 3804 8498 3832 9114
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 3698 6352 3754 6361
rect 3698 6287 3754 6296
rect 3608 5160 3660 5166
rect 3608 5102 3660 5108
rect 3620 4826 3648 5102
rect 3700 5024 3752 5030
rect 3700 4966 3752 4972
rect 3608 4820 3660 4826
rect 3608 4762 3660 4768
rect 3712 2990 3740 4966
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3804 3058 3832 3674
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 3700 2984 3752 2990
rect 3896 2938 3924 10474
rect 3988 8566 4016 12271
rect 3976 8560 4028 8566
rect 4172 8514 4200 15098
rect 4540 15026 4568 15642
rect 4896 15428 4948 15434
rect 4896 15370 4948 15376
rect 4908 15162 4936 15370
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 4344 15020 4396 15026
rect 4344 14962 4396 14968
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 4356 12617 4384 14962
rect 4802 14104 4858 14113
rect 4802 14039 4858 14048
rect 4816 13734 4844 14039
rect 5000 13954 5028 18799
rect 5080 18624 5132 18630
rect 5080 18566 5132 18572
rect 5092 18222 5120 18566
rect 5368 18426 5396 19071
rect 6932 18630 6960 19110
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 5956 18524 6252 18544
rect 6012 18522 6036 18524
rect 6092 18522 6116 18524
rect 6172 18522 6196 18524
rect 6034 18470 6036 18522
rect 6098 18470 6110 18522
rect 6172 18470 6174 18522
rect 6012 18468 6036 18470
rect 6092 18468 6116 18470
rect 6172 18468 6196 18470
rect 5956 18448 6252 18468
rect 5356 18420 5408 18426
rect 5356 18362 5408 18368
rect 5080 18216 5132 18222
rect 5080 18158 5132 18164
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 5184 17678 5212 18022
rect 6368 17740 6420 17746
rect 6368 17682 6420 17688
rect 5172 17672 5224 17678
rect 5170 17640 5172 17649
rect 5724 17672 5776 17678
rect 5224 17640 5226 17649
rect 5724 17614 5776 17620
rect 5170 17575 5226 17584
rect 5736 16998 5764 17614
rect 5956 17436 6252 17456
rect 6012 17434 6036 17436
rect 6092 17434 6116 17436
rect 6172 17434 6196 17436
rect 6034 17382 6036 17434
rect 6098 17382 6110 17434
rect 6172 17382 6174 17434
rect 6012 17380 6036 17382
rect 6092 17380 6116 17382
rect 6172 17380 6196 17382
rect 5956 17360 6252 17380
rect 6380 17338 6408 17682
rect 6368 17332 6420 17338
rect 6368 17274 6420 17280
rect 5814 17232 5870 17241
rect 5814 17167 5870 17176
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 5078 16688 5134 16697
rect 5078 16623 5080 16632
rect 5132 16623 5134 16632
rect 5080 16594 5132 16600
rect 5092 16250 5120 16594
rect 5080 16244 5132 16250
rect 5080 16186 5132 16192
rect 5736 15502 5764 16934
rect 5828 16726 5856 17167
rect 7012 16992 7064 16998
rect 7012 16934 7064 16940
rect 6826 16824 6882 16833
rect 6826 16759 6828 16768
rect 6880 16759 6882 16768
rect 6828 16730 6880 16736
rect 5816 16720 5868 16726
rect 5816 16662 5868 16668
rect 6840 16674 6868 16730
rect 5828 16250 5856 16662
rect 6840 16646 6960 16674
rect 7024 16658 7052 16934
rect 6460 16516 6512 16522
rect 6460 16458 6512 16464
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 5956 16348 6252 16368
rect 6012 16346 6036 16348
rect 6092 16346 6116 16348
rect 6172 16346 6196 16348
rect 6034 16294 6036 16346
rect 6098 16294 6110 16346
rect 6172 16294 6174 16346
rect 6012 16292 6036 16294
rect 6092 16292 6116 16294
rect 6172 16292 6196 16294
rect 5956 16272 6252 16292
rect 5816 16244 5868 16250
rect 5816 16186 5868 16192
rect 5816 15564 5868 15570
rect 5816 15506 5868 15512
rect 5724 15496 5776 15502
rect 5724 15438 5776 15444
rect 5736 15366 5764 15438
rect 5724 15360 5776 15366
rect 5538 15328 5594 15337
rect 5724 15302 5776 15308
rect 5538 15263 5594 15272
rect 5080 14272 5132 14278
rect 5080 14214 5132 14220
rect 4908 13926 5028 13954
rect 5092 13938 5120 14214
rect 5080 13932 5132 13938
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 4540 12782 4568 13126
rect 4816 12918 4844 13670
rect 4908 13462 4936 13926
rect 5080 13874 5132 13880
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 4896 13456 4948 13462
rect 4896 13398 4948 13404
rect 4908 12986 4936 13398
rect 5000 13326 5028 13806
rect 5172 13796 5224 13802
rect 5172 13738 5224 13744
rect 4988 13320 5040 13326
rect 4988 13262 5040 13268
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 4804 12912 4856 12918
rect 4804 12854 4856 12860
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 4342 12608 4398 12617
rect 4342 12543 4398 12552
rect 4816 10538 4844 12854
rect 4908 12617 4936 12922
rect 4894 12608 4950 12617
rect 4894 12543 4950 12552
rect 5000 12442 5028 13262
rect 5184 12986 5212 13738
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5264 12640 5316 12646
rect 5264 12582 5316 12588
rect 4988 12436 5040 12442
rect 4988 12378 5040 12384
rect 5276 12102 5304 12582
rect 5368 12458 5396 13874
rect 5552 13326 5580 15263
rect 5736 15162 5764 15302
rect 5828 15162 5856 15506
rect 5956 15260 6252 15280
rect 6012 15258 6036 15260
rect 6092 15258 6116 15260
rect 6172 15258 6196 15260
rect 6034 15206 6036 15258
rect 6098 15206 6110 15258
rect 6172 15206 6174 15258
rect 6012 15204 6036 15206
rect 6092 15204 6116 15206
rect 6172 15204 6196 15206
rect 5956 15184 6252 15204
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5816 15156 5868 15162
rect 5816 15098 5868 15104
rect 5632 14476 5684 14482
rect 5736 14464 5764 15098
rect 5816 14544 5868 14550
rect 5816 14486 5868 14492
rect 5684 14436 5764 14464
rect 5632 14418 5684 14424
rect 5736 14006 5764 14436
rect 5828 14074 5856 14486
rect 5956 14172 6252 14192
rect 6012 14170 6036 14172
rect 6092 14170 6116 14172
rect 6172 14170 6196 14172
rect 6034 14118 6036 14170
rect 6098 14118 6110 14170
rect 6172 14118 6174 14170
rect 6012 14116 6036 14118
rect 6092 14116 6116 14118
rect 6172 14116 6196 14118
rect 5956 14096 6252 14116
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5724 14000 5776 14006
rect 5724 13942 5776 13948
rect 5724 13728 5776 13734
rect 5724 13670 5776 13676
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5368 12442 5580 12458
rect 5368 12436 5592 12442
rect 5368 12430 5540 12436
rect 5540 12378 5592 12384
rect 5552 12347 5580 12378
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 5448 12096 5500 12102
rect 5500 12044 5580 12050
rect 5448 12038 5580 12044
rect 5460 12022 5580 12038
rect 5552 11393 5580 12022
rect 5644 11898 5672 12242
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5538 11384 5594 11393
rect 5538 11319 5594 11328
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 5184 10742 5212 11086
rect 5276 10810 5304 11154
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5172 10736 5224 10742
rect 5172 10678 5224 10684
rect 4804 10532 4856 10538
rect 4804 10474 4856 10480
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4264 8974 4292 9318
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 3976 8502 4028 8508
rect 4080 8486 4200 8514
rect 4080 8430 4108 8486
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 4264 8294 4292 8910
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4344 8560 4396 8566
rect 4344 8502 4396 8508
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4264 7886 4292 8230
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3988 7154 4016 7686
rect 4264 7410 4292 7822
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 4068 7336 4120 7342
rect 4356 7290 4384 8502
rect 4908 8430 4936 8774
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4120 7284 4384 7290
rect 4068 7278 4384 7284
rect 4080 7262 4384 7278
rect 4068 7200 4120 7206
rect 3988 7148 4068 7154
rect 3988 7142 4120 7148
rect 3988 7126 4108 7142
rect 4080 6934 4108 7126
rect 4068 6928 4120 6934
rect 4068 6870 4120 6876
rect 4356 6866 4384 7262
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 4080 3942 4108 4626
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 4066 3632 4122 3641
rect 4066 3567 4068 3576
rect 4120 3567 4122 3576
rect 4068 3538 4120 3544
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 3976 3120 4028 3126
rect 3976 3062 4028 3068
rect 3700 2926 3752 2932
rect 3804 2910 3924 2938
rect 3804 2854 3832 2910
rect 3792 2848 3844 2854
rect 3792 2790 3844 2796
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3896 2650 3924 2790
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 2134 1456 2190 1465
rect 2134 1391 2190 1400
rect 3528 480 3556 2382
rect 662 0 718 480
rect 2042 0 2098 480
rect 3514 0 3570 480
rect 3988 377 4016 3062
rect 4080 2689 4108 3334
rect 4066 2680 4122 2689
rect 4066 2615 4122 2624
rect 4172 2530 4200 4422
rect 4540 4026 4568 8366
rect 4620 8356 4672 8362
rect 4620 8298 4672 8304
rect 4632 7041 4660 8298
rect 4618 7032 4674 7041
rect 4618 6967 4674 6976
rect 4908 6730 4936 8366
rect 5184 7954 5212 10678
rect 5276 9994 5304 10746
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 5552 9382 5580 11319
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5276 8090 5304 8230
rect 5460 8106 5488 8434
rect 5460 8090 5580 8106
rect 5264 8084 5316 8090
rect 5460 8084 5592 8090
rect 5460 8078 5540 8084
rect 5264 8026 5316 8032
rect 5540 8026 5592 8032
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 4986 7576 5042 7585
rect 4986 7511 4988 7520
rect 5040 7511 5042 7520
rect 4988 7482 5040 7488
rect 5000 7206 5028 7482
rect 5184 7342 5212 7890
rect 5276 7546 5304 8026
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5644 7426 5672 10610
rect 5552 7398 5672 7426
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 4896 6724 4948 6730
rect 4896 6666 4948 6672
rect 5184 5846 5212 7278
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5460 6497 5488 6802
rect 5446 6488 5502 6497
rect 5446 6423 5448 6432
rect 5500 6423 5502 6432
rect 5448 6394 5500 6400
rect 5460 6363 5488 6394
rect 4804 5840 4856 5846
rect 4804 5782 4856 5788
rect 5172 5840 5224 5846
rect 5172 5782 5224 5788
rect 4816 5030 4844 5782
rect 5184 5370 5212 5782
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4816 4282 4844 4966
rect 5184 4826 5212 5306
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 5552 4162 5580 7398
rect 5630 7304 5686 7313
rect 5630 7239 5632 7248
rect 5684 7239 5686 7248
rect 5632 7210 5684 7216
rect 5644 6934 5672 7210
rect 5632 6928 5684 6934
rect 5630 6896 5632 6905
rect 5684 6896 5686 6905
rect 5630 6831 5686 6840
rect 5736 4758 5764 13670
rect 5828 13462 5856 14010
rect 6380 13734 6408 16390
rect 6472 16250 6500 16458
rect 6932 16250 6960 16646
rect 7012 16652 7064 16658
rect 7012 16594 7064 16600
rect 6460 16244 6512 16250
rect 6460 16186 6512 16192
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 6552 15564 6604 15570
rect 6552 15506 6604 15512
rect 6564 14890 6592 15506
rect 6552 14884 6604 14890
rect 6552 14826 6604 14832
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 5816 13456 5868 13462
rect 5816 13398 5868 13404
rect 5828 12850 5856 13398
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 5956 13084 6252 13104
rect 6012 13082 6036 13084
rect 6092 13082 6116 13084
rect 6172 13082 6196 13084
rect 6034 13030 6036 13082
rect 6098 13030 6110 13082
rect 6172 13030 6174 13082
rect 6012 13028 6036 13030
rect 6092 13028 6116 13030
rect 6172 13028 6196 13030
rect 5956 13008 6252 13028
rect 6380 12986 6408 13262
rect 6368 12980 6420 12986
rect 6368 12922 6420 12928
rect 5816 12844 5868 12850
rect 5816 12786 5868 12792
rect 5828 12238 5856 12786
rect 6380 12753 6408 12922
rect 6366 12744 6422 12753
rect 6366 12679 6422 12688
rect 5998 12336 6054 12345
rect 5998 12271 6000 12280
rect 6052 12271 6054 12280
rect 6274 12336 6330 12345
rect 6274 12271 6330 12280
rect 6000 12242 6052 12248
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 5956 11996 6252 12016
rect 6012 11994 6036 11996
rect 6092 11994 6116 11996
rect 6172 11994 6196 11996
rect 6034 11942 6036 11994
rect 6098 11942 6110 11994
rect 6172 11942 6174 11994
rect 6012 11940 6036 11942
rect 6092 11940 6116 11942
rect 6172 11940 6196 11942
rect 5956 11920 6252 11940
rect 6288 11830 6316 12271
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6380 11898 6408 12174
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 6276 11824 6328 11830
rect 6276 11766 6328 11772
rect 6564 11354 6592 14826
rect 7116 14634 7144 19654
rect 7196 18624 7248 18630
rect 7196 18566 7248 18572
rect 7208 17134 7236 18566
rect 7196 17128 7248 17134
rect 7196 17070 7248 17076
rect 7208 16794 7236 17070
rect 7196 16788 7248 16794
rect 7196 16730 7248 16736
rect 6840 14606 7144 14634
rect 6840 14550 6868 14606
rect 6828 14544 6880 14550
rect 7300 14498 7328 21247
rect 8312 20618 8340 23520
rect 10956 21244 11252 21264
rect 11012 21242 11036 21244
rect 11092 21242 11116 21244
rect 11172 21242 11196 21244
rect 11034 21190 11036 21242
rect 11098 21190 11110 21242
rect 11172 21190 11174 21242
rect 11012 21188 11036 21190
rect 11092 21188 11116 21190
rect 11172 21188 11196 21190
rect 10956 21168 11252 21188
rect 10508 21004 10560 21010
rect 10508 20946 10560 20952
rect 10140 20936 10192 20942
rect 10140 20878 10192 20884
rect 10232 20936 10284 20942
rect 10232 20878 10284 20884
rect 9956 20868 10008 20874
rect 9956 20810 10008 20816
rect 8760 20800 8812 20806
rect 8760 20742 8812 20748
rect 8852 20800 8904 20806
rect 8852 20742 8904 20748
rect 8220 20602 8340 20618
rect 8208 20596 8340 20602
rect 8260 20590 8340 20596
rect 8208 20538 8260 20544
rect 8772 20505 8800 20742
rect 8758 20496 8814 20505
rect 8758 20431 8760 20440
rect 8812 20431 8814 20440
rect 8760 20402 8812 20408
rect 8864 20058 8892 20742
rect 9312 20324 9364 20330
rect 9312 20266 9364 20272
rect 8024 20052 8076 20058
rect 8024 19994 8076 20000
rect 8484 20052 8536 20058
rect 8484 19994 8536 20000
rect 8852 20052 8904 20058
rect 8852 19994 8904 20000
rect 8036 19961 8064 19994
rect 8022 19952 8078 19961
rect 8022 19887 8078 19896
rect 8024 19236 8076 19242
rect 8024 19178 8076 19184
rect 8036 18154 8064 19178
rect 8496 18970 8524 19994
rect 8852 19916 8904 19922
rect 8852 19858 8904 19864
rect 8576 19848 8628 19854
rect 8576 19790 8628 19796
rect 8588 19174 8616 19790
rect 8864 19174 8892 19858
rect 9324 19378 9352 20266
rect 9680 20256 9732 20262
rect 9680 20198 9732 20204
rect 9312 19372 9364 19378
rect 9312 19314 9364 19320
rect 8576 19168 8628 19174
rect 8576 19110 8628 19116
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8392 18692 8444 18698
rect 8392 18634 8444 18640
rect 8208 18284 8260 18290
rect 8208 18226 8260 18232
rect 8024 18148 8076 18154
rect 8024 18090 8076 18096
rect 8220 17882 8248 18226
rect 8404 18222 8432 18634
rect 8864 18426 8892 19110
rect 8852 18420 8904 18426
rect 8852 18362 8904 18368
rect 9692 18306 9720 20198
rect 9968 19310 9996 20810
rect 10152 20602 10180 20878
rect 10140 20596 10192 20602
rect 10140 20538 10192 20544
rect 10152 19514 10180 20538
rect 10244 20262 10272 20878
rect 10520 20330 10548 20946
rect 11624 20534 11652 23520
rect 12532 22228 12584 22234
rect 12532 22170 12584 22176
rect 11612 20528 11664 20534
rect 11612 20470 11664 20476
rect 12438 20496 12494 20505
rect 12438 20431 12440 20440
rect 12492 20431 12494 20440
rect 12440 20402 12492 20408
rect 10784 20392 10836 20398
rect 10784 20334 10836 20340
rect 10508 20324 10560 20330
rect 10508 20266 10560 20272
rect 10232 20256 10284 20262
rect 10232 20198 10284 20204
rect 10520 20058 10548 20266
rect 10508 20052 10560 20058
rect 10508 19994 10560 20000
rect 10796 19922 10824 20334
rect 10956 20156 11252 20176
rect 11012 20154 11036 20156
rect 11092 20154 11116 20156
rect 11172 20154 11196 20156
rect 11034 20102 11036 20154
rect 11098 20102 11110 20154
rect 11172 20102 11174 20154
rect 11012 20100 11036 20102
rect 11092 20100 11116 20102
rect 11172 20100 11196 20102
rect 10956 20080 11252 20100
rect 12452 20058 12480 20402
rect 12440 20052 12492 20058
rect 12440 19994 12492 20000
rect 10784 19916 10836 19922
rect 10784 19858 10836 19864
rect 12440 19916 12492 19922
rect 12440 19858 12492 19864
rect 10600 19712 10652 19718
rect 10600 19654 10652 19660
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 10048 19440 10100 19446
rect 10048 19382 10100 19388
rect 9956 19304 10008 19310
rect 9956 19246 10008 19252
rect 9772 18828 9824 18834
rect 9772 18770 9824 18776
rect 9600 18290 9720 18306
rect 9588 18284 9720 18290
rect 9640 18278 9720 18284
rect 9588 18226 9640 18232
rect 8392 18216 8444 18222
rect 9784 18204 9812 18770
rect 10060 18329 10088 19382
rect 10508 19304 10560 19310
rect 10506 19272 10508 19281
rect 10560 19272 10562 19281
rect 10506 19207 10562 19216
rect 10612 19174 10640 19654
rect 10600 19168 10652 19174
rect 10598 19136 10600 19145
rect 10652 19136 10654 19145
rect 10598 19071 10654 19080
rect 10796 18970 10824 19858
rect 10968 19848 11020 19854
rect 10874 19816 10930 19825
rect 10968 19790 11020 19796
rect 10874 19751 10876 19760
rect 10928 19751 10930 19760
rect 10876 19722 10928 19728
rect 10888 19378 10916 19722
rect 10980 19446 11008 19790
rect 10968 19440 11020 19446
rect 10968 19382 11020 19388
rect 10876 19372 10928 19378
rect 10876 19314 10928 19320
rect 10784 18964 10836 18970
rect 10784 18906 10836 18912
rect 10888 18766 10916 19314
rect 12452 19174 12480 19858
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 10956 19068 11252 19088
rect 11012 19066 11036 19068
rect 11092 19066 11116 19068
rect 11172 19066 11196 19068
rect 11034 19014 11036 19066
rect 11098 19014 11110 19066
rect 11172 19014 11174 19066
rect 11012 19012 11036 19014
rect 11092 19012 11116 19014
rect 11172 19012 11196 19014
rect 10956 18992 11252 19012
rect 10140 18760 10192 18766
rect 10140 18702 10192 18708
rect 10876 18760 10928 18766
rect 10876 18702 10928 18708
rect 10046 18320 10102 18329
rect 10046 18255 10102 18264
rect 8392 18158 8444 18164
rect 9692 18176 9812 18204
rect 9692 18086 9720 18176
rect 9680 18080 9732 18086
rect 9678 18048 9680 18057
rect 9732 18048 9734 18057
rect 9678 17983 9734 17992
rect 8208 17876 8260 17882
rect 8208 17818 8260 17824
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 7484 17066 7512 17478
rect 9588 17264 9640 17270
rect 9692 17241 9720 17983
rect 9588 17206 9640 17212
rect 9678 17232 9734 17241
rect 7472 17060 7524 17066
rect 7472 17002 7524 17008
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 8220 15162 8248 15982
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8404 15366 8432 15846
rect 8392 15360 8444 15366
rect 8392 15302 8444 15308
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8220 14618 8248 15098
rect 8404 15026 8432 15302
rect 8588 15162 8616 16934
rect 9600 16697 9628 17206
rect 10060 17218 10088 18255
rect 10152 17746 10180 18702
rect 10888 18426 10916 18702
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10232 18148 10284 18154
rect 10232 18090 10284 18096
rect 10244 17882 10272 18090
rect 10232 17876 10284 17882
rect 10232 17818 10284 17824
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 10152 17338 10180 17682
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 10060 17190 10180 17218
rect 9678 17167 9734 17176
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9586 16688 9642 16697
rect 9586 16623 9642 16632
rect 8760 15972 8812 15978
rect 8760 15914 8812 15920
rect 8576 15156 8628 15162
rect 8576 15098 8628 15104
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8588 14890 8616 15098
rect 8576 14884 8628 14890
rect 8628 14844 8708 14872
rect 8576 14826 8628 14832
rect 8208 14612 8260 14618
rect 8208 14554 8260 14560
rect 6828 14486 6880 14492
rect 7116 14470 7328 14498
rect 8300 14476 8352 14482
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6932 13938 6960 14214
rect 6920 13932 6972 13938
rect 6920 13874 6972 13880
rect 6734 13696 6790 13705
rect 6734 13631 6790 13640
rect 6644 13524 6696 13530
rect 6644 13466 6696 13472
rect 6656 12646 6684 13466
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6656 12481 6684 12582
rect 6642 12472 6698 12481
rect 6642 12407 6698 12416
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 5956 10908 6252 10928
rect 6012 10906 6036 10908
rect 6092 10906 6116 10908
rect 6172 10906 6196 10908
rect 6034 10854 6036 10906
rect 6098 10854 6110 10906
rect 6172 10854 6174 10906
rect 6012 10852 6036 10854
rect 6092 10852 6116 10854
rect 6172 10852 6196 10854
rect 5956 10832 6252 10852
rect 6564 10810 6592 11290
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 5816 10736 5868 10742
rect 5816 10678 5868 10684
rect 5828 9722 5856 10678
rect 6564 10606 6592 10746
rect 6656 10674 6684 12407
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6552 10600 6604 10606
rect 6274 10568 6330 10577
rect 6748 10577 6776 13631
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 7024 12986 7052 13262
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 7116 12356 7144 14470
rect 8300 14418 8352 14424
rect 8312 13938 8340 14418
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 8036 13530 8064 13806
rect 8312 13705 8340 13874
rect 8576 13728 8628 13734
rect 8298 13696 8354 13705
rect 8576 13670 8628 13676
rect 8298 13631 8354 13640
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 8036 12646 8064 13262
rect 8024 12640 8076 12646
rect 8024 12582 8076 12588
rect 8036 12374 8064 12582
rect 8024 12368 8076 12374
rect 7116 12328 7236 12356
rect 6552 10542 6604 10548
rect 6734 10568 6790 10577
rect 6274 10503 6330 10512
rect 6368 10532 6420 10538
rect 5956 9820 6252 9840
rect 6012 9818 6036 9820
rect 6092 9818 6116 9820
rect 6172 9818 6196 9820
rect 6034 9766 6036 9818
rect 6098 9766 6110 9818
rect 6172 9766 6174 9818
rect 6012 9764 6036 9766
rect 6092 9764 6116 9766
rect 6172 9764 6196 9766
rect 5956 9744 6252 9764
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 6092 9512 6144 9518
rect 6092 9454 6144 9460
rect 6104 9178 6132 9454
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 5956 8732 6252 8752
rect 6012 8730 6036 8732
rect 6092 8730 6116 8732
rect 6172 8730 6196 8732
rect 6034 8678 6036 8730
rect 6098 8678 6110 8730
rect 6172 8678 6174 8730
rect 6012 8676 6036 8678
rect 6092 8676 6116 8678
rect 6172 8676 6196 8678
rect 5956 8656 6252 8676
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5828 7410 5856 7890
rect 6288 7834 6316 10503
rect 6734 10503 6790 10512
rect 6368 10474 6420 10480
rect 6380 10266 6408 10474
rect 6644 10464 6696 10470
rect 6458 10432 6514 10441
rect 6644 10406 6696 10412
rect 6458 10367 6514 10376
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6472 9994 6500 10367
rect 6460 9988 6512 9994
rect 6460 9930 6512 9936
rect 6472 9178 6500 9930
rect 6552 9512 6604 9518
rect 6550 9480 6552 9489
rect 6604 9480 6606 9489
rect 6550 9415 6606 9424
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 6472 8362 6500 8978
rect 6460 8356 6512 8362
rect 6460 8298 6512 8304
rect 6288 7806 6408 7834
rect 5956 7644 6252 7664
rect 6012 7642 6036 7644
rect 6092 7642 6116 7644
rect 6172 7642 6196 7644
rect 6034 7590 6036 7642
rect 6098 7590 6110 7642
rect 6172 7590 6174 7642
rect 6012 7588 6036 7590
rect 6092 7588 6116 7590
rect 6172 7588 6196 7590
rect 5956 7568 6252 7588
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6288 7206 6316 7346
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5828 6458 5856 6938
rect 5998 6896 6054 6905
rect 5998 6831 6000 6840
rect 6052 6831 6054 6840
rect 6000 6802 6052 6808
rect 6288 6798 6316 7142
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 5956 6556 6252 6576
rect 6012 6554 6036 6556
rect 6092 6554 6116 6556
rect 6172 6554 6196 6556
rect 6034 6502 6036 6554
rect 6098 6502 6110 6554
rect 6172 6502 6174 6554
rect 6012 6500 6036 6502
rect 6092 6500 6116 6502
rect 6172 6500 6196 6502
rect 5956 6480 6252 6500
rect 6288 6458 6316 6734
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 5956 5468 6252 5488
rect 6012 5466 6036 5468
rect 6092 5466 6116 5468
rect 6172 5466 6196 5468
rect 6034 5414 6036 5466
rect 6098 5414 6110 5466
rect 6172 5414 6174 5466
rect 6012 5412 6036 5414
rect 6092 5412 6116 5414
rect 6172 5412 6196 5414
rect 5956 5392 6252 5412
rect 6288 5370 6316 5510
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6380 4826 6408 7806
rect 6472 5273 6500 8298
rect 6564 6458 6592 9415
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6458 5264 6514 5273
rect 6458 5199 6514 5208
rect 6564 5114 6592 6258
rect 6656 5352 6684 10406
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 6748 9654 6776 10066
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6736 9648 6788 9654
rect 6736 9590 6788 9596
rect 6840 9450 6868 9998
rect 7208 9636 7236 12328
rect 8024 12310 8076 12316
rect 7380 11280 7432 11286
rect 7380 11222 7432 11228
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 7300 10674 7328 10950
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7392 10470 7420 11222
rect 7748 11008 7800 11014
rect 7748 10950 7800 10956
rect 7760 10810 7788 10950
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 7392 9926 7420 10406
rect 7760 10266 7788 10746
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 8208 10124 8260 10130
rect 8312 10112 8340 13631
rect 8392 13388 8444 13394
rect 8392 13330 8444 13336
rect 8404 12646 8432 13330
rect 8588 12850 8616 13670
rect 8680 13326 8708 14844
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 8680 12918 8708 13262
rect 8772 12918 8800 15914
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 9692 15570 9720 15846
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9692 15162 9720 15506
rect 9770 15464 9826 15473
rect 9770 15399 9826 15408
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 9232 14278 9260 14758
rect 9784 14498 9812 15399
rect 9876 14657 9904 16934
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9968 14822 9996 15506
rect 9956 14816 10008 14822
rect 9956 14758 10008 14764
rect 9862 14648 9918 14657
rect 9862 14583 9918 14592
rect 9784 14470 9904 14498
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 9232 13938 9260 14214
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 8668 12912 8720 12918
rect 8668 12854 8720 12860
rect 8760 12912 8812 12918
rect 8760 12854 8812 12860
rect 8576 12844 8628 12850
rect 8576 12786 8628 12792
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8392 12640 8444 12646
rect 8392 12582 8444 12588
rect 8404 12345 8432 12582
rect 8680 12442 8708 12718
rect 8864 12442 8892 12786
rect 9140 12714 9168 13126
rect 9128 12708 9180 12714
rect 9128 12650 9180 12656
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8390 12336 8446 12345
rect 8390 12271 8446 12280
rect 9232 11354 9260 13874
rect 9404 13796 9456 13802
rect 9404 13738 9456 13744
rect 9416 12968 9444 13738
rect 9496 13252 9548 13258
rect 9496 13194 9548 13200
rect 9508 13138 9536 13194
rect 9586 13152 9642 13161
rect 9508 13110 9586 13138
rect 9586 13087 9642 13096
rect 9586 13016 9642 13025
rect 9416 12960 9586 12968
rect 9416 12951 9642 12960
rect 9416 12940 9628 12951
rect 9772 12912 9824 12918
rect 9586 12880 9642 12889
rect 9772 12854 9824 12860
rect 9586 12815 9588 12824
rect 9640 12815 9642 12824
rect 9588 12786 9640 12792
rect 9496 12776 9548 12782
rect 9310 12744 9366 12753
rect 9310 12679 9366 12688
rect 9494 12744 9496 12753
rect 9548 12744 9550 12753
rect 9494 12679 9550 12688
rect 9588 12708 9640 12714
rect 9324 11626 9352 12679
rect 9588 12650 9640 12656
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9600 12594 9628 12650
rect 9312 11620 9364 11626
rect 9312 11562 9364 11568
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8404 10674 8432 10950
rect 9508 10674 9536 12582
rect 9600 12566 9720 12594
rect 9692 12442 9720 12566
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9678 12336 9734 12345
rect 9678 12271 9734 12280
rect 9692 12238 9720 12271
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9692 11393 9720 12174
rect 9678 11384 9734 11393
rect 9678 11319 9734 11328
rect 9692 11286 9720 11319
rect 9680 11280 9732 11286
rect 9680 11222 9732 11228
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 8404 10470 8432 10610
rect 9600 10606 9628 10950
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 8392 10464 8444 10470
rect 8390 10432 8392 10441
rect 8444 10432 8446 10441
rect 8390 10367 8446 10376
rect 8588 10266 8616 10542
rect 8852 10532 8904 10538
rect 8852 10474 8904 10480
rect 8864 10266 8892 10474
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9508 10266 9536 10406
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 8260 10084 8340 10112
rect 8208 10066 8260 10072
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 7288 9648 7340 9654
rect 7208 9608 7288 9636
rect 7288 9590 7340 9596
rect 7392 9586 7420 9862
rect 8024 9716 8076 9722
rect 8128 9704 8156 9862
rect 8220 9722 8248 10066
rect 8076 9676 8156 9704
rect 8024 9658 8076 9664
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7746 9616 7802 9625
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 6828 9444 6880 9450
rect 6828 9386 6880 9392
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6748 6322 6776 9318
rect 6840 9178 6868 9386
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6932 8498 6960 9386
rect 7288 9104 7340 9110
rect 7286 9072 7288 9081
rect 7340 9072 7342 9081
rect 7286 9007 7342 9016
rect 7392 8974 7420 9522
rect 7484 9042 7512 9590
rect 7746 9551 7802 9560
rect 7760 9518 7788 9551
rect 7748 9512 7800 9518
rect 7748 9454 7800 9460
rect 8128 9042 8156 9676
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 9692 9518 9720 11222
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 7472 9036 7524 9042
rect 7472 8978 7524 8984
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7392 8090 7420 8910
rect 7484 8294 7512 8978
rect 8588 8634 8616 8978
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 9048 8430 9076 8774
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7932 8288 7984 8294
rect 7932 8230 7984 8236
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6840 7002 6868 7142
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 7208 6254 7236 6734
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6656 5324 6776 5352
rect 6642 5264 6698 5273
rect 6642 5199 6644 5208
rect 6696 5199 6698 5208
rect 6644 5170 6696 5176
rect 6472 5086 6592 5114
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 5724 4752 5776 4758
rect 5724 4694 5776 4700
rect 6276 4480 6328 4486
rect 6276 4422 6328 4428
rect 5956 4380 6252 4400
rect 6012 4378 6036 4380
rect 6092 4378 6116 4380
rect 6172 4378 6196 4380
rect 6034 4326 6036 4378
rect 6098 4326 6110 4378
rect 6172 4326 6174 4378
rect 6012 4324 6036 4326
rect 6092 4324 6116 4326
rect 6172 4324 6196 4326
rect 5956 4304 6252 4324
rect 5460 4146 5580 4162
rect 5448 4140 5580 4146
rect 5500 4134 5580 4140
rect 5448 4082 5500 4088
rect 4618 4040 4674 4049
rect 4540 3998 4618 4026
rect 4618 3975 4674 3984
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 4528 3936 4580 3942
rect 4528 3878 4580 3884
rect 4264 3505 4292 3878
rect 4434 3632 4490 3641
rect 4434 3567 4490 3576
rect 4250 3496 4306 3505
rect 4250 3431 4306 3440
rect 4448 3194 4476 3567
rect 4540 3369 4568 3878
rect 4526 3360 4582 3369
rect 4526 3295 4582 3304
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4632 2990 4660 3975
rect 5814 3904 5870 3913
rect 5814 3839 5870 3848
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 4816 3194 4844 3538
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4080 2502 4200 2530
rect 5368 2514 5396 3334
rect 5460 2650 5488 3674
rect 5828 3534 5856 3839
rect 6288 3670 6316 4422
rect 6380 4214 6408 4762
rect 6472 4622 6500 5086
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6368 4208 6420 4214
rect 6368 4150 6420 4156
rect 6472 3942 6500 4558
rect 6564 4282 6592 4558
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6276 3664 6328 3670
rect 6276 3606 6328 3612
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 5828 3194 5856 3470
rect 5956 3292 6252 3312
rect 6012 3290 6036 3292
rect 6092 3290 6116 3292
rect 6172 3290 6196 3292
rect 6034 3238 6036 3290
rect 6098 3238 6110 3290
rect 6172 3238 6174 3290
rect 6012 3236 6036 3238
rect 6092 3236 6116 3238
rect 6172 3236 6196 3238
rect 5956 3216 6252 3236
rect 6288 3194 6316 3606
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 6472 2650 6500 3878
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6564 3097 6592 3470
rect 6550 3088 6606 3097
rect 6550 3023 6552 3032
rect 6604 3023 6606 3032
rect 6552 2994 6604 3000
rect 6748 2990 6776 5324
rect 6840 5250 6868 6054
rect 7208 5914 7236 6190
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7576 5710 7604 6258
rect 7944 5846 7972 8230
rect 9048 7750 9076 8366
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 8312 7342 8340 7686
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8312 6934 8340 7278
rect 9600 7154 9628 8298
rect 9680 7200 9732 7206
rect 9600 7148 9680 7154
rect 9600 7142 9732 7148
rect 9600 7126 9720 7142
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 9128 6724 9180 6730
rect 9128 6666 9180 6672
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 7932 5840 7984 5846
rect 7930 5808 7932 5817
rect 7984 5808 7986 5817
rect 7656 5772 7708 5778
rect 7930 5743 7986 5752
rect 7656 5714 7708 5720
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6840 5222 6960 5250
rect 7024 5234 7052 5510
rect 6932 5166 6960 5222
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6840 3602 6868 4966
rect 7024 4826 7052 5170
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 7484 4282 7512 5170
rect 7576 4622 7604 5646
rect 7668 5273 7696 5714
rect 7944 5370 7972 5743
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 7654 5264 7710 5273
rect 7654 5199 7710 5208
rect 8116 4752 8168 4758
rect 8116 4694 8168 4700
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 7484 3534 7512 4218
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7484 3194 7512 3470
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 7748 2916 7800 2922
rect 7748 2858 7800 2864
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 5356 2508 5408 2514
rect 4080 921 4108 2502
rect 5356 2450 5408 2456
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 4066 912 4122 921
rect 4066 847 4122 856
rect 4908 480 4936 2382
rect 5816 2304 5868 2310
rect 5816 2246 5868 2252
rect 5828 2145 5856 2246
rect 5956 2204 6252 2224
rect 6012 2202 6036 2204
rect 6092 2202 6116 2204
rect 6172 2202 6196 2204
rect 6034 2150 6036 2202
rect 6098 2150 6110 2202
rect 6172 2150 6174 2202
rect 6012 2148 6036 2150
rect 6092 2148 6116 2150
rect 6172 2148 6196 2150
rect 5814 2136 5870 2145
rect 5956 2128 6252 2148
rect 5814 2071 5870 2080
rect 6380 480 6408 2382
rect 7760 480 7788 2858
rect 8128 2514 8156 4694
rect 8312 4434 8340 6326
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8864 5914 8892 6258
rect 9140 6186 9168 6666
rect 9600 6322 9628 7126
rect 9680 6928 9732 6934
rect 9680 6870 9732 6876
rect 9588 6316 9640 6322
rect 9588 6258 9640 6264
rect 9128 6180 9180 6186
rect 9128 6122 9180 6128
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 8220 4406 8340 4434
rect 8220 2650 8248 4406
rect 9692 4078 9720 6870
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9036 3936 9088 3942
rect 9034 3904 9036 3913
rect 9088 3904 9090 3913
rect 9034 3839 9090 3848
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 9784 2514 9812 12854
rect 9876 11150 9904 14470
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 10060 12986 10088 13126
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 10046 12608 10102 12617
rect 10046 12543 10102 12552
rect 10060 12306 10088 12543
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10060 11898 10088 12242
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 10152 11642 10180 17190
rect 10336 16794 10364 18158
rect 10956 17980 11252 18000
rect 11012 17978 11036 17980
rect 11092 17978 11116 17980
rect 11172 17978 11196 17980
rect 11034 17926 11036 17978
rect 11098 17926 11110 17978
rect 11172 17926 11174 17978
rect 11012 17924 11036 17926
rect 11092 17924 11116 17926
rect 11172 17924 11196 17926
rect 10956 17904 11252 17924
rect 10600 17740 10652 17746
rect 10600 17682 10652 17688
rect 10784 17740 10836 17746
rect 10784 17682 10836 17688
rect 10416 17536 10468 17542
rect 10612 17513 10640 17682
rect 10416 17478 10468 17484
rect 10598 17504 10654 17513
rect 10428 16998 10456 17478
rect 10598 17439 10654 17448
rect 10612 17270 10640 17439
rect 10600 17264 10652 17270
rect 10600 17206 10652 17212
rect 10796 16998 10824 17682
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 10888 17270 10916 17614
rect 10876 17264 10928 17270
rect 10876 17206 10928 17212
rect 12348 17264 12400 17270
rect 12452 17252 12480 19110
rect 12400 17224 12480 17252
rect 12348 17206 12400 17212
rect 10416 16992 10468 16998
rect 10416 16934 10468 16940
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10324 16788 10376 16794
rect 10324 16730 10376 16736
rect 10428 16697 10456 16934
rect 10414 16688 10470 16697
rect 10414 16623 10470 16632
rect 10508 16652 10560 16658
rect 10508 16594 10560 16600
rect 10520 16250 10548 16594
rect 10600 16584 10652 16590
rect 10598 16552 10600 16561
rect 10652 16552 10654 16561
rect 10598 16487 10654 16496
rect 10508 16244 10560 16250
rect 10508 16186 10560 16192
rect 10520 15745 10548 16186
rect 10612 16182 10640 16487
rect 10600 16176 10652 16182
rect 10600 16118 10652 16124
rect 10796 16017 10824 16934
rect 10888 16590 10916 17206
rect 11610 17096 11666 17105
rect 11610 17031 11612 17040
rect 11664 17031 11666 17040
rect 12070 17096 12126 17105
rect 12070 17031 12126 17040
rect 11612 17002 11664 17008
rect 10956 16892 11252 16912
rect 11012 16890 11036 16892
rect 11092 16890 11116 16892
rect 11172 16890 11196 16892
rect 11034 16838 11036 16890
rect 11098 16838 11110 16890
rect 11172 16838 11174 16890
rect 11012 16836 11036 16838
rect 11092 16836 11116 16838
rect 11172 16836 11196 16838
rect 10956 16816 11252 16836
rect 11978 16688 12034 16697
rect 11978 16623 12034 16632
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 10888 16250 10916 16526
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 10782 16008 10838 16017
rect 10782 15943 10838 15952
rect 10956 15804 11252 15824
rect 11012 15802 11036 15804
rect 11092 15802 11116 15804
rect 11172 15802 11196 15804
rect 11034 15750 11036 15802
rect 11098 15750 11110 15802
rect 11172 15750 11174 15802
rect 11012 15748 11036 15750
rect 11092 15748 11116 15750
rect 11172 15748 11196 15750
rect 10506 15736 10562 15745
rect 10956 15728 11252 15748
rect 10506 15671 10562 15680
rect 11888 15632 11940 15638
rect 11888 15574 11940 15580
rect 10692 15496 10744 15502
rect 10692 15438 10744 15444
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 10600 15156 10652 15162
rect 10704 15144 10732 15438
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 10652 15116 10732 15144
rect 10600 15098 10652 15104
rect 10612 14482 10640 15098
rect 11072 14872 11100 15302
rect 11808 15162 11836 15438
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 10796 14844 11100 14872
rect 10796 14550 10824 14844
rect 11900 14822 11928 15574
rect 11992 15065 12020 16623
rect 11978 15056 12034 15065
rect 11978 14991 12034 15000
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 10956 14716 11252 14736
rect 11012 14714 11036 14716
rect 11092 14714 11116 14716
rect 11172 14714 11196 14716
rect 11034 14662 11036 14714
rect 11098 14662 11110 14714
rect 11172 14662 11174 14714
rect 11012 14660 11036 14662
rect 11092 14660 11116 14662
rect 11172 14660 11196 14662
rect 10956 14640 11252 14660
rect 10784 14544 10836 14550
rect 10784 14486 10836 14492
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10612 14074 10640 14418
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 10796 13870 10824 14486
rect 11900 14278 11928 14758
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10796 13394 10824 13806
rect 10784 13388 10836 13394
rect 10784 13330 10836 13336
rect 10782 13288 10838 13297
rect 10782 13223 10838 13232
rect 10508 13184 10560 13190
rect 10508 13126 10560 13132
rect 10690 13152 10746 13161
rect 10520 12782 10548 13126
rect 10690 13087 10746 13096
rect 10508 12776 10560 12782
rect 10508 12718 10560 12724
rect 10600 12640 10652 12646
rect 10598 12608 10600 12617
rect 10652 12608 10654 12617
rect 10598 12543 10654 12552
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 9968 11614 10180 11642
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9864 10736 9916 10742
rect 9862 10704 9864 10713
rect 9916 10704 9918 10713
rect 9862 10639 9918 10648
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9876 10198 9904 10542
rect 9968 10305 9996 11614
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 10152 10674 10180 11494
rect 10244 11354 10272 12174
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10048 10600 10100 10606
rect 10048 10542 10100 10548
rect 9954 10296 10010 10305
rect 10060 10266 10088 10542
rect 9954 10231 10010 10240
rect 10048 10260 10100 10266
rect 10048 10202 10100 10208
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9876 9722 9904 10134
rect 9864 9716 9916 9722
rect 9916 9676 9996 9704
rect 9864 9658 9916 9664
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9876 6458 9904 7210
rect 9864 6452 9916 6458
rect 9864 6394 9916 6400
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9876 3738 9904 4014
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9968 3505 9996 9676
rect 10244 5846 10272 11086
rect 10324 10736 10376 10742
rect 10324 10678 10376 10684
rect 10336 10538 10364 10678
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 10428 10266 10456 11698
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10520 10810 10548 11086
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10520 10266 10548 10746
rect 10612 10674 10640 11086
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10704 10266 10732 13087
rect 10796 12918 10824 13223
rect 10784 12912 10836 12918
rect 10784 12854 10836 12860
rect 10888 12850 10916 14214
rect 10956 13628 11252 13648
rect 11012 13626 11036 13628
rect 11092 13626 11116 13628
rect 11172 13626 11196 13628
rect 11034 13574 11036 13626
rect 11098 13574 11110 13626
rect 11172 13574 11174 13626
rect 11012 13572 11036 13574
rect 11092 13572 11116 13574
rect 11172 13572 11196 13574
rect 10956 13552 11252 13572
rect 11336 13456 11388 13462
rect 11336 13398 11388 13404
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 11058 13288 11114 13297
rect 10980 13246 11058 13274
rect 10980 13025 11008 13246
rect 11058 13223 11114 13232
rect 10966 13016 11022 13025
rect 10966 12951 11022 12960
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 11164 12782 11192 13330
rect 11152 12776 11204 12782
rect 11150 12744 11152 12753
rect 11204 12744 11206 12753
rect 10784 12708 10836 12714
rect 11150 12679 11206 12688
rect 10784 12650 10836 12656
rect 10796 12481 10824 12650
rect 10956 12540 11252 12560
rect 11012 12538 11036 12540
rect 11092 12538 11116 12540
rect 11172 12538 11196 12540
rect 11034 12486 11036 12538
rect 11098 12486 11110 12538
rect 11172 12486 11174 12538
rect 11012 12484 11036 12486
rect 11092 12484 11116 12486
rect 11172 12484 11196 12486
rect 10782 12472 10838 12481
rect 10956 12464 11252 12484
rect 11348 12442 11376 13398
rect 11520 13252 11572 13258
rect 11520 13194 11572 13200
rect 11532 12986 11560 13194
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11426 12744 11482 12753
rect 11426 12679 11482 12688
rect 11440 12646 11468 12679
rect 11428 12640 11480 12646
rect 11428 12582 11480 12588
rect 10782 12407 10784 12416
rect 10836 12407 10838 12416
rect 11336 12436 11388 12442
rect 10784 12378 10836 12384
rect 11336 12378 11388 12384
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 10796 11694 10824 12378
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11334 11792 11390 11801
rect 11334 11727 11390 11736
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10416 10260 10468 10266
rect 10416 10202 10468 10208
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10428 10062 10456 10202
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10428 9110 10456 9998
rect 10704 9722 10732 10202
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10416 9104 10468 9110
rect 10416 9046 10468 9052
rect 10428 8634 10456 9046
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10796 8430 10824 11494
rect 10956 11452 11252 11472
rect 11012 11450 11036 11452
rect 11092 11450 11116 11452
rect 11172 11450 11196 11452
rect 11034 11398 11036 11450
rect 11098 11398 11110 11450
rect 11172 11398 11174 11450
rect 11012 11396 11036 11398
rect 11092 11396 11116 11398
rect 11172 11396 11196 11398
rect 10956 11376 11252 11396
rect 11348 11393 11376 11727
rect 11440 11558 11468 12174
rect 11900 11898 11928 12378
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11428 11552 11480 11558
rect 11428 11494 11480 11500
rect 11518 11520 11574 11529
rect 11334 11384 11390 11393
rect 11334 11319 11390 11328
rect 11440 11257 11468 11494
rect 11518 11455 11574 11464
rect 11426 11248 11482 11257
rect 10968 11212 11020 11218
rect 11426 11183 11482 11192
rect 10968 11154 11020 11160
rect 10980 10826 11008 11154
rect 10888 10798 11100 10826
rect 10888 9654 10916 10798
rect 11072 10674 11100 10798
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 11336 10600 11388 10606
rect 11336 10542 11388 10548
rect 10956 10364 11252 10384
rect 11012 10362 11036 10364
rect 11092 10362 11116 10364
rect 11172 10362 11196 10364
rect 11034 10310 11036 10362
rect 11098 10310 11110 10362
rect 11172 10310 11174 10362
rect 11012 10308 11036 10310
rect 11092 10308 11116 10310
rect 11172 10308 11196 10310
rect 10956 10288 11252 10308
rect 10968 9988 11020 9994
rect 10968 9930 11020 9936
rect 10876 9648 10928 9654
rect 10876 9590 10928 9596
rect 10980 9586 11008 9930
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10956 9276 11252 9296
rect 11012 9274 11036 9276
rect 11092 9274 11116 9276
rect 11172 9274 11196 9276
rect 11034 9222 11036 9274
rect 11098 9222 11110 9274
rect 11172 9222 11174 9274
rect 11012 9220 11036 9222
rect 11092 9220 11116 9222
rect 11172 9220 11196 9222
rect 10956 9200 11252 9220
rect 11348 9178 11376 10542
rect 11532 10198 11560 11455
rect 11520 10192 11572 10198
rect 11520 10134 11572 10140
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10796 7886 10824 8230
rect 10956 8188 11252 8208
rect 11012 8186 11036 8188
rect 11092 8186 11116 8188
rect 11172 8186 11196 8188
rect 11034 8134 11036 8186
rect 11098 8134 11110 8186
rect 11172 8134 11174 8186
rect 11012 8132 11036 8134
rect 11092 8132 11116 8134
rect 11172 8132 11196 8134
rect 10956 8112 11252 8132
rect 11336 8016 11388 8022
rect 11336 7958 11388 7964
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10796 7206 10824 7822
rect 11348 7206 11376 7958
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 11336 7200 11388 7206
rect 11336 7142 11388 7148
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11794 7168 11850 7177
rect 10796 6934 10824 7142
rect 10956 7100 11252 7120
rect 11012 7098 11036 7100
rect 11092 7098 11116 7100
rect 11172 7098 11196 7100
rect 11034 7046 11036 7098
rect 11098 7046 11110 7098
rect 11172 7046 11174 7098
rect 11012 7044 11036 7046
rect 11092 7044 11116 7046
rect 11172 7044 11196 7046
rect 10956 7024 11252 7044
rect 11348 7002 11376 7142
rect 11336 6996 11388 7002
rect 11336 6938 11388 6944
rect 10784 6928 10836 6934
rect 10784 6870 10836 6876
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10428 6322 10456 6598
rect 10416 6316 10468 6322
rect 10416 6258 10468 6264
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10416 6180 10468 6186
rect 10416 6122 10468 6128
rect 10428 5914 10456 6122
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 10508 5908 10560 5914
rect 10508 5850 10560 5856
rect 10232 5840 10284 5846
rect 10232 5782 10284 5788
rect 10244 5302 10272 5782
rect 10520 5370 10548 5850
rect 10704 5370 10732 6258
rect 10956 6012 11252 6032
rect 11012 6010 11036 6012
rect 11092 6010 11116 6012
rect 11172 6010 11196 6012
rect 11034 5958 11036 6010
rect 11098 5958 11110 6010
rect 11172 5958 11174 6010
rect 11012 5956 11036 5958
rect 11092 5956 11116 5958
rect 11172 5956 11196 5958
rect 10956 5936 11252 5956
rect 11348 5710 11376 6938
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10232 5296 10284 5302
rect 10232 5238 10284 5244
rect 10244 5137 10272 5238
rect 11348 5234 11376 5646
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 10230 5128 10286 5137
rect 10230 5063 10286 5072
rect 10796 4826 10824 5170
rect 11440 5098 11468 5510
rect 11428 5092 11480 5098
rect 11428 5034 11480 5040
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 10956 4924 11252 4944
rect 11012 4922 11036 4924
rect 11092 4922 11116 4924
rect 11172 4922 11196 4924
rect 11034 4870 11036 4922
rect 11098 4870 11110 4922
rect 11172 4870 11174 4922
rect 11012 4868 11036 4870
rect 11092 4868 11116 4870
rect 11172 4868 11196 4870
rect 10956 4848 11252 4868
rect 11348 4826 11376 4966
rect 11440 4826 11468 5034
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11624 4690 11652 4966
rect 11716 4729 11744 7142
rect 11794 7103 11850 7112
rect 11808 4758 11836 7103
rect 11992 5778 12020 14991
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 12084 5710 12112 17031
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12360 12442 12388 13262
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12452 12442 12480 12922
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12544 12306 12572 22170
rect 13820 20256 13872 20262
rect 14936 20233 14964 23520
rect 15956 21788 16252 21808
rect 16012 21786 16036 21788
rect 16092 21786 16116 21788
rect 16172 21786 16196 21788
rect 16034 21734 16036 21786
rect 16098 21734 16110 21786
rect 16172 21734 16174 21786
rect 16012 21732 16036 21734
rect 16092 21732 16116 21734
rect 16172 21732 16196 21734
rect 15956 21712 16252 21732
rect 15956 20700 16252 20720
rect 16012 20698 16036 20700
rect 16092 20698 16116 20700
rect 16172 20698 16196 20700
rect 16034 20646 16036 20698
rect 16098 20646 16110 20698
rect 16172 20646 16174 20698
rect 16012 20644 16036 20646
rect 16092 20644 16116 20646
rect 16172 20644 16196 20646
rect 15956 20624 16252 20644
rect 18340 20505 18368 23520
rect 21456 22160 21508 22166
rect 21456 22102 21508 22108
rect 20956 21244 21252 21264
rect 21012 21242 21036 21244
rect 21092 21242 21116 21244
rect 21172 21242 21196 21244
rect 21034 21190 21036 21242
rect 21098 21190 21110 21242
rect 21172 21190 21174 21242
rect 21012 21188 21036 21190
rect 21092 21188 21116 21190
rect 21172 21188 21196 21190
rect 20956 21168 21252 21188
rect 19708 20936 19760 20942
rect 19708 20878 19760 20884
rect 16118 20496 16174 20505
rect 16118 20431 16120 20440
rect 16172 20431 16174 20440
rect 18326 20496 18382 20505
rect 19720 20466 19748 20878
rect 18326 20431 18382 20440
rect 19708 20460 19760 20466
rect 16120 20402 16172 20408
rect 19708 20402 19760 20408
rect 15844 20392 15896 20398
rect 15844 20334 15896 20340
rect 13820 20198 13872 20204
rect 14922 20224 14978 20233
rect 13832 19922 13860 20198
rect 14922 20159 14978 20168
rect 15856 19961 15884 20334
rect 20720 20324 20772 20330
rect 20720 20266 20772 20272
rect 15842 19952 15898 19961
rect 13820 19916 13872 19922
rect 15842 19887 15898 19896
rect 13820 19858 13872 19864
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 14186 19816 14242 19825
rect 12636 19242 12664 19790
rect 14186 19751 14188 19760
rect 14240 19751 14242 19760
rect 14188 19722 14240 19728
rect 16488 19712 16540 19718
rect 13910 19680 13966 19689
rect 16488 19654 16540 19660
rect 19616 19712 19668 19718
rect 19616 19654 19668 19660
rect 13910 19615 13966 19624
rect 12624 19236 12676 19242
rect 12624 19178 12676 19184
rect 12636 18630 12664 19178
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12636 18222 12664 18566
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12636 15162 12664 18158
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13266 17912 13322 17921
rect 13266 17847 13268 17856
rect 13320 17847 13322 17856
rect 13268 17818 13320 17824
rect 12716 17536 12768 17542
rect 12716 17478 12768 17484
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 12452 11558 12480 12106
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12452 11354 12480 11494
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 12162 7440 12218 7449
rect 12162 7375 12164 7384
rect 12216 7375 12218 7384
rect 12164 7346 12216 7352
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12268 6934 12296 7142
rect 12256 6928 12308 6934
rect 12256 6870 12308 6876
rect 12268 6458 12296 6870
rect 12360 6798 12388 7686
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12360 6390 12388 6734
rect 12348 6384 12400 6390
rect 12348 6326 12400 6332
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 12084 5370 12112 5646
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 11796 4752 11848 4758
rect 11702 4720 11758 4729
rect 11612 4684 11664 4690
rect 11796 4694 11848 4700
rect 11702 4655 11758 4664
rect 11612 4626 11664 4632
rect 11428 4276 11480 4282
rect 11428 4218 11480 4224
rect 10956 3836 11252 3856
rect 11012 3834 11036 3836
rect 11092 3834 11116 3836
rect 11172 3834 11196 3836
rect 11034 3782 11036 3834
rect 11098 3782 11110 3834
rect 11172 3782 11174 3834
rect 11012 3780 11036 3782
rect 11092 3780 11116 3782
rect 11172 3780 11196 3782
rect 10956 3760 11252 3780
rect 11440 3738 11468 4218
rect 11624 4078 11652 4626
rect 11808 4214 11836 4694
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11992 4282 12020 4558
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 11796 4208 11848 4214
rect 11796 4150 11848 4156
rect 11612 4072 11664 4078
rect 11610 4040 11612 4049
rect 12084 4049 12112 5306
rect 12360 4434 12388 5714
rect 12440 4480 12492 4486
rect 12360 4428 12440 4434
rect 12360 4422 12492 4428
rect 12360 4406 12480 4422
rect 11664 4040 11666 4049
rect 11610 3975 11666 3984
rect 12070 4040 12126 4049
rect 12070 3975 12126 3984
rect 11624 3949 11652 3975
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 12360 3641 12388 4406
rect 12346 3632 12402 3641
rect 12346 3567 12402 3576
rect 9954 3496 10010 3505
rect 9954 3431 10010 3440
rect 10956 2748 11252 2768
rect 11012 2746 11036 2748
rect 11092 2746 11116 2748
rect 11172 2746 11196 2748
rect 11034 2694 11036 2746
rect 11098 2694 11110 2746
rect 11172 2694 11174 2746
rect 11012 2692 11036 2694
rect 11092 2692 11116 2694
rect 11172 2692 11196 2694
rect 10956 2672 11252 2692
rect 12728 2514 12756 17478
rect 13280 17202 13308 17818
rect 13832 17762 13860 18022
rect 13740 17734 13860 17762
rect 13740 17678 13768 17734
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13372 17338 13400 17614
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 13372 16726 13400 17274
rect 13740 17270 13768 17614
rect 13820 17536 13872 17542
rect 13820 17478 13872 17484
rect 13728 17264 13780 17270
rect 13728 17206 13780 17212
rect 13452 17060 13504 17066
rect 13452 17002 13504 17008
rect 13464 16794 13492 17002
rect 13452 16788 13504 16794
rect 13452 16730 13504 16736
rect 13360 16720 13412 16726
rect 13360 16662 13412 16668
rect 13636 16720 13688 16726
rect 13636 16662 13688 16668
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12820 15473 12848 15846
rect 13280 15706 13308 16050
rect 13372 15910 13400 16526
rect 13648 16250 13676 16662
rect 13636 16244 13688 16250
rect 13636 16186 13688 16192
rect 13740 16130 13768 17206
rect 13832 16998 13860 17478
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13832 16250 13860 16934
rect 13924 16726 13952 19615
rect 15956 19612 16252 19632
rect 16012 19610 16036 19612
rect 16092 19610 16116 19612
rect 16172 19610 16196 19612
rect 16034 19558 16036 19610
rect 16098 19558 16110 19610
rect 16172 19558 16174 19610
rect 16012 19556 16036 19558
rect 16092 19556 16116 19558
rect 16172 19556 16196 19558
rect 15956 19536 16252 19556
rect 16394 19408 16450 19417
rect 16500 19394 16528 19654
rect 16450 19366 16528 19394
rect 19628 19378 19656 19654
rect 16394 19343 16450 19352
rect 15844 19236 15896 19242
rect 15844 19178 15896 19184
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 15752 19168 15804 19174
rect 15752 19110 15804 19116
rect 15212 18834 15240 19110
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 14476 17338 14504 18158
rect 15212 18086 15240 18770
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 15212 17649 15240 18022
rect 15198 17640 15254 17649
rect 15198 17575 15254 17584
rect 14464 17332 14516 17338
rect 14464 17274 14516 17280
rect 13912 16720 13964 16726
rect 13912 16662 13964 16668
rect 14464 16720 14516 16726
rect 14464 16662 14516 16668
rect 14004 16584 14056 16590
rect 14004 16526 14056 16532
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13740 16102 13860 16130
rect 13360 15904 13412 15910
rect 13360 15846 13412 15852
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 13372 15706 13400 15846
rect 13268 15700 13320 15706
rect 13268 15642 13320 15648
rect 13360 15700 13412 15706
rect 13360 15642 13412 15648
rect 13648 15609 13676 15846
rect 13634 15600 13690 15609
rect 13176 15564 13228 15570
rect 13634 15535 13636 15544
rect 13176 15506 13228 15512
rect 13688 15535 13690 15544
rect 13636 15506 13688 15512
rect 12806 15464 12862 15473
rect 12806 15399 12862 15408
rect 12808 12300 12860 12306
rect 12808 12242 12860 12248
rect 12820 11830 12848 12242
rect 12900 12232 12952 12238
rect 12898 12200 12900 12209
rect 12952 12200 12954 12209
rect 12898 12135 12954 12144
rect 12912 11898 12940 12135
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12808 11824 12860 11830
rect 12808 11766 12860 11772
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12820 9926 12848 11086
rect 12912 10810 12940 11154
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12820 9518 12848 9862
rect 13188 9722 13216 15506
rect 13832 15162 13860 16102
rect 14016 16046 14044 16526
rect 14004 16040 14056 16046
rect 14004 15982 14056 15988
rect 14016 15638 14044 15982
rect 14004 15632 14056 15638
rect 14004 15574 14056 15580
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13832 14958 13860 15098
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13728 14884 13780 14890
rect 13728 14826 13780 14832
rect 13740 14278 13768 14826
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13740 13841 13768 14214
rect 13726 13832 13782 13841
rect 13726 13767 13782 13776
rect 14188 13728 14240 13734
rect 14188 13670 14240 13676
rect 13912 13388 13964 13394
rect 13912 13330 13964 13336
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 13820 13184 13872 13190
rect 13820 13126 13872 13132
rect 13452 12640 13504 12646
rect 13450 12608 13452 12617
rect 13504 12608 13506 12617
rect 13450 12543 13506 12552
rect 13634 12336 13690 12345
rect 13832 12306 13860 13126
rect 13924 12481 13952 13330
rect 14108 13297 14136 13330
rect 14200 13326 14228 13670
rect 14188 13320 14240 13326
rect 14094 13288 14150 13297
rect 14188 13262 14240 13268
rect 14278 13288 14334 13297
rect 14094 13223 14150 13232
rect 14108 12617 14136 13223
rect 14094 12608 14150 12617
rect 14094 12543 14150 12552
rect 13910 12472 13966 12481
rect 14200 12442 14228 13262
rect 14278 13223 14334 13232
rect 14292 12714 14320 13223
rect 14280 12708 14332 12714
rect 14280 12650 14332 12656
rect 13910 12407 13966 12416
rect 14188 12436 14240 12442
rect 13924 12345 13952 12407
rect 14188 12378 14240 12384
rect 13910 12336 13966 12345
rect 13634 12271 13636 12280
rect 13688 12271 13690 12280
rect 13820 12300 13872 12306
rect 13636 12242 13688 12248
rect 13910 12271 13966 12280
rect 14096 12300 14148 12306
rect 13820 12242 13872 12248
rect 14096 12242 14148 12248
rect 13820 11688 13872 11694
rect 13740 11636 13820 11642
rect 13740 11630 13872 11636
rect 13740 11614 13860 11630
rect 13912 11620 13964 11626
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13556 10452 13584 11494
rect 13740 10810 13768 11614
rect 13912 11562 13964 11568
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13832 11218 13860 11494
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13924 10826 13952 11562
rect 14004 11552 14056 11558
rect 14004 11494 14056 11500
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13832 10798 13952 10826
rect 13832 10690 13860 10798
rect 13740 10674 13860 10690
rect 13728 10668 13860 10674
rect 13780 10662 13860 10668
rect 13728 10610 13780 10616
rect 13820 10464 13872 10470
rect 13556 10424 13820 10452
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13464 9518 13492 9658
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 13452 9512 13504 9518
rect 13452 9454 13504 9460
rect 12820 8838 12848 9454
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12806 7440 12862 7449
rect 12806 7375 12862 7384
rect 12820 7206 12848 7375
rect 12912 7274 12940 9454
rect 13556 9450 13584 10424
rect 13820 10406 13872 10412
rect 14016 10130 14044 11494
rect 14108 10810 14136 12242
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14200 11014 14228 11698
rect 14292 11694 14320 12038
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14384 11626 14412 12038
rect 14372 11620 14424 11626
rect 14372 11562 14424 11568
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 14200 10674 14228 10950
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 14200 10470 14228 10610
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 13636 9920 13688 9926
rect 13636 9862 13688 9868
rect 13544 9444 13596 9450
rect 13544 9386 13596 9392
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 13280 8634 13308 8774
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 12900 7268 12952 7274
rect 12900 7210 12952 7216
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 13096 7002 13124 7346
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 13096 6730 13124 6938
rect 13084 6724 13136 6730
rect 13084 6666 13136 6672
rect 13280 6338 13308 8570
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13372 7002 13400 7822
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13450 6760 13506 6769
rect 13450 6695 13506 6704
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13372 6458 13400 6598
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13280 6310 13400 6338
rect 13372 5574 13400 6310
rect 12900 5568 12952 5574
rect 12900 5510 12952 5516
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 12912 5098 12940 5510
rect 13372 5166 13400 5510
rect 13360 5160 13412 5166
rect 13360 5102 13412 5108
rect 12900 5092 12952 5098
rect 12900 5034 12952 5040
rect 12912 4622 12940 5034
rect 13266 4856 13322 4865
rect 13464 4826 13492 6695
rect 13266 4791 13268 4800
rect 13320 4791 13322 4800
rect 13452 4820 13504 4826
rect 13268 4762 13320 4768
rect 13452 4762 13504 4768
rect 12900 4616 12952 4622
rect 12900 4558 12952 4564
rect 13280 4282 13308 4762
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 13280 4185 13308 4218
rect 13464 4214 13492 4762
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13556 4282 13584 4558
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 13452 4208 13504 4214
rect 13266 4176 13322 4185
rect 13452 4150 13504 4156
rect 13266 4111 13322 4120
rect 13648 3194 13676 9862
rect 13740 9178 13768 10066
rect 14108 9178 14136 10202
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14200 9722 14228 9998
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 14476 8129 14504 16662
rect 15212 15978 15240 17575
rect 15304 17542 15332 18702
rect 15764 18193 15792 19110
rect 15856 18290 15884 19178
rect 16500 19174 16528 19366
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 16488 19168 16540 19174
rect 16488 19110 16540 19116
rect 16856 19168 16908 19174
rect 16856 19110 16908 19116
rect 16672 18624 16724 18630
rect 16672 18566 16724 18572
rect 15956 18524 16252 18544
rect 16012 18522 16036 18524
rect 16092 18522 16116 18524
rect 16172 18522 16196 18524
rect 16034 18470 16036 18522
rect 16098 18470 16110 18522
rect 16172 18470 16174 18522
rect 16012 18468 16036 18470
rect 16092 18468 16116 18470
rect 16172 18468 16196 18470
rect 15956 18448 16252 18468
rect 16684 18290 16712 18566
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 16672 18284 16724 18290
rect 16672 18226 16724 18232
rect 15750 18184 15806 18193
rect 15750 18119 15806 18128
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 15396 17921 15424 18022
rect 15382 17912 15438 17921
rect 16224 17882 16252 18022
rect 15382 17847 15438 17856
rect 16212 17876 16264 17882
rect 16212 17818 16264 17824
rect 16672 17808 16724 17814
rect 16670 17776 16672 17785
rect 16724 17776 16726 17785
rect 16670 17711 16726 17720
rect 16396 17604 16448 17610
rect 16396 17546 16448 17552
rect 15292 17536 15344 17542
rect 16304 17536 16356 17542
rect 15292 17478 15344 17484
rect 15750 17504 15806 17513
rect 16304 17478 16356 17484
rect 15750 17439 15806 17448
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15396 16561 15424 16934
rect 15382 16552 15438 16561
rect 15382 16487 15438 16496
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 15396 16046 15424 16390
rect 15488 16114 15516 16934
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 15200 15972 15252 15978
rect 15200 15914 15252 15920
rect 15396 15706 15424 15982
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 15488 15638 15516 16050
rect 15764 15881 15792 17439
rect 15956 17436 16252 17456
rect 16012 17434 16036 17436
rect 16092 17434 16116 17436
rect 16172 17434 16196 17436
rect 16034 17382 16036 17434
rect 16098 17382 16110 17434
rect 16172 17382 16174 17434
rect 16012 17380 16036 17382
rect 16092 17380 16116 17382
rect 16172 17380 16196 17382
rect 15956 17360 16252 17380
rect 15844 16992 15896 16998
rect 15844 16934 15896 16940
rect 15856 16658 15884 16934
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 16212 16652 16264 16658
rect 16212 16594 16264 16600
rect 15856 16454 15884 16594
rect 16224 16538 16252 16594
rect 16316 16538 16344 17478
rect 16408 17202 16436 17546
rect 16684 17338 16712 17711
rect 16764 17672 16816 17678
rect 16762 17640 16764 17649
rect 16816 17640 16818 17649
rect 16762 17575 16818 17584
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16776 17270 16804 17575
rect 16764 17264 16816 17270
rect 16764 17206 16816 17212
rect 16396 17196 16448 17202
rect 16396 17138 16448 17144
rect 16408 16658 16436 17138
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 16224 16510 16344 16538
rect 15844 16448 15896 16454
rect 15844 16390 15896 16396
rect 15956 16348 16252 16368
rect 16012 16346 16036 16348
rect 16092 16346 16116 16348
rect 16172 16346 16196 16348
rect 16034 16294 16036 16346
rect 16098 16294 16110 16346
rect 16172 16294 16174 16346
rect 16012 16292 16036 16294
rect 16092 16292 16116 16294
rect 16172 16292 16196 16294
rect 15956 16272 16252 16292
rect 16120 16176 16172 16182
rect 16120 16118 16172 16124
rect 16026 16008 16082 16017
rect 16026 15943 16082 15952
rect 15750 15872 15806 15881
rect 15750 15807 15806 15816
rect 15764 15706 15792 15807
rect 16040 15706 16068 15943
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 16028 15700 16080 15706
rect 16028 15642 16080 15648
rect 15476 15632 15528 15638
rect 15476 15574 15528 15580
rect 15764 15162 15792 15642
rect 16040 15450 16068 15642
rect 16132 15502 16160 16118
rect 16316 15910 16344 16510
rect 16408 16182 16436 16594
rect 16396 16176 16448 16182
rect 16396 16118 16448 16124
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 15856 15422 16068 15450
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 16304 15496 16356 15502
rect 16304 15438 16356 15444
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15856 15094 15884 15422
rect 15956 15260 16252 15280
rect 16012 15258 16036 15260
rect 16092 15258 16116 15260
rect 16172 15258 16196 15260
rect 16034 15206 16036 15258
rect 16098 15206 16110 15258
rect 16172 15206 16174 15258
rect 16012 15204 16036 15206
rect 16092 15204 16116 15206
rect 16172 15204 16196 15206
rect 15956 15184 16252 15204
rect 16316 15162 16344 15438
rect 16304 15156 16356 15162
rect 16304 15098 16356 15104
rect 15292 15088 15344 15094
rect 15292 15030 15344 15036
rect 15844 15088 15896 15094
rect 15844 15030 15896 15036
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 14936 13802 14964 14758
rect 15200 14544 15252 14550
rect 15200 14486 15252 14492
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 15014 13832 15070 13841
rect 14924 13796 14976 13802
rect 15014 13767 15070 13776
rect 14924 13738 14976 13744
rect 14830 13696 14886 13705
rect 14830 13631 14886 13640
rect 14844 12986 14872 13631
rect 15028 13530 15056 13767
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 14832 12980 14884 12986
rect 14832 12922 14884 12928
rect 15120 12306 15148 14214
rect 15212 13870 15240 14486
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15212 13569 15240 13806
rect 15198 13560 15254 13569
rect 15198 13495 15254 13504
rect 15212 13161 15240 13495
rect 15198 13152 15254 13161
rect 15198 13087 15254 13096
rect 15304 13002 15332 15030
rect 16304 14476 16356 14482
rect 16304 14418 16356 14424
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15384 13864 15436 13870
rect 15382 13832 15384 13841
rect 15436 13832 15438 13841
rect 15856 13802 15884 14350
rect 15956 14172 16252 14192
rect 16012 14170 16036 14172
rect 16092 14170 16116 14172
rect 16172 14170 16196 14172
rect 16034 14118 16036 14170
rect 16098 14118 16110 14170
rect 16172 14118 16174 14170
rect 16012 14116 16036 14118
rect 16092 14116 16116 14118
rect 16172 14116 16196 14118
rect 15956 14096 16252 14116
rect 16316 14074 16344 14418
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 15382 13767 15438 13776
rect 15844 13796 15896 13802
rect 15844 13738 15896 13744
rect 15752 13456 15804 13462
rect 15752 13398 15804 13404
rect 15660 13184 15712 13190
rect 15660 13126 15712 13132
rect 15212 12974 15332 13002
rect 15568 12980 15620 12986
rect 15108 12300 15160 12306
rect 15108 12242 15160 12248
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 14568 11354 14596 12174
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14936 11218 14964 12174
rect 14924 11212 14976 11218
rect 14924 11154 14976 11160
rect 15108 11008 15160 11014
rect 15108 10950 15160 10956
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14568 10266 14596 10406
rect 14752 10266 14780 10542
rect 15120 10538 15148 10950
rect 15108 10532 15160 10538
rect 15108 10474 15160 10480
rect 15120 10266 15148 10474
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 15016 9512 15068 9518
rect 15016 9454 15068 9460
rect 15028 9042 15056 9454
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14462 8120 14518 8129
rect 14462 8055 14518 8064
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 14660 7002 14688 7346
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 13726 6896 13782 6905
rect 13726 6831 13728 6840
rect 13780 6831 13782 6840
rect 13728 6802 13780 6808
rect 13740 6390 13768 6802
rect 13832 6458 13860 6938
rect 14004 6792 14056 6798
rect 14004 6734 14056 6740
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13728 6384 13780 6390
rect 13728 6326 13780 6332
rect 14016 6118 14044 6734
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 14016 5370 14044 6054
rect 14004 5364 14056 5370
rect 14004 5306 14056 5312
rect 14660 5234 14688 6938
rect 14648 5228 14700 5234
rect 14648 5170 14700 5176
rect 14660 4826 14688 5170
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14936 4729 14964 8366
rect 15028 7546 15056 8978
rect 15212 8362 15240 12974
rect 15568 12922 15620 12928
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15396 11665 15424 11834
rect 15382 11656 15438 11665
rect 15292 11620 15344 11626
rect 15382 11591 15438 11600
rect 15292 11562 15344 11568
rect 15304 9489 15332 11562
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15396 10606 15424 11494
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15488 10266 15516 11154
rect 15580 10713 15608 12922
rect 15672 12866 15700 13126
rect 15764 12986 15792 13398
rect 15856 13326 15884 13738
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15856 12986 15884 13262
rect 15956 13084 16252 13104
rect 16012 13082 16036 13084
rect 16092 13082 16116 13084
rect 16172 13082 16196 13084
rect 16034 13030 16036 13082
rect 16098 13030 16110 13082
rect 16172 13030 16174 13082
rect 16012 13028 16036 13030
rect 16092 13028 16116 13030
rect 16172 13028 16196 13030
rect 15956 13008 16252 13028
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15672 12838 15792 12866
rect 15660 12776 15712 12782
rect 15660 12718 15712 12724
rect 15566 10704 15622 10713
rect 15566 10639 15622 10648
rect 15476 10260 15528 10266
rect 15476 10202 15528 10208
rect 15290 9480 15346 9489
rect 15290 9415 15346 9424
rect 15200 8356 15252 8362
rect 15200 8298 15252 8304
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 15580 6225 15608 10639
rect 15672 9081 15700 12718
rect 15764 12306 15792 12838
rect 15844 12368 15896 12374
rect 15842 12336 15844 12345
rect 15896 12336 15898 12345
rect 15752 12300 15804 12306
rect 15842 12271 15898 12280
rect 15752 12242 15804 12248
rect 15856 11898 15884 12271
rect 15956 11996 16252 12016
rect 16012 11994 16036 11996
rect 16092 11994 16116 11996
rect 16172 11994 16196 11996
rect 16034 11942 16036 11994
rect 16098 11942 16110 11994
rect 16172 11942 16174 11994
rect 16012 11940 16036 11942
rect 16092 11940 16116 11942
rect 16172 11940 16196 11942
rect 15956 11920 16252 11940
rect 15844 11892 15896 11898
rect 15844 11834 15896 11840
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 15936 11280 15988 11286
rect 15856 11257 15936 11268
rect 15842 11248 15936 11257
rect 15752 11212 15804 11218
rect 15898 11240 15936 11248
rect 15936 11222 15988 11228
rect 15842 11183 15898 11192
rect 15752 11154 15804 11160
rect 15764 10810 15792 11154
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 15856 10742 15884 11183
rect 16132 11150 16160 11698
rect 16316 11529 16344 14010
rect 16580 14000 16632 14006
rect 16580 13942 16632 13948
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16408 13161 16436 13330
rect 16394 13152 16450 13161
rect 16394 13087 16450 13096
rect 16408 12918 16436 13087
rect 16396 12912 16448 12918
rect 16396 12854 16448 12860
rect 16592 12238 16620 13942
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16408 11665 16436 12038
rect 16672 11824 16724 11830
rect 16670 11792 16672 11801
rect 16724 11792 16726 11801
rect 16670 11727 16726 11736
rect 16394 11656 16450 11665
rect 16394 11591 16396 11600
rect 16448 11591 16450 11600
rect 16396 11562 16448 11568
rect 16408 11531 16436 11562
rect 16302 11520 16358 11529
rect 16302 11455 16358 11464
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 15956 10908 16252 10928
rect 16012 10906 16036 10908
rect 16092 10906 16116 10908
rect 16172 10906 16196 10908
rect 16034 10854 16036 10906
rect 16098 10854 16110 10906
rect 16172 10854 16174 10906
rect 16012 10852 16036 10854
rect 16092 10852 16116 10854
rect 16172 10852 16196 10854
rect 15956 10832 16252 10852
rect 15844 10736 15896 10742
rect 15844 10678 15896 10684
rect 15956 9820 16252 9840
rect 16012 9818 16036 9820
rect 16092 9818 16116 9820
rect 16172 9818 16196 9820
rect 16034 9766 16036 9818
rect 16098 9766 16110 9818
rect 16172 9766 16174 9818
rect 16012 9764 16036 9766
rect 16092 9764 16116 9766
rect 16172 9764 16196 9766
rect 15956 9744 16252 9764
rect 16868 9722 16896 19110
rect 18878 18864 18934 18873
rect 18878 18799 18934 18808
rect 18892 18426 18920 18799
rect 18880 18420 18932 18426
rect 18880 18362 18932 18368
rect 19340 18216 19392 18222
rect 19338 18184 19340 18193
rect 19392 18184 19394 18193
rect 18604 18148 18656 18154
rect 19338 18119 19394 18128
rect 18604 18090 18656 18096
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 16960 17746 16988 18022
rect 16948 17740 17000 17746
rect 16948 17682 17000 17688
rect 16960 17338 16988 17682
rect 16948 17332 17000 17338
rect 16948 17274 17000 17280
rect 17500 17264 17552 17270
rect 17500 17206 17552 17212
rect 18236 17264 18288 17270
rect 18236 17206 18288 17212
rect 17512 16794 17540 17206
rect 17500 16788 17552 16794
rect 17500 16730 17552 16736
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17788 15366 17816 15846
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17776 15360 17828 15366
rect 17776 15302 17828 15308
rect 17788 15026 17816 15302
rect 17972 15178 18000 15506
rect 17880 15162 18000 15178
rect 17868 15156 18000 15162
rect 17920 15150 18000 15156
rect 17868 15098 17920 15104
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 17776 15020 17828 15026
rect 17776 14962 17828 14968
rect 17788 13841 17816 14962
rect 17774 13832 17830 13841
rect 17774 13767 17830 13776
rect 17788 13394 17816 13767
rect 17776 13388 17828 13394
rect 17776 13330 17828 13336
rect 17314 12880 17370 12889
rect 17314 12815 17370 12824
rect 17328 12306 17356 12815
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17420 12442 17448 12582
rect 17788 12442 17816 13330
rect 17972 12730 18000 15030
rect 18144 14476 18196 14482
rect 18144 14418 18196 14424
rect 18156 13734 18184 14418
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 18156 13530 18184 13670
rect 18144 13524 18196 13530
rect 18144 13466 18196 13472
rect 18052 13388 18104 13394
rect 18052 13330 18104 13336
rect 18064 12850 18092 13330
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 17972 12702 18092 12730
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 17776 12436 17828 12442
rect 17776 12378 17828 12384
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 17052 11354 17080 12242
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 17144 11898 17172 12174
rect 17420 11898 17448 12378
rect 17684 12096 17736 12102
rect 17684 12038 17736 12044
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 15658 9072 15714 9081
rect 15658 9007 15714 9016
rect 16210 8936 16266 8945
rect 16316 8922 16344 9522
rect 16396 9376 16448 9382
rect 16396 9318 16448 9324
rect 16408 9110 16436 9318
rect 16396 9104 16448 9110
rect 16396 9046 16448 9052
rect 17408 9104 17460 9110
rect 17408 9046 17460 9052
rect 16266 8894 16344 8922
rect 16210 8871 16266 8880
rect 15956 8732 16252 8752
rect 16012 8730 16036 8732
rect 16092 8730 16116 8732
rect 16172 8730 16196 8732
rect 16034 8678 16036 8730
rect 16098 8678 16110 8730
rect 16172 8678 16174 8730
rect 16012 8676 16036 8678
rect 16092 8676 16116 8678
rect 16172 8676 16196 8678
rect 15956 8656 16252 8676
rect 16316 8537 16344 8894
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16302 8528 16358 8537
rect 16500 8498 16528 8774
rect 17420 8634 17448 9046
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 16302 8463 16358 8472
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16304 8356 16356 8362
rect 16304 8298 16356 8304
rect 15956 7644 16252 7664
rect 16012 7642 16036 7644
rect 16092 7642 16116 7644
rect 16172 7642 16196 7644
rect 16034 7590 16036 7642
rect 16098 7590 16110 7642
rect 16172 7590 16174 7642
rect 16012 7588 16036 7590
rect 16092 7588 16116 7590
rect 16172 7588 16196 7590
rect 15956 7568 16252 7588
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 15856 6254 15884 7142
rect 16316 6769 16344 8298
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16408 6866 16436 8230
rect 16592 8106 16620 8366
rect 16500 8090 16620 8106
rect 16868 8090 16896 8434
rect 17420 8344 17448 8570
rect 17420 8316 17540 8344
rect 16488 8084 16620 8090
rect 16540 8078 16620 8084
rect 16856 8084 16908 8090
rect 16488 8026 16540 8032
rect 16856 8026 16908 8032
rect 16500 7342 16528 8026
rect 17406 7984 17462 7993
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 17316 7948 17368 7954
rect 17406 7919 17462 7928
rect 17316 7890 17368 7896
rect 16960 7585 16988 7890
rect 16946 7576 17002 7585
rect 16946 7511 17002 7520
rect 16488 7336 16540 7342
rect 16488 7278 16540 7284
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 16302 6760 16358 6769
rect 16302 6695 16358 6704
rect 15956 6556 16252 6576
rect 16012 6554 16036 6556
rect 16092 6554 16116 6556
rect 16172 6554 16196 6556
rect 16034 6502 16036 6554
rect 16098 6502 16110 6554
rect 16172 6502 16174 6554
rect 16012 6500 16036 6502
rect 16092 6500 16116 6502
rect 16172 6500 16196 6502
rect 15956 6480 16252 6500
rect 16408 6322 16436 6802
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 15844 6248 15896 6254
rect 15566 6216 15622 6225
rect 15844 6190 15896 6196
rect 15566 6151 15622 6160
rect 15200 6112 15252 6118
rect 15120 6060 15200 6066
rect 15120 6054 15252 6060
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 15120 6038 15240 6054
rect 15120 5098 15148 6038
rect 16132 5914 16160 6054
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15108 5092 15160 5098
rect 15108 5034 15160 5040
rect 14922 4720 14978 4729
rect 14922 4655 14978 4664
rect 15488 3194 15516 5510
rect 15856 4826 15884 5850
rect 16488 5772 16540 5778
rect 16592 5760 16620 6598
rect 16540 5732 16620 5760
rect 16488 5714 16540 5720
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 15956 5468 16252 5488
rect 16012 5466 16036 5468
rect 16092 5466 16116 5468
rect 16172 5466 16196 5468
rect 16034 5414 16036 5466
rect 16098 5414 16110 5466
rect 16172 5414 16174 5466
rect 16012 5412 16036 5414
rect 16092 5412 16116 5414
rect 16172 5412 16196 5414
rect 15956 5392 16252 5412
rect 16316 5370 16344 5646
rect 16592 5370 16620 5732
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 16316 4758 16344 5306
rect 16684 5030 16712 7210
rect 16960 7206 16988 7511
rect 17328 7274 17356 7890
rect 17316 7268 17368 7274
rect 17316 7210 17368 7216
rect 16948 7200 17000 7206
rect 16946 7168 16948 7177
rect 17420 7177 17448 7919
rect 17512 7886 17540 8316
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 17512 7546 17540 7822
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17000 7168 17002 7177
rect 16946 7103 17002 7112
rect 17406 7168 17462 7177
rect 17406 7103 17462 7112
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 16856 6724 16908 6730
rect 16856 6666 16908 6672
rect 16868 5914 16896 6666
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16960 5846 16988 6802
rect 17132 6792 17184 6798
rect 17132 6734 17184 6740
rect 17144 6254 17172 6734
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17040 6180 17092 6186
rect 17040 6122 17092 6128
rect 17052 5914 17080 6122
rect 17420 5914 17448 7103
rect 17592 6384 17644 6390
rect 17592 6326 17644 6332
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 16948 5840 17000 5846
rect 16948 5782 17000 5788
rect 17420 5302 17448 5850
rect 17604 5710 17632 6326
rect 17500 5704 17552 5710
rect 17498 5672 17500 5681
rect 17592 5704 17644 5710
rect 17552 5672 17554 5681
rect 17592 5646 17644 5652
rect 17696 5658 17724 12038
rect 17868 9036 17920 9042
rect 17868 8978 17920 8984
rect 17880 8673 17908 8978
rect 17866 8664 17922 8673
rect 17866 8599 17868 8608
rect 17920 8599 17922 8608
rect 17868 8570 17920 8576
rect 18064 8022 18092 12702
rect 18156 12238 18184 13466
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 18052 8016 18104 8022
rect 18052 7958 18104 7964
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 18064 7313 18092 7686
rect 18050 7304 18106 7313
rect 18106 7274 18184 7290
rect 18106 7268 18196 7274
rect 18106 7262 18144 7268
rect 18050 7239 18106 7248
rect 18144 7210 18196 7216
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17880 6866 17908 7142
rect 17868 6860 17920 6866
rect 17868 6802 17920 6808
rect 17498 5607 17554 5616
rect 17512 5370 17540 5607
rect 17604 5370 17632 5646
rect 17696 5630 18000 5658
rect 17500 5364 17552 5370
rect 17500 5306 17552 5312
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17408 5296 17460 5302
rect 17408 5238 17460 5244
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 17512 4865 17540 5306
rect 17498 4856 17554 4865
rect 17498 4791 17554 4800
rect 16304 4752 16356 4758
rect 16304 4694 16356 4700
rect 16396 4752 16448 4758
rect 16396 4694 16448 4700
rect 15956 4380 16252 4400
rect 16012 4378 16036 4380
rect 16092 4378 16116 4380
rect 16172 4378 16196 4380
rect 16034 4326 16036 4378
rect 16098 4326 16110 4378
rect 16172 4326 16174 4378
rect 16012 4324 16036 4326
rect 16092 4324 16116 4326
rect 16172 4324 16196 4326
rect 15956 4304 16252 4324
rect 16316 4214 16344 4694
rect 16408 4282 16436 4694
rect 17776 4480 17828 4486
rect 17776 4422 17828 4428
rect 17788 4282 17816 4422
rect 16396 4276 16448 4282
rect 16396 4218 16448 4224
rect 17776 4276 17828 4282
rect 17776 4218 17828 4224
rect 16304 4208 16356 4214
rect 15658 4176 15714 4185
rect 16304 4150 16356 4156
rect 15658 4111 15714 4120
rect 15672 3602 15700 4111
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 15672 3194 15700 3538
rect 16304 3528 16356 3534
rect 17328 3505 17356 3538
rect 16304 3470 16356 3476
rect 17314 3496 17370 3505
rect 15956 3292 16252 3312
rect 16012 3290 16036 3292
rect 16092 3290 16116 3292
rect 16172 3290 16196 3292
rect 16034 3238 16036 3290
rect 16098 3238 16110 3290
rect 16172 3238 16174 3290
rect 16012 3236 16036 3238
rect 16092 3236 16116 3238
rect 16172 3236 16196 3238
rect 15956 3216 16252 3236
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 13648 2990 13676 3130
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 13452 2916 13504 2922
rect 13452 2858 13504 2864
rect 14924 2916 14976 2922
rect 14924 2858 14976 2864
rect 8116 2508 8168 2514
rect 8116 2450 8168 2456
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 12716 2508 12768 2514
rect 12716 2450 12768 2456
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 12072 2440 12124 2446
rect 12072 2382 12124 2388
rect 9232 480 9260 2382
rect 10612 480 10640 2382
rect 12084 480 12112 2382
rect 13464 480 13492 2858
rect 14936 480 14964 2858
rect 15956 2204 16252 2224
rect 16012 2202 16036 2204
rect 16092 2202 16116 2204
rect 16172 2202 16196 2204
rect 16034 2150 16036 2202
rect 16098 2150 16110 2202
rect 16172 2150 16174 2202
rect 16012 2148 16036 2150
rect 16092 2148 16116 2150
rect 16172 2148 16196 2150
rect 15956 2128 16252 2148
rect 16316 480 16344 3470
rect 17314 3431 17370 3440
rect 17328 3194 17356 3431
rect 17316 3188 17368 3194
rect 17316 3130 17368 3136
rect 16854 2680 16910 2689
rect 17788 2650 17816 4218
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17880 3126 17908 3470
rect 17868 3120 17920 3126
rect 17866 3088 17868 3097
rect 17920 3088 17922 3097
rect 17866 3023 17922 3032
rect 17972 2990 18000 5630
rect 18052 4684 18104 4690
rect 18052 4626 18104 4632
rect 18064 4078 18092 4626
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 16854 2615 16856 2624
rect 16908 2615 16910 2624
rect 17776 2644 17828 2650
rect 16856 2586 16908 2592
rect 17776 2586 17828 2592
rect 18248 2514 18276 17206
rect 18328 16992 18380 16998
rect 18328 16934 18380 16940
rect 18340 16794 18368 16934
rect 18328 16788 18380 16794
rect 18328 16730 18380 16736
rect 18616 16250 18644 18090
rect 19524 17536 19576 17542
rect 19524 17478 19576 17484
rect 19338 17232 19394 17241
rect 19338 17167 19394 17176
rect 18788 16448 18840 16454
rect 18788 16390 18840 16396
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 18800 15484 18828 16390
rect 19352 16182 19380 17167
rect 19536 17134 19564 17478
rect 19628 17218 19656 19314
rect 20732 19310 20760 20266
rect 20812 20256 20864 20262
rect 20810 20224 20812 20233
rect 20864 20224 20866 20233
rect 20810 20159 20866 20168
rect 20824 19922 20852 20159
rect 20956 20156 21252 20176
rect 21012 20154 21036 20156
rect 21092 20154 21116 20156
rect 21172 20154 21196 20156
rect 21034 20102 21036 20154
rect 21098 20102 21110 20154
rect 21172 20102 21174 20154
rect 21012 20100 21036 20102
rect 21092 20100 21116 20102
rect 21172 20100 21196 20102
rect 20956 20080 21252 20100
rect 20812 19916 20864 19922
rect 20812 19858 20864 19864
rect 20824 19514 20852 19858
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20720 19304 20772 19310
rect 20720 19246 20772 19252
rect 19984 19236 20036 19242
rect 19984 19178 20036 19184
rect 19996 18290 20024 19178
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 20956 19068 21252 19088
rect 21012 19066 21036 19068
rect 21092 19066 21116 19068
rect 21172 19066 21196 19068
rect 21034 19014 21036 19066
rect 21098 19014 21110 19066
rect 21172 19014 21174 19066
rect 21012 19012 21036 19014
rect 21092 19012 21116 19014
rect 21172 19012 21196 19014
rect 20956 18992 21252 19012
rect 20444 18760 20496 18766
rect 20444 18702 20496 18708
rect 20456 18426 20484 18702
rect 20444 18420 20496 18426
rect 20444 18362 20496 18368
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 20456 18222 20484 18362
rect 20720 18352 20772 18358
rect 20720 18294 20772 18300
rect 20444 18216 20496 18222
rect 20444 18158 20496 18164
rect 19708 18080 19760 18086
rect 19708 18022 19760 18028
rect 19720 17882 19748 18022
rect 19708 17876 19760 17882
rect 19708 17818 19760 17824
rect 19720 17338 19748 17818
rect 20732 17762 20760 18294
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20824 17882 20852 18226
rect 20956 17980 21252 18000
rect 21012 17978 21036 17980
rect 21092 17978 21116 17980
rect 21172 17978 21196 17980
rect 21034 17926 21036 17978
rect 21098 17926 21110 17978
rect 21172 17926 21174 17978
rect 21012 17924 21036 17926
rect 21092 17924 21116 17926
rect 21172 17924 21196 17926
rect 20956 17904 21252 17924
rect 20812 17876 20864 17882
rect 20812 17818 20864 17824
rect 20640 17746 20760 17762
rect 20628 17740 20760 17746
rect 20680 17734 20760 17740
rect 20628 17682 20680 17688
rect 19800 17672 19852 17678
rect 19800 17614 19852 17620
rect 19708 17332 19760 17338
rect 19708 17274 19760 17280
rect 19628 17190 19748 17218
rect 19524 17128 19576 17134
rect 19524 17070 19576 17076
rect 19616 16992 19668 16998
rect 19616 16934 19668 16940
rect 19628 16794 19656 16934
rect 19616 16788 19668 16794
rect 19616 16730 19668 16736
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 19340 16176 19392 16182
rect 19154 16144 19210 16153
rect 19340 16118 19392 16124
rect 19154 16079 19210 16088
rect 18880 15904 18932 15910
rect 18878 15872 18880 15881
rect 18932 15872 18934 15881
rect 18878 15807 18934 15816
rect 19168 15722 19196 16079
rect 19444 15910 19472 16594
rect 19614 16008 19670 16017
rect 19614 15943 19670 15952
rect 19628 15910 19656 15943
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 19616 15904 19668 15910
rect 19616 15846 19668 15852
rect 19168 15694 19380 15722
rect 19444 15706 19472 15846
rect 18880 15496 18932 15502
rect 18800 15456 18880 15484
rect 18880 15438 18932 15444
rect 18892 15162 18920 15438
rect 19168 15162 19196 15694
rect 19352 15586 19380 15694
rect 19432 15700 19484 15706
rect 19432 15642 19484 15648
rect 19524 15700 19576 15706
rect 19524 15642 19576 15648
rect 19536 15586 19564 15642
rect 19248 15564 19300 15570
rect 19352 15558 19564 15586
rect 19616 15564 19668 15570
rect 19248 15506 19300 15512
rect 19616 15506 19668 15512
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 19156 15156 19208 15162
rect 19156 15098 19208 15104
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 18788 14272 18840 14278
rect 18892 14226 18920 14962
rect 18840 14220 18920 14226
rect 18788 14214 18920 14220
rect 18800 14198 18920 14214
rect 18892 14074 18920 14198
rect 19260 14074 19288 15506
rect 19628 15473 19656 15506
rect 19614 15464 19670 15473
rect 19614 15399 19670 15408
rect 19720 15162 19748 17190
rect 19812 17066 19840 17614
rect 20628 17264 20680 17270
rect 20732 17252 20760 17734
rect 21284 17678 21312 19110
rect 21468 18442 21496 22102
rect 21652 20058 21680 23520
rect 24964 23474 24992 23520
rect 24964 23446 25268 23474
rect 25134 22400 25190 22409
rect 25134 22335 25190 22344
rect 22376 21004 22428 21010
rect 22376 20946 22428 20952
rect 22284 20936 22336 20942
rect 22284 20878 22336 20884
rect 22296 20534 22324 20878
rect 22388 20602 22416 20946
rect 22652 20800 22704 20806
rect 22652 20742 22704 20748
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 22284 20528 22336 20534
rect 22284 20470 22336 20476
rect 21730 20088 21786 20097
rect 21640 20052 21692 20058
rect 21730 20023 21786 20032
rect 21640 19994 21692 20000
rect 21744 19394 21772 20023
rect 22296 19922 22324 20470
rect 22284 19916 22336 19922
rect 22284 19858 22336 19864
rect 22100 19712 22152 19718
rect 22100 19654 22152 19660
rect 21376 18414 21496 18442
rect 21652 19366 21772 19394
rect 21376 18086 21404 18414
rect 21364 18080 21416 18086
rect 21364 18022 21416 18028
rect 21376 17785 21404 18022
rect 21362 17776 21418 17785
rect 21362 17711 21418 17720
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21284 17270 21312 17614
rect 20680 17224 20760 17252
rect 21272 17264 21324 17270
rect 20628 17206 20680 17212
rect 21272 17206 21324 17212
rect 21364 17128 21416 17134
rect 21364 17070 21416 17076
rect 19800 17060 19852 17066
rect 19800 17002 19852 17008
rect 19812 16590 19840 17002
rect 20956 16892 21252 16912
rect 21012 16890 21036 16892
rect 21092 16890 21116 16892
rect 21172 16890 21196 16892
rect 21034 16838 21036 16890
rect 21098 16838 21110 16890
rect 21172 16838 21174 16890
rect 21012 16836 21036 16838
rect 21092 16836 21116 16838
rect 21172 16836 21196 16838
rect 20956 16816 21252 16836
rect 21376 16794 21404 17070
rect 21364 16788 21416 16794
rect 21364 16730 21416 16736
rect 19800 16584 19852 16590
rect 19800 16526 19852 16532
rect 20996 16584 21048 16590
rect 20996 16526 21048 16532
rect 19812 15638 19840 16526
rect 21008 16250 21036 16526
rect 20996 16244 21048 16250
rect 20996 16186 21048 16192
rect 20720 16108 20772 16114
rect 20720 16050 20772 16056
rect 20074 16008 20130 16017
rect 19892 15972 19944 15978
rect 20074 15943 20130 15952
rect 19892 15914 19944 15920
rect 19800 15632 19852 15638
rect 19800 15574 19852 15580
rect 19800 15496 19852 15502
rect 19800 15438 19852 15444
rect 19708 15156 19760 15162
rect 19708 15098 19760 15104
rect 19812 14890 19840 15438
rect 19904 15337 19932 15914
rect 19890 15328 19946 15337
rect 19890 15263 19946 15272
rect 19800 14884 19852 14890
rect 19800 14826 19852 14832
rect 19812 14618 19840 14826
rect 19800 14612 19852 14618
rect 19800 14554 19852 14560
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19708 13864 19760 13870
rect 19708 13806 19760 13812
rect 19720 13705 19748 13806
rect 18694 13696 18750 13705
rect 18694 13631 18750 13640
rect 19706 13696 19762 13705
rect 19706 13631 19762 13640
rect 18512 12708 18564 12714
rect 18512 12650 18564 12656
rect 18524 12442 18552 12650
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18512 12436 18564 12442
rect 18512 12378 18564 12384
rect 18420 12368 18472 12374
rect 18418 12336 18420 12345
rect 18472 12336 18474 12345
rect 18418 12271 18474 12280
rect 18432 11558 18460 12271
rect 18616 11898 18644 12582
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18420 11552 18472 11558
rect 18420 11494 18472 11500
rect 18512 11552 18564 11558
rect 18512 11494 18564 11500
rect 18432 10713 18460 11494
rect 18524 11014 18552 11494
rect 18512 11008 18564 11014
rect 18512 10950 18564 10956
rect 18418 10704 18474 10713
rect 18418 10639 18474 10648
rect 18418 10568 18474 10577
rect 18418 10503 18420 10512
rect 18472 10503 18474 10512
rect 18420 10474 18472 10480
rect 18524 10266 18552 10950
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 18708 10130 18736 13631
rect 19706 13424 19762 13433
rect 19706 13359 19762 13368
rect 18786 13016 18842 13025
rect 18786 12951 18842 12960
rect 18800 12850 18828 12951
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 19616 12708 19668 12714
rect 19616 12650 19668 12656
rect 18972 12232 19024 12238
rect 18972 12174 19024 12180
rect 19156 12232 19208 12238
rect 19156 12174 19208 12180
rect 18984 11354 19012 12174
rect 19168 11762 19196 12174
rect 19628 11830 19656 12650
rect 19720 12481 19748 13359
rect 19706 12472 19762 12481
rect 19706 12407 19762 12416
rect 19616 11824 19668 11830
rect 19616 11766 19668 11772
rect 19156 11756 19208 11762
rect 19156 11698 19208 11704
rect 19064 11620 19116 11626
rect 19064 11562 19116 11568
rect 18972 11348 19024 11354
rect 18972 11290 19024 11296
rect 19076 10810 19104 11562
rect 19338 11520 19394 11529
rect 19338 11455 19394 11464
rect 19352 11121 19380 11455
rect 19524 11144 19576 11150
rect 19338 11112 19394 11121
rect 19524 11086 19576 11092
rect 19338 11047 19394 11056
rect 19064 10804 19116 10810
rect 19064 10746 19116 10752
rect 19352 10606 19380 11047
rect 19340 10600 19392 10606
rect 19536 10577 19564 11086
rect 19616 11008 19668 11014
rect 19616 10950 19668 10956
rect 19628 10674 19656 10950
rect 19616 10668 19668 10674
rect 19616 10610 19668 10616
rect 19340 10542 19392 10548
rect 19522 10568 19578 10577
rect 19522 10503 19578 10512
rect 18880 10464 18932 10470
rect 18880 10406 18932 10412
rect 18696 10124 18748 10130
rect 18696 10066 18748 10072
rect 18708 9722 18736 10066
rect 18696 9716 18748 9722
rect 18696 9658 18748 9664
rect 18512 8832 18564 8838
rect 18512 8774 18564 8780
rect 18524 8498 18552 8774
rect 18512 8492 18564 8498
rect 18512 8434 18564 8440
rect 18524 8090 18552 8434
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18418 7984 18474 7993
rect 18418 7919 18474 7928
rect 18432 7342 18460 7919
rect 18524 7392 18552 8026
rect 18604 7404 18656 7410
rect 18524 7364 18604 7392
rect 18604 7346 18656 7352
rect 18420 7336 18472 7342
rect 18420 7278 18472 7284
rect 18510 6896 18566 6905
rect 18420 6860 18472 6866
rect 18510 6831 18512 6840
rect 18420 6802 18472 6808
rect 18564 6831 18566 6840
rect 18512 6802 18564 6808
rect 18432 6322 18460 6802
rect 18524 6458 18552 6802
rect 18616 6798 18644 7346
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 18512 6452 18564 6458
rect 18512 6394 18564 6400
rect 18616 6390 18644 6734
rect 18604 6384 18656 6390
rect 18604 6326 18656 6332
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 18340 3534 18368 4014
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18892 3097 18920 10406
rect 19340 10124 19392 10130
rect 19340 10066 19392 10072
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19260 9058 19288 9862
rect 19352 9586 19380 10066
rect 19628 10062 19656 10610
rect 19720 10130 19748 12407
rect 20088 11218 20116 15943
rect 20732 15162 20760 16050
rect 20956 15804 21252 15824
rect 21012 15802 21036 15804
rect 21092 15802 21116 15804
rect 21172 15802 21196 15804
rect 21034 15750 21036 15802
rect 21098 15750 21110 15802
rect 21172 15750 21174 15802
rect 21012 15748 21036 15750
rect 21092 15748 21116 15750
rect 21172 15748 21196 15750
rect 20956 15728 21252 15748
rect 21376 15706 21404 16730
rect 21456 15904 21508 15910
rect 21456 15846 21508 15852
rect 21364 15700 21416 15706
rect 21364 15642 21416 15648
rect 21376 15366 21404 15642
rect 21468 15434 21496 15846
rect 21456 15428 21508 15434
rect 21456 15370 21508 15376
rect 21364 15360 21416 15366
rect 21364 15302 21416 15308
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20534 15056 20590 15065
rect 20534 14991 20590 15000
rect 20350 13832 20406 13841
rect 20350 13767 20406 13776
rect 20364 12850 20392 13767
rect 20442 13560 20498 13569
rect 20442 13495 20498 13504
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20166 12608 20222 12617
rect 20166 12543 20222 12552
rect 20180 12345 20208 12543
rect 20364 12442 20392 12786
rect 20456 12782 20484 13495
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 20166 12336 20222 12345
rect 20166 12271 20222 12280
rect 20076 11212 20128 11218
rect 20076 11154 20128 11160
rect 19708 10124 19760 10130
rect 19708 10066 19760 10072
rect 19432 10056 19484 10062
rect 19432 9998 19484 10004
rect 19616 10056 19668 10062
rect 19616 9998 19668 10004
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19444 9450 19472 9998
rect 19628 9722 19656 9998
rect 20180 9994 20208 12271
rect 20260 11212 20312 11218
rect 20260 11154 20312 11160
rect 20272 10470 20300 11154
rect 20456 10538 20484 12718
rect 20548 11898 20576 14991
rect 20956 14716 21252 14736
rect 21012 14714 21036 14716
rect 21092 14714 21116 14716
rect 21172 14714 21196 14716
rect 21034 14662 21036 14714
rect 21098 14662 21110 14714
rect 21172 14662 21174 14714
rect 21012 14660 21036 14662
rect 21092 14660 21116 14662
rect 21172 14660 21196 14662
rect 20956 14640 21252 14660
rect 20956 13628 21252 13648
rect 21012 13626 21036 13628
rect 21092 13626 21116 13628
rect 21172 13626 21196 13628
rect 21034 13574 21036 13626
rect 21098 13574 21110 13626
rect 21172 13574 21174 13626
rect 21012 13572 21036 13574
rect 21092 13572 21116 13574
rect 21172 13572 21196 13574
rect 20956 13552 21252 13572
rect 21272 13388 21324 13394
rect 21272 13330 21324 13336
rect 20904 13184 20956 13190
rect 20904 13126 20956 13132
rect 20810 13016 20866 13025
rect 20810 12951 20866 12960
rect 20824 12646 20852 12951
rect 20916 12889 20944 13126
rect 21284 12986 21312 13330
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21456 13320 21508 13326
rect 21456 13262 21508 13268
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 20902 12880 20958 12889
rect 20902 12815 20958 12824
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20824 12442 20852 12582
rect 20956 12540 21252 12560
rect 21012 12538 21036 12540
rect 21092 12538 21116 12540
rect 21172 12538 21196 12540
rect 21034 12486 21036 12538
rect 21098 12486 21110 12538
rect 21172 12486 21174 12538
rect 21012 12484 21036 12486
rect 21092 12484 21116 12486
rect 21172 12484 21196 12486
rect 20956 12464 21252 12484
rect 20812 12436 20864 12442
rect 20812 12378 20864 12384
rect 21284 11898 21312 12922
rect 21376 12918 21404 13262
rect 21364 12912 21416 12918
rect 21364 12854 21416 12860
rect 21376 12442 21404 12854
rect 21468 12646 21496 13262
rect 21456 12640 21508 12646
rect 21456 12582 21508 12588
rect 21652 12442 21680 19366
rect 22112 19310 22140 19654
rect 22388 19514 22416 20538
rect 22376 19508 22428 19514
rect 22376 19450 22428 19456
rect 22664 19378 22692 20742
rect 25042 20496 25098 20505
rect 25042 20431 25098 20440
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 23112 19916 23164 19922
rect 23112 19858 23164 19864
rect 22652 19372 22704 19378
rect 22652 19314 22704 19320
rect 22100 19304 22152 19310
rect 22100 19246 22152 19252
rect 21732 19168 21784 19174
rect 21732 19110 21784 19116
rect 22468 19168 22520 19174
rect 22468 19110 22520 19116
rect 21364 12436 21416 12442
rect 21364 12378 21416 12384
rect 21640 12436 21692 12442
rect 21640 12378 21692 12384
rect 21640 12300 21692 12306
rect 21640 12242 21692 12248
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 21652 11558 21680 12242
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 20824 11393 20852 11494
rect 20956 11452 21252 11472
rect 21012 11450 21036 11452
rect 21092 11450 21116 11452
rect 21172 11450 21196 11452
rect 21034 11398 21036 11450
rect 21098 11398 21110 11450
rect 21172 11398 21174 11450
rect 21012 11396 21036 11398
rect 21092 11396 21116 11398
rect 21172 11396 21196 11398
rect 20810 11384 20866 11393
rect 20956 11376 21252 11396
rect 20810 11319 20866 11328
rect 21652 10577 21680 11494
rect 21638 10568 21694 10577
rect 20444 10532 20496 10538
rect 21638 10503 21694 10512
rect 20444 10474 20496 10480
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 21638 10432 21694 10441
rect 20168 9988 20220 9994
rect 20168 9930 20220 9936
rect 19616 9716 19668 9722
rect 19616 9658 19668 9664
rect 19432 9444 19484 9450
rect 19432 9386 19484 9392
rect 19260 9042 19380 9058
rect 19260 9036 19392 9042
rect 19260 9030 19340 9036
rect 19340 8978 19392 8984
rect 19352 8634 19380 8978
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 19708 8832 19760 8838
rect 19708 8774 19760 8780
rect 19444 8673 19472 8774
rect 19430 8664 19486 8673
rect 19340 8628 19392 8634
rect 19430 8599 19486 8608
rect 19340 8570 19392 8576
rect 19720 8430 19748 8774
rect 19708 8424 19760 8430
rect 19708 8366 19760 8372
rect 19720 7750 19748 8366
rect 19708 7744 19760 7750
rect 19708 7686 19760 7692
rect 19720 6254 19748 7686
rect 19708 6248 19760 6254
rect 19708 6190 19760 6196
rect 19720 5846 19748 6190
rect 19708 5840 19760 5846
rect 19708 5782 19760 5788
rect 19708 4820 19760 4826
rect 19708 4762 19760 4768
rect 19616 4616 19668 4622
rect 19616 4558 19668 4564
rect 19248 4480 19300 4486
rect 19248 4422 19300 4428
rect 19260 4185 19288 4422
rect 19246 4176 19302 4185
rect 19246 4111 19302 4120
rect 19628 3534 19656 4558
rect 19720 3738 19748 4762
rect 19892 4616 19944 4622
rect 19890 4584 19892 4593
rect 19944 4584 19946 4593
rect 19890 4519 19946 4528
rect 19904 4282 19932 4519
rect 19892 4276 19944 4282
rect 19892 4218 19944 4224
rect 20180 4146 20208 9930
rect 20272 5710 20300 10406
rect 20956 10364 21252 10384
rect 21638 10367 21694 10376
rect 21012 10362 21036 10364
rect 21092 10362 21116 10364
rect 21172 10362 21196 10364
rect 21034 10310 21036 10362
rect 21098 10310 21110 10362
rect 21172 10310 21174 10362
rect 21012 10308 21036 10310
rect 21092 10308 21116 10310
rect 21172 10308 21196 10310
rect 20956 10288 21252 10308
rect 21270 9616 21326 9625
rect 20628 9580 20680 9586
rect 21270 9551 21326 9560
rect 20628 9522 20680 9528
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 20456 8838 20484 9318
rect 20536 9036 20588 9042
rect 20536 8978 20588 8984
rect 20444 8832 20496 8838
rect 20444 8774 20496 8780
rect 20548 8090 20576 8978
rect 20536 8084 20588 8090
rect 20536 8026 20588 8032
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 20272 5302 20300 5646
rect 20640 5302 20668 9522
rect 20956 9276 21252 9296
rect 21012 9274 21036 9276
rect 21092 9274 21116 9276
rect 21172 9274 21196 9276
rect 21034 9222 21036 9274
rect 21098 9222 21110 9274
rect 21172 9222 21174 9274
rect 21012 9220 21036 9222
rect 21092 9220 21116 9222
rect 21172 9220 21196 9222
rect 20956 9200 21252 9220
rect 20812 8832 20864 8838
rect 20812 8774 20864 8780
rect 20718 8120 20774 8129
rect 20718 8055 20774 8064
rect 20732 7954 20760 8055
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20260 5296 20312 5302
rect 20258 5264 20260 5273
rect 20628 5296 20680 5302
rect 20312 5264 20314 5273
rect 20628 5238 20680 5244
rect 20258 5199 20314 5208
rect 20732 5166 20760 6598
rect 20720 5160 20772 5166
rect 20720 5102 20772 5108
rect 20444 5024 20496 5030
rect 20444 4966 20496 4972
rect 20456 4826 20484 4966
rect 20444 4820 20496 4826
rect 20444 4762 20496 4768
rect 20352 4208 20404 4214
rect 20352 4150 20404 4156
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 19708 3732 19760 3738
rect 19708 3674 19760 3680
rect 20272 3670 20300 3878
rect 20364 3738 20392 4150
rect 20628 4072 20680 4078
rect 20628 4014 20680 4020
rect 20352 3732 20404 3738
rect 20352 3674 20404 3680
rect 20260 3664 20312 3670
rect 20640 3641 20668 4014
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 20260 3606 20312 3612
rect 20626 3632 20682 3641
rect 20626 3567 20682 3576
rect 19616 3528 19668 3534
rect 19616 3470 19668 3476
rect 20732 3466 20760 3878
rect 20720 3460 20772 3466
rect 20720 3402 20772 3408
rect 18878 3088 18934 3097
rect 18878 3023 18934 3032
rect 19156 2916 19208 2922
rect 19156 2858 19208 2864
rect 18236 2508 18288 2514
rect 18236 2450 18288 2456
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 17788 480 17816 2382
rect 19168 480 19196 2858
rect 20824 2689 20852 8774
rect 20956 8188 21252 8208
rect 21012 8186 21036 8188
rect 21092 8186 21116 8188
rect 21172 8186 21196 8188
rect 21034 8134 21036 8186
rect 21098 8134 21110 8186
rect 21172 8134 21174 8186
rect 21012 8132 21036 8134
rect 21092 8132 21116 8134
rect 21172 8132 21196 8134
rect 20956 8112 21252 8132
rect 21284 7970 21312 9551
rect 21456 9444 21508 9450
rect 21456 9386 21508 9392
rect 21364 9172 21416 9178
rect 21364 9114 21416 9120
rect 21376 8974 21404 9114
rect 21468 8974 21496 9386
rect 21548 9104 21600 9110
rect 21548 9046 21600 9052
rect 21364 8968 21416 8974
rect 21364 8910 21416 8916
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21376 8090 21404 8910
rect 21468 8634 21496 8910
rect 21456 8628 21508 8634
rect 21456 8570 21508 8576
rect 21560 8090 21588 9046
rect 21364 8084 21416 8090
rect 21364 8026 21416 8032
rect 21548 8084 21600 8090
rect 21548 8026 21600 8032
rect 21284 7942 21404 7970
rect 20956 7100 21252 7120
rect 21012 7098 21036 7100
rect 21092 7098 21116 7100
rect 21172 7098 21196 7100
rect 21034 7046 21036 7098
rect 21098 7046 21110 7098
rect 21172 7046 21174 7098
rect 21012 7044 21036 7046
rect 21092 7044 21116 7046
rect 21172 7044 21196 7046
rect 20956 7024 21252 7044
rect 21272 6928 21324 6934
rect 21272 6870 21324 6876
rect 21284 6458 21312 6870
rect 21376 6866 21404 7942
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 21272 6452 21324 6458
rect 21272 6394 21324 6400
rect 21376 6390 21404 6802
rect 21364 6384 21416 6390
rect 21364 6326 21416 6332
rect 21272 6112 21324 6118
rect 21272 6054 21324 6060
rect 20956 6012 21252 6032
rect 21012 6010 21036 6012
rect 21092 6010 21116 6012
rect 21172 6010 21196 6012
rect 21034 5958 21036 6010
rect 21098 5958 21110 6010
rect 21172 5958 21174 6010
rect 21012 5956 21036 5958
rect 21092 5956 21116 5958
rect 21172 5956 21196 5958
rect 20956 5936 21252 5956
rect 21178 5808 21234 5817
rect 21178 5743 21180 5752
rect 21232 5743 21234 5752
rect 21180 5714 21232 5720
rect 20904 5568 20956 5574
rect 20904 5510 20956 5516
rect 20916 5234 20944 5510
rect 21192 5370 21220 5714
rect 21180 5364 21232 5370
rect 21180 5306 21232 5312
rect 21284 5234 21312 6054
rect 21364 5296 21416 5302
rect 21364 5238 21416 5244
rect 20904 5228 20956 5234
rect 20904 5170 20956 5176
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 20956 4924 21252 4944
rect 21012 4922 21036 4924
rect 21092 4922 21116 4924
rect 21172 4922 21196 4924
rect 21034 4870 21036 4922
rect 21098 4870 21110 4922
rect 21172 4870 21174 4922
rect 21012 4868 21036 4870
rect 21092 4868 21116 4870
rect 21172 4868 21196 4870
rect 20956 4848 21252 4868
rect 21284 4826 21312 5170
rect 21376 4826 21404 5238
rect 21272 4820 21324 4826
rect 21272 4762 21324 4768
rect 21364 4820 21416 4826
rect 21364 4762 21416 4768
rect 20956 3836 21252 3856
rect 21012 3834 21036 3836
rect 21092 3834 21116 3836
rect 21172 3834 21196 3836
rect 21034 3782 21036 3834
rect 21098 3782 21110 3834
rect 21172 3782 21174 3834
rect 21012 3780 21036 3782
rect 21092 3780 21116 3782
rect 21172 3780 21196 3782
rect 20956 3760 21252 3780
rect 21284 3534 21312 4762
rect 21364 4684 21416 4690
rect 21364 4626 21416 4632
rect 21376 4214 21404 4626
rect 21652 4282 21680 10367
rect 21640 4276 21692 4282
rect 21640 4218 21692 4224
rect 21364 4208 21416 4214
rect 21364 4150 21416 4156
rect 21652 4078 21680 4218
rect 21640 4072 21692 4078
rect 21640 4014 21692 4020
rect 21364 3664 21416 3670
rect 21364 3606 21416 3612
rect 21272 3528 21324 3534
rect 21272 3470 21324 3476
rect 21284 3126 21312 3470
rect 21376 3194 21404 3606
rect 21364 3188 21416 3194
rect 21364 3130 21416 3136
rect 21272 3120 21324 3126
rect 21272 3062 21324 3068
rect 21744 2922 21772 19110
rect 22480 18970 22508 19110
rect 22468 18964 22520 18970
rect 22468 18906 22520 18912
rect 22848 18902 22876 19858
rect 23124 19174 23152 19858
rect 24216 19712 24268 19718
rect 24216 19654 24268 19660
rect 24228 19514 24256 19654
rect 23572 19508 23624 19514
rect 23572 19450 23624 19456
rect 24216 19508 24268 19514
rect 24216 19450 24268 19456
rect 23112 19168 23164 19174
rect 23112 19110 23164 19116
rect 22836 18896 22888 18902
rect 22836 18838 22888 18844
rect 22744 17332 22796 17338
rect 22744 17274 22796 17280
rect 22652 16244 22704 16250
rect 22652 16186 22704 16192
rect 21916 15700 21968 15706
rect 21916 15642 21968 15648
rect 21824 15564 21876 15570
rect 21824 15506 21876 15512
rect 21836 15162 21864 15506
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 21836 14074 21864 15098
rect 21928 15065 21956 15642
rect 22664 15570 22692 16186
rect 22756 15638 22784 17274
rect 22848 16250 22876 18838
rect 23124 17610 23152 19110
rect 23296 18828 23348 18834
rect 23296 18770 23348 18776
rect 23480 18828 23532 18834
rect 23480 18770 23532 18776
rect 23308 18154 23336 18770
rect 23296 18148 23348 18154
rect 23296 18090 23348 18096
rect 23308 17882 23336 18090
rect 23492 18086 23520 18770
rect 23584 18766 23612 19450
rect 24952 19372 25004 19378
rect 24952 19314 25004 19320
rect 24584 19304 24636 19310
rect 24584 19246 24636 19252
rect 24124 19236 24176 19242
rect 24124 19178 24176 19184
rect 24136 18970 24164 19178
rect 24596 18970 24624 19246
rect 24124 18964 24176 18970
rect 24124 18906 24176 18912
rect 24584 18964 24636 18970
rect 24584 18906 24636 18912
rect 23572 18760 23624 18766
rect 23572 18702 23624 18708
rect 23584 18426 23612 18702
rect 23572 18420 23624 18426
rect 23572 18362 23624 18368
rect 23480 18080 23532 18086
rect 23480 18022 23532 18028
rect 24768 18080 24820 18086
rect 24820 18028 24900 18034
rect 24768 18022 24900 18028
rect 24780 18006 24900 18022
rect 24872 17882 24900 18006
rect 23296 17876 23348 17882
rect 23296 17818 23348 17824
rect 24860 17876 24912 17882
rect 24860 17818 24912 17824
rect 24676 17808 24728 17814
rect 24676 17750 24728 17756
rect 23204 17740 23256 17746
rect 23204 17682 23256 17688
rect 23112 17604 23164 17610
rect 23112 17546 23164 17552
rect 23124 17270 23152 17546
rect 23112 17264 23164 17270
rect 23216 17241 23244 17682
rect 23480 17672 23532 17678
rect 23480 17614 23532 17620
rect 23492 17338 23520 17614
rect 23480 17332 23532 17338
rect 23480 17274 23532 17280
rect 23112 17206 23164 17212
rect 23202 17232 23258 17241
rect 23124 16794 23152 17206
rect 23202 17167 23258 17176
rect 24216 17196 24268 17202
rect 23216 16998 23244 17167
rect 24216 17138 24268 17144
rect 23478 17096 23534 17105
rect 23478 17031 23480 17040
rect 23532 17031 23534 17040
rect 23480 17002 23532 17008
rect 23204 16992 23256 16998
rect 23202 16960 23204 16969
rect 23664 16992 23716 16998
rect 23256 16960 23258 16969
rect 23664 16934 23716 16940
rect 23202 16895 23258 16904
rect 23112 16788 23164 16794
rect 23112 16730 23164 16736
rect 23676 16658 23704 16934
rect 24228 16794 24256 17138
rect 24216 16788 24268 16794
rect 24216 16730 24268 16736
rect 23664 16652 23716 16658
rect 23664 16594 23716 16600
rect 24400 16652 24452 16658
rect 24400 16594 24452 16600
rect 22836 16244 22888 16250
rect 22836 16186 22888 16192
rect 22744 15632 22796 15638
rect 22744 15574 22796 15580
rect 22652 15564 22704 15570
rect 22652 15506 22704 15512
rect 22664 15366 22692 15506
rect 22652 15360 22704 15366
rect 22652 15302 22704 15308
rect 22664 15094 22692 15302
rect 22756 15162 22784 15574
rect 23676 15201 23704 16594
rect 23756 15904 23808 15910
rect 23756 15846 23808 15852
rect 23662 15192 23718 15201
rect 22744 15156 22796 15162
rect 23662 15127 23718 15136
rect 22744 15098 22796 15104
rect 22652 15088 22704 15094
rect 21914 15056 21970 15065
rect 22652 15030 22704 15036
rect 21914 14991 21970 15000
rect 22664 14550 22692 15030
rect 22652 14544 22704 14550
rect 22652 14486 22704 14492
rect 22376 14476 22428 14482
rect 22376 14418 22428 14424
rect 22388 14074 22416 14418
rect 22664 14074 22692 14486
rect 23768 14278 23796 15846
rect 24412 15434 24440 16594
rect 24688 16454 24716 17750
rect 24860 17740 24912 17746
rect 24860 17682 24912 17688
rect 24768 17128 24820 17134
rect 24768 17070 24820 17076
rect 24676 16448 24728 16454
rect 24676 16390 24728 16396
rect 24688 16182 24716 16390
rect 24780 16250 24808 17070
rect 24872 16794 24900 17682
rect 24860 16788 24912 16794
rect 24860 16730 24912 16736
rect 24858 16688 24914 16697
rect 24858 16623 24914 16632
rect 24768 16244 24820 16250
rect 24768 16186 24820 16192
rect 24676 16176 24728 16182
rect 24676 16118 24728 16124
rect 24872 15450 24900 16623
rect 24400 15428 24452 15434
rect 24400 15370 24452 15376
rect 24688 15422 24900 15450
rect 24412 15337 24440 15370
rect 24398 15328 24454 15337
rect 24398 15263 24454 15272
rect 23756 14272 23808 14278
rect 23756 14214 23808 14220
rect 21824 14068 21876 14074
rect 21824 14010 21876 14016
rect 22376 14068 22428 14074
rect 22376 14010 22428 14016
rect 22652 14068 22704 14074
rect 22652 14010 22704 14016
rect 22664 13841 22692 14010
rect 22650 13832 22706 13841
rect 22650 13767 22706 13776
rect 22928 13456 22980 13462
rect 21822 13424 21878 13433
rect 22928 13398 22980 13404
rect 23664 13456 23716 13462
rect 23664 13398 23716 13404
rect 21822 13359 21878 13368
rect 21836 13025 21864 13359
rect 22560 13184 22612 13190
rect 22560 13126 22612 13132
rect 21822 13016 21878 13025
rect 21822 12951 21878 12960
rect 22100 12708 22152 12714
rect 22100 12650 22152 12656
rect 21824 12436 21876 12442
rect 21824 12378 21876 12384
rect 21836 11665 21864 12378
rect 22112 12238 22140 12650
rect 22100 12232 22152 12238
rect 22100 12174 22152 12180
rect 22112 11762 22140 12174
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 21822 11656 21878 11665
rect 21822 11591 21878 11600
rect 21836 11354 21864 11591
rect 21824 11348 21876 11354
rect 21824 11290 21876 11296
rect 22100 11280 22152 11286
rect 22100 11222 22152 11228
rect 21916 11144 21968 11150
rect 21916 11086 21968 11092
rect 21928 10538 21956 11086
rect 22112 10962 22140 11222
rect 22020 10934 22140 10962
rect 22020 10810 22048 10934
rect 22008 10804 22060 10810
rect 22008 10746 22060 10752
rect 21916 10532 21968 10538
rect 21916 10474 21968 10480
rect 22020 9722 22048 10746
rect 22100 10532 22152 10538
rect 22100 10474 22152 10480
rect 22008 9716 22060 9722
rect 22008 9658 22060 9664
rect 22112 9518 22140 10474
rect 22100 9512 22152 9518
rect 22100 9454 22152 9460
rect 22100 8356 22152 8362
rect 22020 8316 22100 8344
rect 22020 8090 22048 8316
rect 22100 8298 22152 8304
rect 22008 8084 22060 8090
rect 22008 8026 22060 8032
rect 21824 7948 21876 7954
rect 21824 7890 21876 7896
rect 22376 7948 22428 7954
rect 22376 7890 22428 7896
rect 21836 7546 21864 7890
rect 21824 7540 21876 7546
rect 21824 7482 21876 7488
rect 22284 7404 22336 7410
rect 22284 7346 22336 7352
rect 22008 7336 22060 7342
rect 22008 7278 22060 7284
rect 22020 7002 22048 7278
rect 22296 7274 22324 7346
rect 22284 7268 22336 7274
rect 22284 7210 22336 7216
rect 22008 6996 22060 7002
rect 22008 6938 22060 6944
rect 21824 6792 21876 6798
rect 21916 6792 21968 6798
rect 21824 6734 21876 6740
rect 21914 6760 21916 6769
rect 21968 6760 21970 6769
rect 21836 6458 21864 6734
rect 22296 6730 22324 7210
rect 22388 6769 22416 7890
rect 22468 7404 22520 7410
rect 22468 7346 22520 7352
rect 22480 7002 22508 7346
rect 22468 6996 22520 7002
rect 22468 6938 22520 6944
rect 22374 6760 22430 6769
rect 21914 6695 21970 6704
rect 22284 6724 22336 6730
rect 22374 6695 22430 6704
rect 22284 6666 22336 6672
rect 21824 6452 21876 6458
rect 21824 6394 21876 6400
rect 21836 6186 21864 6394
rect 21824 6180 21876 6186
rect 21824 6122 21876 6128
rect 21836 5710 21864 6122
rect 22192 5840 22244 5846
rect 22192 5782 22244 5788
rect 21824 5704 21876 5710
rect 21824 5646 21876 5652
rect 21836 4690 21864 5646
rect 22204 5234 22232 5782
rect 22192 5228 22244 5234
rect 22192 5170 22244 5176
rect 22100 4820 22152 4826
rect 22100 4762 22152 4768
rect 21824 4684 21876 4690
rect 21824 4626 21876 4632
rect 22112 4146 22140 4762
rect 22204 4622 22232 5170
rect 22376 5160 22428 5166
rect 22376 5102 22428 5108
rect 22388 4758 22416 5102
rect 22376 4752 22428 4758
rect 22376 4694 22428 4700
rect 22192 4616 22244 4622
rect 22244 4564 22324 4570
rect 22192 4558 22324 4564
rect 22204 4542 22324 4558
rect 22100 4140 22152 4146
rect 22100 4082 22152 4088
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 21836 3738 21864 3878
rect 22296 3738 22324 4542
rect 22388 4282 22416 4694
rect 22376 4276 22428 4282
rect 22376 4218 22428 4224
rect 21824 3732 21876 3738
rect 21824 3674 21876 3680
rect 22284 3732 22336 3738
rect 22284 3674 22336 3680
rect 21836 3194 21864 3674
rect 21824 3188 21876 3194
rect 21824 3130 21876 3136
rect 21732 2916 21784 2922
rect 21732 2858 21784 2864
rect 20956 2748 21252 2768
rect 21012 2746 21036 2748
rect 21092 2746 21116 2748
rect 21172 2746 21196 2748
rect 21034 2694 21036 2746
rect 21098 2694 21110 2746
rect 21172 2694 21174 2746
rect 21012 2692 21036 2694
rect 21092 2692 21116 2694
rect 21172 2692 21196 2694
rect 20810 2680 20866 2689
rect 20956 2672 21252 2692
rect 22572 2650 22600 13126
rect 22940 12986 22968 13398
rect 23572 13388 23624 13394
rect 23572 13330 23624 13336
rect 23584 12986 23612 13330
rect 22928 12980 22980 12986
rect 22928 12922 22980 12928
rect 23572 12980 23624 12986
rect 23572 12922 23624 12928
rect 23584 12442 23612 12922
rect 23676 12442 23704 13398
rect 23768 13326 23796 14214
rect 24412 13569 24440 15263
rect 24492 15156 24544 15162
rect 24492 15098 24544 15104
rect 24398 13560 24454 13569
rect 24398 13495 24454 13504
rect 23756 13320 23808 13326
rect 23756 13262 23808 13268
rect 23768 12918 23796 13262
rect 24308 13184 24360 13190
rect 24308 13126 24360 13132
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 24320 12646 24348 13126
rect 24412 12889 24440 13495
rect 24398 12880 24454 12889
rect 24398 12815 24454 12824
rect 24400 12776 24452 12782
rect 24400 12718 24452 12724
rect 24308 12640 24360 12646
rect 24308 12582 24360 12588
rect 23572 12436 23624 12442
rect 23572 12378 23624 12384
rect 23664 12436 23716 12442
rect 24412 12424 24440 12718
rect 23664 12378 23716 12384
rect 24320 12396 24440 12424
rect 24124 12368 24176 12374
rect 24124 12310 24176 12316
rect 23020 12232 23072 12238
rect 23020 12174 23072 12180
rect 23032 11626 23060 12174
rect 24136 11898 24164 12310
rect 24320 12102 24348 12396
rect 24504 12356 24532 15098
rect 24584 14816 24636 14822
rect 24584 14758 24636 14764
rect 24596 14482 24624 14758
rect 24584 14476 24636 14482
rect 24584 14418 24636 14424
rect 24596 12850 24624 14418
rect 24688 13161 24716 15422
rect 24768 15360 24820 15366
rect 24820 15308 24900 15314
rect 24768 15302 24900 15308
rect 24780 15286 24900 15302
rect 24872 14074 24900 15286
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 24860 13932 24912 13938
rect 24860 13874 24912 13880
rect 24872 13274 24900 13874
rect 24780 13246 24900 13274
rect 24674 13152 24730 13161
rect 24674 13087 24730 13096
rect 24674 12880 24730 12889
rect 24584 12844 24636 12850
rect 24674 12815 24730 12824
rect 24584 12786 24636 12792
rect 24596 12374 24624 12786
rect 24412 12328 24532 12356
rect 24584 12368 24636 12374
rect 24308 12096 24360 12102
rect 24308 12038 24360 12044
rect 24124 11892 24176 11898
rect 24124 11834 24176 11840
rect 24320 11665 24348 12038
rect 24306 11656 24362 11665
rect 23020 11620 23072 11626
rect 24306 11591 24362 11600
rect 23020 11562 23072 11568
rect 22928 11552 22980 11558
rect 22928 11494 22980 11500
rect 22940 11354 22968 11494
rect 22928 11348 22980 11354
rect 22928 11290 22980 11296
rect 24412 9625 24440 12328
rect 24584 12310 24636 12316
rect 24584 12232 24636 12238
rect 24584 12174 24636 12180
rect 24596 11354 24624 12174
rect 24584 11348 24636 11354
rect 24584 11290 24636 11296
rect 24688 10010 24716 12815
rect 24780 12782 24808 13246
rect 24860 13184 24912 13190
rect 24860 13126 24912 13132
rect 24768 12776 24820 12782
rect 24768 12718 24820 12724
rect 24768 12436 24820 12442
rect 24872 12424 24900 13126
rect 24820 12396 24900 12424
rect 24768 12378 24820 12384
rect 24766 12336 24822 12345
rect 24766 12271 24822 12280
rect 24596 9982 24716 10010
rect 24398 9616 24454 9625
rect 24398 9551 24454 9560
rect 23664 9512 23716 9518
rect 23664 9454 23716 9460
rect 23480 9376 23532 9382
rect 23480 9318 23532 9324
rect 22744 9172 22796 9178
rect 22744 9114 22796 9120
rect 22756 8498 22784 9114
rect 22836 9036 22888 9042
rect 22836 8978 22888 8984
rect 22744 8492 22796 8498
rect 22744 8434 22796 8440
rect 22652 7880 22704 7886
rect 22652 7822 22704 7828
rect 22664 7410 22692 7822
rect 22756 7546 22784 8434
rect 22848 8362 22876 8978
rect 23020 8968 23072 8974
rect 23020 8910 23072 8916
rect 22836 8356 22888 8362
rect 22836 8298 22888 8304
rect 23032 8294 23060 8910
rect 23020 8288 23072 8294
rect 23492 8242 23520 9318
rect 23676 8838 23704 9454
rect 23664 8832 23716 8838
rect 23664 8774 23716 8780
rect 23020 8230 23072 8236
rect 23400 8214 23520 8242
rect 22836 8084 22888 8090
rect 22836 8026 22888 8032
rect 22744 7540 22796 7546
rect 22744 7482 22796 7488
rect 22652 7404 22704 7410
rect 22652 7346 22704 7352
rect 22848 6934 22876 8026
rect 23400 7886 23428 8214
rect 23388 7880 23440 7886
rect 23388 7822 23440 7828
rect 23478 7576 23534 7585
rect 23112 7540 23164 7546
rect 23478 7511 23534 7520
rect 23112 7482 23164 7488
rect 23124 7313 23152 7482
rect 23492 7410 23520 7511
rect 23480 7404 23532 7410
rect 23480 7346 23532 7352
rect 23676 7313 23704 8774
rect 23848 7948 23900 7954
rect 23848 7890 23900 7896
rect 23860 7449 23888 7890
rect 24032 7880 24084 7886
rect 24032 7822 24084 7828
rect 24308 7880 24360 7886
rect 24308 7822 24360 7828
rect 24044 7546 24072 7822
rect 24032 7540 24084 7546
rect 24032 7482 24084 7488
rect 24044 7449 24072 7482
rect 23846 7440 23902 7449
rect 23846 7375 23902 7384
rect 24030 7440 24086 7449
rect 24320 7410 24348 7822
rect 24030 7375 24086 7384
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 24308 7404 24360 7410
rect 24308 7346 24360 7352
rect 23110 7304 23166 7313
rect 23110 7239 23166 7248
rect 23662 7304 23718 7313
rect 23662 7239 23718 7248
rect 22836 6928 22888 6934
rect 22836 6870 22888 6876
rect 23572 6316 23624 6322
rect 23572 6258 23624 6264
rect 23584 5681 23612 6258
rect 23570 5672 23626 5681
rect 23570 5607 23626 5616
rect 23676 5574 23704 7239
rect 24136 7041 24164 7346
rect 24122 7032 24178 7041
rect 24122 6967 24178 6976
rect 24320 6798 24348 7346
rect 24596 7002 24624 9982
rect 24676 9920 24728 9926
rect 24676 9862 24728 9868
rect 24688 9450 24716 9862
rect 24676 9444 24728 9450
rect 24676 9386 24728 9392
rect 24676 9104 24728 9110
rect 24676 9046 24728 9052
rect 24688 8634 24716 9046
rect 24676 8628 24728 8634
rect 24676 8570 24728 8576
rect 24780 7546 24808 12271
rect 24964 12186 24992 19314
rect 25056 13190 25084 20431
rect 25148 15706 25176 22335
rect 25240 19378 25268 23446
rect 25778 23080 25834 23089
rect 25778 23015 25834 23024
rect 25792 22166 25820 23015
rect 25780 22160 25832 22166
rect 25780 22102 25832 22108
rect 25884 21434 25912 23559
rect 28262 23520 28318 24000
rect 27526 21856 27582 21865
rect 25956 21788 26252 21808
rect 27526 21791 27582 21800
rect 26012 21786 26036 21788
rect 26092 21786 26116 21788
rect 26172 21786 26196 21788
rect 26034 21734 26036 21786
rect 26098 21734 26110 21786
rect 26172 21734 26174 21786
rect 26012 21732 26036 21734
rect 26092 21732 26116 21734
rect 26172 21732 26196 21734
rect 25956 21712 26252 21732
rect 25608 21406 25912 21434
rect 25412 19712 25464 19718
rect 25412 19654 25464 19660
rect 25424 19378 25452 19654
rect 25504 19440 25556 19446
rect 25504 19382 25556 19388
rect 25228 19372 25280 19378
rect 25228 19314 25280 19320
rect 25412 19372 25464 19378
rect 25412 19314 25464 19320
rect 25318 19272 25374 19281
rect 25318 19207 25374 19216
rect 25332 19174 25360 19207
rect 25320 19168 25372 19174
rect 25320 19110 25372 19116
rect 25226 18728 25282 18737
rect 25226 18663 25282 18672
rect 25136 15700 25188 15706
rect 25136 15642 25188 15648
rect 25240 13938 25268 18663
rect 25424 17678 25452 19314
rect 25516 19242 25544 19382
rect 25504 19236 25556 19242
rect 25504 19178 25556 19184
rect 25502 19000 25558 19009
rect 25502 18935 25558 18944
rect 25516 18329 25544 18935
rect 25502 18320 25558 18329
rect 25502 18255 25558 18264
rect 25412 17672 25464 17678
rect 25412 17614 25464 17620
rect 25424 17338 25452 17614
rect 25412 17332 25464 17338
rect 25412 17274 25464 17280
rect 25412 17196 25464 17202
rect 25412 17138 25464 17144
rect 25320 16584 25372 16590
rect 25320 16526 25372 16532
rect 25332 16046 25360 16526
rect 25424 16522 25452 17138
rect 25502 17096 25558 17105
rect 25502 17031 25558 17040
rect 25412 16516 25464 16522
rect 25412 16458 25464 16464
rect 25424 16250 25452 16458
rect 25412 16244 25464 16250
rect 25412 16186 25464 16192
rect 25424 16046 25452 16186
rect 25320 16040 25372 16046
rect 25320 15982 25372 15988
rect 25412 16040 25464 16046
rect 25412 15982 25464 15988
rect 25318 15872 25374 15881
rect 25318 15807 25374 15816
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 25332 13410 25360 15807
rect 25424 15706 25452 15982
rect 25412 15700 25464 15706
rect 25412 15642 25464 15648
rect 25516 15609 25544 17031
rect 25502 15600 25558 15609
rect 25502 15535 25558 15544
rect 25410 15464 25466 15473
rect 25410 15399 25466 15408
rect 25424 15366 25452 15399
rect 25412 15360 25464 15366
rect 25412 15302 25464 15308
rect 25412 15020 25464 15026
rect 25412 14962 25464 14968
rect 25424 14618 25452 14962
rect 25504 14884 25556 14890
rect 25504 14826 25556 14832
rect 25412 14612 25464 14618
rect 25412 14554 25464 14560
rect 25424 13870 25452 14554
rect 25412 13864 25464 13870
rect 25412 13806 25464 13812
rect 25136 13388 25188 13394
rect 25332 13382 25452 13410
rect 25136 13330 25188 13336
rect 25044 13184 25096 13190
rect 25044 13126 25096 13132
rect 25044 12708 25096 12714
rect 25044 12650 25096 12656
rect 24872 12158 24992 12186
rect 24872 11234 24900 12158
rect 24952 12096 25004 12102
rect 24952 12038 25004 12044
rect 24964 11354 24992 12038
rect 25056 11898 25084 12650
rect 25148 12646 25176 13330
rect 25320 13320 25372 13326
rect 25320 13262 25372 13268
rect 25332 12986 25360 13262
rect 25320 12980 25372 12986
rect 25320 12922 25372 12928
rect 25424 12866 25452 13382
rect 25516 13326 25544 14826
rect 25504 13320 25556 13326
rect 25504 13262 25556 13268
rect 25504 13184 25556 13190
rect 25504 13126 25556 13132
rect 25332 12838 25452 12866
rect 25228 12708 25280 12714
rect 25228 12650 25280 12656
rect 25136 12640 25188 12646
rect 25136 12582 25188 12588
rect 25148 12481 25176 12582
rect 25134 12472 25190 12481
rect 25134 12407 25190 12416
rect 25240 12209 25268 12650
rect 25226 12200 25282 12209
rect 25226 12135 25282 12144
rect 25044 11892 25096 11898
rect 25044 11834 25096 11840
rect 25240 11830 25268 12135
rect 25228 11824 25280 11830
rect 25134 11792 25190 11801
rect 25228 11766 25280 11772
rect 25134 11727 25136 11736
rect 25188 11727 25190 11736
rect 25136 11698 25188 11704
rect 24952 11348 25004 11354
rect 24952 11290 25004 11296
rect 24872 11206 24992 11234
rect 24860 9920 24912 9926
rect 24860 9862 24912 9868
rect 24872 9178 24900 9862
rect 24860 9172 24912 9178
rect 24860 9114 24912 9120
rect 24872 8634 24900 9114
rect 24860 8628 24912 8634
rect 24860 8570 24912 8576
rect 24768 7540 24820 7546
rect 24768 7482 24820 7488
rect 24780 7342 24808 7482
rect 24768 7336 24820 7342
rect 24768 7278 24820 7284
rect 24584 6996 24636 7002
rect 24584 6938 24636 6944
rect 23940 6792 23992 6798
rect 23940 6734 23992 6740
rect 24308 6792 24360 6798
rect 24308 6734 24360 6740
rect 23952 6390 23980 6734
rect 24320 6458 24348 6734
rect 24308 6452 24360 6458
rect 24308 6394 24360 6400
rect 23940 6384 23992 6390
rect 23940 6326 23992 6332
rect 23664 5568 23716 5574
rect 23664 5510 23716 5516
rect 23676 5234 23704 5510
rect 23664 5228 23716 5234
rect 23664 5170 23716 5176
rect 23572 5024 23624 5030
rect 23572 4966 23624 4972
rect 23584 4593 23612 4966
rect 23570 4584 23626 4593
rect 23570 4519 23572 4528
rect 23624 4519 23626 4528
rect 23572 4490 23624 4496
rect 23952 3602 23980 6326
rect 24596 6322 24624 6938
rect 24584 6316 24636 6322
rect 24584 6258 24636 6264
rect 24858 3768 24914 3777
rect 24858 3703 24914 3712
rect 23940 3596 23992 3602
rect 23940 3538 23992 3544
rect 23846 2952 23902 2961
rect 23846 2887 23902 2896
rect 24032 2916 24084 2922
rect 23860 2854 23888 2887
rect 24032 2858 24084 2864
rect 23848 2848 23900 2854
rect 23848 2790 23900 2796
rect 20810 2615 20866 2624
rect 22560 2644 22612 2650
rect 22560 2586 22612 2592
rect 24044 2514 24072 2858
rect 24032 2508 24084 2514
rect 24032 2450 24084 2456
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 22008 2440 22060 2446
rect 22008 2382 22060 2388
rect 23480 2440 23532 2446
rect 23480 2382 23532 2388
rect 20640 480 20668 2382
rect 22020 480 22048 2382
rect 23492 480 23520 2382
rect 24872 480 24900 3703
rect 24964 2990 24992 11206
rect 25228 10464 25280 10470
rect 25228 10406 25280 10412
rect 25240 10130 25268 10406
rect 25228 10124 25280 10130
rect 25228 10066 25280 10072
rect 25044 9376 25096 9382
rect 25044 9318 25096 9324
rect 25056 8974 25084 9318
rect 25240 9178 25268 10066
rect 25228 9172 25280 9178
rect 25228 9114 25280 9120
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 25332 7970 25360 12838
rect 25412 12776 25464 12782
rect 25412 12718 25464 12724
rect 25424 12102 25452 12718
rect 25516 12594 25544 13126
rect 25608 12714 25636 21406
rect 25870 21312 25926 21321
rect 25870 21247 25926 21256
rect 25688 19236 25740 19242
rect 25688 19178 25740 19184
rect 25700 18873 25728 19178
rect 25686 18864 25742 18873
rect 25686 18799 25742 18808
rect 25700 18630 25728 18799
rect 25688 18624 25740 18630
rect 25688 18566 25740 18572
rect 25700 18329 25728 18566
rect 25686 18320 25742 18329
rect 25686 18255 25742 18264
rect 25686 17640 25742 17649
rect 25686 17575 25742 17584
rect 25700 16697 25728 17575
rect 25780 17536 25832 17542
rect 25780 17478 25832 17484
rect 25792 17066 25820 17478
rect 25780 17060 25832 17066
rect 25780 17002 25832 17008
rect 25780 16788 25832 16794
rect 25780 16730 25832 16736
rect 25686 16688 25742 16697
rect 25686 16623 25742 16632
rect 25686 16280 25742 16289
rect 25686 16215 25688 16224
rect 25740 16215 25742 16224
rect 25688 16186 25740 16192
rect 25686 15464 25742 15473
rect 25686 15399 25742 15408
rect 25700 13297 25728 15399
rect 25792 14498 25820 16730
rect 25884 15162 25912 21247
rect 25956 20700 26252 20720
rect 26012 20698 26036 20700
rect 26092 20698 26116 20700
rect 26172 20698 26196 20700
rect 26034 20646 26036 20698
rect 26098 20646 26110 20698
rect 26172 20646 26174 20698
rect 26012 20644 26036 20646
rect 26092 20644 26116 20646
rect 26172 20644 26196 20646
rect 25956 20624 26252 20644
rect 26054 20360 26110 20369
rect 26054 20295 26110 20304
rect 26068 20262 26096 20295
rect 26056 20256 26108 20262
rect 26056 20198 26108 20204
rect 27252 20256 27304 20262
rect 27252 20198 27304 20204
rect 27436 20256 27488 20262
rect 27436 20198 27488 20204
rect 25956 19612 26252 19632
rect 26012 19610 26036 19612
rect 26092 19610 26116 19612
rect 26172 19610 26196 19612
rect 26034 19558 26036 19610
rect 26098 19558 26110 19610
rect 26172 19558 26174 19610
rect 26012 19556 26036 19558
rect 26092 19556 26116 19558
rect 26172 19556 26196 19558
rect 25956 19536 26252 19556
rect 26976 19236 27028 19242
rect 26976 19178 27028 19184
rect 26424 19168 26476 19174
rect 26424 19110 26476 19116
rect 25956 18524 26252 18544
rect 26012 18522 26036 18524
rect 26092 18522 26116 18524
rect 26172 18522 26196 18524
rect 26034 18470 26036 18522
rect 26098 18470 26110 18522
rect 26172 18470 26174 18522
rect 26012 18468 26036 18470
rect 26092 18468 26116 18470
rect 26172 18468 26196 18470
rect 25956 18448 26252 18468
rect 25956 17436 26252 17456
rect 26012 17434 26036 17436
rect 26092 17434 26116 17436
rect 26172 17434 26196 17436
rect 26034 17382 26036 17434
rect 26098 17382 26110 17434
rect 26172 17382 26174 17434
rect 26012 17380 26036 17382
rect 26092 17380 26116 17382
rect 26172 17380 26196 17382
rect 25956 17360 26252 17380
rect 26330 16960 26386 16969
rect 26330 16895 26386 16904
rect 25956 16348 26252 16368
rect 26012 16346 26036 16348
rect 26092 16346 26116 16348
rect 26172 16346 26196 16348
rect 26034 16294 26036 16346
rect 26098 16294 26110 16346
rect 26172 16294 26174 16346
rect 26012 16292 26036 16294
rect 26092 16292 26116 16294
rect 26172 16292 26196 16294
rect 25956 16272 26252 16292
rect 26240 15904 26292 15910
rect 26240 15846 26292 15852
rect 26252 15348 26280 15846
rect 26344 15570 26372 16895
rect 26332 15564 26384 15570
rect 26332 15506 26384 15512
rect 26332 15360 26384 15366
rect 26252 15320 26332 15348
rect 26332 15302 26384 15308
rect 25956 15260 26252 15280
rect 26012 15258 26036 15260
rect 26092 15258 26116 15260
rect 26172 15258 26196 15260
rect 26034 15206 26036 15258
rect 26098 15206 26110 15258
rect 26172 15206 26174 15258
rect 26012 15204 26036 15206
rect 26092 15204 26116 15206
rect 26172 15204 26196 15206
rect 25956 15184 26252 15204
rect 25872 15156 25924 15162
rect 25872 15098 25924 15104
rect 25792 14470 25912 14498
rect 25780 13864 25832 13870
rect 25780 13806 25832 13812
rect 25686 13288 25742 13297
rect 25686 13223 25742 13232
rect 25792 12850 25820 13806
rect 25780 12844 25832 12850
rect 25780 12786 25832 12792
rect 25596 12708 25648 12714
rect 25596 12650 25648 12656
rect 25516 12566 25636 12594
rect 25502 12472 25558 12481
rect 25502 12407 25558 12416
rect 25412 12096 25464 12102
rect 25412 12038 25464 12044
rect 25424 11121 25452 12038
rect 25410 11112 25466 11121
rect 25410 11047 25466 11056
rect 25516 10266 25544 12407
rect 25504 10260 25556 10266
rect 25504 10202 25556 10208
rect 25516 9722 25544 10202
rect 25504 9716 25556 9722
rect 25504 9658 25556 9664
rect 25240 7954 25360 7970
rect 25228 7948 25360 7954
rect 25280 7942 25360 7948
rect 25228 7890 25280 7896
rect 25240 7546 25268 7890
rect 25320 7744 25372 7750
rect 25320 7686 25372 7692
rect 25228 7540 25280 7546
rect 25228 7482 25280 7488
rect 25332 7342 25360 7686
rect 25320 7336 25372 7342
rect 25318 7304 25320 7313
rect 25372 7304 25374 7313
rect 25318 7239 25374 7248
rect 25608 6905 25636 12566
rect 25792 12442 25820 12786
rect 25780 12436 25832 12442
rect 25780 12378 25832 12384
rect 25780 12096 25832 12102
rect 25780 12038 25832 12044
rect 25688 11688 25740 11694
rect 25688 11630 25740 11636
rect 25700 11218 25728 11630
rect 25688 11212 25740 11218
rect 25688 11154 25740 11160
rect 25792 6905 25820 12038
rect 25884 11121 25912 14470
rect 25956 14172 26252 14192
rect 26012 14170 26036 14172
rect 26092 14170 26116 14172
rect 26172 14170 26196 14172
rect 26034 14118 26036 14170
rect 26098 14118 26110 14170
rect 26172 14118 26174 14170
rect 26012 14116 26036 14118
rect 26092 14116 26116 14118
rect 26172 14116 26196 14118
rect 25956 14096 26252 14116
rect 25956 13084 26252 13104
rect 26012 13082 26036 13084
rect 26092 13082 26116 13084
rect 26172 13082 26196 13084
rect 26034 13030 26036 13082
rect 26098 13030 26110 13082
rect 26172 13030 26174 13082
rect 26012 13028 26036 13030
rect 26092 13028 26116 13030
rect 26172 13028 26196 13030
rect 25956 13008 26252 13028
rect 26148 12912 26200 12918
rect 25962 12880 26018 12889
rect 26148 12854 26200 12860
rect 25962 12815 26018 12824
rect 25976 12782 26004 12815
rect 25964 12776 26016 12782
rect 25964 12718 26016 12724
rect 26160 12374 26188 12854
rect 26148 12368 26200 12374
rect 26344 12345 26372 15302
rect 26436 12866 26464 19110
rect 26988 19009 27016 19178
rect 27160 19168 27212 19174
rect 27160 19110 27212 19116
rect 26974 19000 27030 19009
rect 27172 18970 27200 19110
rect 26974 18935 27030 18944
rect 27160 18964 27212 18970
rect 27160 18906 27212 18912
rect 26514 18184 26570 18193
rect 26514 18119 26570 18128
rect 26528 16658 26556 18119
rect 26516 16652 26568 16658
rect 26516 16594 26568 16600
rect 26528 16250 26556 16594
rect 26516 16244 26568 16250
rect 26516 16186 26568 16192
rect 26792 15360 26844 15366
rect 26792 15302 26844 15308
rect 26516 13728 26568 13734
rect 26516 13670 26568 13676
rect 26528 13326 26556 13670
rect 26516 13320 26568 13326
rect 26516 13262 26568 13268
rect 26528 12986 26556 13262
rect 26516 12980 26568 12986
rect 26516 12922 26568 12928
rect 26436 12838 26556 12866
rect 26424 12708 26476 12714
rect 26424 12650 26476 12656
rect 26148 12310 26200 12316
rect 26330 12336 26386 12345
rect 26330 12271 26386 12280
rect 25956 11996 26252 12016
rect 26012 11994 26036 11996
rect 26092 11994 26116 11996
rect 26172 11994 26196 11996
rect 26034 11942 26036 11994
rect 26098 11942 26110 11994
rect 26172 11942 26174 11994
rect 26012 11940 26036 11942
rect 26092 11940 26116 11942
rect 26172 11940 26196 11942
rect 25956 11920 26252 11940
rect 26238 11656 26294 11665
rect 26238 11591 26294 11600
rect 26252 11558 26280 11591
rect 26240 11552 26292 11558
rect 26240 11494 26292 11500
rect 26436 11286 26464 12650
rect 26424 11280 26476 11286
rect 26422 11248 26424 11257
rect 26476 11248 26478 11257
rect 26422 11183 26478 11192
rect 26436 11157 26464 11183
rect 25870 11112 25926 11121
rect 25870 11047 25926 11056
rect 25956 10908 26252 10928
rect 26012 10906 26036 10908
rect 26092 10906 26116 10908
rect 26172 10906 26196 10908
rect 26034 10854 26036 10906
rect 26098 10854 26110 10906
rect 26172 10854 26174 10906
rect 26012 10852 26036 10854
rect 26092 10852 26116 10854
rect 26172 10852 26196 10854
rect 25956 10832 26252 10852
rect 26424 10600 26476 10606
rect 26422 10568 26424 10577
rect 26476 10568 26478 10577
rect 26422 10503 26478 10512
rect 26528 10130 26556 12838
rect 26698 11656 26754 11665
rect 26698 11591 26754 11600
rect 26712 11082 26740 11591
rect 26700 11076 26752 11082
rect 26700 11018 26752 11024
rect 26608 10464 26660 10470
rect 26606 10432 26608 10441
rect 26660 10432 26662 10441
rect 26606 10367 26662 10376
rect 26516 10124 26568 10130
rect 26516 10066 26568 10072
rect 25872 10056 25924 10062
rect 25872 9998 25924 10004
rect 25884 9586 25912 9998
rect 25956 9820 26252 9840
rect 26012 9818 26036 9820
rect 26092 9818 26116 9820
rect 26172 9818 26196 9820
rect 26034 9766 26036 9818
rect 26098 9766 26110 9818
rect 26172 9766 26174 9818
rect 26012 9764 26036 9766
rect 26092 9764 26116 9766
rect 26172 9764 26196 9766
rect 25956 9744 26252 9764
rect 26528 9722 26556 10066
rect 26700 9920 26752 9926
rect 26698 9888 26700 9897
rect 26752 9888 26754 9897
rect 26698 9823 26754 9832
rect 26516 9716 26568 9722
rect 26516 9658 26568 9664
rect 25872 9580 25924 9586
rect 25872 9522 25924 9528
rect 26332 9580 26384 9586
rect 26332 9522 26384 9528
rect 25964 9444 26016 9450
rect 25964 9386 26016 9392
rect 25872 9376 25924 9382
rect 25872 9318 25924 9324
rect 25884 9110 25912 9318
rect 25872 9104 25924 9110
rect 25872 9046 25924 9052
rect 25872 8968 25924 8974
rect 25870 8936 25872 8945
rect 25924 8936 25926 8945
rect 25976 8922 26004 9386
rect 25926 8894 26004 8922
rect 25870 8871 25926 8880
rect 25956 8732 26252 8752
rect 26012 8730 26036 8732
rect 26092 8730 26116 8732
rect 26172 8730 26196 8732
rect 26034 8678 26036 8730
rect 26098 8678 26110 8730
rect 26172 8678 26174 8730
rect 26012 8676 26036 8678
rect 26092 8676 26116 8678
rect 26172 8676 26196 8678
rect 25956 8656 26252 8676
rect 25956 7644 26252 7664
rect 26012 7642 26036 7644
rect 26092 7642 26116 7644
rect 26172 7642 26196 7644
rect 26034 7590 26036 7642
rect 26098 7590 26110 7642
rect 26172 7590 26174 7642
rect 26012 7588 26036 7590
rect 26092 7588 26116 7590
rect 26172 7588 26196 7590
rect 25956 7568 26252 7588
rect 26344 7478 26372 9522
rect 26528 9518 26556 9658
rect 26516 9512 26568 9518
rect 26516 9454 26568 9460
rect 26606 9344 26662 9353
rect 26606 9279 26662 9288
rect 26620 8634 26648 9279
rect 26698 8664 26754 8673
rect 26608 8628 26660 8634
rect 26698 8599 26754 8608
rect 26608 8570 26660 8576
rect 26424 8424 26476 8430
rect 26424 8366 26476 8372
rect 26332 7472 26384 7478
rect 26332 7414 26384 7420
rect 26330 7032 26386 7041
rect 26330 6967 26386 6976
rect 25594 6896 25650 6905
rect 25594 6831 25650 6840
rect 25778 6896 25834 6905
rect 25778 6831 25834 6840
rect 25044 6656 25096 6662
rect 25044 6598 25096 6604
rect 25056 5370 25084 6598
rect 25956 6556 26252 6576
rect 26012 6554 26036 6556
rect 26092 6554 26116 6556
rect 26172 6554 26196 6556
rect 26034 6502 26036 6554
rect 26098 6502 26110 6554
rect 26172 6502 26174 6554
rect 26012 6500 26036 6502
rect 26092 6500 26116 6502
rect 26172 6500 26196 6502
rect 25956 6480 26252 6500
rect 26238 6216 26294 6225
rect 26238 6151 26240 6160
rect 26292 6151 26294 6160
rect 26240 6122 26292 6128
rect 25956 5468 26252 5488
rect 26012 5466 26036 5468
rect 26092 5466 26116 5468
rect 26172 5466 26196 5468
rect 26034 5414 26036 5466
rect 26098 5414 26110 5466
rect 26172 5414 26174 5466
rect 26012 5412 26036 5414
rect 26092 5412 26116 5414
rect 26172 5412 26196 5414
rect 25956 5392 26252 5412
rect 25044 5364 25096 5370
rect 25044 5306 25096 5312
rect 26238 5128 26294 5137
rect 26238 5063 26240 5072
rect 26292 5063 26294 5072
rect 26240 5034 26292 5040
rect 25956 4380 26252 4400
rect 26012 4378 26036 4380
rect 26092 4378 26116 4380
rect 26172 4378 26196 4380
rect 26034 4326 26036 4378
rect 26098 4326 26110 4378
rect 26172 4326 26174 4378
rect 26012 4324 26036 4326
rect 26092 4324 26116 4326
rect 26172 4324 26196 4326
rect 25956 4304 26252 4324
rect 26344 3924 26372 6967
rect 26436 5817 26464 8366
rect 26712 8090 26740 8599
rect 26700 8084 26752 8090
rect 26700 8026 26752 8032
rect 26514 7984 26570 7993
rect 26514 7919 26516 7928
rect 26568 7919 26570 7928
rect 26516 7890 26568 7896
rect 26528 7546 26556 7890
rect 26516 7540 26568 7546
rect 26516 7482 26568 7488
rect 26514 7440 26570 7449
rect 26514 7375 26570 7384
rect 26698 7440 26754 7449
rect 26698 7375 26754 7384
rect 26422 5808 26478 5817
rect 26528 5778 26556 7375
rect 26712 6730 26740 7375
rect 26700 6724 26752 6730
rect 26700 6666 26752 6672
rect 26804 6361 26832 15302
rect 26882 12744 26938 12753
rect 26882 12679 26938 12688
rect 26896 12646 26924 12679
rect 26884 12640 26936 12646
rect 26884 12582 26936 12588
rect 26896 12306 26924 12582
rect 26884 12300 26936 12306
rect 26884 12242 26936 12248
rect 26896 11898 26924 12242
rect 26884 11892 26936 11898
rect 26884 11834 26936 11840
rect 27068 11688 27120 11694
rect 27068 11630 27120 11636
rect 27264 11642 27292 20198
rect 27344 15564 27396 15570
rect 27344 15506 27396 15512
rect 27356 15162 27384 15506
rect 27344 15156 27396 15162
rect 27344 15098 27396 15104
rect 27344 12980 27396 12986
rect 27344 12922 27396 12928
rect 27356 11778 27384 12922
rect 27448 11914 27476 20198
rect 27540 19310 27568 21791
rect 28276 20602 28304 23520
rect 28264 20596 28316 20602
rect 28264 20538 28316 20544
rect 27528 19304 27580 19310
rect 27528 19246 27580 19252
rect 27526 14104 27582 14113
rect 27526 14039 27582 14048
rect 27540 13297 27568 14039
rect 27526 13288 27582 13297
rect 27526 13223 27582 13232
rect 27540 12782 27568 13223
rect 27528 12776 27580 12782
rect 27528 12718 27580 12724
rect 27540 12442 27568 12718
rect 27528 12436 27580 12442
rect 27528 12378 27580 12384
rect 27448 11886 27568 11914
rect 27356 11762 27476 11778
rect 27356 11756 27488 11762
rect 27356 11750 27436 11756
rect 27436 11698 27488 11704
rect 27080 11286 27108 11630
rect 27264 11614 27384 11642
rect 27252 11552 27304 11558
rect 27252 11494 27304 11500
rect 27264 11354 27292 11494
rect 27252 11348 27304 11354
rect 27252 11290 27304 11296
rect 27068 11280 27120 11286
rect 27068 11222 27120 11228
rect 27252 11212 27304 11218
rect 27252 11154 27304 11160
rect 27264 10810 27292 11154
rect 27252 10804 27304 10810
rect 27252 10746 27304 10752
rect 26976 6860 27028 6866
rect 26976 6802 27028 6808
rect 26988 6769 27016 6802
rect 26974 6760 27030 6769
rect 26974 6695 27030 6704
rect 26988 6458 27016 6695
rect 26976 6452 27028 6458
rect 26976 6394 27028 6400
rect 26790 6352 26846 6361
rect 26790 6287 26846 6296
rect 26608 6112 26660 6118
rect 26608 6054 26660 6060
rect 26422 5743 26478 5752
rect 26516 5772 26568 5778
rect 26516 5714 26568 5720
rect 26620 5681 26648 6054
rect 26976 5772 27028 5778
rect 26976 5714 27028 5720
rect 26606 5672 26662 5681
rect 26606 5607 26662 5616
rect 26792 5568 26844 5574
rect 26792 5510 26844 5516
rect 26606 5128 26662 5137
rect 26606 5063 26662 5072
rect 26620 5030 26648 5063
rect 26608 5024 26660 5030
rect 26608 4966 26660 4972
rect 26514 4720 26570 4729
rect 26514 4655 26516 4664
rect 26568 4655 26570 4664
rect 26516 4626 26568 4632
rect 26528 4282 26556 4626
rect 26516 4276 26568 4282
rect 26516 4218 26568 4224
rect 26424 4072 26476 4078
rect 26422 4040 26424 4049
rect 26476 4040 26478 4049
rect 26422 3975 26478 3984
rect 26700 3936 26752 3942
rect 26344 3896 26464 3924
rect 25956 3292 26252 3312
rect 26012 3290 26036 3292
rect 26092 3290 26116 3292
rect 26172 3290 26196 3292
rect 26034 3238 26036 3290
rect 26098 3238 26110 3290
rect 26172 3238 26174 3290
rect 26012 3236 26036 3238
rect 26092 3236 26116 3238
rect 26172 3236 26196 3238
rect 25956 3216 26252 3236
rect 26332 3120 26384 3126
rect 25686 3088 25742 3097
rect 26332 3062 26384 3068
rect 25686 3023 25742 3032
rect 24952 2984 25004 2990
rect 24952 2926 25004 2932
rect 25700 2514 25728 3023
rect 25688 2508 25740 2514
rect 25688 2450 25740 2456
rect 25872 2304 25924 2310
rect 25872 2246 25924 2252
rect 25884 921 25912 2246
rect 25956 2204 26252 2224
rect 26012 2202 26036 2204
rect 26092 2202 26116 2204
rect 26172 2202 26196 2204
rect 26034 2150 26036 2202
rect 26098 2150 26110 2202
rect 26172 2150 26174 2202
rect 26012 2148 26036 2150
rect 26092 2148 26116 2150
rect 26172 2148 26196 2150
rect 25956 2128 26252 2148
rect 25870 912 25926 921
rect 25870 847 25926 856
rect 26344 480 26372 3062
rect 26436 2990 26464 3896
rect 26804 3913 26832 5510
rect 26988 5370 27016 5714
rect 26976 5364 27028 5370
rect 26976 5306 27028 5312
rect 27356 4826 27384 11614
rect 27448 11354 27476 11698
rect 27436 11348 27488 11354
rect 27436 11290 27488 11296
rect 27540 10792 27568 11886
rect 27448 10764 27568 10792
rect 27344 4820 27396 4826
rect 27344 4762 27396 4768
rect 26884 4480 26936 4486
rect 26884 4422 26936 4428
rect 26700 3878 26752 3884
rect 26790 3904 26846 3913
rect 26424 2984 26476 2990
rect 26424 2926 26476 2932
rect 26608 2848 26660 2854
rect 26712 2825 26740 3878
rect 26790 3839 26846 3848
rect 26792 3392 26844 3398
rect 26896 3369 26924 4422
rect 27448 3777 27476 10764
rect 27526 10704 27582 10713
rect 27526 10639 27582 10648
rect 27540 10606 27568 10639
rect 27528 10600 27580 10606
rect 27528 10542 27580 10548
rect 27712 10464 27764 10470
rect 27712 10406 27764 10412
rect 27724 8129 27752 10406
rect 27710 8120 27766 8129
rect 27710 8055 27766 8064
rect 27804 4820 27856 4826
rect 27804 4762 27856 4768
rect 27710 4448 27766 4457
rect 27710 4383 27766 4392
rect 27724 3942 27752 4383
rect 27712 3936 27764 3942
rect 27712 3878 27764 3884
rect 27434 3768 27490 3777
rect 27434 3703 27490 3712
rect 27526 3632 27582 3641
rect 27344 3596 27396 3602
rect 27526 3567 27582 3576
rect 27344 3538 27396 3544
rect 26792 3334 26844 3340
rect 26882 3360 26938 3369
rect 26608 2790 26660 2796
rect 26698 2816 26754 2825
rect 3974 368 4030 377
rect 3974 303 4030 312
rect 4894 0 4950 480
rect 6366 0 6422 480
rect 7746 0 7802 480
rect 9218 0 9274 480
rect 10598 0 10654 480
rect 12070 0 12126 480
rect 13450 0 13506 480
rect 14922 0 14978 480
rect 16302 0 16358 480
rect 17774 0 17830 480
rect 19154 0 19210 480
rect 20626 0 20682 480
rect 22006 0 22062 480
rect 23478 0 23534 480
rect 24858 0 24914 480
rect 26330 0 26386 480
rect 26620 377 26648 2790
rect 26698 2751 26754 2760
rect 26804 1465 26832 3334
rect 26882 3295 26938 3304
rect 27356 3194 27384 3538
rect 27344 3188 27396 3194
rect 27344 3130 27396 3136
rect 27540 2990 27568 3567
rect 27528 2984 27580 2990
rect 27528 2926 27580 2932
rect 27712 2848 27764 2854
rect 27712 2790 27764 2796
rect 27724 2145 27752 2790
rect 27710 2136 27766 2145
rect 27710 2071 27766 2080
rect 27816 1986 27844 4762
rect 29184 2304 29236 2310
rect 29184 2246 29236 2252
rect 27724 1958 27844 1986
rect 26790 1456 26846 1465
rect 26790 1391 26846 1400
rect 27724 480 27752 1958
rect 29196 480 29224 2246
rect 26606 368 26662 377
rect 26606 303 26662 312
rect 27710 0 27766 480
rect 29182 0 29238 480
<< via2 >>
rect 3974 23568 4030 23624
rect 2870 22344 2926 22400
rect 2042 17992 2098 18048
rect 1398 17740 1454 17776
rect 1398 17720 1400 17740
rect 1400 17720 1452 17740
rect 1452 17720 1454 17740
rect 2778 15816 2834 15872
rect 1490 12144 1546 12200
rect 1398 11056 1454 11112
rect 1582 10376 1638 10432
rect 1674 9424 1730 9480
rect 1582 9288 1638 9344
rect 1490 8608 1546 8664
rect 1398 8064 1454 8120
rect 1582 7384 1638 7440
rect 1766 6840 1822 6896
rect 1582 5616 1638 5672
rect 1582 5072 1638 5128
rect 1858 5072 1914 5128
rect 1582 4392 1638 4448
rect 25870 23568 25926 23624
rect 4250 23024 4306 23080
rect 4066 21800 4122 21856
rect 3238 20576 3294 20632
rect 3330 20032 3386 20088
rect 5956 21786 6012 21788
rect 6036 21786 6092 21788
rect 6116 21786 6172 21788
rect 6196 21786 6252 21788
rect 5956 21734 5982 21786
rect 5982 21734 6012 21786
rect 6036 21734 6046 21786
rect 6046 21734 6092 21786
rect 6116 21734 6162 21786
rect 6162 21734 6172 21786
rect 6196 21734 6226 21786
rect 6226 21734 6252 21786
rect 5956 21732 6012 21734
rect 6036 21732 6092 21734
rect 6116 21732 6172 21734
rect 6196 21732 6252 21734
rect 7286 21256 7342 21312
rect 5956 20698 6012 20700
rect 6036 20698 6092 20700
rect 6116 20698 6172 20700
rect 6196 20698 6252 20700
rect 5956 20646 5982 20698
rect 5982 20646 6012 20698
rect 6036 20646 6046 20698
rect 6046 20646 6092 20698
rect 6116 20646 6162 20698
rect 6162 20646 6172 20698
rect 6196 20646 6226 20698
rect 6226 20646 6252 20698
rect 5956 20644 6012 20646
rect 6036 20644 6092 20646
rect 6116 20644 6172 20646
rect 6196 20644 6252 20646
rect 4986 20304 5042 20360
rect 5956 19610 6012 19612
rect 6036 19610 6092 19612
rect 6116 19610 6172 19612
rect 6196 19610 6252 19612
rect 5956 19558 5982 19610
rect 5982 19558 6012 19610
rect 6036 19558 6046 19610
rect 6046 19558 6092 19610
rect 6116 19558 6162 19610
rect 6162 19558 6172 19610
rect 6196 19558 6226 19610
rect 6226 19558 6252 19610
rect 5956 19556 6012 19558
rect 6036 19556 6092 19558
rect 6116 19556 6172 19558
rect 6196 19556 6252 19558
rect 5354 19080 5410 19136
rect 4986 18808 5042 18864
rect 4250 18148 4306 18184
rect 4250 18128 4252 18148
rect 4252 18128 4304 18148
rect 4304 18128 4306 18148
rect 4710 18264 4766 18320
rect 3422 17584 3478 17640
rect 3146 17040 3202 17096
rect 3238 16768 3294 16824
rect 3146 15408 3202 15464
rect 3238 14864 3294 14920
rect 2870 12144 2926 12200
rect 3238 12552 3294 12608
rect 2686 11600 2742 11656
rect 2686 11212 2742 11248
rect 2686 11192 2688 11212
rect 2688 11192 2740 11212
rect 2740 11192 2742 11212
rect 2502 10240 2558 10296
rect 2686 9868 2688 9888
rect 2688 9868 2740 9888
rect 2740 9868 2742 9888
rect 2686 9832 2742 9868
rect 2042 9580 2098 9616
rect 2042 9560 2044 9580
rect 2044 9560 2096 9580
rect 2096 9560 2098 9580
rect 2502 6840 2558 6896
rect 2042 6452 2098 6488
rect 2042 6432 2044 6452
rect 2044 6432 2096 6452
rect 2096 6432 2098 6452
rect 2042 5228 2098 5264
rect 2042 5208 2044 5228
rect 2044 5208 2096 5228
rect 2096 5208 2098 5228
rect 2042 4684 2098 4720
rect 2962 11736 3018 11792
rect 2870 8492 2926 8528
rect 2870 8472 2872 8492
rect 2872 8472 2924 8492
rect 2924 8472 2926 8492
rect 2778 7964 2780 7984
rect 2780 7964 2832 7984
rect 2832 7964 2834 7984
rect 2778 7928 2834 7964
rect 2962 6976 3018 7032
rect 2042 4664 2044 4684
rect 2044 4664 2096 4684
rect 2096 4664 2098 4684
rect 1950 4120 2006 4176
rect 3422 11600 3478 11656
rect 3606 15952 3662 16008
rect 3606 13368 3662 13424
rect 3514 10648 3570 10704
rect 4526 17992 4582 18048
rect 4710 17992 4766 18048
rect 4066 17176 4122 17232
rect 4526 16496 4582 16552
rect 3882 16360 3938 16416
rect 4434 15700 4490 15736
rect 4434 15680 4436 15700
rect 4436 15680 4488 15700
rect 4488 15680 4490 15700
rect 3882 13640 3938 13696
rect 3974 12552 4030 12608
rect 3974 12280 4030 12336
rect 3330 7520 3386 7576
rect 3422 4120 3478 4176
rect 2686 3848 2742 3904
rect 662 2896 718 2952
rect 3330 3068 3332 3088
rect 3332 3068 3384 3088
rect 3384 3068 3386 3088
rect 3330 3032 3386 3068
rect 3698 6296 3754 6352
rect 4802 14048 4858 14104
rect 5956 18522 6012 18524
rect 6036 18522 6092 18524
rect 6116 18522 6172 18524
rect 6196 18522 6252 18524
rect 5956 18470 5982 18522
rect 5982 18470 6012 18522
rect 6036 18470 6046 18522
rect 6046 18470 6092 18522
rect 6116 18470 6162 18522
rect 6162 18470 6172 18522
rect 6196 18470 6226 18522
rect 6226 18470 6252 18522
rect 5956 18468 6012 18470
rect 6036 18468 6092 18470
rect 6116 18468 6172 18470
rect 6196 18468 6252 18470
rect 5170 17620 5172 17640
rect 5172 17620 5224 17640
rect 5224 17620 5226 17640
rect 5170 17584 5226 17620
rect 5956 17434 6012 17436
rect 6036 17434 6092 17436
rect 6116 17434 6172 17436
rect 6196 17434 6252 17436
rect 5956 17382 5982 17434
rect 5982 17382 6012 17434
rect 6036 17382 6046 17434
rect 6046 17382 6092 17434
rect 6116 17382 6162 17434
rect 6162 17382 6172 17434
rect 6196 17382 6226 17434
rect 6226 17382 6252 17434
rect 5956 17380 6012 17382
rect 6036 17380 6092 17382
rect 6116 17380 6172 17382
rect 6196 17380 6252 17382
rect 5814 17176 5870 17232
rect 5078 16652 5134 16688
rect 5078 16632 5080 16652
rect 5080 16632 5132 16652
rect 5132 16632 5134 16652
rect 6826 16788 6882 16824
rect 6826 16768 6828 16788
rect 6828 16768 6880 16788
rect 6880 16768 6882 16788
rect 5956 16346 6012 16348
rect 6036 16346 6092 16348
rect 6116 16346 6172 16348
rect 6196 16346 6252 16348
rect 5956 16294 5982 16346
rect 5982 16294 6012 16346
rect 6036 16294 6046 16346
rect 6046 16294 6092 16346
rect 6116 16294 6162 16346
rect 6162 16294 6172 16346
rect 6196 16294 6226 16346
rect 6226 16294 6252 16346
rect 5956 16292 6012 16294
rect 6036 16292 6092 16294
rect 6116 16292 6172 16294
rect 6196 16292 6252 16294
rect 5538 15272 5594 15328
rect 4342 12552 4398 12608
rect 4894 12552 4950 12608
rect 5956 15258 6012 15260
rect 6036 15258 6092 15260
rect 6116 15258 6172 15260
rect 6196 15258 6252 15260
rect 5956 15206 5982 15258
rect 5982 15206 6012 15258
rect 6036 15206 6046 15258
rect 6046 15206 6092 15258
rect 6116 15206 6162 15258
rect 6162 15206 6172 15258
rect 6196 15206 6226 15258
rect 6226 15206 6252 15258
rect 5956 15204 6012 15206
rect 6036 15204 6092 15206
rect 6116 15204 6172 15206
rect 6196 15204 6252 15206
rect 5956 14170 6012 14172
rect 6036 14170 6092 14172
rect 6116 14170 6172 14172
rect 6196 14170 6252 14172
rect 5956 14118 5982 14170
rect 5982 14118 6012 14170
rect 6036 14118 6046 14170
rect 6046 14118 6092 14170
rect 6116 14118 6162 14170
rect 6162 14118 6172 14170
rect 6196 14118 6226 14170
rect 6226 14118 6252 14170
rect 5956 14116 6012 14118
rect 6036 14116 6092 14118
rect 6116 14116 6172 14118
rect 6196 14116 6252 14118
rect 5538 11328 5594 11384
rect 4066 3596 4122 3632
rect 4066 3576 4068 3596
rect 4068 3576 4120 3596
rect 4120 3576 4122 3596
rect 2134 1400 2190 1456
rect 4066 2624 4122 2680
rect 4618 6976 4674 7032
rect 4986 7540 5042 7576
rect 4986 7520 4988 7540
rect 4988 7520 5040 7540
rect 5040 7520 5042 7540
rect 5446 6452 5502 6488
rect 5446 6432 5448 6452
rect 5448 6432 5500 6452
rect 5500 6432 5502 6452
rect 5630 7268 5686 7304
rect 5630 7248 5632 7268
rect 5632 7248 5684 7268
rect 5684 7248 5686 7268
rect 5630 6876 5632 6896
rect 5632 6876 5684 6896
rect 5684 6876 5686 6896
rect 5630 6840 5686 6876
rect 5956 13082 6012 13084
rect 6036 13082 6092 13084
rect 6116 13082 6172 13084
rect 6196 13082 6252 13084
rect 5956 13030 5982 13082
rect 5982 13030 6012 13082
rect 6036 13030 6046 13082
rect 6046 13030 6092 13082
rect 6116 13030 6162 13082
rect 6162 13030 6172 13082
rect 6196 13030 6226 13082
rect 6226 13030 6252 13082
rect 5956 13028 6012 13030
rect 6036 13028 6092 13030
rect 6116 13028 6172 13030
rect 6196 13028 6252 13030
rect 6366 12688 6422 12744
rect 5998 12300 6054 12336
rect 5998 12280 6000 12300
rect 6000 12280 6052 12300
rect 6052 12280 6054 12300
rect 6274 12280 6330 12336
rect 5956 11994 6012 11996
rect 6036 11994 6092 11996
rect 6116 11994 6172 11996
rect 6196 11994 6252 11996
rect 5956 11942 5982 11994
rect 5982 11942 6012 11994
rect 6036 11942 6046 11994
rect 6046 11942 6092 11994
rect 6116 11942 6162 11994
rect 6162 11942 6172 11994
rect 6196 11942 6226 11994
rect 6226 11942 6252 11994
rect 5956 11940 6012 11942
rect 6036 11940 6092 11942
rect 6116 11940 6172 11942
rect 6196 11940 6252 11942
rect 10956 21242 11012 21244
rect 11036 21242 11092 21244
rect 11116 21242 11172 21244
rect 11196 21242 11252 21244
rect 10956 21190 10982 21242
rect 10982 21190 11012 21242
rect 11036 21190 11046 21242
rect 11046 21190 11092 21242
rect 11116 21190 11162 21242
rect 11162 21190 11172 21242
rect 11196 21190 11226 21242
rect 11226 21190 11252 21242
rect 10956 21188 11012 21190
rect 11036 21188 11092 21190
rect 11116 21188 11172 21190
rect 11196 21188 11252 21190
rect 8758 20460 8814 20496
rect 8758 20440 8760 20460
rect 8760 20440 8812 20460
rect 8812 20440 8814 20460
rect 8022 19896 8078 19952
rect 12438 20460 12494 20496
rect 12438 20440 12440 20460
rect 12440 20440 12492 20460
rect 12492 20440 12494 20460
rect 10956 20154 11012 20156
rect 11036 20154 11092 20156
rect 11116 20154 11172 20156
rect 11196 20154 11252 20156
rect 10956 20102 10982 20154
rect 10982 20102 11012 20154
rect 11036 20102 11046 20154
rect 11046 20102 11092 20154
rect 11116 20102 11162 20154
rect 11162 20102 11172 20154
rect 11196 20102 11226 20154
rect 11226 20102 11252 20154
rect 10956 20100 11012 20102
rect 11036 20100 11092 20102
rect 11116 20100 11172 20102
rect 11196 20100 11252 20102
rect 10506 19252 10508 19272
rect 10508 19252 10560 19272
rect 10560 19252 10562 19272
rect 10506 19216 10562 19252
rect 10598 19116 10600 19136
rect 10600 19116 10652 19136
rect 10652 19116 10654 19136
rect 10598 19080 10654 19116
rect 10874 19780 10930 19816
rect 10874 19760 10876 19780
rect 10876 19760 10928 19780
rect 10928 19760 10930 19780
rect 10956 19066 11012 19068
rect 11036 19066 11092 19068
rect 11116 19066 11172 19068
rect 11196 19066 11252 19068
rect 10956 19014 10982 19066
rect 10982 19014 11012 19066
rect 11036 19014 11046 19066
rect 11046 19014 11092 19066
rect 11116 19014 11162 19066
rect 11162 19014 11172 19066
rect 11196 19014 11226 19066
rect 11226 19014 11252 19066
rect 10956 19012 11012 19014
rect 11036 19012 11092 19014
rect 11116 19012 11172 19014
rect 11196 19012 11252 19014
rect 10046 18264 10102 18320
rect 9678 18028 9680 18048
rect 9680 18028 9732 18048
rect 9732 18028 9734 18048
rect 9678 17992 9734 18028
rect 9678 17176 9734 17232
rect 9586 16632 9642 16688
rect 6734 13640 6790 13696
rect 6642 12416 6698 12472
rect 5956 10906 6012 10908
rect 6036 10906 6092 10908
rect 6116 10906 6172 10908
rect 6196 10906 6252 10908
rect 5956 10854 5982 10906
rect 5982 10854 6012 10906
rect 6036 10854 6046 10906
rect 6046 10854 6092 10906
rect 6116 10854 6162 10906
rect 6162 10854 6172 10906
rect 6196 10854 6226 10906
rect 6226 10854 6252 10906
rect 5956 10852 6012 10854
rect 6036 10852 6092 10854
rect 6116 10852 6172 10854
rect 6196 10852 6252 10854
rect 6274 10512 6330 10568
rect 8298 13640 8354 13696
rect 5956 9818 6012 9820
rect 6036 9818 6092 9820
rect 6116 9818 6172 9820
rect 6196 9818 6252 9820
rect 5956 9766 5982 9818
rect 5982 9766 6012 9818
rect 6036 9766 6046 9818
rect 6046 9766 6092 9818
rect 6116 9766 6162 9818
rect 6162 9766 6172 9818
rect 6196 9766 6226 9818
rect 6226 9766 6252 9818
rect 5956 9764 6012 9766
rect 6036 9764 6092 9766
rect 6116 9764 6172 9766
rect 6196 9764 6252 9766
rect 5956 8730 6012 8732
rect 6036 8730 6092 8732
rect 6116 8730 6172 8732
rect 6196 8730 6252 8732
rect 5956 8678 5982 8730
rect 5982 8678 6012 8730
rect 6036 8678 6046 8730
rect 6046 8678 6092 8730
rect 6116 8678 6162 8730
rect 6162 8678 6172 8730
rect 6196 8678 6226 8730
rect 6226 8678 6252 8730
rect 5956 8676 6012 8678
rect 6036 8676 6092 8678
rect 6116 8676 6172 8678
rect 6196 8676 6252 8678
rect 6734 10512 6790 10568
rect 6458 10376 6514 10432
rect 6550 9460 6552 9480
rect 6552 9460 6604 9480
rect 6604 9460 6606 9480
rect 6550 9424 6606 9460
rect 5956 7642 6012 7644
rect 6036 7642 6092 7644
rect 6116 7642 6172 7644
rect 6196 7642 6252 7644
rect 5956 7590 5982 7642
rect 5982 7590 6012 7642
rect 6036 7590 6046 7642
rect 6046 7590 6092 7642
rect 6116 7590 6162 7642
rect 6162 7590 6172 7642
rect 6196 7590 6226 7642
rect 6226 7590 6252 7642
rect 5956 7588 6012 7590
rect 6036 7588 6092 7590
rect 6116 7588 6172 7590
rect 6196 7588 6252 7590
rect 5998 6860 6054 6896
rect 5998 6840 6000 6860
rect 6000 6840 6052 6860
rect 6052 6840 6054 6860
rect 5956 6554 6012 6556
rect 6036 6554 6092 6556
rect 6116 6554 6172 6556
rect 6196 6554 6252 6556
rect 5956 6502 5982 6554
rect 5982 6502 6012 6554
rect 6036 6502 6046 6554
rect 6046 6502 6092 6554
rect 6116 6502 6162 6554
rect 6162 6502 6172 6554
rect 6196 6502 6226 6554
rect 6226 6502 6252 6554
rect 5956 6500 6012 6502
rect 6036 6500 6092 6502
rect 6116 6500 6172 6502
rect 6196 6500 6252 6502
rect 5956 5466 6012 5468
rect 6036 5466 6092 5468
rect 6116 5466 6172 5468
rect 6196 5466 6252 5468
rect 5956 5414 5982 5466
rect 5982 5414 6012 5466
rect 6036 5414 6046 5466
rect 6046 5414 6092 5466
rect 6116 5414 6162 5466
rect 6162 5414 6172 5466
rect 6196 5414 6226 5466
rect 6226 5414 6252 5466
rect 5956 5412 6012 5414
rect 6036 5412 6092 5414
rect 6116 5412 6172 5414
rect 6196 5412 6252 5414
rect 6458 5208 6514 5264
rect 9770 15408 9826 15464
rect 9862 14592 9918 14648
rect 8390 12280 8446 12336
rect 9586 13096 9642 13152
rect 9586 12960 9642 13016
rect 9586 12844 9642 12880
rect 9586 12824 9588 12844
rect 9588 12824 9640 12844
rect 9640 12824 9642 12844
rect 9310 12688 9366 12744
rect 9494 12724 9496 12744
rect 9496 12724 9548 12744
rect 9548 12724 9550 12744
rect 9494 12688 9550 12724
rect 9678 12280 9734 12336
rect 9678 11328 9734 11384
rect 8390 10412 8392 10432
rect 8392 10412 8444 10432
rect 8444 10412 8446 10432
rect 8390 10376 8446 10412
rect 7286 9052 7288 9072
rect 7288 9052 7340 9072
rect 7340 9052 7342 9072
rect 7286 9016 7342 9052
rect 7746 9560 7802 9616
rect 6642 5228 6698 5264
rect 6642 5208 6644 5228
rect 6644 5208 6696 5228
rect 6696 5208 6698 5228
rect 5956 4378 6012 4380
rect 6036 4378 6092 4380
rect 6116 4378 6172 4380
rect 6196 4378 6252 4380
rect 5956 4326 5982 4378
rect 5982 4326 6012 4378
rect 6036 4326 6046 4378
rect 6046 4326 6092 4378
rect 6116 4326 6162 4378
rect 6162 4326 6172 4378
rect 6196 4326 6226 4378
rect 6226 4326 6252 4378
rect 5956 4324 6012 4326
rect 6036 4324 6092 4326
rect 6116 4324 6172 4326
rect 6196 4324 6252 4326
rect 4618 3984 4674 4040
rect 4434 3576 4490 3632
rect 4250 3440 4306 3496
rect 4526 3304 4582 3360
rect 5814 3848 5870 3904
rect 5956 3290 6012 3292
rect 6036 3290 6092 3292
rect 6116 3290 6172 3292
rect 6196 3290 6252 3292
rect 5956 3238 5982 3290
rect 5982 3238 6012 3290
rect 6036 3238 6046 3290
rect 6046 3238 6092 3290
rect 6116 3238 6162 3290
rect 6162 3238 6172 3290
rect 6196 3238 6226 3290
rect 6226 3238 6252 3290
rect 5956 3236 6012 3238
rect 6036 3236 6092 3238
rect 6116 3236 6172 3238
rect 6196 3236 6252 3238
rect 6550 3052 6606 3088
rect 6550 3032 6552 3052
rect 6552 3032 6604 3052
rect 6604 3032 6606 3052
rect 7930 5788 7932 5808
rect 7932 5788 7984 5808
rect 7984 5788 7986 5808
rect 7930 5752 7986 5788
rect 7654 5208 7710 5264
rect 4066 856 4122 912
rect 5956 2202 6012 2204
rect 6036 2202 6092 2204
rect 6116 2202 6172 2204
rect 6196 2202 6252 2204
rect 5956 2150 5982 2202
rect 5982 2150 6012 2202
rect 6036 2150 6046 2202
rect 6046 2150 6092 2202
rect 6116 2150 6162 2202
rect 6162 2150 6172 2202
rect 6196 2150 6226 2202
rect 6226 2150 6252 2202
rect 5956 2148 6012 2150
rect 6036 2148 6092 2150
rect 6116 2148 6172 2150
rect 6196 2148 6252 2150
rect 5814 2080 5870 2136
rect 9034 3884 9036 3904
rect 9036 3884 9088 3904
rect 9088 3884 9090 3904
rect 9034 3848 9090 3884
rect 10046 12552 10102 12608
rect 10956 17978 11012 17980
rect 11036 17978 11092 17980
rect 11116 17978 11172 17980
rect 11196 17978 11252 17980
rect 10956 17926 10982 17978
rect 10982 17926 11012 17978
rect 11036 17926 11046 17978
rect 11046 17926 11092 17978
rect 11116 17926 11162 17978
rect 11162 17926 11172 17978
rect 11196 17926 11226 17978
rect 11226 17926 11252 17978
rect 10956 17924 11012 17926
rect 11036 17924 11092 17926
rect 11116 17924 11172 17926
rect 11196 17924 11252 17926
rect 10598 17448 10654 17504
rect 10414 16632 10470 16688
rect 10598 16532 10600 16552
rect 10600 16532 10652 16552
rect 10652 16532 10654 16552
rect 10598 16496 10654 16532
rect 11610 17060 11666 17096
rect 11610 17040 11612 17060
rect 11612 17040 11664 17060
rect 11664 17040 11666 17060
rect 12070 17040 12126 17096
rect 10956 16890 11012 16892
rect 11036 16890 11092 16892
rect 11116 16890 11172 16892
rect 11196 16890 11252 16892
rect 10956 16838 10982 16890
rect 10982 16838 11012 16890
rect 11036 16838 11046 16890
rect 11046 16838 11092 16890
rect 11116 16838 11162 16890
rect 11162 16838 11172 16890
rect 11196 16838 11226 16890
rect 11226 16838 11252 16890
rect 10956 16836 11012 16838
rect 11036 16836 11092 16838
rect 11116 16836 11172 16838
rect 11196 16836 11252 16838
rect 11978 16632 12034 16688
rect 10782 15952 10838 16008
rect 10956 15802 11012 15804
rect 11036 15802 11092 15804
rect 11116 15802 11172 15804
rect 11196 15802 11252 15804
rect 10956 15750 10982 15802
rect 10982 15750 11012 15802
rect 11036 15750 11046 15802
rect 11046 15750 11092 15802
rect 11116 15750 11162 15802
rect 11162 15750 11172 15802
rect 11196 15750 11226 15802
rect 11226 15750 11252 15802
rect 10956 15748 11012 15750
rect 11036 15748 11092 15750
rect 11116 15748 11172 15750
rect 11196 15748 11252 15750
rect 10506 15680 10562 15736
rect 11978 15000 12034 15056
rect 10956 14714 11012 14716
rect 11036 14714 11092 14716
rect 11116 14714 11172 14716
rect 11196 14714 11252 14716
rect 10956 14662 10982 14714
rect 10982 14662 11012 14714
rect 11036 14662 11046 14714
rect 11046 14662 11092 14714
rect 11116 14662 11162 14714
rect 11162 14662 11172 14714
rect 11196 14662 11226 14714
rect 11226 14662 11252 14714
rect 10956 14660 11012 14662
rect 11036 14660 11092 14662
rect 11116 14660 11172 14662
rect 11196 14660 11252 14662
rect 10782 13232 10838 13288
rect 10690 13096 10746 13152
rect 10598 12588 10600 12608
rect 10600 12588 10652 12608
rect 10652 12588 10654 12608
rect 10598 12552 10654 12588
rect 9862 10684 9864 10704
rect 9864 10684 9916 10704
rect 9916 10684 9918 10704
rect 9862 10648 9918 10684
rect 9954 10240 10010 10296
rect 10956 13626 11012 13628
rect 11036 13626 11092 13628
rect 11116 13626 11172 13628
rect 11196 13626 11252 13628
rect 10956 13574 10982 13626
rect 10982 13574 11012 13626
rect 11036 13574 11046 13626
rect 11046 13574 11092 13626
rect 11116 13574 11162 13626
rect 11162 13574 11172 13626
rect 11196 13574 11226 13626
rect 11226 13574 11252 13626
rect 10956 13572 11012 13574
rect 11036 13572 11092 13574
rect 11116 13572 11172 13574
rect 11196 13572 11252 13574
rect 11058 13232 11114 13288
rect 10966 12960 11022 13016
rect 11150 12724 11152 12744
rect 11152 12724 11204 12744
rect 11204 12724 11206 12744
rect 11150 12688 11206 12724
rect 10956 12538 11012 12540
rect 11036 12538 11092 12540
rect 11116 12538 11172 12540
rect 11196 12538 11252 12540
rect 10956 12486 10982 12538
rect 10982 12486 11012 12538
rect 11036 12486 11046 12538
rect 11046 12486 11092 12538
rect 11116 12486 11162 12538
rect 11162 12486 11172 12538
rect 11196 12486 11226 12538
rect 11226 12486 11252 12538
rect 10956 12484 11012 12486
rect 11036 12484 11092 12486
rect 11116 12484 11172 12486
rect 11196 12484 11252 12486
rect 10782 12436 10838 12472
rect 11426 12688 11482 12744
rect 10782 12416 10784 12436
rect 10784 12416 10836 12436
rect 10836 12416 10838 12436
rect 11334 11736 11390 11792
rect 10956 11450 11012 11452
rect 11036 11450 11092 11452
rect 11116 11450 11172 11452
rect 11196 11450 11252 11452
rect 10956 11398 10982 11450
rect 10982 11398 11012 11450
rect 11036 11398 11046 11450
rect 11046 11398 11092 11450
rect 11116 11398 11162 11450
rect 11162 11398 11172 11450
rect 11196 11398 11226 11450
rect 11226 11398 11252 11450
rect 10956 11396 11012 11398
rect 11036 11396 11092 11398
rect 11116 11396 11172 11398
rect 11196 11396 11252 11398
rect 11334 11328 11390 11384
rect 11518 11464 11574 11520
rect 11426 11192 11482 11248
rect 10956 10362 11012 10364
rect 11036 10362 11092 10364
rect 11116 10362 11172 10364
rect 11196 10362 11252 10364
rect 10956 10310 10982 10362
rect 10982 10310 11012 10362
rect 11036 10310 11046 10362
rect 11046 10310 11092 10362
rect 11116 10310 11162 10362
rect 11162 10310 11172 10362
rect 11196 10310 11226 10362
rect 11226 10310 11252 10362
rect 10956 10308 11012 10310
rect 11036 10308 11092 10310
rect 11116 10308 11172 10310
rect 11196 10308 11252 10310
rect 10956 9274 11012 9276
rect 11036 9274 11092 9276
rect 11116 9274 11172 9276
rect 11196 9274 11252 9276
rect 10956 9222 10982 9274
rect 10982 9222 11012 9274
rect 11036 9222 11046 9274
rect 11046 9222 11092 9274
rect 11116 9222 11162 9274
rect 11162 9222 11172 9274
rect 11196 9222 11226 9274
rect 11226 9222 11252 9274
rect 10956 9220 11012 9222
rect 11036 9220 11092 9222
rect 11116 9220 11172 9222
rect 11196 9220 11252 9222
rect 10956 8186 11012 8188
rect 11036 8186 11092 8188
rect 11116 8186 11172 8188
rect 11196 8186 11252 8188
rect 10956 8134 10982 8186
rect 10982 8134 11012 8186
rect 11036 8134 11046 8186
rect 11046 8134 11092 8186
rect 11116 8134 11162 8186
rect 11162 8134 11172 8186
rect 11196 8134 11226 8186
rect 11226 8134 11252 8186
rect 10956 8132 11012 8134
rect 11036 8132 11092 8134
rect 11116 8132 11172 8134
rect 11196 8132 11252 8134
rect 10956 7098 11012 7100
rect 11036 7098 11092 7100
rect 11116 7098 11172 7100
rect 11196 7098 11252 7100
rect 10956 7046 10982 7098
rect 10982 7046 11012 7098
rect 11036 7046 11046 7098
rect 11046 7046 11092 7098
rect 11116 7046 11162 7098
rect 11162 7046 11172 7098
rect 11196 7046 11226 7098
rect 11226 7046 11252 7098
rect 10956 7044 11012 7046
rect 11036 7044 11092 7046
rect 11116 7044 11172 7046
rect 11196 7044 11252 7046
rect 10956 6010 11012 6012
rect 11036 6010 11092 6012
rect 11116 6010 11172 6012
rect 11196 6010 11252 6012
rect 10956 5958 10982 6010
rect 10982 5958 11012 6010
rect 11036 5958 11046 6010
rect 11046 5958 11092 6010
rect 11116 5958 11162 6010
rect 11162 5958 11172 6010
rect 11196 5958 11226 6010
rect 11226 5958 11252 6010
rect 10956 5956 11012 5958
rect 11036 5956 11092 5958
rect 11116 5956 11172 5958
rect 11196 5956 11252 5958
rect 10230 5072 10286 5128
rect 10956 4922 11012 4924
rect 11036 4922 11092 4924
rect 11116 4922 11172 4924
rect 11196 4922 11252 4924
rect 10956 4870 10982 4922
rect 10982 4870 11012 4922
rect 11036 4870 11046 4922
rect 11046 4870 11092 4922
rect 11116 4870 11162 4922
rect 11162 4870 11172 4922
rect 11196 4870 11226 4922
rect 11226 4870 11252 4922
rect 10956 4868 11012 4870
rect 11036 4868 11092 4870
rect 11116 4868 11172 4870
rect 11196 4868 11252 4870
rect 11794 7112 11850 7168
rect 15956 21786 16012 21788
rect 16036 21786 16092 21788
rect 16116 21786 16172 21788
rect 16196 21786 16252 21788
rect 15956 21734 15982 21786
rect 15982 21734 16012 21786
rect 16036 21734 16046 21786
rect 16046 21734 16092 21786
rect 16116 21734 16162 21786
rect 16162 21734 16172 21786
rect 16196 21734 16226 21786
rect 16226 21734 16252 21786
rect 15956 21732 16012 21734
rect 16036 21732 16092 21734
rect 16116 21732 16172 21734
rect 16196 21732 16252 21734
rect 15956 20698 16012 20700
rect 16036 20698 16092 20700
rect 16116 20698 16172 20700
rect 16196 20698 16252 20700
rect 15956 20646 15982 20698
rect 15982 20646 16012 20698
rect 16036 20646 16046 20698
rect 16046 20646 16092 20698
rect 16116 20646 16162 20698
rect 16162 20646 16172 20698
rect 16196 20646 16226 20698
rect 16226 20646 16252 20698
rect 15956 20644 16012 20646
rect 16036 20644 16092 20646
rect 16116 20644 16172 20646
rect 16196 20644 16252 20646
rect 20956 21242 21012 21244
rect 21036 21242 21092 21244
rect 21116 21242 21172 21244
rect 21196 21242 21252 21244
rect 20956 21190 20982 21242
rect 20982 21190 21012 21242
rect 21036 21190 21046 21242
rect 21046 21190 21092 21242
rect 21116 21190 21162 21242
rect 21162 21190 21172 21242
rect 21196 21190 21226 21242
rect 21226 21190 21252 21242
rect 20956 21188 21012 21190
rect 21036 21188 21092 21190
rect 21116 21188 21172 21190
rect 21196 21188 21252 21190
rect 16118 20460 16174 20496
rect 16118 20440 16120 20460
rect 16120 20440 16172 20460
rect 16172 20440 16174 20460
rect 18326 20440 18382 20496
rect 14922 20168 14978 20224
rect 15842 19896 15898 19952
rect 14186 19780 14242 19816
rect 14186 19760 14188 19780
rect 14188 19760 14240 19780
rect 14240 19760 14242 19780
rect 13910 19624 13966 19680
rect 13266 17876 13322 17912
rect 13266 17856 13268 17876
rect 13268 17856 13320 17876
rect 13320 17856 13322 17876
rect 12162 7404 12218 7440
rect 12162 7384 12164 7404
rect 12164 7384 12216 7404
rect 12216 7384 12218 7404
rect 11702 4664 11758 4720
rect 10956 3834 11012 3836
rect 11036 3834 11092 3836
rect 11116 3834 11172 3836
rect 11196 3834 11252 3836
rect 10956 3782 10982 3834
rect 10982 3782 11012 3834
rect 11036 3782 11046 3834
rect 11046 3782 11092 3834
rect 11116 3782 11162 3834
rect 11162 3782 11172 3834
rect 11196 3782 11226 3834
rect 11226 3782 11252 3834
rect 10956 3780 11012 3782
rect 11036 3780 11092 3782
rect 11116 3780 11172 3782
rect 11196 3780 11252 3782
rect 11610 4020 11612 4040
rect 11612 4020 11664 4040
rect 11664 4020 11666 4040
rect 11610 3984 11666 4020
rect 12070 3984 12126 4040
rect 12346 3576 12402 3632
rect 9954 3440 10010 3496
rect 10956 2746 11012 2748
rect 11036 2746 11092 2748
rect 11116 2746 11172 2748
rect 11196 2746 11252 2748
rect 10956 2694 10982 2746
rect 10982 2694 11012 2746
rect 11036 2694 11046 2746
rect 11046 2694 11092 2746
rect 11116 2694 11162 2746
rect 11162 2694 11172 2746
rect 11196 2694 11226 2746
rect 11226 2694 11252 2746
rect 10956 2692 11012 2694
rect 11036 2692 11092 2694
rect 11116 2692 11172 2694
rect 11196 2692 11252 2694
rect 15956 19610 16012 19612
rect 16036 19610 16092 19612
rect 16116 19610 16172 19612
rect 16196 19610 16252 19612
rect 15956 19558 15982 19610
rect 15982 19558 16012 19610
rect 16036 19558 16046 19610
rect 16046 19558 16092 19610
rect 16116 19558 16162 19610
rect 16162 19558 16172 19610
rect 16196 19558 16226 19610
rect 16226 19558 16252 19610
rect 15956 19556 16012 19558
rect 16036 19556 16092 19558
rect 16116 19556 16172 19558
rect 16196 19556 16252 19558
rect 16394 19352 16450 19408
rect 15198 17584 15254 17640
rect 13634 15564 13690 15600
rect 13634 15544 13636 15564
rect 13636 15544 13688 15564
rect 13688 15544 13690 15564
rect 12806 15408 12862 15464
rect 12898 12180 12900 12200
rect 12900 12180 12952 12200
rect 12952 12180 12954 12200
rect 12898 12144 12954 12180
rect 13726 13776 13782 13832
rect 13450 12588 13452 12608
rect 13452 12588 13504 12608
rect 13504 12588 13506 12608
rect 13450 12552 13506 12588
rect 13634 12300 13690 12336
rect 14094 13232 14150 13288
rect 14094 12552 14150 12608
rect 13910 12416 13966 12472
rect 14278 13232 14334 13288
rect 13634 12280 13636 12300
rect 13636 12280 13688 12300
rect 13688 12280 13690 12300
rect 13910 12280 13966 12336
rect 12806 7384 12862 7440
rect 13450 6704 13506 6760
rect 13266 4820 13322 4856
rect 13266 4800 13268 4820
rect 13268 4800 13320 4820
rect 13320 4800 13322 4820
rect 13266 4120 13322 4176
rect 15956 18522 16012 18524
rect 16036 18522 16092 18524
rect 16116 18522 16172 18524
rect 16196 18522 16252 18524
rect 15956 18470 15982 18522
rect 15982 18470 16012 18522
rect 16036 18470 16046 18522
rect 16046 18470 16092 18522
rect 16116 18470 16162 18522
rect 16162 18470 16172 18522
rect 16196 18470 16226 18522
rect 16226 18470 16252 18522
rect 15956 18468 16012 18470
rect 16036 18468 16092 18470
rect 16116 18468 16172 18470
rect 16196 18468 16252 18470
rect 15750 18128 15806 18184
rect 15382 17856 15438 17912
rect 16670 17756 16672 17776
rect 16672 17756 16724 17776
rect 16724 17756 16726 17776
rect 16670 17720 16726 17756
rect 15750 17448 15806 17504
rect 15382 16496 15438 16552
rect 15956 17434 16012 17436
rect 16036 17434 16092 17436
rect 16116 17434 16172 17436
rect 16196 17434 16252 17436
rect 15956 17382 15982 17434
rect 15982 17382 16012 17434
rect 16036 17382 16046 17434
rect 16046 17382 16092 17434
rect 16116 17382 16162 17434
rect 16162 17382 16172 17434
rect 16196 17382 16226 17434
rect 16226 17382 16252 17434
rect 15956 17380 16012 17382
rect 16036 17380 16092 17382
rect 16116 17380 16172 17382
rect 16196 17380 16252 17382
rect 16762 17620 16764 17640
rect 16764 17620 16816 17640
rect 16816 17620 16818 17640
rect 16762 17584 16818 17620
rect 15956 16346 16012 16348
rect 16036 16346 16092 16348
rect 16116 16346 16172 16348
rect 16196 16346 16252 16348
rect 15956 16294 15982 16346
rect 15982 16294 16012 16346
rect 16036 16294 16046 16346
rect 16046 16294 16092 16346
rect 16116 16294 16162 16346
rect 16162 16294 16172 16346
rect 16196 16294 16226 16346
rect 16226 16294 16252 16346
rect 15956 16292 16012 16294
rect 16036 16292 16092 16294
rect 16116 16292 16172 16294
rect 16196 16292 16252 16294
rect 16026 15952 16082 16008
rect 15750 15816 15806 15872
rect 15956 15258 16012 15260
rect 16036 15258 16092 15260
rect 16116 15258 16172 15260
rect 16196 15258 16252 15260
rect 15956 15206 15982 15258
rect 15982 15206 16012 15258
rect 16036 15206 16046 15258
rect 16046 15206 16092 15258
rect 16116 15206 16162 15258
rect 16162 15206 16172 15258
rect 16196 15206 16226 15258
rect 16226 15206 16252 15258
rect 15956 15204 16012 15206
rect 16036 15204 16092 15206
rect 16116 15204 16172 15206
rect 16196 15204 16252 15206
rect 15014 13776 15070 13832
rect 14830 13640 14886 13696
rect 15198 13504 15254 13560
rect 15198 13096 15254 13152
rect 15382 13812 15384 13832
rect 15384 13812 15436 13832
rect 15436 13812 15438 13832
rect 15382 13776 15438 13812
rect 15956 14170 16012 14172
rect 16036 14170 16092 14172
rect 16116 14170 16172 14172
rect 16196 14170 16252 14172
rect 15956 14118 15982 14170
rect 15982 14118 16012 14170
rect 16036 14118 16046 14170
rect 16046 14118 16092 14170
rect 16116 14118 16162 14170
rect 16162 14118 16172 14170
rect 16196 14118 16226 14170
rect 16226 14118 16252 14170
rect 15956 14116 16012 14118
rect 16036 14116 16092 14118
rect 16116 14116 16172 14118
rect 16196 14116 16252 14118
rect 14462 8064 14518 8120
rect 13726 6860 13782 6896
rect 13726 6840 13728 6860
rect 13728 6840 13780 6860
rect 13780 6840 13782 6860
rect 15382 11600 15438 11656
rect 15956 13082 16012 13084
rect 16036 13082 16092 13084
rect 16116 13082 16172 13084
rect 16196 13082 16252 13084
rect 15956 13030 15982 13082
rect 15982 13030 16012 13082
rect 16036 13030 16046 13082
rect 16046 13030 16092 13082
rect 16116 13030 16162 13082
rect 16162 13030 16172 13082
rect 16196 13030 16226 13082
rect 16226 13030 16252 13082
rect 15956 13028 16012 13030
rect 16036 13028 16092 13030
rect 16116 13028 16172 13030
rect 16196 13028 16252 13030
rect 15566 10648 15622 10704
rect 15290 9424 15346 9480
rect 15842 12316 15844 12336
rect 15844 12316 15896 12336
rect 15896 12316 15898 12336
rect 15842 12280 15898 12316
rect 15956 11994 16012 11996
rect 16036 11994 16092 11996
rect 16116 11994 16172 11996
rect 16196 11994 16252 11996
rect 15956 11942 15982 11994
rect 15982 11942 16012 11994
rect 16036 11942 16046 11994
rect 16046 11942 16092 11994
rect 16116 11942 16162 11994
rect 16162 11942 16172 11994
rect 16196 11942 16226 11994
rect 16226 11942 16252 11994
rect 15956 11940 16012 11942
rect 16036 11940 16092 11942
rect 16116 11940 16172 11942
rect 16196 11940 16252 11942
rect 15842 11192 15898 11248
rect 16394 13096 16450 13152
rect 16670 11772 16672 11792
rect 16672 11772 16724 11792
rect 16724 11772 16726 11792
rect 16670 11736 16726 11772
rect 16394 11620 16450 11656
rect 16394 11600 16396 11620
rect 16396 11600 16448 11620
rect 16448 11600 16450 11620
rect 16302 11464 16358 11520
rect 15956 10906 16012 10908
rect 16036 10906 16092 10908
rect 16116 10906 16172 10908
rect 16196 10906 16252 10908
rect 15956 10854 15982 10906
rect 15982 10854 16012 10906
rect 16036 10854 16046 10906
rect 16046 10854 16092 10906
rect 16116 10854 16162 10906
rect 16162 10854 16172 10906
rect 16196 10854 16226 10906
rect 16226 10854 16252 10906
rect 15956 10852 16012 10854
rect 16036 10852 16092 10854
rect 16116 10852 16172 10854
rect 16196 10852 16252 10854
rect 15956 9818 16012 9820
rect 16036 9818 16092 9820
rect 16116 9818 16172 9820
rect 16196 9818 16252 9820
rect 15956 9766 15982 9818
rect 15982 9766 16012 9818
rect 16036 9766 16046 9818
rect 16046 9766 16092 9818
rect 16116 9766 16162 9818
rect 16162 9766 16172 9818
rect 16196 9766 16226 9818
rect 16226 9766 16252 9818
rect 15956 9764 16012 9766
rect 16036 9764 16092 9766
rect 16116 9764 16172 9766
rect 16196 9764 16252 9766
rect 18878 18808 18934 18864
rect 19338 18164 19340 18184
rect 19340 18164 19392 18184
rect 19392 18164 19394 18184
rect 19338 18128 19394 18164
rect 17774 13776 17830 13832
rect 17314 12824 17370 12880
rect 15658 9016 15714 9072
rect 16210 8880 16266 8936
rect 15956 8730 16012 8732
rect 16036 8730 16092 8732
rect 16116 8730 16172 8732
rect 16196 8730 16252 8732
rect 15956 8678 15982 8730
rect 15982 8678 16012 8730
rect 16036 8678 16046 8730
rect 16046 8678 16092 8730
rect 16116 8678 16162 8730
rect 16162 8678 16172 8730
rect 16196 8678 16226 8730
rect 16226 8678 16252 8730
rect 15956 8676 16012 8678
rect 16036 8676 16092 8678
rect 16116 8676 16172 8678
rect 16196 8676 16252 8678
rect 16302 8472 16358 8528
rect 15956 7642 16012 7644
rect 16036 7642 16092 7644
rect 16116 7642 16172 7644
rect 16196 7642 16252 7644
rect 15956 7590 15982 7642
rect 15982 7590 16012 7642
rect 16036 7590 16046 7642
rect 16046 7590 16092 7642
rect 16116 7590 16162 7642
rect 16162 7590 16172 7642
rect 16196 7590 16226 7642
rect 16226 7590 16252 7642
rect 15956 7588 16012 7590
rect 16036 7588 16092 7590
rect 16116 7588 16172 7590
rect 16196 7588 16252 7590
rect 17406 7928 17462 7984
rect 16946 7520 17002 7576
rect 16302 6704 16358 6760
rect 15956 6554 16012 6556
rect 16036 6554 16092 6556
rect 16116 6554 16172 6556
rect 16196 6554 16252 6556
rect 15956 6502 15982 6554
rect 15982 6502 16012 6554
rect 16036 6502 16046 6554
rect 16046 6502 16092 6554
rect 16116 6502 16162 6554
rect 16162 6502 16172 6554
rect 16196 6502 16226 6554
rect 16226 6502 16252 6554
rect 15956 6500 16012 6502
rect 16036 6500 16092 6502
rect 16116 6500 16172 6502
rect 16196 6500 16252 6502
rect 15566 6160 15622 6216
rect 14922 4664 14978 4720
rect 15956 5466 16012 5468
rect 16036 5466 16092 5468
rect 16116 5466 16172 5468
rect 16196 5466 16252 5468
rect 15956 5414 15982 5466
rect 15982 5414 16012 5466
rect 16036 5414 16046 5466
rect 16046 5414 16092 5466
rect 16116 5414 16162 5466
rect 16162 5414 16172 5466
rect 16196 5414 16226 5466
rect 16226 5414 16252 5466
rect 15956 5412 16012 5414
rect 16036 5412 16092 5414
rect 16116 5412 16172 5414
rect 16196 5412 16252 5414
rect 16946 7148 16948 7168
rect 16948 7148 17000 7168
rect 17000 7148 17002 7168
rect 16946 7112 17002 7148
rect 17406 7112 17462 7168
rect 17498 5652 17500 5672
rect 17500 5652 17552 5672
rect 17552 5652 17554 5672
rect 17498 5616 17554 5652
rect 17866 8628 17922 8664
rect 17866 8608 17868 8628
rect 17868 8608 17920 8628
rect 17920 8608 17922 8628
rect 18050 7248 18106 7304
rect 17498 4800 17554 4856
rect 15956 4378 16012 4380
rect 16036 4378 16092 4380
rect 16116 4378 16172 4380
rect 16196 4378 16252 4380
rect 15956 4326 15982 4378
rect 15982 4326 16012 4378
rect 16036 4326 16046 4378
rect 16046 4326 16092 4378
rect 16116 4326 16162 4378
rect 16162 4326 16172 4378
rect 16196 4326 16226 4378
rect 16226 4326 16252 4378
rect 15956 4324 16012 4326
rect 16036 4324 16092 4326
rect 16116 4324 16172 4326
rect 16196 4324 16252 4326
rect 15658 4120 15714 4176
rect 15956 3290 16012 3292
rect 16036 3290 16092 3292
rect 16116 3290 16172 3292
rect 16196 3290 16252 3292
rect 15956 3238 15982 3290
rect 15982 3238 16012 3290
rect 16036 3238 16046 3290
rect 16046 3238 16092 3290
rect 16116 3238 16162 3290
rect 16162 3238 16172 3290
rect 16196 3238 16226 3290
rect 16226 3238 16252 3290
rect 15956 3236 16012 3238
rect 16036 3236 16092 3238
rect 16116 3236 16172 3238
rect 16196 3236 16252 3238
rect 15956 2202 16012 2204
rect 16036 2202 16092 2204
rect 16116 2202 16172 2204
rect 16196 2202 16252 2204
rect 15956 2150 15982 2202
rect 15982 2150 16012 2202
rect 16036 2150 16046 2202
rect 16046 2150 16092 2202
rect 16116 2150 16162 2202
rect 16162 2150 16172 2202
rect 16196 2150 16226 2202
rect 16226 2150 16252 2202
rect 15956 2148 16012 2150
rect 16036 2148 16092 2150
rect 16116 2148 16172 2150
rect 16196 2148 16252 2150
rect 17314 3440 17370 3496
rect 16854 2644 16910 2680
rect 17866 3068 17868 3088
rect 17868 3068 17920 3088
rect 17920 3068 17922 3088
rect 17866 3032 17922 3068
rect 16854 2624 16856 2644
rect 16856 2624 16908 2644
rect 16908 2624 16910 2644
rect 19338 17176 19394 17232
rect 20810 20204 20812 20224
rect 20812 20204 20864 20224
rect 20864 20204 20866 20224
rect 20810 20168 20866 20204
rect 20956 20154 21012 20156
rect 21036 20154 21092 20156
rect 21116 20154 21172 20156
rect 21196 20154 21252 20156
rect 20956 20102 20982 20154
rect 20982 20102 21012 20154
rect 21036 20102 21046 20154
rect 21046 20102 21092 20154
rect 21116 20102 21162 20154
rect 21162 20102 21172 20154
rect 21196 20102 21226 20154
rect 21226 20102 21252 20154
rect 20956 20100 21012 20102
rect 21036 20100 21092 20102
rect 21116 20100 21172 20102
rect 21196 20100 21252 20102
rect 20956 19066 21012 19068
rect 21036 19066 21092 19068
rect 21116 19066 21172 19068
rect 21196 19066 21252 19068
rect 20956 19014 20982 19066
rect 20982 19014 21012 19066
rect 21036 19014 21046 19066
rect 21046 19014 21092 19066
rect 21116 19014 21162 19066
rect 21162 19014 21172 19066
rect 21196 19014 21226 19066
rect 21226 19014 21252 19066
rect 20956 19012 21012 19014
rect 21036 19012 21092 19014
rect 21116 19012 21172 19014
rect 21196 19012 21252 19014
rect 20956 17978 21012 17980
rect 21036 17978 21092 17980
rect 21116 17978 21172 17980
rect 21196 17978 21252 17980
rect 20956 17926 20982 17978
rect 20982 17926 21012 17978
rect 21036 17926 21046 17978
rect 21046 17926 21092 17978
rect 21116 17926 21162 17978
rect 21162 17926 21172 17978
rect 21196 17926 21226 17978
rect 21226 17926 21252 17978
rect 20956 17924 21012 17926
rect 21036 17924 21092 17926
rect 21116 17924 21172 17926
rect 21196 17924 21252 17926
rect 19154 16088 19210 16144
rect 18878 15852 18880 15872
rect 18880 15852 18932 15872
rect 18932 15852 18934 15872
rect 18878 15816 18934 15852
rect 19614 15952 19670 16008
rect 19614 15408 19670 15464
rect 25134 22344 25190 22400
rect 21730 20032 21786 20088
rect 21362 17720 21418 17776
rect 20956 16890 21012 16892
rect 21036 16890 21092 16892
rect 21116 16890 21172 16892
rect 21196 16890 21252 16892
rect 20956 16838 20982 16890
rect 20982 16838 21012 16890
rect 21036 16838 21046 16890
rect 21046 16838 21092 16890
rect 21116 16838 21162 16890
rect 21162 16838 21172 16890
rect 21196 16838 21226 16890
rect 21226 16838 21252 16890
rect 20956 16836 21012 16838
rect 21036 16836 21092 16838
rect 21116 16836 21172 16838
rect 21196 16836 21252 16838
rect 20074 15952 20130 16008
rect 19890 15272 19946 15328
rect 18694 13640 18750 13696
rect 19706 13640 19762 13696
rect 18418 12316 18420 12336
rect 18420 12316 18472 12336
rect 18472 12316 18474 12336
rect 18418 12280 18474 12316
rect 18418 10648 18474 10704
rect 18418 10532 18474 10568
rect 18418 10512 18420 10532
rect 18420 10512 18472 10532
rect 18472 10512 18474 10532
rect 19706 13368 19762 13424
rect 18786 12960 18842 13016
rect 19706 12416 19762 12472
rect 19338 11464 19394 11520
rect 19338 11056 19394 11112
rect 19522 10512 19578 10568
rect 18418 7928 18474 7984
rect 18510 6860 18566 6896
rect 18510 6840 18512 6860
rect 18512 6840 18564 6860
rect 18564 6840 18566 6860
rect 20956 15802 21012 15804
rect 21036 15802 21092 15804
rect 21116 15802 21172 15804
rect 21196 15802 21252 15804
rect 20956 15750 20982 15802
rect 20982 15750 21012 15802
rect 21036 15750 21046 15802
rect 21046 15750 21092 15802
rect 21116 15750 21162 15802
rect 21162 15750 21172 15802
rect 21196 15750 21226 15802
rect 21226 15750 21252 15802
rect 20956 15748 21012 15750
rect 21036 15748 21092 15750
rect 21116 15748 21172 15750
rect 21196 15748 21252 15750
rect 20534 15000 20590 15056
rect 20350 13776 20406 13832
rect 20442 13504 20498 13560
rect 20166 12552 20222 12608
rect 20166 12280 20222 12336
rect 20956 14714 21012 14716
rect 21036 14714 21092 14716
rect 21116 14714 21172 14716
rect 21196 14714 21252 14716
rect 20956 14662 20982 14714
rect 20982 14662 21012 14714
rect 21036 14662 21046 14714
rect 21046 14662 21092 14714
rect 21116 14662 21162 14714
rect 21162 14662 21172 14714
rect 21196 14662 21226 14714
rect 21226 14662 21252 14714
rect 20956 14660 21012 14662
rect 21036 14660 21092 14662
rect 21116 14660 21172 14662
rect 21196 14660 21252 14662
rect 20956 13626 21012 13628
rect 21036 13626 21092 13628
rect 21116 13626 21172 13628
rect 21196 13626 21252 13628
rect 20956 13574 20982 13626
rect 20982 13574 21012 13626
rect 21036 13574 21046 13626
rect 21046 13574 21092 13626
rect 21116 13574 21162 13626
rect 21162 13574 21172 13626
rect 21196 13574 21226 13626
rect 21226 13574 21252 13626
rect 20956 13572 21012 13574
rect 21036 13572 21092 13574
rect 21116 13572 21172 13574
rect 21196 13572 21252 13574
rect 20810 12960 20866 13016
rect 20902 12824 20958 12880
rect 20956 12538 21012 12540
rect 21036 12538 21092 12540
rect 21116 12538 21172 12540
rect 21196 12538 21252 12540
rect 20956 12486 20982 12538
rect 20982 12486 21012 12538
rect 21036 12486 21046 12538
rect 21046 12486 21092 12538
rect 21116 12486 21162 12538
rect 21162 12486 21172 12538
rect 21196 12486 21226 12538
rect 21226 12486 21252 12538
rect 20956 12484 21012 12486
rect 21036 12484 21092 12486
rect 21116 12484 21172 12486
rect 21196 12484 21252 12486
rect 25042 20440 25098 20496
rect 20956 11450 21012 11452
rect 21036 11450 21092 11452
rect 21116 11450 21172 11452
rect 21196 11450 21252 11452
rect 20956 11398 20982 11450
rect 20982 11398 21012 11450
rect 21036 11398 21046 11450
rect 21046 11398 21092 11450
rect 21116 11398 21162 11450
rect 21162 11398 21172 11450
rect 21196 11398 21226 11450
rect 21226 11398 21252 11450
rect 20956 11396 21012 11398
rect 21036 11396 21092 11398
rect 21116 11396 21172 11398
rect 21196 11396 21252 11398
rect 20810 11328 20866 11384
rect 21638 10512 21694 10568
rect 19430 8608 19486 8664
rect 19246 4120 19302 4176
rect 19890 4564 19892 4584
rect 19892 4564 19944 4584
rect 19944 4564 19946 4584
rect 19890 4528 19946 4564
rect 21638 10376 21694 10432
rect 20956 10362 21012 10364
rect 21036 10362 21092 10364
rect 21116 10362 21172 10364
rect 21196 10362 21252 10364
rect 20956 10310 20982 10362
rect 20982 10310 21012 10362
rect 21036 10310 21046 10362
rect 21046 10310 21092 10362
rect 21116 10310 21162 10362
rect 21162 10310 21172 10362
rect 21196 10310 21226 10362
rect 21226 10310 21252 10362
rect 20956 10308 21012 10310
rect 21036 10308 21092 10310
rect 21116 10308 21172 10310
rect 21196 10308 21252 10310
rect 21270 9560 21326 9616
rect 20956 9274 21012 9276
rect 21036 9274 21092 9276
rect 21116 9274 21172 9276
rect 21196 9274 21252 9276
rect 20956 9222 20982 9274
rect 20982 9222 21012 9274
rect 21036 9222 21046 9274
rect 21046 9222 21092 9274
rect 21116 9222 21162 9274
rect 21162 9222 21172 9274
rect 21196 9222 21226 9274
rect 21226 9222 21252 9274
rect 20956 9220 21012 9222
rect 21036 9220 21092 9222
rect 21116 9220 21172 9222
rect 21196 9220 21252 9222
rect 20718 8064 20774 8120
rect 20258 5244 20260 5264
rect 20260 5244 20312 5264
rect 20312 5244 20314 5264
rect 20258 5208 20314 5244
rect 20626 3576 20682 3632
rect 18878 3032 18934 3088
rect 20956 8186 21012 8188
rect 21036 8186 21092 8188
rect 21116 8186 21172 8188
rect 21196 8186 21252 8188
rect 20956 8134 20982 8186
rect 20982 8134 21012 8186
rect 21036 8134 21046 8186
rect 21046 8134 21092 8186
rect 21116 8134 21162 8186
rect 21162 8134 21172 8186
rect 21196 8134 21226 8186
rect 21226 8134 21252 8186
rect 20956 8132 21012 8134
rect 21036 8132 21092 8134
rect 21116 8132 21172 8134
rect 21196 8132 21252 8134
rect 20956 7098 21012 7100
rect 21036 7098 21092 7100
rect 21116 7098 21172 7100
rect 21196 7098 21252 7100
rect 20956 7046 20982 7098
rect 20982 7046 21012 7098
rect 21036 7046 21046 7098
rect 21046 7046 21092 7098
rect 21116 7046 21162 7098
rect 21162 7046 21172 7098
rect 21196 7046 21226 7098
rect 21226 7046 21252 7098
rect 20956 7044 21012 7046
rect 21036 7044 21092 7046
rect 21116 7044 21172 7046
rect 21196 7044 21252 7046
rect 20956 6010 21012 6012
rect 21036 6010 21092 6012
rect 21116 6010 21172 6012
rect 21196 6010 21252 6012
rect 20956 5958 20982 6010
rect 20982 5958 21012 6010
rect 21036 5958 21046 6010
rect 21046 5958 21092 6010
rect 21116 5958 21162 6010
rect 21162 5958 21172 6010
rect 21196 5958 21226 6010
rect 21226 5958 21252 6010
rect 20956 5956 21012 5958
rect 21036 5956 21092 5958
rect 21116 5956 21172 5958
rect 21196 5956 21252 5958
rect 21178 5772 21234 5808
rect 21178 5752 21180 5772
rect 21180 5752 21232 5772
rect 21232 5752 21234 5772
rect 20956 4922 21012 4924
rect 21036 4922 21092 4924
rect 21116 4922 21172 4924
rect 21196 4922 21252 4924
rect 20956 4870 20982 4922
rect 20982 4870 21012 4922
rect 21036 4870 21046 4922
rect 21046 4870 21092 4922
rect 21116 4870 21162 4922
rect 21162 4870 21172 4922
rect 21196 4870 21226 4922
rect 21226 4870 21252 4922
rect 20956 4868 21012 4870
rect 21036 4868 21092 4870
rect 21116 4868 21172 4870
rect 21196 4868 21252 4870
rect 20956 3834 21012 3836
rect 21036 3834 21092 3836
rect 21116 3834 21172 3836
rect 21196 3834 21252 3836
rect 20956 3782 20982 3834
rect 20982 3782 21012 3834
rect 21036 3782 21046 3834
rect 21046 3782 21092 3834
rect 21116 3782 21162 3834
rect 21162 3782 21172 3834
rect 21196 3782 21226 3834
rect 21226 3782 21252 3834
rect 20956 3780 21012 3782
rect 21036 3780 21092 3782
rect 21116 3780 21172 3782
rect 21196 3780 21252 3782
rect 23202 17176 23258 17232
rect 23478 17060 23534 17096
rect 23478 17040 23480 17060
rect 23480 17040 23532 17060
rect 23532 17040 23534 17060
rect 23202 16940 23204 16960
rect 23204 16940 23256 16960
rect 23256 16940 23258 16960
rect 23202 16904 23258 16940
rect 23662 15136 23718 15192
rect 21914 15000 21970 15056
rect 24858 16632 24914 16688
rect 24398 15272 24454 15328
rect 22650 13776 22706 13832
rect 21822 13368 21878 13424
rect 21822 12960 21878 13016
rect 21822 11600 21878 11656
rect 21914 6740 21916 6760
rect 21916 6740 21968 6760
rect 21968 6740 21970 6760
rect 21914 6704 21970 6740
rect 22374 6704 22430 6760
rect 20956 2746 21012 2748
rect 21036 2746 21092 2748
rect 21116 2746 21172 2748
rect 21196 2746 21252 2748
rect 20956 2694 20982 2746
rect 20982 2694 21012 2746
rect 21036 2694 21046 2746
rect 21046 2694 21092 2746
rect 21116 2694 21162 2746
rect 21162 2694 21172 2746
rect 21196 2694 21226 2746
rect 21226 2694 21252 2746
rect 20956 2692 21012 2694
rect 21036 2692 21092 2694
rect 21116 2692 21172 2694
rect 21196 2692 21252 2694
rect 20810 2624 20866 2680
rect 24398 13504 24454 13560
rect 24398 12824 24454 12880
rect 24674 13096 24730 13152
rect 24674 12824 24730 12880
rect 24306 11600 24362 11656
rect 24766 12280 24822 12336
rect 24398 9560 24454 9616
rect 23478 7520 23534 7576
rect 23846 7384 23902 7440
rect 24030 7384 24086 7440
rect 23110 7248 23166 7304
rect 23662 7248 23718 7304
rect 23570 5616 23626 5672
rect 24122 6976 24178 7032
rect 25778 23024 25834 23080
rect 27526 21800 27582 21856
rect 25956 21786 26012 21788
rect 26036 21786 26092 21788
rect 26116 21786 26172 21788
rect 26196 21786 26252 21788
rect 25956 21734 25982 21786
rect 25982 21734 26012 21786
rect 26036 21734 26046 21786
rect 26046 21734 26092 21786
rect 26116 21734 26162 21786
rect 26162 21734 26172 21786
rect 26196 21734 26226 21786
rect 26226 21734 26252 21786
rect 25956 21732 26012 21734
rect 26036 21732 26092 21734
rect 26116 21732 26172 21734
rect 26196 21732 26252 21734
rect 25318 19216 25374 19272
rect 25226 18672 25282 18728
rect 25502 18944 25558 19000
rect 25502 18264 25558 18320
rect 25502 17040 25558 17096
rect 25318 15816 25374 15872
rect 25502 15544 25558 15600
rect 25410 15408 25466 15464
rect 25134 12416 25190 12472
rect 25226 12144 25282 12200
rect 25134 11756 25190 11792
rect 25134 11736 25136 11756
rect 25136 11736 25188 11756
rect 25188 11736 25190 11756
rect 23570 4548 23626 4584
rect 23570 4528 23572 4548
rect 23572 4528 23624 4548
rect 23624 4528 23626 4548
rect 24858 3712 24914 3768
rect 23846 2896 23902 2952
rect 25870 21256 25926 21312
rect 25686 18808 25742 18864
rect 25686 18264 25742 18320
rect 25686 17584 25742 17640
rect 25686 16632 25742 16688
rect 25686 16244 25742 16280
rect 25686 16224 25688 16244
rect 25688 16224 25740 16244
rect 25740 16224 25742 16244
rect 25686 15408 25742 15464
rect 25956 20698 26012 20700
rect 26036 20698 26092 20700
rect 26116 20698 26172 20700
rect 26196 20698 26252 20700
rect 25956 20646 25982 20698
rect 25982 20646 26012 20698
rect 26036 20646 26046 20698
rect 26046 20646 26092 20698
rect 26116 20646 26162 20698
rect 26162 20646 26172 20698
rect 26196 20646 26226 20698
rect 26226 20646 26252 20698
rect 25956 20644 26012 20646
rect 26036 20644 26092 20646
rect 26116 20644 26172 20646
rect 26196 20644 26252 20646
rect 26054 20304 26110 20360
rect 25956 19610 26012 19612
rect 26036 19610 26092 19612
rect 26116 19610 26172 19612
rect 26196 19610 26252 19612
rect 25956 19558 25982 19610
rect 25982 19558 26012 19610
rect 26036 19558 26046 19610
rect 26046 19558 26092 19610
rect 26116 19558 26162 19610
rect 26162 19558 26172 19610
rect 26196 19558 26226 19610
rect 26226 19558 26252 19610
rect 25956 19556 26012 19558
rect 26036 19556 26092 19558
rect 26116 19556 26172 19558
rect 26196 19556 26252 19558
rect 25956 18522 26012 18524
rect 26036 18522 26092 18524
rect 26116 18522 26172 18524
rect 26196 18522 26252 18524
rect 25956 18470 25982 18522
rect 25982 18470 26012 18522
rect 26036 18470 26046 18522
rect 26046 18470 26092 18522
rect 26116 18470 26162 18522
rect 26162 18470 26172 18522
rect 26196 18470 26226 18522
rect 26226 18470 26252 18522
rect 25956 18468 26012 18470
rect 26036 18468 26092 18470
rect 26116 18468 26172 18470
rect 26196 18468 26252 18470
rect 25956 17434 26012 17436
rect 26036 17434 26092 17436
rect 26116 17434 26172 17436
rect 26196 17434 26252 17436
rect 25956 17382 25982 17434
rect 25982 17382 26012 17434
rect 26036 17382 26046 17434
rect 26046 17382 26092 17434
rect 26116 17382 26162 17434
rect 26162 17382 26172 17434
rect 26196 17382 26226 17434
rect 26226 17382 26252 17434
rect 25956 17380 26012 17382
rect 26036 17380 26092 17382
rect 26116 17380 26172 17382
rect 26196 17380 26252 17382
rect 26330 16904 26386 16960
rect 25956 16346 26012 16348
rect 26036 16346 26092 16348
rect 26116 16346 26172 16348
rect 26196 16346 26252 16348
rect 25956 16294 25982 16346
rect 25982 16294 26012 16346
rect 26036 16294 26046 16346
rect 26046 16294 26092 16346
rect 26116 16294 26162 16346
rect 26162 16294 26172 16346
rect 26196 16294 26226 16346
rect 26226 16294 26252 16346
rect 25956 16292 26012 16294
rect 26036 16292 26092 16294
rect 26116 16292 26172 16294
rect 26196 16292 26252 16294
rect 25956 15258 26012 15260
rect 26036 15258 26092 15260
rect 26116 15258 26172 15260
rect 26196 15258 26252 15260
rect 25956 15206 25982 15258
rect 25982 15206 26012 15258
rect 26036 15206 26046 15258
rect 26046 15206 26092 15258
rect 26116 15206 26162 15258
rect 26162 15206 26172 15258
rect 26196 15206 26226 15258
rect 26226 15206 26252 15258
rect 25956 15204 26012 15206
rect 26036 15204 26092 15206
rect 26116 15204 26172 15206
rect 26196 15204 26252 15206
rect 25686 13232 25742 13288
rect 25502 12416 25558 12472
rect 25410 11056 25466 11112
rect 25318 7284 25320 7304
rect 25320 7284 25372 7304
rect 25372 7284 25374 7304
rect 25318 7248 25374 7284
rect 25956 14170 26012 14172
rect 26036 14170 26092 14172
rect 26116 14170 26172 14172
rect 26196 14170 26252 14172
rect 25956 14118 25982 14170
rect 25982 14118 26012 14170
rect 26036 14118 26046 14170
rect 26046 14118 26092 14170
rect 26116 14118 26162 14170
rect 26162 14118 26172 14170
rect 26196 14118 26226 14170
rect 26226 14118 26252 14170
rect 25956 14116 26012 14118
rect 26036 14116 26092 14118
rect 26116 14116 26172 14118
rect 26196 14116 26252 14118
rect 25956 13082 26012 13084
rect 26036 13082 26092 13084
rect 26116 13082 26172 13084
rect 26196 13082 26252 13084
rect 25956 13030 25982 13082
rect 25982 13030 26012 13082
rect 26036 13030 26046 13082
rect 26046 13030 26092 13082
rect 26116 13030 26162 13082
rect 26162 13030 26172 13082
rect 26196 13030 26226 13082
rect 26226 13030 26252 13082
rect 25956 13028 26012 13030
rect 26036 13028 26092 13030
rect 26116 13028 26172 13030
rect 26196 13028 26252 13030
rect 25962 12824 26018 12880
rect 26974 18944 27030 19000
rect 26514 18128 26570 18184
rect 26330 12280 26386 12336
rect 25956 11994 26012 11996
rect 26036 11994 26092 11996
rect 26116 11994 26172 11996
rect 26196 11994 26252 11996
rect 25956 11942 25982 11994
rect 25982 11942 26012 11994
rect 26036 11942 26046 11994
rect 26046 11942 26092 11994
rect 26116 11942 26162 11994
rect 26162 11942 26172 11994
rect 26196 11942 26226 11994
rect 26226 11942 26252 11994
rect 25956 11940 26012 11942
rect 26036 11940 26092 11942
rect 26116 11940 26172 11942
rect 26196 11940 26252 11942
rect 26238 11600 26294 11656
rect 26422 11228 26424 11248
rect 26424 11228 26476 11248
rect 26476 11228 26478 11248
rect 26422 11192 26478 11228
rect 25870 11056 25926 11112
rect 25956 10906 26012 10908
rect 26036 10906 26092 10908
rect 26116 10906 26172 10908
rect 26196 10906 26252 10908
rect 25956 10854 25982 10906
rect 25982 10854 26012 10906
rect 26036 10854 26046 10906
rect 26046 10854 26092 10906
rect 26116 10854 26162 10906
rect 26162 10854 26172 10906
rect 26196 10854 26226 10906
rect 26226 10854 26252 10906
rect 25956 10852 26012 10854
rect 26036 10852 26092 10854
rect 26116 10852 26172 10854
rect 26196 10852 26252 10854
rect 26422 10548 26424 10568
rect 26424 10548 26476 10568
rect 26476 10548 26478 10568
rect 26422 10512 26478 10548
rect 26698 11600 26754 11656
rect 26606 10412 26608 10432
rect 26608 10412 26660 10432
rect 26660 10412 26662 10432
rect 26606 10376 26662 10412
rect 25956 9818 26012 9820
rect 26036 9818 26092 9820
rect 26116 9818 26172 9820
rect 26196 9818 26252 9820
rect 25956 9766 25982 9818
rect 25982 9766 26012 9818
rect 26036 9766 26046 9818
rect 26046 9766 26092 9818
rect 26116 9766 26162 9818
rect 26162 9766 26172 9818
rect 26196 9766 26226 9818
rect 26226 9766 26252 9818
rect 25956 9764 26012 9766
rect 26036 9764 26092 9766
rect 26116 9764 26172 9766
rect 26196 9764 26252 9766
rect 26698 9868 26700 9888
rect 26700 9868 26752 9888
rect 26752 9868 26754 9888
rect 26698 9832 26754 9868
rect 25870 8916 25872 8936
rect 25872 8916 25924 8936
rect 25924 8916 25926 8936
rect 25870 8880 25926 8916
rect 25956 8730 26012 8732
rect 26036 8730 26092 8732
rect 26116 8730 26172 8732
rect 26196 8730 26252 8732
rect 25956 8678 25982 8730
rect 25982 8678 26012 8730
rect 26036 8678 26046 8730
rect 26046 8678 26092 8730
rect 26116 8678 26162 8730
rect 26162 8678 26172 8730
rect 26196 8678 26226 8730
rect 26226 8678 26252 8730
rect 25956 8676 26012 8678
rect 26036 8676 26092 8678
rect 26116 8676 26172 8678
rect 26196 8676 26252 8678
rect 25956 7642 26012 7644
rect 26036 7642 26092 7644
rect 26116 7642 26172 7644
rect 26196 7642 26252 7644
rect 25956 7590 25982 7642
rect 25982 7590 26012 7642
rect 26036 7590 26046 7642
rect 26046 7590 26092 7642
rect 26116 7590 26162 7642
rect 26162 7590 26172 7642
rect 26196 7590 26226 7642
rect 26226 7590 26252 7642
rect 25956 7588 26012 7590
rect 26036 7588 26092 7590
rect 26116 7588 26172 7590
rect 26196 7588 26252 7590
rect 26606 9288 26662 9344
rect 26698 8608 26754 8664
rect 26330 6976 26386 7032
rect 25594 6840 25650 6896
rect 25778 6840 25834 6896
rect 25956 6554 26012 6556
rect 26036 6554 26092 6556
rect 26116 6554 26172 6556
rect 26196 6554 26252 6556
rect 25956 6502 25982 6554
rect 25982 6502 26012 6554
rect 26036 6502 26046 6554
rect 26046 6502 26092 6554
rect 26116 6502 26162 6554
rect 26162 6502 26172 6554
rect 26196 6502 26226 6554
rect 26226 6502 26252 6554
rect 25956 6500 26012 6502
rect 26036 6500 26092 6502
rect 26116 6500 26172 6502
rect 26196 6500 26252 6502
rect 26238 6180 26294 6216
rect 26238 6160 26240 6180
rect 26240 6160 26292 6180
rect 26292 6160 26294 6180
rect 25956 5466 26012 5468
rect 26036 5466 26092 5468
rect 26116 5466 26172 5468
rect 26196 5466 26252 5468
rect 25956 5414 25982 5466
rect 25982 5414 26012 5466
rect 26036 5414 26046 5466
rect 26046 5414 26092 5466
rect 26116 5414 26162 5466
rect 26162 5414 26172 5466
rect 26196 5414 26226 5466
rect 26226 5414 26252 5466
rect 25956 5412 26012 5414
rect 26036 5412 26092 5414
rect 26116 5412 26172 5414
rect 26196 5412 26252 5414
rect 26238 5092 26294 5128
rect 26238 5072 26240 5092
rect 26240 5072 26292 5092
rect 26292 5072 26294 5092
rect 25956 4378 26012 4380
rect 26036 4378 26092 4380
rect 26116 4378 26172 4380
rect 26196 4378 26252 4380
rect 25956 4326 25982 4378
rect 25982 4326 26012 4378
rect 26036 4326 26046 4378
rect 26046 4326 26092 4378
rect 26116 4326 26162 4378
rect 26162 4326 26172 4378
rect 26196 4326 26226 4378
rect 26226 4326 26252 4378
rect 25956 4324 26012 4326
rect 26036 4324 26092 4326
rect 26116 4324 26172 4326
rect 26196 4324 26252 4326
rect 26514 7948 26570 7984
rect 26514 7928 26516 7948
rect 26516 7928 26568 7948
rect 26568 7928 26570 7948
rect 26514 7384 26570 7440
rect 26698 7384 26754 7440
rect 26422 5752 26478 5808
rect 26882 12688 26938 12744
rect 27526 14048 27582 14104
rect 27526 13232 27582 13288
rect 26974 6704 27030 6760
rect 26790 6296 26846 6352
rect 26606 5616 26662 5672
rect 26606 5072 26662 5128
rect 26514 4684 26570 4720
rect 26514 4664 26516 4684
rect 26516 4664 26568 4684
rect 26568 4664 26570 4684
rect 26422 4020 26424 4040
rect 26424 4020 26476 4040
rect 26476 4020 26478 4040
rect 26422 3984 26478 4020
rect 25956 3290 26012 3292
rect 26036 3290 26092 3292
rect 26116 3290 26172 3292
rect 26196 3290 26252 3292
rect 25956 3238 25982 3290
rect 25982 3238 26012 3290
rect 26036 3238 26046 3290
rect 26046 3238 26092 3290
rect 26116 3238 26162 3290
rect 26162 3238 26172 3290
rect 26196 3238 26226 3290
rect 26226 3238 26252 3290
rect 25956 3236 26012 3238
rect 26036 3236 26092 3238
rect 26116 3236 26172 3238
rect 26196 3236 26252 3238
rect 25686 3032 25742 3088
rect 25956 2202 26012 2204
rect 26036 2202 26092 2204
rect 26116 2202 26172 2204
rect 26196 2202 26252 2204
rect 25956 2150 25982 2202
rect 25982 2150 26012 2202
rect 26036 2150 26046 2202
rect 26046 2150 26092 2202
rect 26116 2150 26162 2202
rect 26162 2150 26172 2202
rect 26196 2150 26226 2202
rect 26226 2150 26252 2202
rect 25956 2148 26012 2150
rect 26036 2148 26092 2150
rect 26116 2148 26172 2150
rect 26196 2148 26252 2150
rect 25870 856 25926 912
rect 26790 3848 26846 3904
rect 27526 10648 27582 10704
rect 27710 8064 27766 8120
rect 27710 4392 27766 4448
rect 27434 3712 27490 3768
rect 27526 3576 27582 3632
rect 3974 312 4030 368
rect 26698 2760 26754 2816
rect 26882 3304 26938 3360
rect 27710 2080 27766 2136
rect 26790 1400 26846 1456
rect 26606 312 26662 368
<< metal3 >>
rect 0 23626 480 23656
rect 3969 23626 4035 23629
rect 0 23624 4035 23626
rect 0 23568 3974 23624
rect 4030 23568 4035 23624
rect 0 23566 4035 23568
rect 0 23536 480 23566
rect 3969 23563 4035 23566
rect 25865 23626 25931 23629
rect 29520 23626 30000 23656
rect 25865 23624 30000 23626
rect 25865 23568 25870 23624
rect 25926 23568 30000 23624
rect 25865 23566 30000 23568
rect 25865 23563 25931 23566
rect 29520 23536 30000 23566
rect 0 23082 480 23112
rect 4245 23082 4311 23085
rect 0 23080 4311 23082
rect 0 23024 4250 23080
rect 4306 23024 4311 23080
rect 0 23022 4311 23024
rect 0 22992 480 23022
rect 4245 23019 4311 23022
rect 25773 23082 25839 23085
rect 29520 23082 30000 23112
rect 25773 23080 30000 23082
rect 25773 23024 25778 23080
rect 25834 23024 30000 23080
rect 25773 23022 30000 23024
rect 25773 23019 25839 23022
rect 29520 22992 30000 23022
rect 0 22402 480 22432
rect 2865 22402 2931 22405
rect 0 22400 2931 22402
rect 0 22344 2870 22400
rect 2926 22344 2931 22400
rect 0 22342 2931 22344
rect 0 22312 480 22342
rect 2865 22339 2931 22342
rect 25129 22402 25195 22405
rect 29520 22402 30000 22432
rect 25129 22400 30000 22402
rect 25129 22344 25134 22400
rect 25190 22344 30000 22400
rect 25129 22342 30000 22344
rect 25129 22339 25195 22342
rect 29520 22312 30000 22342
rect 0 21858 480 21888
rect 4061 21858 4127 21861
rect 0 21856 4127 21858
rect 0 21800 4066 21856
rect 4122 21800 4127 21856
rect 0 21798 4127 21800
rect 0 21768 480 21798
rect 4061 21795 4127 21798
rect 27521 21858 27587 21861
rect 29520 21858 30000 21888
rect 27521 21856 30000 21858
rect 27521 21800 27526 21856
rect 27582 21800 30000 21856
rect 27521 21798 30000 21800
rect 27521 21795 27587 21798
rect 5944 21792 6264 21793
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 21727 6264 21728
rect 15944 21792 16264 21793
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 21727 16264 21728
rect 25944 21792 26264 21793
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 29520 21768 30000 21798
rect 25944 21727 26264 21728
rect 0 21314 480 21344
rect 7281 21314 7347 21317
rect 0 21312 7347 21314
rect 0 21256 7286 21312
rect 7342 21256 7347 21312
rect 0 21254 7347 21256
rect 0 21224 480 21254
rect 7281 21251 7347 21254
rect 25865 21314 25931 21317
rect 29520 21314 30000 21344
rect 25865 21312 30000 21314
rect 25865 21256 25870 21312
rect 25926 21256 30000 21312
rect 25865 21254 30000 21256
rect 25865 21251 25931 21254
rect 10944 21248 11264 21249
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 21183 11264 21184
rect 20944 21248 21264 21249
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 29520 21224 30000 21254
rect 20944 21183 21264 21184
rect 5944 20704 6264 20705
rect 0 20634 480 20664
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 20639 6264 20640
rect 15944 20704 16264 20705
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 20639 16264 20640
rect 25944 20704 26264 20705
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 20639 26264 20640
rect 3233 20634 3299 20637
rect 29520 20634 30000 20664
rect 0 20632 3299 20634
rect 0 20576 3238 20632
rect 3294 20576 3299 20632
rect 0 20574 3299 20576
rect 0 20544 480 20574
rect 3233 20571 3299 20574
rect 26374 20574 30000 20634
rect 8753 20498 8819 20501
rect 12433 20498 12499 20501
rect 8753 20496 12499 20498
rect 8753 20440 8758 20496
rect 8814 20440 12438 20496
rect 12494 20440 12499 20496
rect 8753 20438 12499 20440
rect 8753 20435 8819 20438
rect 12433 20435 12499 20438
rect 16113 20498 16179 20501
rect 18321 20498 18387 20501
rect 16113 20496 18387 20498
rect 16113 20440 16118 20496
rect 16174 20440 18326 20496
rect 18382 20440 18387 20496
rect 16113 20438 18387 20440
rect 16113 20435 16179 20438
rect 18321 20435 18387 20438
rect 25037 20498 25103 20501
rect 26374 20498 26434 20574
rect 29520 20544 30000 20574
rect 25037 20496 26434 20498
rect 25037 20440 25042 20496
rect 25098 20440 26434 20496
rect 25037 20438 26434 20440
rect 25037 20435 25103 20438
rect 4981 20362 5047 20365
rect 26049 20362 26115 20365
rect 4981 20360 26115 20362
rect 4981 20304 4986 20360
rect 5042 20304 26054 20360
rect 26110 20304 26115 20360
rect 4981 20302 26115 20304
rect 4981 20299 5047 20302
rect 26049 20299 26115 20302
rect 14917 20226 14983 20229
rect 20805 20226 20871 20229
rect 14917 20224 20871 20226
rect 14917 20168 14922 20224
rect 14978 20168 20810 20224
rect 20866 20168 20871 20224
rect 14917 20166 20871 20168
rect 14917 20163 14983 20166
rect 20805 20163 20871 20166
rect 10944 20160 11264 20161
rect 0 20090 480 20120
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 20095 11264 20096
rect 20944 20160 21264 20161
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 20095 21264 20096
rect 3325 20090 3391 20093
rect 0 20088 3391 20090
rect 0 20032 3330 20088
rect 3386 20032 3391 20088
rect 0 20030 3391 20032
rect 0 20000 480 20030
rect 3325 20027 3391 20030
rect 21725 20090 21791 20093
rect 29520 20090 30000 20120
rect 21725 20088 30000 20090
rect 21725 20032 21730 20088
rect 21786 20032 30000 20088
rect 21725 20030 30000 20032
rect 21725 20027 21791 20030
rect 29520 20000 30000 20030
rect 8017 19954 8083 19957
rect 15837 19954 15903 19957
rect 614 19894 7666 19954
rect 0 19410 480 19440
rect 614 19410 674 19894
rect 7606 19682 7666 19894
rect 8017 19952 15903 19954
rect 8017 19896 8022 19952
rect 8078 19896 15842 19952
rect 15898 19896 15903 19952
rect 8017 19894 15903 19896
rect 8017 19891 8083 19894
rect 15837 19891 15903 19894
rect 10869 19818 10935 19821
rect 14181 19818 14247 19821
rect 10869 19816 14247 19818
rect 10869 19760 10874 19816
rect 10930 19760 14186 19816
rect 14242 19760 14247 19816
rect 10869 19758 14247 19760
rect 10869 19755 10935 19758
rect 14181 19755 14247 19758
rect 13905 19682 13971 19685
rect 7606 19680 13971 19682
rect 7606 19624 13910 19680
rect 13966 19624 13971 19680
rect 7606 19622 13971 19624
rect 13905 19619 13971 19622
rect 5944 19616 6264 19617
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 19551 6264 19552
rect 15944 19616 16264 19617
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 19551 16264 19552
rect 25944 19616 26264 19617
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 19551 26264 19552
rect 0 19350 674 19410
rect 16389 19410 16455 19413
rect 29520 19410 30000 19440
rect 16389 19408 30000 19410
rect 16389 19352 16394 19408
rect 16450 19352 30000 19408
rect 16389 19350 30000 19352
rect 0 19320 480 19350
rect 16389 19347 16455 19350
rect 29520 19320 30000 19350
rect 10501 19274 10567 19277
rect 25313 19274 25379 19277
rect 10501 19272 25379 19274
rect 10501 19216 10506 19272
rect 10562 19216 25318 19272
rect 25374 19216 25379 19272
rect 10501 19214 25379 19216
rect 10501 19211 10567 19214
rect 25313 19211 25379 19214
rect 5349 19138 5415 19141
rect 10593 19138 10659 19141
rect 5349 19136 10794 19138
rect 5349 19080 5354 19136
rect 5410 19080 10598 19136
rect 10654 19080 10794 19136
rect 5349 19078 10794 19080
rect 5349 19075 5415 19078
rect 10593 19075 10659 19078
rect 0 18866 480 18896
rect 4981 18866 5047 18869
rect 0 18864 5047 18866
rect 0 18808 4986 18864
rect 5042 18808 5047 18864
rect 0 18806 5047 18808
rect 10734 18866 10794 19078
rect 10944 19072 11264 19073
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 19007 11264 19008
rect 20944 19072 21264 19073
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 19007 21264 19008
rect 25497 19002 25563 19005
rect 26969 19002 27035 19005
rect 25497 19000 27035 19002
rect 25497 18944 25502 19000
rect 25558 18944 26974 19000
rect 27030 18944 27035 19000
rect 25497 18942 27035 18944
rect 25497 18939 25563 18942
rect 26969 18939 27035 18942
rect 18873 18866 18939 18869
rect 25681 18866 25747 18869
rect 29520 18866 30000 18896
rect 10734 18864 25747 18866
rect 10734 18808 18878 18864
rect 18934 18808 25686 18864
rect 25742 18808 25747 18864
rect 10734 18806 25747 18808
rect 0 18776 480 18806
rect 4981 18803 5047 18806
rect 18873 18803 18939 18806
rect 25681 18803 25747 18806
rect 26742 18806 30000 18866
rect 25221 18730 25287 18733
rect 26742 18730 26802 18806
rect 29520 18776 30000 18806
rect 25221 18728 26802 18730
rect 25221 18672 25226 18728
rect 25282 18672 26802 18728
rect 25221 18670 26802 18672
rect 25221 18667 25287 18670
rect 5944 18528 6264 18529
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 18463 6264 18464
rect 15944 18528 16264 18529
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 18463 16264 18464
rect 25944 18528 26264 18529
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 18463 26264 18464
rect 0 18322 480 18352
rect 4705 18322 4771 18325
rect 0 18320 4771 18322
rect 0 18264 4710 18320
rect 4766 18264 4771 18320
rect 0 18262 4771 18264
rect 0 18232 480 18262
rect 4705 18259 4771 18262
rect 10041 18322 10107 18325
rect 25497 18324 25563 18325
rect 25446 18322 25452 18324
rect 10041 18320 25452 18322
rect 25516 18320 25563 18324
rect 10041 18264 10046 18320
rect 10102 18264 25452 18320
rect 25558 18264 25563 18320
rect 10041 18262 25452 18264
rect 10041 18259 10107 18262
rect 25446 18260 25452 18262
rect 25516 18260 25563 18264
rect 25497 18259 25563 18260
rect 25681 18322 25747 18325
rect 29520 18322 30000 18352
rect 25681 18320 30000 18322
rect 25681 18264 25686 18320
rect 25742 18264 30000 18320
rect 25681 18262 30000 18264
rect 25681 18259 25747 18262
rect 29520 18232 30000 18262
rect 4245 18186 4311 18189
rect 15745 18186 15811 18189
rect 19333 18186 19399 18189
rect 26509 18186 26575 18189
rect 4245 18184 26575 18186
rect 4245 18128 4250 18184
rect 4306 18128 15750 18184
rect 15806 18128 19338 18184
rect 19394 18128 26514 18184
rect 26570 18128 26575 18184
rect 4245 18126 26575 18128
rect 4245 18123 4311 18126
rect 15745 18123 15811 18126
rect 19333 18123 19399 18126
rect 26509 18123 26575 18126
rect 2037 18050 2103 18053
rect 4521 18050 4587 18053
rect 2037 18048 4587 18050
rect 2037 17992 2042 18048
rect 2098 17992 4526 18048
rect 4582 17992 4587 18048
rect 2037 17990 4587 17992
rect 2037 17987 2103 17990
rect 4521 17987 4587 17990
rect 4705 18050 4771 18053
rect 9673 18050 9739 18053
rect 4705 18048 9739 18050
rect 4705 17992 4710 18048
rect 4766 17992 9678 18048
rect 9734 17992 9739 18048
rect 4705 17990 9739 17992
rect 4705 17987 4771 17990
rect 9673 17987 9739 17990
rect 10944 17984 11264 17985
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 17919 11264 17920
rect 20944 17984 21264 17985
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 17919 21264 17920
rect 13261 17914 13327 17917
rect 15377 17914 15443 17917
rect 13261 17912 15443 17914
rect 13261 17856 13266 17912
rect 13322 17856 15382 17912
rect 15438 17856 15443 17912
rect 13261 17854 15443 17856
rect 13261 17851 13327 17854
rect 15377 17851 15443 17854
rect 1393 17778 1459 17781
rect 16665 17778 16731 17781
rect 21357 17778 21423 17781
rect 1393 17776 5090 17778
rect 1393 17720 1398 17776
rect 1454 17720 5090 17776
rect 1393 17718 5090 17720
rect 1393 17715 1459 17718
rect 0 17642 480 17672
rect 3417 17642 3483 17645
rect 0 17640 3483 17642
rect 0 17584 3422 17640
rect 3478 17584 3483 17640
rect 0 17582 3483 17584
rect 5030 17642 5090 17718
rect 14966 17776 21423 17778
rect 14966 17720 16670 17776
rect 16726 17720 21362 17776
rect 21418 17720 21423 17776
rect 14966 17718 21423 17720
rect 5165 17642 5231 17645
rect 14966 17642 15026 17718
rect 16665 17715 16731 17718
rect 21357 17715 21423 17718
rect 5030 17640 15026 17642
rect 5030 17584 5170 17640
rect 5226 17584 15026 17640
rect 5030 17582 15026 17584
rect 15193 17642 15259 17645
rect 16757 17642 16823 17645
rect 15193 17640 16823 17642
rect 15193 17584 15198 17640
rect 15254 17584 16762 17640
rect 16818 17584 16823 17640
rect 15193 17582 16823 17584
rect 0 17552 480 17582
rect 3417 17579 3483 17582
rect 5165 17579 5231 17582
rect 15193 17579 15259 17582
rect 16757 17579 16823 17582
rect 25681 17642 25747 17645
rect 29520 17642 30000 17672
rect 25681 17640 30000 17642
rect 25681 17584 25686 17640
rect 25742 17584 30000 17640
rect 25681 17582 30000 17584
rect 25681 17579 25747 17582
rect 29520 17552 30000 17582
rect 10593 17506 10659 17509
rect 15745 17506 15811 17509
rect 10593 17504 15811 17506
rect 10593 17448 10598 17504
rect 10654 17448 15750 17504
rect 15806 17448 15811 17504
rect 10593 17446 15811 17448
rect 10593 17443 10659 17446
rect 15745 17443 15811 17446
rect 5944 17440 6264 17441
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 17375 6264 17376
rect 15944 17440 16264 17441
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 17375 16264 17376
rect 25944 17440 26264 17441
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 17375 26264 17376
rect 4061 17234 4127 17237
rect 5809 17234 5875 17237
rect 4061 17232 5875 17234
rect 4061 17176 4066 17232
rect 4122 17176 5814 17232
rect 5870 17176 5875 17232
rect 4061 17174 5875 17176
rect 4061 17171 4127 17174
rect 5809 17171 5875 17174
rect 9673 17234 9739 17237
rect 19333 17234 19399 17237
rect 23197 17234 23263 17237
rect 9673 17232 23263 17234
rect 9673 17176 9678 17232
rect 9734 17176 19338 17232
rect 19394 17176 23202 17232
rect 23258 17176 23263 17232
rect 9673 17174 23263 17176
rect 9673 17171 9739 17174
rect 19333 17171 19399 17174
rect 23197 17171 23263 17174
rect 0 17098 480 17128
rect 3141 17098 3207 17101
rect 0 17096 3207 17098
rect 0 17040 3146 17096
rect 3202 17040 3207 17096
rect 0 17038 3207 17040
rect 0 17008 480 17038
rect 3141 17035 3207 17038
rect 11605 17098 11671 17101
rect 12065 17098 12131 17101
rect 23473 17098 23539 17101
rect 11605 17096 23539 17098
rect 11605 17040 11610 17096
rect 11666 17040 12070 17096
rect 12126 17040 23478 17096
rect 23534 17040 23539 17096
rect 11605 17038 23539 17040
rect 11605 17035 11671 17038
rect 12065 17035 12131 17038
rect 23473 17035 23539 17038
rect 25497 17098 25563 17101
rect 29520 17098 30000 17128
rect 25497 17096 30000 17098
rect 25497 17040 25502 17096
rect 25558 17040 30000 17096
rect 25497 17038 30000 17040
rect 25497 17035 25563 17038
rect 29520 17008 30000 17038
rect 23197 16962 23263 16965
rect 26325 16962 26391 16965
rect 23197 16960 26391 16962
rect 23197 16904 23202 16960
rect 23258 16904 26330 16960
rect 26386 16904 26391 16960
rect 23197 16902 26391 16904
rect 23197 16899 23263 16902
rect 26325 16899 26391 16902
rect 10944 16896 11264 16897
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 16831 11264 16832
rect 20944 16896 21264 16897
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 16831 21264 16832
rect 3233 16826 3299 16829
rect 6821 16826 6887 16829
rect 3233 16824 6887 16826
rect 3233 16768 3238 16824
rect 3294 16768 6826 16824
rect 6882 16768 6887 16824
rect 3233 16766 6887 16768
rect 3233 16763 3299 16766
rect 6821 16763 6887 16766
rect 5073 16690 5139 16693
rect 9581 16690 9647 16693
rect 5073 16688 9647 16690
rect 5073 16632 5078 16688
rect 5134 16632 9586 16688
rect 9642 16632 9647 16688
rect 5073 16630 9647 16632
rect 5073 16627 5139 16630
rect 9581 16627 9647 16630
rect 10409 16690 10475 16693
rect 11973 16690 12039 16693
rect 10409 16688 12039 16690
rect 10409 16632 10414 16688
rect 10470 16632 11978 16688
rect 12034 16632 12039 16688
rect 10409 16630 12039 16632
rect 10409 16627 10475 16630
rect 11973 16627 12039 16630
rect 24853 16690 24919 16693
rect 25681 16690 25747 16693
rect 24853 16688 25747 16690
rect 24853 16632 24858 16688
rect 24914 16632 25686 16688
rect 25742 16632 25747 16688
rect 24853 16630 25747 16632
rect 24853 16627 24919 16630
rect 25681 16627 25747 16630
rect 4521 16554 4587 16557
rect 10593 16554 10659 16557
rect 15377 16554 15443 16557
rect 4521 16552 15762 16554
rect 4521 16496 4526 16552
rect 4582 16496 10598 16552
rect 10654 16496 15382 16552
rect 15438 16496 15762 16552
rect 4521 16494 15762 16496
rect 4521 16491 4587 16494
rect 10593 16491 10659 16494
rect 15377 16491 15443 16494
rect 0 16418 480 16448
rect 3877 16418 3943 16421
rect 0 16416 3943 16418
rect 0 16360 3882 16416
rect 3938 16360 3943 16416
rect 0 16358 3943 16360
rect 0 16328 480 16358
rect 3877 16355 3943 16358
rect 5944 16352 6264 16353
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 16287 6264 16288
rect 15702 16146 15762 16494
rect 29520 16418 30000 16448
rect 26374 16358 30000 16418
rect 15944 16352 16264 16353
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 16287 16264 16288
rect 25944 16352 26264 16353
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 16287 26264 16288
rect 25681 16282 25747 16285
rect 19198 16280 25747 16282
rect 19198 16224 25686 16280
rect 25742 16224 25747 16280
rect 19198 16222 25747 16224
rect 19198 16149 19258 16222
rect 25681 16219 25747 16222
rect 19149 16146 19258 16149
rect 15702 16144 19258 16146
rect 15702 16088 19154 16144
rect 19210 16088 19258 16144
rect 15702 16086 19258 16088
rect 19149 16083 19215 16086
rect 3601 16010 3667 16013
rect 10777 16010 10843 16013
rect 16021 16010 16087 16013
rect 19609 16010 19675 16013
rect 3601 16008 19675 16010
rect 3601 15952 3606 16008
rect 3662 15952 10782 16008
rect 10838 15952 16026 16008
rect 16082 15952 19614 16008
rect 19670 15952 19675 16008
rect 3601 15950 19675 15952
rect 3601 15947 3667 15950
rect 10777 15947 10843 15950
rect 16021 15947 16087 15950
rect 19609 15947 19675 15950
rect 20069 16010 20135 16013
rect 26374 16010 26434 16358
rect 29520 16328 30000 16358
rect 20069 16008 26434 16010
rect 20069 15952 20074 16008
rect 20130 15952 26434 16008
rect 20069 15950 26434 15952
rect 20069 15947 20135 15950
rect 0 15874 480 15904
rect 2773 15874 2839 15877
rect 0 15872 2839 15874
rect 0 15816 2778 15872
rect 2834 15816 2839 15872
rect 0 15814 2839 15816
rect 0 15784 480 15814
rect 2773 15811 2839 15814
rect 15745 15874 15811 15877
rect 18873 15874 18939 15877
rect 15745 15872 18939 15874
rect 15745 15816 15750 15872
rect 15806 15816 18878 15872
rect 18934 15816 18939 15872
rect 15745 15814 18939 15816
rect 15745 15811 15811 15814
rect 18873 15811 18939 15814
rect 25313 15874 25379 15877
rect 29520 15874 30000 15904
rect 25313 15872 30000 15874
rect 25313 15816 25318 15872
rect 25374 15816 30000 15872
rect 25313 15814 30000 15816
rect 25313 15811 25379 15814
rect 10944 15808 11264 15809
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 15743 11264 15744
rect 20944 15808 21264 15809
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 29520 15784 30000 15814
rect 20944 15743 21264 15744
rect 4429 15738 4495 15741
rect 10501 15738 10567 15741
rect 4429 15736 10567 15738
rect 4429 15680 4434 15736
rect 4490 15680 10506 15736
rect 10562 15680 10567 15736
rect 4429 15678 10567 15680
rect 4429 15675 4495 15678
rect 10501 15675 10567 15678
rect 13629 15602 13695 15605
rect 25497 15602 25563 15605
rect 13629 15600 25563 15602
rect 13629 15544 13634 15600
rect 13690 15544 25502 15600
rect 25558 15544 25563 15600
rect 13629 15542 25563 15544
rect 13629 15539 13695 15542
rect 25497 15539 25563 15542
rect 3141 15466 3207 15469
rect 9765 15466 9831 15469
rect 12801 15466 12867 15469
rect 3141 15464 12867 15466
rect 3141 15408 3146 15464
rect 3202 15408 9770 15464
rect 9826 15408 12806 15464
rect 12862 15408 12867 15464
rect 3141 15406 12867 15408
rect 3141 15403 3207 15406
rect 9765 15403 9831 15406
rect 12801 15403 12867 15406
rect 19609 15466 19675 15469
rect 25405 15466 25471 15469
rect 19609 15464 25471 15466
rect 19609 15408 19614 15464
rect 19670 15408 25410 15464
rect 25466 15408 25471 15464
rect 19609 15406 25471 15408
rect 19609 15403 19675 15406
rect 25405 15403 25471 15406
rect 25681 15466 25747 15469
rect 25681 15464 26434 15466
rect 25681 15408 25686 15464
rect 25742 15408 26434 15464
rect 25681 15406 26434 15408
rect 25681 15403 25747 15406
rect 0 15330 480 15360
rect 5533 15330 5599 15333
rect 0 15328 5599 15330
rect 0 15272 5538 15328
rect 5594 15272 5599 15328
rect 0 15270 5599 15272
rect 0 15240 480 15270
rect 5533 15267 5599 15270
rect 19885 15330 19951 15333
rect 24393 15330 24459 15333
rect 19885 15328 24459 15330
rect 19885 15272 19890 15328
rect 19946 15272 24398 15328
rect 24454 15272 24459 15328
rect 19885 15270 24459 15272
rect 26374 15330 26434 15406
rect 29520 15330 30000 15360
rect 26374 15270 30000 15330
rect 19885 15267 19951 15270
rect 24393 15267 24459 15270
rect 5944 15264 6264 15265
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 15199 6264 15200
rect 15944 15264 16264 15265
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 15199 16264 15200
rect 25944 15264 26264 15265
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 29520 15240 30000 15270
rect 25944 15199 26264 15200
rect 23657 15194 23723 15197
rect 17174 15192 24916 15194
rect 17174 15136 23662 15192
rect 23718 15136 24916 15192
rect 17174 15134 24916 15136
rect 11973 15058 12039 15061
rect 17174 15058 17234 15134
rect 23657 15131 23723 15134
rect 20529 15058 20595 15061
rect 21909 15058 21975 15061
rect 11973 15056 17234 15058
rect 11973 15000 11978 15056
rect 12034 15000 17234 15056
rect 19336 15056 21975 15058
rect 19336 15024 20534 15056
rect 11973 14998 17234 15000
rect 19152 15000 20534 15024
rect 20590 15000 21914 15056
rect 21970 15000 21975 15056
rect 19152 14998 21975 15000
rect 11973 14995 12039 14998
rect 19152 14964 19396 14998
rect 20529 14995 20595 14998
rect 21909 14995 21975 14998
rect 3233 14922 3299 14925
rect 19152 14922 19212 14964
rect 3233 14920 19212 14922
rect 3233 14864 3238 14920
rect 3294 14864 19212 14920
rect 3233 14862 19212 14864
rect 3233 14859 3299 14862
rect 10944 14720 11264 14721
rect 0 14650 480 14680
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 14655 11264 14656
rect 20944 14720 21264 14721
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 14655 21264 14656
rect 9857 14650 9923 14653
rect 0 14648 9923 14650
rect 0 14592 9862 14648
rect 9918 14592 9923 14648
rect 0 14590 9923 14592
rect 24856 14650 24916 15134
rect 29520 14650 30000 14680
rect 24856 14590 30000 14650
rect 0 14560 480 14590
rect 9857 14587 9923 14590
rect 29520 14560 30000 14590
rect 5944 14176 6264 14177
rect 0 14106 480 14136
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 14111 6264 14112
rect 15944 14176 16264 14177
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 14111 16264 14112
rect 25944 14176 26264 14177
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 14111 26264 14112
rect 4797 14106 4863 14109
rect 0 14104 4863 14106
rect 0 14048 4802 14104
rect 4858 14048 4863 14104
rect 0 14046 4863 14048
rect 0 14016 480 14046
rect 4797 14043 4863 14046
rect 27521 14106 27587 14109
rect 29520 14106 30000 14136
rect 27521 14104 30000 14106
rect 27521 14048 27526 14104
rect 27582 14048 30000 14104
rect 27521 14046 30000 14048
rect 27521 14043 27587 14046
rect 29520 14016 30000 14046
rect 13721 13834 13787 13837
rect 15009 13834 15075 13837
rect 15377 13834 15443 13837
rect 17769 13834 17835 13837
rect 10734 13774 11530 13834
rect 3877 13698 3943 13701
rect 6729 13698 6795 13701
rect 3877 13696 6795 13698
rect 3877 13640 3882 13696
rect 3938 13640 6734 13696
rect 6790 13640 6795 13696
rect 3877 13638 6795 13640
rect 3877 13635 3943 13638
rect 6729 13635 6795 13638
rect 8293 13698 8359 13701
rect 10734 13698 10794 13774
rect 8293 13696 10794 13698
rect 8293 13640 8298 13696
rect 8354 13640 10794 13696
rect 8293 13638 10794 13640
rect 11470 13698 11530 13774
rect 13721 13832 17835 13834
rect 13721 13776 13726 13832
rect 13782 13776 15014 13832
rect 15070 13776 15382 13832
rect 15438 13776 17774 13832
rect 17830 13776 17835 13832
rect 13721 13774 17835 13776
rect 13721 13771 13787 13774
rect 15009 13771 15075 13774
rect 15377 13771 15443 13774
rect 17769 13771 17835 13774
rect 20345 13834 20411 13837
rect 22645 13834 22711 13837
rect 20345 13832 22711 13834
rect 20345 13776 20350 13832
rect 20406 13776 22650 13832
rect 22706 13776 22711 13832
rect 20345 13774 22711 13776
rect 20345 13771 20411 13774
rect 22645 13771 22711 13774
rect 14825 13698 14891 13701
rect 18689 13698 18755 13701
rect 19701 13698 19767 13701
rect 11470 13696 19767 13698
rect 11470 13640 14830 13696
rect 14886 13640 18694 13696
rect 18750 13640 19706 13696
rect 19762 13640 19767 13696
rect 11470 13638 19767 13640
rect 8293 13635 8359 13638
rect 14825 13635 14891 13638
rect 18689 13635 18755 13638
rect 19701 13635 19767 13638
rect 10944 13632 11264 13633
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 13567 11264 13568
rect 20944 13632 21264 13633
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 13567 21264 13568
rect 15193 13562 15259 13565
rect 20437 13562 20503 13565
rect 15193 13560 20503 13562
rect 15193 13504 15198 13560
rect 15254 13504 20442 13560
rect 20498 13504 20503 13560
rect 15193 13502 20503 13504
rect 15193 13499 15259 13502
rect 20437 13499 20503 13502
rect 24393 13562 24459 13565
rect 24393 13560 25514 13562
rect 24393 13504 24398 13560
rect 24454 13504 25514 13560
rect 24393 13502 25514 13504
rect 24393 13499 24459 13502
rect 0 13426 480 13456
rect 3601 13426 3667 13429
rect 0 13424 3667 13426
rect 0 13368 3606 13424
rect 3662 13368 3667 13424
rect 0 13366 3667 13368
rect 0 13336 480 13366
rect 3601 13363 3667 13366
rect 19701 13426 19767 13429
rect 21817 13426 21883 13429
rect 19701 13424 21883 13426
rect 19701 13368 19706 13424
rect 19762 13368 21822 13424
rect 21878 13368 21883 13424
rect 19701 13366 21883 13368
rect 25454 13426 25514 13502
rect 29520 13426 30000 13456
rect 25454 13366 30000 13426
rect 19701 13363 19767 13366
rect 21817 13363 21883 13366
rect 29520 13336 30000 13366
rect 9622 13228 9628 13292
rect 9692 13290 9698 13292
rect 10777 13290 10843 13293
rect 9692 13288 10843 13290
rect 9692 13232 10782 13288
rect 10838 13232 10843 13288
rect 9692 13230 10843 13232
rect 9692 13228 9698 13230
rect 10777 13227 10843 13230
rect 11053 13290 11119 13293
rect 14089 13290 14155 13293
rect 11053 13288 14155 13290
rect 11053 13232 11058 13288
rect 11114 13232 14094 13288
rect 14150 13232 14155 13288
rect 11053 13230 14155 13232
rect 11053 13227 11119 13230
rect 14089 13227 14155 13230
rect 14273 13290 14339 13293
rect 25681 13290 25747 13293
rect 27521 13290 27587 13293
rect 14273 13288 25747 13290
rect 14273 13232 14278 13288
rect 14334 13232 25686 13288
rect 25742 13232 25747 13288
rect 14273 13230 25747 13232
rect 14273 13227 14339 13230
rect 25681 13227 25747 13230
rect 25822 13288 27587 13290
rect 25822 13232 27526 13288
rect 27582 13232 27587 13288
rect 25822 13230 27587 13232
rect 9581 13154 9647 13157
rect 10685 13154 10751 13157
rect 15193 13154 15259 13157
rect 9581 13152 15259 13154
rect 9581 13096 9586 13152
rect 9642 13096 10690 13152
rect 10746 13096 15198 13152
rect 15254 13096 15259 13152
rect 9581 13094 15259 13096
rect 9581 13091 9647 13094
rect 10685 13091 10751 13094
rect 15193 13091 15259 13094
rect 16389 13154 16455 13157
rect 24669 13154 24735 13157
rect 16389 13152 24735 13154
rect 16389 13096 16394 13152
rect 16450 13096 24674 13152
rect 24730 13096 24735 13152
rect 16389 13094 24735 13096
rect 16389 13091 16455 13094
rect 24669 13091 24735 13094
rect 5944 13088 6264 13089
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 13023 6264 13024
rect 15944 13088 16264 13089
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 13023 16264 13024
rect 9581 13018 9647 13021
rect 10961 13018 11027 13021
rect 9581 13016 11027 13018
rect 9581 12960 9586 13016
rect 9642 12960 10966 13016
rect 11022 12960 11027 13016
rect 9581 12958 11027 12960
rect 9581 12955 9647 12958
rect 10961 12955 11027 12958
rect 18781 13018 18847 13021
rect 20805 13018 20871 13021
rect 18781 13016 20871 13018
rect 18781 12960 18786 13016
rect 18842 12960 20810 13016
rect 20866 12960 20871 13016
rect 18781 12958 20871 12960
rect 18781 12955 18847 12958
rect 20805 12955 20871 12958
rect 21817 13018 21883 13021
rect 25822 13018 25882 13230
rect 27521 13227 27587 13230
rect 25944 13088 26264 13089
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 13023 26264 13024
rect 21817 13016 25882 13018
rect 21817 12960 21822 13016
rect 21878 12960 25882 13016
rect 21817 12958 25882 12960
rect 21817 12955 21883 12958
rect 0 12882 480 12912
rect 9581 12884 9647 12885
rect 0 12822 2698 12882
rect 0 12792 480 12822
rect 2638 12610 2698 12822
rect 9581 12880 9628 12884
rect 9692 12882 9698 12884
rect 17309 12882 17375 12885
rect 20897 12882 20963 12885
rect 9581 12824 9586 12880
rect 9581 12820 9628 12824
rect 9692 12822 9774 12882
rect 17309 12880 20963 12882
rect 17309 12824 17314 12880
rect 17370 12824 20902 12880
rect 20958 12824 20963 12880
rect 17309 12822 20963 12824
rect 9692 12820 9698 12822
rect 9581 12819 9647 12820
rect 17309 12819 17375 12822
rect 20897 12819 20963 12822
rect 24393 12882 24459 12885
rect 24669 12882 24735 12885
rect 24393 12880 24735 12882
rect 24393 12824 24398 12880
rect 24454 12824 24674 12880
rect 24730 12824 24735 12880
rect 24393 12822 24735 12824
rect 24393 12819 24459 12822
rect 24669 12819 24735 12822
rect 25957 12882 26023 12885
rect 29520 12882 30000 12912
rect 25957 12880 30000 12882
rect 25957 12824 25962 12880
rect 26018 12824 30000 12880
rect 25957 12822 30000 12824
rect 25957 12819 26023 12822
rect 29520 12792 30000 12822
rect 6361 12746 6427 12749
rect 9305 12746 9371 12749
rect 6361 12744 9371 12746
rect 6361 12688 6366 12744
rect 6422 12688 9310 12744
rect 9366 12688 9371 12744
rect 6361 12686 9371 12688
rect 6361 12683 6427 12686
rect 9305 12683 9371 12686
rect 9489 12746 9555 12749
rect 11145 12746 11211 12749
rect 9489 12744 11211 12746
rect 9489 12688 9494 12744
rect 9550 12688 11150 12744
rect 11206 12688 11211 12744
rect 9489 12686 11211 12688
rect 9489 12683 9555 12686
rect 11145 12683 11211 12686
rect 11421 12746 11487 12749
rect 26877 12746 26943 12749
rect 11421 12744 26943 12746
rect 11421 12688 11426 12744
rect 11482 12688 26882 12744
rect 26938 12688 26943 12744
rect 11421 12686 26943 12688
rect 11421 12683 11487 12686
rect 26877 12683 26943 12686
rect 3233 12610 3299 12613
rect 2638 12608 3299 12610
rect 2638 12552 3238 12608
rect 3294 12552 3299 12608
rect 2638 12550 3299 12552
rect 3233 12547 3299 12550
rect 3969 12610 4035 12613
rect 4337 12610 4403 12613
rect 3969 12608 4403 12610
rect 3969 12552 3974 12608
rect 4030 12552 4342 12608
rect 4398 12552 4403 12608
rect 3969 12550 4403 12552
rect 3969 12547 4035 12550
rect 4337 12547 4403 12550
rect 4889 12610 4955 12613
rect 10041 12610 10107 12613
rect 10593 12610 10659 12613
rect 4889 12608 10659 12610
rect 4889 12552 4894 12608
rect 4950 12552 10046 12608
rect 10102 12552 10598 12608
rect 10654 12552 10659 12608
rect 4889 12550 10659 12552
rect 4889 12547 4955 12550
rect 10041 12547 10107 12550
rect 10593 12547 10659 12550
rect 13445 12610 13511 12613
rect 14089 12610 14155 12613
rect 20161 12610 20227 12613
rect 13445 12608 20227 12610
rect 13445 12552 13450 12608
rect 13506 12552 14094 12608
rect 14150 12552 20166 12608
rect 20222 12552 20227 12608
rect 13445 12550 20227 12552
rect 13445 12547 13511 12550
rect 14089 12547 14155 12550
rect 20161 12547 20227 12550
rect 10944 12544 11264 12545
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 12479 11264 12480
rect 20944 12544 21264 12545
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 12479 21264 12480
rect 6637 12474 6703 12477
rect 10777 12474 10843 12477
rect 6637 12472 10843 12474
rect 6637 12416 6642 12472
rect 6698 12416 10782 12472
rect 10838 12416 10843 12472
rect 6637 12414 10843 12416
rect 6637 12411 6703 12414
rect 10777 12411 10843 12414
rect 13905 12474 13971 12477
rect 19701 12474 19767 12477
rect 25129 12474 25195 12477
rect 25497 12476 25563 12477
rect 13905 12472 19767 12474
rect 13905 12416 13910 12472
rect 13966 12416 19706 12472
rect 19762 12416 19767 12472
rect 13905 12414 19767 12416
rect 13905 12411 13971 12414
rect 19701 12411 19767 12414
rect 21406 12472 25195 12474
rect 21406 12416 25134 12472
rect 25190 12416 25195 12472
rect 21406 12414 25195 12416
rect 0 12338 480 12368
rect 3969 12338 4035 12341
rect 0 12336 4035 12338
rect 0 12280 3974 12336
rect 4030 12280 4035 12336
rect 0 12278 4035 12280
rect 0 12248 480 12278
rect 3969 12275 4035 12278
rect 5993 12338 6059 12341
rect 6269 12338 6335 12341
rect 8385 12338 8451 12341
rect 5993 12336 8451 12338
rect 5993 12280 5998 12336
rect 6054 12280 6274 12336
rect 6330 12280 8390 12336
rect 8446 12280 8451 12336
rect 5993 12278 8451 12280
rect 5993 12275 6059 12278
rect 6269 12275 6335 12278
rect 8385 12275 8451 12278
rect 9673 12338 9739 12341
rect 13629 12338 13695 12341
rect 13905 12338 13971 12341
rect 9673 12336 13971 12338
rect 9673 12280 9678 12336
rect 9734 12280 13634 12336
rect 13690 12280 13910 12336
rect 13966 12280 13971 12336
rect 9673 12278 13971 12280
rect 9673 12275 9739 12278
rect 13629 12275 13695 12278
rect 13905 12275 13971 12278
rect 15837 12338 15903 12341
rect 18413 12338 18479 12341
rect 15837 12336 18479 12338
rect 15837 12280 15842 12336
rect 15898 12280 18418 12336
rect 18474 12280 18479 12336
rect 15837 12278 18479 12280
rect 15837 12275 15903 12278
rect 18413 12275 18479 12278
rect 20161 12338 20227 12341
rect 21406 12338 21466 12414
rect 25129 12411 25195 12414
rect 25446 12412 25452 12476
rect 25516 12474 25563 12476
rect 25516 12472 25608 12474
rect 25558 12416 25608 12472
rect 25516 12414 25608 12416
rect 25516 12412 25563 12414
rect 25497 12411 25563 12412
rect 20161 12336 21466 12338
rect 20161 12280 20166 12336
rect 20222 12280 21466 12336
rect 20161 12278 21466 12280
rect 24761 12338 24827 12341
rect 26325 12338 26391 12341
rect 29520 12338 30000 12368
rect 24761 12336 30000 12338
rect 24761 12280 24766 12336
rect 24822 12280 26330 12336
rect 26386 12280 30000 12336
rect 24761 12278 30000 12280
rect 20161 12275 20227 12278
rect 24761 12275 24827 12278
rect 26325 12275 26391 12278
rect 29520 12248 30000 12278
rect 1485 12202 1551 12205
rect 2865 12202 2931 12205
rect 12893 12202 12959 12205
rect 25221 12202 25287 12205
rect 1485 12200 25287 12202
rect 1485 12144 1490 12200
rect 1546 12144 2870 12200
rect 2926 12144 12898 12200
rect 12954 12144 25226 12200
rect 25282 12144 25287 12200
rect 1485 12142 25287 12144
rect 1485 12139 1551 12142
rect 2865 12139 2931 12142
rect 12893 12139 12959 12142
rect 25221 12139 25287 12142
rect 5944 12000 6264 12001
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 11935 6264 11936
rect 15944 12000 16264 12001
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 11935 16264 11936
rect 25944 12000 26264 12001
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 11935 26264 11936
rect 2957 11794 3023 11797
rect 11329 11794 11395 11797
rect 2957 11792 11395 11794
rect 2957 11736 2962 11792
rect 3018 11736 11334 11792
rect 11390 11736 11395 11792
rect 2957 11734 11395 11736
rect 2957 11731 3023 11734
rect 11329 11731 11395 11734
rect 16665 11794 16731 11797
rect 25129 11794 25195 11797
rect 16665 11792 25195 11794
rect 16665 11736 16670 11792
rect 16726 11736 25134 11792
rect 25190 11736 25195 11792
rect 16665 11734 25195 11736
rect 16665 11731 16731 11734
rect 25129 11731 25195 11734
rect 0 11658 480 11688
rect 2681 11658 2747 11661
rect 0 11656 2747 11658
rect 0 11600 2686 11656
rect 2742 11600 2747 11656
rect 0 11598 2747 11600
rect 0 11568 480 11598
rect 2681 11595 2747 11598
rect 3417 11658 3483 11661
rect 15377 11658 15443 11661
rect 3417 11656 15443 11658
rect 3417 11600 3422 11656
rect 3478 11600 15382 11656
rect 15438 11600 15443 11656
rect 3417 11598 15443 11600
rect 3417 11595 3483 11598
rect 15377 11595 15443 11598
rect 16389 11658 16455 11661
rect 21817 11658 21883 11661
rect 16389 11656 21883 11658
rect 16389 11600 16394 11656
rect 16450 11600 21822 11656
rect 21878 11600 21883 11656
rect 16389 11598 21883 11600
rect 16389 11595 16455 11598
rect 21817 11595 21883 11598
rect 24301 11658 24367 11661
rect 26233 11658 26299 11661
rect 24301 11656 26299 11658
rect 24301 11600 24306 11656
rect 24362 11600 26238 11656
rect 26294 11600 26299 11656
rect 24301 11598 26299 11600
rect 24301 11595 24367 11598
rect 26233 11595 26299 11598
rect 26693 11658 26759 11661
rect 29520 11658 30000 11688
rect 26693 11656 30000 11658
rect 26693 11600 26698 11656
rect 26754 11600 30000 11656
rect 26693 11598 30000 11600
rect 26693 11595 26759 11598
rect 29520 11568 30000 11598
rect 11513 11522 11579 11525
rect 16297 11522 16363 11525
rect 19333 11522 19399 11525
rect 11513 11520 19399 11522
rect 11513 11464 11518 11520
rect 11574 11464 16302 11520
rect 16358 11464 19338 11520
rect 19394 11464 19399 11520
rect 11513 11462 19399 11464
rect 11513 11459 11579 11462
rect 16297 11459 16363 11462
rect 19333 11459 19399 11462
rect 10944 11456 11264 11457
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 11391 11264 11392
rect 20944 11456 21264 11457
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 11391 21264 11392
rect 5533 11386 5599 11389
rect 9673 11386 9739 11389
rect 5533 11384 9739 11386
rect 5533 11328 5538 11384
rect 5594 11328 9678 11384
rect 9734 11328 9739 11384
rect 5533 11326 9739 11328
rect 5533 11323 5599 11326
rect 9673 11323 9739 11326
rect 11329 11386 11395 11389
rect 20805 11386 20871 11389
rect 11329 11384 20871 11386
rect 11329 11328 11334 11384
rect 11390 11328 20810 11384
rect 20866 11328 20871 11384
rect 11329 11326 20871 11328
rect 11329 11323 11395 11326
rect 20805 11323 20871 11326
rect 2681 11250 2747 11253
rect 11421 11250 11487 11253
rect 15837 11250 15903 11253
rect 26417 11250 26483 11253
rect 2681 11248 26483 11250
rect 2681 11192 2686 11248
rect 2742 11192 11426 11248
rect 11482 11192 15842 11248
rect 15898 11192 26422 11248
rect 26478 11192 26483 11248
rect 2681 11190 26483 11192
rect 2681 11187 2747 11190
rect 11421 11187 11487 11190
rect 15837 11187 15903 11190
rect 26417 11187 26483 11190
rect 0 11114 480 11144
rect 1393 11114 1459 11117
rect 0 11112 1459 11114
rect 0 11056 1398 11112
rect 1454 11056 1459 11112
rect 0 11054 1459 11056
rect 0 11024 480 11054
rect 1393 11051 1459 11054
rect 19333 11114 19399 11117
rect 25405 11114 25471 11117
rect 19333 11112 25471 11114
rect 19333 11056 19338 11112
rect 19394 11056 25410 11112
rect 25466 11056 25471 11112
rect 19333 11054 25471 11056
rect 19333 11051 19399 11054
rect 25405 11051 25471 11054
rect 25865 11114 25931 11117
rect 29520 11114 30000 11144
rect 25865 11112 30000 11114
rect 25865 11056 25870 11112
rect 25926 11056 30000 11112
rect 25865 11054 30000 11056
rect 25865 11051 25931 11054
rect 29520 11024 30000 11054
rect 5944 10912 6264 10913
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 10847 6264 10848
rect 15944 10912 16264 10913
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 10847 16264 10848
rect 25944 10912 26264 10913
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 10847 26264 10848
rect 3509 10706 3575 10709
rect 9857 10706 9923 10709
rect 15561 10706 15627 10709
rect 3509 10704 15627 10706
rect 3509 10648 3514 10704
rect 3570 10648 9862 10704
rect 9918 10648 15566 10704
rect 15622 10648 15627 10704
rect 3509 10646 15627 10648
rect 3509 10643 3575 10646
rect 9857 10643 9923 10646
rect 15561 10643 15627 10646
rect 18413 10706 18479 10709
rect 27521 10706 27587 10709
rect 18413 10704 27587 10706
rect 18413 10648 18418 10704
rect 18474 10648 27526 10704
rect 27582 10648 27587 10704
rect 18413 10646 27587 10648
rect 18413 10643 18479 10646
rect 27521 10643 27587 10646
rect 6269 10570 6335 10573
rect 6729 10570 6795 10573
rect 18413 10570 18479 10573
rect 19517 10570 19583 10573
rect 21633 10570 21699 10573
rect 26417 10570 26483 10573
rect 6269 10568 21466 10570
rect 6269 10512 6274 10568
rect 6330 10512 6734 10568
rect 6790 10512 18418 10568
rect 18474 10512 19522 10568
rect 19578 10512 21466 10568
rect 6269 10510 21466 10512
rect 6269 10507 6335 10510
rect 6729 10507 6795 10510
rect 18413 10507 18479 10510
rect 19517 10507 19583 10510
rect 0 10434 480 10464
rect 1577 10434 1643 10437
rect 0 10432 1643 10434
rect 0 10376 1582 10432
rect 1638 10376 1643 10432
rect 0 10374 1643 10376
rect 0 10344 480 10374
rect 1577 10371 1643 10374
rect 6453 10434 6519 10437
rect 8385 10434 8451 10437
rect 6453 10432 8451 10434
rect 6453 10376 6458 10432
rect 6514 10376 8390 10432
rect 8446 10376 8451 10432
rect 6453 10374 8451 10376
rect 21406 10434 21466 10510
rect 21633 10568 26483 10570
rect 21633 10512 21638 10568
rect 21694 10512 26422 10568
rect 26478 10512 26483 10568
rect 21633 10510 26483 10512
rect 21633 10507 21699 10510
rect 26417 10507 26483 10510
rect 21633 10434 21699 10437
rect 21406 10432 21699 10434
rect 21406 10376 21638 10432
rect 21694 10376 21699 10432
rect 21406 10374 21699 10376
rect 6453 10371 6519 10374
rect 8385 10371 8451 10374
rect 21633 10371 21699 10374
rect 26601 10434 26667 10437
rect 29520 10434 30000 10464
rect 26601 10432 30000 10434
rect 26601 10376 26606 10432
rect 26662 10376 30000 10432
rect 26601 10374 30000 10376
rect 26601 10371 26667 10374
rect 10944 10368 11264 10369
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 10303 11264 10304
rect 20944 10368 21264 10369
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 29520 10344 30000 10374
rect 20944 10303 21264 10304
rect 2497 10298 2563 10301
rect 9949 10298 10015 10301
rect 2497 10296 10015 10298
rect 2497 10240 2502 10296
rect 2558 10240 9954 10296
rect 10010 10240 10015 10296
rect 2497 10238 10015 10240
rect 2497 10235 2563 10238
rect 9949 10235 10015 10238
rect 0 9890 480 9920
rect 2681 9890 2747 9893
rect 0 9888 2747 9890
rect 0 9832 2686 9888
rect 2742 9832 2747 9888
rect 0 9830 2747 9832
rect 0 9800 480 9830
rect 2681 9827 2747 9830
rect 26693 9890 26759 9893
rect 29520 9890 30000 9920
rect 26693 9888 30000 9890
rect 26693 9832 26698 9888
rect 26754 9832 30000 9888
rect 26693 9830 30000 9832
rect 26693 9827 26759 9830
rect 5944 9824 6264 9825
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 9759 6264 9760
rect 15944 9824 16264 9825
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 9759 16264 9760
rect 25944 9824 26264 9825
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 29520 9800 30000 9830
rect 25944 9759 26264 9760
rect 2037 9618 2103 9621
rect 7741 9618 7807 9621
rect 21265 9618 21331 9621
rect 24393 9618 24459 9621
rect 2037 9616 7666 9618
rect 2037 9560 2042 9616
rect 2098 9560 7666 9616
rect 2037 9558 7666 9560
rect 2037 9555 2103 9558
rect 1669 9482 1735 9485
rect 6545 9482 6611 9485
rect 1669 9480 6611 9482
rect 1669 9424 1674 9480
rect 1730 9424 6550 9480
rect 6606 9424 6611 9480
rect 1669 9422 6611 9424
rect 7606 9482 7666 9558
rect 7741 9616 24459 9618
rect 7741 9560 7746 9616
rect 7802 9560 21270 9616
rect 21326 9560 24398 9616
rect 24454 9560 24459 9616
rect 7741 9558 24459 9560
rect 7741 9555 7807 9558
rect 21265 9555 21331 9558
rect 24393 9555 24459 9558
rect 15285 9482 15351 9485
rect 7606 9480 15351 9482
rect 7606 9424 15290 9480
rect 15346 9424 15351 9480
rect 7606 9422 15351 9424
rect 1669 9419 1735 9422
rect 6545 9419 6611 9422
rect 15285 9419 15351 9422
rect 0 9346 480 9376
rect 1577 9346 1643 9349
rect 0 9344 1643 9346
rect 0 9288 1582 9344
rect 1638 9288 1643 9344
rect 0 9286 1643 9288
rect 0 9256 480 9286
rect 1577 9283 1643 9286
rect 26601 9346 26667 9349
rect 29520 9346 30000 9376
rect 26601 9344 30000 9346
rect 26601 9288 26606 9344
rect 26662 9288 30000 9344
rect 26601 9286 30000 9288
rect 26601 9283 26667 9286
rect 10944 9280 11264 9281
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 9215 11264 9216
rect 20944 9280 21264 9281
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 29520 9256 30000 9286
rect 20944 9215 21264 9216
rect 7281 9074 7347 9077
rect 15653 9074 15719 9077
rect 7281 9072 15719 9074
rect 7281 9016 7286 9072
rect 7342 9016 15658 9072
rect 15714 9016 15719 9072
rect 7281 9014 15719 9016
rect 7281 9011 7347 9014
rect 15653 9011 15719 9014
rect 16205 8938 16271 8941
rect 25865 8938 25931 8941
rect 16205 8936 25931 8938
rect 16205 8880 16210 8936
rect 16266 8880 25870 8936
rect 25926 8880 25931 8936
rect 16205 8878 25931 8880
rect 16205 8875 16271 8878
rect 25865 8875 25931 8878
rect 5944 8736 6264 8737
rect 0 8666 480 8696
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 8671 6264 8672
rect 15944 8736 16264 8737
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 8671 16264 8672
rect 25944 8736 26264 8737
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 8671 26264 8672
rect 1485 8666 1551 8669
rect 0 8664 1551 8666
rect 0 8608 1490 8664
rect 1546 8608 1551 8664
rect 0 8606 1551 8608
rect 0 8576 480 8606
rect 1485 8603 1551 8606
rect 17861 8666 17927 8669
rect 19425 8666 19491 8669
rect 17861 8664 19491 8666
rect 17861 8608 17866 8664
rect 17922 8608 19430 8664
rect 19486 8608 19491 8664
rect 17861 8606 19491 8608
rect 17861 8603 17927 8606
rect 19425 8603 19491 8606
rect 26693 8666 26759 8669
rect 29520 8666 30000 8696
rect 26693 8664 30000 8666
rect 26693 8608 26698 8664
rect 26754 8608 30000 8664
rect 26693 8606 30000 8608
rect 26693 8603 26759 8606
rect 29520 8576 30000 8606
rect 2865 8530 2931 8533
rect 16297 8530 16363 8533
rect 2865 8528 16363 8530
rect 2865 8472 2870 8528
rect 2926 8472 16302 8528
rect 16358 8472 16363 8528
rect 2865 8470 16363 8472
rect 2865 8467 2931 8470
rect 16297 8467 16363 8470
rect 10944 8192 11264 8193
rect 0 8122 480 8152
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 8127 11264 8128
rect 20944 8192 21264 8193
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 8127 21264 8128
rect 1393 8122 1459 8125
rect 0 8120 1459 8122
rect 0 8064 1398 8120
rect 1454 8064 1459 8120
rect 0 8062 1459 8064
rect 0 8032 480 8062
rect 1393 8059 1459 8062
rect 14457 8122 14523 8125
rect 20713 8122 20779 8125
rect 14457 8120 20779 8122
rect 14457 8064 14462 8120
rect 14518 8064 20718 8120
rect 20774 8064 20779 8120
rect 14457 8062 20779 8064
rect 14457 8059 14523 8062
rect 20713 8059 20779 8062
rect 27705 8122 27771 8125
rect 29520 8122 30000 8152
rect 27705 8120 30000 8122
rect 27705 8064 27710 8120
rect 27766 8064 30000 8120
rect 27705 8062 30000 8064
rect 27705 8059 27771 8062
rect 29520 8032 30000 8062
rect 2773 7986 2839 7989
rect 17401 7986 17467 7989
rect 2773 7984 17467 7986
rect 2773 7928 2778 7984
rect 2834 7928 17406 7984
rect 17462 7928 17467 7984
rect 2773 7926 17467 7928
rect 2773 7923 2839 7926
rect 17401 7923 17467 7926
rect 18413 7986 18479 7989
rect 26509 7986 26575 7989
rect 18413 7984 26575 7986
rect 18413 7928 18418 7984
rect 18474 7928 26514 7984
rect 26570 7928 26575 7984
rect 18413 7926 26575 7928
rect 18413 7923 18479 7926
rect 26509 7923 26575 7926
rect 5944 7648 6264 7649
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 7583 6264 7584
rect 15944 7648 16264 7649
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 7583 16264 7584
rect 25944 7648 26264 7649
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 7583 26264 7584
rect 3325 7578 3391 7581
rect 4981 7578 5047 7581
rect 16941 7578 17007 7581
rect 23473 7578 23539 7581
rect 3325 7576 5826 7578
rect 3325 7520 3330 7576
rect 3386 7520 4986 7576
rect 5042 7520 5826 7576
rect 3325 7518 5826 7520
rect 3325 7515 3391 7518
rect 4981 7515 5047 7518
rect 0 7442 480 7472
rect 1577 7442 1643 7445
rect 0 7440 1643 7442
rect 0 7384 1582 7440
rect 1638 7384 1643 7440
rect 0 7382 1643 7384
rect 5766 7442 5826 7518
rect 16941 7576 23539 7578
rect 16941 7520 16946 7576
rect 17002 7520 23478 7576
rect 23534 7520 23539 7576
rect 16941 7518 23539 7520
rect 16941 7515 17007 7518
rect 23473 7515 23539 7518
rect 12157 7442 12223 7445
rect 12801 7442 12867 7445
rect 23841 7442 23907 7445
rect 5766 7440 12867 7442
rect 5766 7384 12162 7440
rect 12218 7384 12806 7440
rect 12862 7384 12867 7440
rect 5766 7382 12867 7384
rect 0 7352 480 7382
rect 1577 7379 1643 7382
rect 12157 7379 12223 7382
rect 12801 7379 12867 7382
rect 18094 7440 23907 7442
rect 18094 7384 23846 7440
rect 23902 7384 23907 7440
rect 18094 7382 23907 7384
rect 18094 7309 18154 7382
rect 23841 7379 23907 7382
rect 24025 7442 24091 7445
rect 26509 7442 26575 7445
rect 24025 7440 26575 7442
rect 24025 7384 24030 7440
rect 24086 7384 26514 7440
rect 26570 7384 26575 7440
rect 24025 7382 26575 7384
rect 24025 7379 24091 7382
rect 26509 7379 26575 7382
rect 26693 7442 26759 7445
rect 29520 7442 30000 7472
rect 26693 7440 30000 7442
rect 26693 7384 26698 7440
rect 26754 7384 30000 7440
rect 26693 7382 30000 7384
rect 26693 7379 26759 7382
rect 29520 7352 30000 7382
rect 5625 7306 5691 7309
rect 18045 7306 18154 7309
rect 23105 7306 23171 7309
rect 5625 7304 18154 7306
rect 5625 7248 5630 7304
rect 5686 7248 18050 7304
rect 18106 7248 18154 7304
rect 5625 7246 18154 7248
rect 18278 7304 23171 7306
rect 18278 7248 23110 7304
rect 23166 7248 23171 7304
rect 18278 7246 23171 7248
rect 5625 7243 5691 7246
rect 18045 7243 18111 7246
rect 11789 7170 11855 7173
rect 16941 7170 17007 7173
rect 11789 7168 17007 7170
rect 11789 7112 11794 7168
rect 11850 7112 16946 7168
rect 17002 7112 17007 7168
rect 11789 7110 17007 7112
rect 11789 7107 11855 7110
rect 16941 7107 17007 7110
rect 17401 7170 17467 7173
rect 18278 7170 18338 7246
rect 23105 7243 23171 7246
rect 23657 7306 23723 7309
rect 25313 7306 25379 7309
rect 23657 7304 25379 7306
rect 23657 7248 23662 7304
rect 23718 7248 25318 7304
rect 25374 7248 25379 7304
rect 23657 7246 25379 7248
rect 23657 7243 23723 7246
rect 25313 7243 25379 7246
rect 17401 7168 18338 7170
rect 17401 7112 17406 7168
rect 17462 7112 18338 7168
rect 17401 7110 18338 7112
rect 17401 7107 17467 7110
rect 10944 7104 11264 7105
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 7039 11264 7040
rect 20944 7104 21264 7105
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 7039 21264 7040
rect 2957 7034 3023 7037
rect 4613 7034 4679 7037
rect 2957 7032 4679 7034
rect 2957 6976 2962 7032
rect 3018 6976 4618 7032
rect 4674 6976 4679 7032
rect 2957 6974 4679 6976
rect 2957 6971 3023 6974
rect 4613 6971 4679 6974
rect 24117 7034 24183 7037
rect 26325 7034 26391 7037
rect 24117 7032 26391 7034
rect 24117 6976 24122 7032
rect 24178 6976 26330 7032
rect 26386 6976 26391 7032
rect 24117 6974 26391 6976
rect 24117 6971 24183 6974
rect 26325 6971 26391 6974
rect 0 6898 480 6928
rect 1761 6898 1827 6901
rect 0 6896 1827 6898
rect 0 6840 1766 6896
rect 1822 6840 1827 6896
rect 0 6838 1827 6840
rect 0 6808 480 6838
rect 1761 6835 1827 6838
rect 2497 6898 2563 6901
rect 5625 6898 5691 6901
rect 2497 6896 5691 6898
rect 2497 6840 2502 6896
rect 2558 6840 5630 6896
rect 5686 6840 5691 6896
rect 2497 6838 5691 6840
rect 2497 6835 2563 6838
rect 5625 6835 5691 6838
rect 5993 6898 6059 6901
rect 13721 6898 13787 6901
rect 18505 6898 18571 6901
rect 25589 6898 25655 6901
rect 5993 6896 25655 6898
rect 5993 6840 5998 6896
rect 6054 6840 13726 6896
rect 13782 6840 18510 6896
rect 18566 6840 25594 6896
rect 25650 6840 25655 6896
rect 5993 6838 25655 6840
rect 5993 6835 6059 6838
rect 13721 6835 13787 6838
rect 18505 6835 18571 6838
rect 25589 6835 25655 6838
rect 25773 6898 25839 6901
rect 29520 6898 30000 6928
rect 25773 6896 30000 6898
rect 25773 6840 25778 6896
rect 25834 6840 30000 6896
rect 25773 6838 30000 6840
rect 25773 6835 25839 6838
rect 29520 6808 30000 6838
rect 13445 6762 13511 6765
rect 16297 6762 16363 6765
rect 21909 6762 21975 6765
rect 13445 6760 21975 6762
rect 13445 6704 13450 6760
rect 13506 6704 16302 6760
rect 16358 6704 21914 6760
rect 21970 6704 21975 6760
rect 13445 6702 21975 6704
rect 13445 6699 13511 6702
rect 16297 6699 16363 6702
rect 21909 6699 21975 6702
rect 22369 6762 22435 6765
rect 26969 6762 27035 6765
rect 22369 6760 27035 6762
rect 22369 6704 22374 6760
rect 22430 6704 26974 6760
rect 27030 6704 27035 6760
rect 22369 6702 27035 6704
rect 22369 6699 22435 6702
rect 26969 6699 27035 6702
rect 5944 6560 6264 6561
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 6495 6264 6496
rect 15944 6560 16264 6561
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 6495 16264 6496
rect 25944 6560 26264 6561
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 6495 26264 6496
rect 2037 6490 2103 6493
rect 5441 6490 5507 6493
rect 2037 6488 5507 6490
rect 2037 6432 2042 6488
rect 2098 6432 5446 6488
rect 5502 6432 5507 6488
rect 2037 6430 5507 6432
rect 2037 6427 2103 6430
rect 5441 6427 5507 6430
rect 0 6354 480 6384
rect 3693 6354 3759 6357
rect 0 6352 3759 6354
rect 0 6296 3698 6352
rect 3754 6296 3759 6352
rect 0 6294 3759 6296
rect 0 6264 480 6294
rect 3693 6291 3759 6294
rect 26785 6354 26851 6357
rect 29520 6354 30000 6384
rect 26785 6352 30000 6354
rect 26785 6296 26790 6352
rect 26846 6296 30000 6352
rect 26785 6294 30000 6296
rect 26785 6291 26851 6294
rect 29520 6264 30000 6294
rect 15561 6218 15627 6221
rect 26233 6218 26299 6221
rect 15561 6216 26299 6218
rect 15561 6160 15566 6216
rect 15622 6160 26238 6216
rect 26294 6160 26299 6216
rect 15561 6158 26299 6160
rect 15561 6155 15627 6158
rect 26233 6155 26299 6158
rect 10944 6016 11264 6017
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 5951 11264 5952
rect 20944 6016 21264 6017
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 5951 21264 5952
rect 7925 5810 7991 5813
rect 21173 5810 21239 5813
rect 26417 5810 26483 5813
rect 7925 5808 26483 5810
rect 7925 5752 7930 5808
rect 7986 5752 21178 5808
rect 21234 5752 26422 5808
rect 26478 5752 26483 5808
rect 7925 5750 26483 5752
rect 7925 5747 7991 5750
rect 21173 5747 21239 5750
rect 26417 5747 26483 5750
rect 0 5674 480 5704
rect 1577 5674 1643 5677
rect 0 5672 1643 5674
rect 0 5616 1582 5672
rect 1638 5616 1643 5672
rect 0 5614 1643 5616
rect 0 5584 480 5614
rect 1577 5611 1643 5614
rect 17493 5674 17559 5677
rect 23565 5674 23631 5677
rect 17493 5672 23631 5674
rect 17493 5616 17498 5672
rect 17554 5616 23570 5672
rect 23626 5616 23631 5672
rect 17493 5614 23631 5616
rect 17493 5611 17559 5614
rect 23565 5611 23631 5614
rect 26601 5674 26667 5677
rect 29520 5674 30000 5704
rect 26601 5672 30000 5674
rect 26601 5616 26606 5672
rect 26662 5616 30000 5672
rect 26601 5614 30000 5616
rect 26601 5611 26667 5614
rect 29520 5584 30000 5614
rect 5944 5472 6264 5473
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 5407 6264 5408
rect 15944 5472 16264 5473
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 5407 16264 5408
rect 25944 5472 26264 5473
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 5407 26264 5408
rect 2037 5266 2103 5269
rect 6453 5266 6519 5269
rect 2037 5264 6519 5266
rect 2037 5208 2042 5264
rect 2098 5208 6458 5264
rect 6514 5208 6519 5264
rect 2037 5206 6519 5208
rect 2037 5203 2103 5206
rect 6453 5203 6519 5206
rect 6637 5266 6703 5269
rect 7649 5266 7715 5269
rect 20253 5266 20319 5269
rect 6637 5264 20319 5266
rect 6637 5208 6642 5264
rect 6698 5208 7654 5264
rect 7710 5208 20258 5264
rect 20314 5208 20319 5264
rect 6637 5206 20319 5208
rect 6637 5203 6703 5206
rect 7649 5203 7715 5206
rect 20253 5203 20319 5206
rect 0 5130 480 5160
rect 1577 5130 1643 5133
rect 0 5128 1643 5130
rect 0 5072 1582 5128
rect 1638 5072 1643 5128
rect 0 5070 1643 5072
rect 0 5040 480 5070
rect 1577 5067 1643 5070
rect 1853 5130 1919 5133
rect 6640 5130 6700 5203
rect 1853 5128 6700 5130
rect 1853 5072 1858 5128
rect 1914 5072 6700 5128
rect 1853 5070 6700 5072
rect 10225 5130 10291 5133
rect 26233 5130 26299 5133
rect 10225 5128 26299 5130
rect 10225 5072 10230 5128
rect 10286 5072 26238 5128
rect 26294 5072 26299 5128
rect 10225 5070 26299 5072
rect 1853 5067 1919 5070
rect 10225 5067 10291 5070
rect 26233 5067 26299 5070
rect 26601 5130 26667 5133
rect 29520 5130 30000 5160
rect 26601 5128 30000 5130
rect 26601 5072 26606 5128
rect 26662 5072 30000 5128
rect 26601 5070 30000 5072
rect 26601 5067 26667 5070
rect 29520 5040 30000 5070
rect 10944 4928 11264 4929
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 4863 11264 4864
rect 20944 4928 21264 4929
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 4863 21264 4864
rect 13261 4858 13327 4861
rect 17493 4858 17559 4861
rect 13261 4856 17559 4858
rect 13261 4800 13266 4856
rect 13322 4800 17498 4856
rect 17554 4800 17559 4856
rect 13261 4798 17559 4800
rect 13261 4795 13327 4798
rect 17493 4795 17559 4798
rect 2037 4722 2103 4725
rect 11697 4722 11763 4725
rect 2037 4720 11763 4722
rect 2037 4664 2042 4720
rect 2098 4664 11702 4720
rect 11758 4664 11763 4720
rect 2037 4662 11763 4664
rect 2037 4659 2103 4662
rect 11697 4659 11763 4662
rect 14917 4722 14983 4725
rect 26509 4722 26575 4725
rect 14917 4720 26575 4722
rect 14917 4664 14922 4720
rect 14978 4664 26514 4720
rect 26570 4664 26575 4720
rect 14917 4662 26575 4664
rect 14917 4659 14983 4662
rect 26509 4659 26575 4662
rect 19885 4586 19951 4589
rect 23565 4586 23631 4589
rect 19885 4584 23631 4586
rect 19885 4528 19890 4584
rect 19946 4528 23570 4584
rect 23626 4528 23631 4584
rect 19885 4526 23631 4528
rect 19885 4523 19951 4526
rect 23565 4523 23631 4526
rect 0 4450 480 4480
rect 1577 4450 1643 4453
rect 0 4448 1643 4450
rect 0 4392 1582 4448
rect 1638 4392 1643 4448
rect 0 4390 1643 4392
rect 0 4360 480 4390
rect 1577 4387 1643 4390
rect 27705 4450 27771 4453
rect 29520 4450 30000 4480
rect 27705 4448 30000 4450
rect 27705 4392 27710 4448
rect 27766 4392 30000 4448
rect 27705 4390 30000 4392
rect 27705 4387 27771 4390
rect 5944 4384 6264 4385
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 4319 6264 4320
rect 15944 4384 16264 4385
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 4319 16264 4320
rect 25944 4384 26264 4385
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 29520 4360 30000 4390
rect 25944 4319 26264 4320
rect 1945 4178 2011 4181
rect 3417 4178 3483 4181
rect 13261 4178 13327 4181
rect 1945 4176 13327 4178
rect 1945 4120 1950 4176
rect 2006 4120 3422 4176
rect 3478 4120 13266 4176
rect 13322 4120 13327 4176
rect 1945 4118 13327 4120
rect 1945 4115 2011 4118
rect 3417 4115 3483 4118
rect 13261 4115 13327 4118
rect 15653 4178 15719 4181
rect 19241 4178 19307 4181
rect 15653 4176 19307 4178
rect 15653 4120 15658 4176
rect 15714 4120 19246 4176
rect 19302 4120 19307 4176
rect 15653 4118 19307 4120
rect 15653 4115 15719 4118
rect 19241 4115 19307 4118
rect 4613 4042 4679 4045
rect 11605 4042 11671 4045
rect 4613 4040 11671 4042
rect 4613 3984 4618 4040
rect 4674 3984 11610 4040
rect 11666 3984 11671 4040
rect 4613 3982 11671 3984
rect 4613 3979 4679 3982
rect 11605 3979 11671 3982
rect 12065 4042 12131 4045
rect 26417 4042 26483 4045
rect 12065 4040 26483 4042
rect 12065 3984 12070 4040
rect 12126 3984 26422 4040
rect 26478 3984 26483 4040
rect 12065 3982 26483 3984
rect 12065 3979 12131 3982
rect 26417 3979 26483 3982
rect 0 3906 480 3936
rect 2681 3906 2747 3909
rect 0 3904 2747 3906
rect 0 3848 2686 3904
rect 2742 3848 2747 3904
rect 0 3846 2747 3848
rect 0 3816 480 3846
rect 2681 3843 2747 3846
rect 5809 3906 5875 3909
rect 9029 3906 9095 3909
rect 5809 3904 9095 3906
rect 5809 3848 5814 3904
rect 5870 3848 9034 3904
rect 9090 3848 9095 3904
rect 5809 3846 9095 3848
rect 5809 3843 5875 3846
rect 9029 3843 9095 3846
rect 26785 3906 26851 3909
rect 29520 3906 30000 3936
rect 26785 3904 30000 3906
rect 26785 3848 26790 3904
rect 26846 3848 30000 3904
rect 26785 3846 30000 3848
rect 26785 3843 26851 3846
rect 10944 3840 11264 3841
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 3775 11264 3776
rect 20944 3840 21264 3841
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 29520 3816 30000 3846
rect 20944 3775 21264 3776
rect 24853 3770 24919 3773
rect 27429 3770 27495 3773
rect 24853 3768 27495 3770
rect 24853 3712 24858 3768
rect 24914 3712 27434 3768
rect 27490 3712 27495 3768
rect 24853 3710 27495 3712
rect 24853 3707 24919 3710
rect 27429 3707 27495 3710
rect 4061 3634 4127 3637
rect 4429 3634 4495 3637
rect 12341 3634 12407 3637
rect 4061 3632 12407 3634
rect 4061 3576 4066 3632
rect 4122 3576 4434 3632
rect 4490 3576 12346 3632
rect 12402 3576 12407 3632
rect 4061 3574 12407 3576
rect 4061 3571 4127 3574
rect 4429 3571 4495 3574
rect 12341 3571 12407 3574
rect 20621 3634 20687 3637
rect 27521 3634 27587 3637
rect 20621 3632 27587 3634
rect 20621 3576 20626 3632
rect 20682 3576 27526 3632
rect 27582 3576 27587 3632
rect 20621 3574 27587 3576
rect 20621 3571 20687 3574
rect 27521 3571 27587 3574
rect 4245 3498 4311 3501
rect 9949 3498 10015 3501
rect 17309 3498 17375 3501
rect 4245 3496 17375 3498
rect 4245 3440 4250 3496
rect 4306 3440 9954 3496
rect 10010 3440 17314 3496
rect 17370 3440 17375 3496
rect 4245 3438 17375 3440
rect 4245 3435 4311 3438
rect 9949 3435 10015 3438
rect 17309 3435 17375 3438
rect 0 3362 480 3392
rect 4521 3362 4587 3365
rect 0 3360 4587 3362
rect 0 3304 4526 3360
rect 4582 3304 4587 3360
rect 0 3302 4587 3304
rect 0 3272 480 3302
rect 4521 3299 4587 3302
rect 26877 3362 26943 3365
rect 29520 3362 30000 3392
rect 26877 3360 30000 3362
rect 26877 3304 26882 3360
rect 26938 3304 30000 3360
rect 26877 3302 30000 3304
rect 26877 3299 26943 3302
rect 5944 3296 6264 3297
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 3231 6264 3232
rect 15944 3296 16264 3297
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 3231 16264 3232
rect 25944 3296 26264 3297
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 29520 3272 30000 3302
rect 25944 3231 26264 3232
rect 3325 3090 3391 3093
rect 6545 3090 6611 3093
rect 3325 3088 6611 3090
rect 3325 3032 3330 3088
rect 3386 3032 6550 3088
rect 6606 3032 6611 3088
rect 3325 3030 6611 3032
rect 3325 3027 3391 3030
rect 6545 3027 6611 3030
rect 17861 3090 17927 3093
rect 18873 3090 18939 3093
rect 25681 3090 25747 3093
rect 17861 3088 25747 3090
rect 17861 3032 17866 3088
rect 17922 3032 18878 3088
rect 18934 3032 25686 3088
rect 25742 3032 25747 3088
rect 17861 3030 25747 3032
rect 17861 3027 17927 3030
rect 18873 3027 18939 3030
rect 25681 3027 25747 3030
rect 657 2954 723 2957
rect 23841 2954 23907 2957
rect 657 2952 23907 2954
rect 657 2896 662 2952
rect 718 2896 23846 2952
rect 23902 2896 23907 2952
rect 657 2894 23907 2896
rect 657 2891 723 2894
rect 23841 2891 23907 2894
rect 26693 2818 26759 2821
rect 26693 2816 26986 2818
rect 26693 2760 26698 2816
rect 26754 2760 26986 2816
rect 26693 2758 26986 2760
rect 26693 2755 26759 2758
rect 10944 2752 11264 2753
rect 0 2682 480 2712
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2687 11264 2688
rect 20944 2752 21264 2753
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2687 21264 2688
rect 4061 2682 4127 2685
rect 0 2680 4127 2682
rect 0 2624 4066 2680
rect 4122 2624 4127 2680
rect 0 2622 4127 2624
rect 0 2592 480 2622
rect 4061 2619 4127 2622
rect 16849 2682 16915 2685
rect 20805 2682 20871 2685
rect 16849 2680 20871 2682
rect 16849 2624 16854 2680
rect 16910 2624 20810 2680
rect 20866 2624 20871 2680
rect 16849 2622 20871 2624
rect 26926 2682 26986 2758
rect 29520 2682 30000 2712
rect 26926 2622 30000 2682
rect 16849 2619 16915 2622
rect 20805 2619 20871 2622
rect 29520 2592 30000 2622
rect 5944 2208 6264 2209
rect 0 2138 480 2168
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2143 6264 2144
rect 15944 2208 16264 2209
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2143 16264 2144
rect 25944 2208 26264 2209
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2143 26264 2144
rect 5809 2138 5875 2141
rect 0 2136 5875 2138
rect 0 2080 5814 2136
rect 5870 2080 5875 2136
rect 0 2078 5875 2080
rect 0 2048 480 2078
rect 5809 2075 5875 2078
rect 27705 2138 27771 2141
rect 29520 2138 30000 2168
rect 27705 2136 30000 2138
rect 27705 2080 27710 2136
rect 27766 2080 30000 2136
rect 27705 2078 30000 2080
rect 27705 2075 27771 2078
rect 29520 2048 30000 2078
rect 0 1458 480 1488
rect 2129 1458 2195 1461
rect 0 1456 2195 1458
rect 0 1400 2134 1456
rect 2190 1400 2195 1456
rect 0 1398 2195 1400
rect 0 1368 480 1398
rect 2129 1395 2195 1398
rect 26785 1458 26851 1461
rect 29520 1458 30000 1488
rect 26785 1456 30000 1458
rect 26785 1400 26790 1456
rect 26846 1400 30000 1456
rect 26785 1398 30000 1400
rect 26785 1395 26851 1398
rect 29520 1368 30000 1398
rect 0 914 480 944
rect 4061 914 4127 917
rect 0 912 4127 914
rect 0 856 4066 912
rect 4122 856 4127 912
rect 0 854 4127 856
rect 0 824 480 854
rect 4061 851 4127 854
rect 25865 914 25931 917
rect 29520 914 30000 944
rect 25865 912 30000 914
rect 25865 856 25870 912
rect 25926 856 30000 912
rect 25865 854 30000 856
rect 25865 851 25931 854
rect 29520 824 30000 854
rect 0 370 480 400
rect 3969 370 4035 373
rect 0 368 4035 370
rect 0 312 3974 368
rect 4030 312 4035 368
rect 0 310 4035 312
rect 0 280 480 310
rect 3969 307 4035 310
rect 26601 370 26667 373
rect 29520 370 30000 400
rect 26601 368 30000 370
rect 26601 312 26606 368
rect 26662 312 30000 368
rect 26601 310 30000 312
rect 26601 307 26667 310
rect 29520 280 30000 310
<< via3 >>
rect 5952 21788 6016 21792
rect 5952 21732 5956 21788
rect 5956 21732 6012 21788
rect 6012 21732 6016 21788
rect 5952 21728 6016 21732
rect 6032 21788 6096 21792
rect 6032 21732 6036 21788
rect 6036 21732 6092 21788
rect 6092 21732 6096 21788
rect 6032 21728 6096 21732
rect 6112 21788 6176 21792
rect 6112 21732 6116 21788
rect 6116 21732 6172 21788
rect 6172 21732 6176 21788
rect 6112 21728 6176 21732
rect 6192 21788 6256 21792
rect 6192 21732 6196 21788
rect 6196 21732 6252 21788
rect 6252 21732 6256 21788
rect 6192 21728 6256 21732
rect 15952 21788 16016 21792
rect 15952 21732 15956 21788
rect 15956 21732 16012 21788
rect 16012 21732 16016 21788
rect 15952 21728 16016 21732
rect 16032 21788 16096 21792
rect 16032 21732 16036 21788
rect 16036 21732 16092 21788
rect 16092 21732 16096 21788
rect 16032 21728 16096 21732
rect 16112 21788 16176 21792
rect 16112 21732 16116 21788
rect 16116 21732 16172 21788
rect 16172 21732 16176 21788
rect 16112 21728 16176 21732
rect 16192 21788 16256 21792
rect 16192 21732 16196 21788
rect 16196 21732 16252 21788
rect 16252 21732 16256 21788
rect 16192 21728 16256 21732
rect 25952 21788 26016 21792
rect 25952 21732 25956 21788
rect 25956 21732 26012 21788
rect 26012 21732 26016 21788
rect 25952 21728 26016 21732
rect 26032 21788 26096 21792
rect 26032 21732 26036 21788
rect 26036 21732 26092 21788
rect 26092 21732 26096 21788
rect 26032 21728 26096 21732
rect 26112 21788 26176 21792
rect 26112 21732 26116 21788
rect 26116 21732 26172 21788
rect 26172 21732 26176 21788
rect 26112 21728 26176 21732
rect 26192 21788 26256 21792
rect 26192 21732 26196 21788
rect 26196 21732 26252 21788
rect 26252 21732 26256 21788
rect 26192 21728 26256 21732
rect 10952 21244 11016 21248
rect 10952 21188 10956 21244
rect 10956 21188 11012 21244
rect 11012 21188 11016 21244
rect 10952 21184 11016 21188
rect 11032 21244 11096 21248
rect 11032 21188 11036 21244
rect 11036 21188 11092 21244
rect 11092 21188 11096 21244
rect 11032 21184 11096 21188
rect 11112 21244 11176 21248
rect 11112 21188 11116 21244
rect 11116 21188 11172 21244
rect 11172 21188 11176 21244
rect 11112 21184 11176 21188
rect 11192 21244 11256 21248
rect 11192 21188 11196 21244
rect 11196 21188 11252 21244
rect 11252 21188 11256 21244
rect 11192 21184 11256 21188
rect 20952 21244 21016 21248
rect 20952 21188 20956 21244
rect 20956 21188 21012 21244
rect 21012 21188 21016 21244
rect 20952 21184 21016 21188
rect 21032 21244 21096 21248
rect 21032 21188 21036 21244
rect 21036 21188 21092 21244
rect 21092 21188 21096 21244
rect 21032 21184 21096 21188
rect 21112 21244 21176 21248
rect 21112 21188 21116 21244
rect 21116 21188 21172 21244
rect 21172 21188 21176 21244
rect 21112 21184 21176 21188
rect 21192 21244 21256 21248
rect 21192 21188 21196 21244
rect 21196 21188 21252 21244
rect 21252 21188 21256 21244
rect 21192 21184 21256 21188
rect 5952 20700 6016 20704
rect 5952 20644 5956 20700
rect 5956 20644 6012 20700
rect 6012 20644 6016 20700
rect 5952 20640 6016 20644
rect 6032 20700 6096 20704
rect 6032 20644 6036 20700
rect 6036 20644 6092 20700
rect 6092 20644 6096 20700
rect 6032 20640 6096 20644
rect 6112 20700 6176 20704
rect 6112 20644 6116 20700
rect 6116 20644 6172 20700
rect 6172 20644 6176 20700
rect 6112 20640 6176 20644
rect 6192 20700 6256 20704
rect 6192 20644 6196 20700
rect 6196 20644 6252 20700
rect 6252 20644 6256 20700
rect 6192 20640 6256 20644
rect 15952 20700 16016 20704
rect 15952 20644 15956 20700
rect 15956 20644 16012 20700
rect 16012 20644 16016 20700
rect 15952 20640 16016 20644
rect 16032 20700 16096 20704
rect 16032 20644 16036 20700
rect 16036 20644 16092 20700
rect 16092 20644 16096 20700
rect 16032 20640 16096 20644
rect 16112 20700 16176 20704
rect 16112 20644 16116 20700
rect 16116 20644 16172 20700
rect 16172 20644 16176 20700
rect 16112 20640 16176 20644
rect 16192 20700 16256 20704
rect 16192 20644 16196 20700
rect 16196 20644 16252 20700
rect 16252 20644 16256 20700
rect 16192 20640 16256 20644
rect 25952 20700 26016 20704
rect 25952 20644 25956 20700
rect 25956 20644 26012 20700
rect 26012 20644 26016 20700
rect 25952 20640 26016 20644
rect 26032 20700 26096 20704
rect 26032 20644 26036 20700
rect 26036 20644 26092 20700
rect 26092 20644 26096 20700
rect 26032 20640 26096 20644
rect 26112 20700 26176 20704
rect 26112 20644 26116 20700
rect 26116 20644 26172 20700
rect 26172 20644 26176 20700
rect 26112 20640 26176 20644
rect 26192 20700 26256 20704
rect 26192 20644 26196 20700
rect 26196 20644 26252 20700
rect 26252 20644 26256 20700
rect 26192 20640 26256 20644
rect 10952 20156 11016 20160
rect 10952 20100 10956 20156
rect 10956 20100 11012 20156
rect 11012 20100 11016 20156
rect 10952 20096 11016 20100
rect 11032 20156 11096 20160
rect 11032 20100 11036 20156
rect 11036 20100 11092 20156
rect 11092 20100 11096 20156
rect 11032 20096 11096 20100
rect 11112 20156 11176 20160
rect 11112 20100 11116 20156
rect 11116 20100 11172 20156
rect 11172 20100 11176 20156
rect 11112 20096 11176 20100
rect 11192 20156 11256 20160
rect 11192 20100 11196 20156
rect 11196 20100 11252 20156
rect 11252 20100 11256 20156
rect 11192 20096 11256 20100
rect 20952 20156 21016 20160
rect 20952 20100 20956 20156
rect 20956 20100 21012 20156
rect 21012 20100 21016 20156
rect 20952 20096 21016 20100
rect 21032 20156 21096 20160
rect 21032 20100 21036 20156
rect 21036 20100 21092 20156
rect 21092 20100 21096 20156
rect 21032 20096 21096 20100
rect 21112 20156 21176 20160
rect 21112 20100 21116 20156
rect 21116 20100 21172 20156
rect 21172 20100 21176 20156
rect 21112 20096 21176 20100
rect 21192 20156 21256 20160
rect 21192 20100 21196 20156
rect 21196 20100 21252 20156
rect 21252 20100 21256 20156
rect 21192 20096 21256 20100
rect 5952 19612 6016 19616
rect 5952 19556 5956 19612
rect 5956 19556 6012 19612
rect 6012 19556 6016 19612
rect 5952 19552 6016 19556
rect 6032 19612 6096 19616
rect 6032 19556 6036 19612
rect 6036 19556 6092 19612
rect 6092 19556 6096 19612
rect 6032 19552 6096 19556
rect 6112 19612 6176 19616
rect 6112 19556 6116 19612
rect 6116 19556 6172 19612
rect 6172 19556 6176 19612
rect 6112 19552 6176 19556
rect 6192 19612 6256 19616
rect 6192 19556 6196 19612
rect 6196 19556 6252 19612
rect 6252 19556 6256 19612
rect 6192 19552 6256 19556
rect 15952 19612 16016 19616
rect 15952 19556 15956 19612
rect 15956 19556 16012 19612
rect 16012 19556 16016 19612
rect 15952 19552 16016 19556
rect 16032 19612 16096 19616
rect 16032 19556 16036 19612
rect 16036 19556 16092 19612
rect 16092 19556 16096 19612
rect 16032 19552 16096 19556
rect 16112 19612 16176 19616
rect 16112 19556 16116 19612
rect 16116 19556 16172 19612
rect 16172 19556 16176 19612
rect 16112 19552 16176 19556
rect 16192 19612 16256 19616
rect 16192 19556 16196 19612
rect 16196 19556 16252 19612
rect 16252 19556 16256 19612
rect 16192 19552 16256 19556
rect 25952 19612 26016 19616
rect 25952 19556 25956 19612
rect 25956 19556 26012 19612
rect 26012 19556 26016 19612
rect 25952 19552 26016 19556
rect 26032 19612 26096 19616
rect 26032 19556 26036 19612
rect 26036 19556 26092 19612
rect 26092 19556 26096 19612
rect 26032 19552 26096 19556
rect 26112 19612 26176 19616
rect 26112 19556 26116 19612
rect 26116 19556 26172 19612
rect 26172 19556 26176 19612
rect 26112 19552 26176 19556
rect 26192 19612 26256 19616
rect 26192 19556 26196 19612
rect 26196 19556 26252 19612
rect 26252 19556 26256 19612
rect 26192 19552 26256 19556
rect 10952 19068 11016 19072
rect 10952 19012 10956 19068
rect 10956 19012 11012 19068
rect 11012 19012 11016 19068
rect 10952 19008 11016 19012
rect 11032 19068 11096 19072
rect 11032 19012 11036 19068
rect 11036 19012 11092 19068
rect 11092 19012 11096 19068
rect 11032 19008 11096 19012
rect 11112 19068 11176 19072
rect 11112 19012 11116 19068
rect 11116 19012 11172 19068
rect 11172 19012 11176 19068
rect 11112 19008 11176 19012
rect 11192 19068 11256 19072
rect 11192 19012 11196 19068
rect 11196 19012 11252 19068
rect 11252 19012 11256 19068
rect 11192 19008 11256 19012
rect 20952 19068 21016 19072
rect 20952 19012 20956 19068
rect 20956 19012 21012 19068
rect 21012 19012 21016 19068
rect 20952 19008 21016 19012
rect 21032 19068 21096 19072
rect 21032 19012 21036 19068
rect 21036 19012 21092 19068
rect 21092 19012 21096 19068
rect 21032 19008 21096 19012
rect 21112 19068 21176 19072
rect 21112 19012 21116 19068
rect 21116 19012 21172 19068
rect 21172 19012 21176 19068
rect 21112 19008 21176 19012
rect 21192 19068 21256 19072
rect 21192 19012 21196 19068
rect 21196 19012 21252 19068
rect 21252 19012 21256 19068
rect 21192 19008 21256 19012
rect 5952 18524 6016 18528
rect 5952 18468 5956 18524
rect 5956 18468 6012 18524
rect 6012 18468 6016 18524
rect 5952 18464 6016 18468
rect 6032 18524 6096 18528
rect 6032 18468 6036 18524
rect 6036 18468 6092 18524
rect 6092 18468 6096 18524
rect 6032 18464 6096 18468
rect 6112 18524 6176 18528
rect 6112 18468 6116 18524
rect 6116 18468 6172 18524
rect 6172 18468 6176 18524
rect 6112 18464 6176 18468
rect 6192 18524 6256 18528
rect 6192 18468 6196 18524
rect 6196 18468 6252 18524
rect 6252 18468 6256 18524
rect 6192 18464 6256 18468
rect 15952 18524 16016 18528
rect 15952 18468 15956 18524
rect 15956 18468 16012 18524
rect 16012 18468 16016 18524
rect 15952 18464 16016 18468
rect 16032 18524 16096 18528
rect 16032 18468 16036 18524
rect 16036 18468 16092 18524
rect 16092 18468 16096 18524
rect 16032 18464 16096 18468
rect 16112 18524 16176 18528
rect 16112 18468 16116 18524
rect 16116 18468 16172 18524
rect 16172 18468 16176 18524
rect 16112 18464 16176 18468
rect 16192 18524 16256 18528
rect 16192 18468 16196 18524
rect 16196 18468 16252 18524
rect 16252 18468 16256 18524
rect 16192 18464 16256 18468
rect 25952 18524 26016 18528
rect 25952 18468 25956 18524
rect 25956 18468 26012 18524
rect 26012 18468 26016 18524
rect 25952 18464 26016 18468
rect 26032 18524 26096 18528
rect 26032 18468 26036 18524
rect 26036 18468 26092 18524
rect 26092 18468 26096 18524
rect 26032 18464 26096 18468
rect 26112 18524 26176 18528
rect 26112 18468 26116 18524
rect 26116 18468 26172 18524
rect 26172 18468 26176 18524
rect 26112 18464 26176 18468
rect 26192 18524 26256 18528
rect 26192 18468 26196 18524
rect 26196 18468 26252 18524
rect 26252 18468 26256 18524
rect 26192 18464 26256 18468
rect 25452 18320 25516 18324
rect 25452 18264 25502 18320
rect 25502 18264 25516 18320
rect 25452 18260 25516 18264
rect 10952 17980 11016 17984
rect 10952 17924 10956 17980
rect 10956 17924 11012 17980
rect 11012 17924 11016 17980
rect 10952 17920 11016 17924
rect 11032 17980 11096 17984
rect 11032 17924 11036 17980
rect 11036 17924 11092 17980
rect 11092 17924 11096 17980
rect 11032 17920 11096 17924
rect 11112 17980 11176 17984
rect 11112 17924 11116 17980
rect 11116 17924 11172 17980
rect 11172 17924 11176 17980
rect 11112 17920 11176 17924
rect 11192 17980 11256 17984
rect 11192 17924 11196 17980
rect 11196 17924 11252 17980
rect 11252 17924 11256 17980
rect 11192 17920 11256 17924
rect 20952 17980 21016 17984
rect 20952 17924 20956 17980
rect 20956 17924 21012 17980
rect 21012 17924 21016 17980
rect 20952 17920 21016 17924
rect 21032 17980 21096 17984
rect 21032 17924 21036 17980
rect 21036 17924 21092 17980
rect 21092 17924 21096 17980
rect 21032 17920 21096 17924
rect 21112 17980 21176 17984
rect 21112 17924 21116 17980
rect 21116 17924 21172 17980
rect 21172 17924 21176 17980
rect 21112 17920 21176 17924
rect 21192 17980 21256 17984
rect 21192 17924 21196 17980
rect 21196 17924 21252 17980
rect 21252 17924 21256 17980
rect 21192 17920 21256 17924
rect 5952 17436 6016 17440
rect 5952 17380 5956 17436
rect 5956 17380 6012 17436
rect 6012 17380 6016 17436
rect 5952 17376 6016 17380
rect 6032 17436 6096 17440
rect 6032 17380 6036 17436
rect 6036 17380 6092 17436
rect 6092 17380 6096 17436
rect 6032 17376 6096 17380
rect 6112 17436 6176 17440
rect 6112 17380 6116 17436
rect 6116 17380 6172 17436
rect 6172 17380 6176 17436
rect 6112 17376 6176 17380
rect 6192 17436 6256 17440
rect 6192 17380 6196 17436
rect 6196 17380 6252 17436
rect 6252 17380 6256 17436
rect 6192 17376 6256 17380
rect 15952 17436 16016 17440
rect 15952 17380 15956 17436
rect 15956 17380 16012 17436
rect 16012 17380 16016 17436
rect 15952 17376 16016 17380
rect 16032 17436 16096 17440
rect 16032 17380 16036 17436
rect 16036 17380 16092 17436
rect 16092 17380 16096 17436
rect 16032 17376 16096 17380
rect 16112 17436 16176 17440
rect 16112 17380 16116 17436
rect 16116 17380 16172 17436
rect 16172 17380 16176 17436
rect 16112 17376 16176 17380
rect 16192 17436 16256 17440
rect 16192 17380 16196 17436
rect 16196 17380 16252 17436
rect 16252 17380 16256 17436
rect 16192 17376 16256 17380
rect 25952 17436 26016 17440
rect 25952 17380 25956 17436
rect 25956 17380 26012 17436
rect 26012 17380 26016 17436
rect 25952 17376 26016 17380
rect 26032 17436 26096 17440
rect 26032 17380 26036 17436
rect 26036 17380 26092 17436
rect 26092 17380 26096 17436
rect 26032 17376 26096 17380
rect 26112 17436 26176 17440
rect 26112 17380 26116 17436
rect 26116 17380 26172 17436
rect 26172 17380 26176 17436
rect 26112 17376 26176 17380
rect 26192 17436 26256 17440
rect 26192 17380 26196 17436
rect 26196 17380 26252 17436
rect 26252 17380 26256 17436
rect 26192 17376 26256 17380
rect 10952 16892 11016 16896
rect 10952 16836 10956 16892
rect 10956 16836 11012 16892
rect 11012 16836 11016 16892
rect 10952 16832 11016 16836
rect 11032 16892 11096 16896
rect 11032 16836 11036 16892
rect 11036 16836 11092 16892
rect 11092 16836 11096 16892
rect 11032 16832 11096 16836
rect 11112 16892 11176 16896
rect 11112 16836 11116 16892
rect 11116 16836 11172 16892
rect 11172 16836 11176 16892
rect 11112 16832 11176 16836
rect 11192 16892 11256 16896
rect 11192 16836 11196 16892
rect 11196 16836 11252 16892
rect 11252 16836 11256 16892
rect 11192 16832 11256 16836
rect 20952 16892 21016 16896
rect 20952 16836 20956 16892
rect 20956 16836 21012 16892
rect 21012 16836 21016 16892
rect 20952 16832 21016 16836
rect 21032 16892 21096 16896
rect 21032 16836 21036 16892
rect 21036 16836 21092 16892
rect 21092 16836 21096 16892
rect 21032 16832 21096 16836
rect 21112 16892 21176 16896
rect 21112 16836 21116 16892
rect 21116 16836 21172 16892
rect 21172 16836 21176 16892
rect 21112 16832 21176 16836
rect 21192 16892 21256 16896
rect 21192 16836 21196 16892
rect 21196 16836 21252 16892
rect 21252 16836 21256 16892
rect 21192 16832 21256 16836
rect 5952 16348 6016 16352
rect 5952 16292 5956 16348
rect 5956 16292 6012 16348
rect 6012 16292 6016 16348
rect 5952 16288 6016 16292
rect 6032 16348 6096 16352
rect 6032 16292 6036 16348
rect 6036 16292 6092 16348
rect 6092 16292 6096 16348
rect 6032 16288 6096 16292
rect 6112 16348 6176 16352
rect 6112 16292 6116 16348
rect 6116 16292 6172 16348
rect 6172 16292 6176 16348
rect 6112 16288 6176 16292
rect 6192 16348 6256 16352
rect 6192 16292 6196 16348
rect 6196 16292 6252 16348
rect 6252 16292 6256 16348
rect 6192 16288 6256 16292
rect 15952 16348 16016 16352
rect 15952 16292 15956 16348
rect 15956 16292 16012 16348
rect 16012 16292 16016 16348
rect 15952 16288 16016 16292
rect 16032 16348 16096 16352
rect 16032 16292 16036 16348
rect 16036 16292 16092 16348
rect 16092 16292 16096 16348
rect 16032 16288 16096 16292
rect 16112 16348 16176 16352
rect 16112 16292 16116 16348
rect 16116 16292 16172 16348
rect 16172 16292 16176 16348
rect 16112 16288 16176 16292
rect 16192 16348 16256 16352
rect 16192 16292 16196 16348
rect 16196 16292 16252 16348
rect 16252 16292 16256 16348
rect 16192 16288 16256 16292
rect 25952 16348 26016 16352
rect 25952 16292 25956 16348
rect 25956 16292 26012 16348
rect 26012 16292 26016 16348
rect 25952 16288 26016 16292
rect 26032 16348 26096 16352
rect 26032 16292 26036 16348
rect 26036 16292 26092 16348
rect 26092 16292 26096 16348
rect 26032 16288 26096 16292
rect 26112 16348 26176 16352
rect 26112 16292 26116 16348
rect 26116 16292 26172 16348
rect 26172 16292 26176 16348
rect 26112 16288 26176 16292
rect 26192 16348 26256 16352
rect 26192 16292 26196 16348
rect 26196 16292 26252 16348
rect 26252 16292 26256 16348
rect 26192 16288 26256 16292
rect 10952 15804 11016 15808
rect 10952 15748 10956 15804
rect 10956 15748 11012 15804
rect 11012 15748 11016 15804
rect 10952 15744 11016 15748
rect 11032 15804 11096 15808
rect 11032 15748 11036 15804
rect 11036 15748 11092 15804
rect 11092 15748 11096 15804
rect 11032 15744 11096 15748
rect 11112 15804 11176 15808
rect 11112 15748 11116 15804
rect 11116 15748 11172 15804
rect 11172 15748 11176 15804
rect 11112 15744 11176 15748
rect 11192 15804 11256 15808
rect 11192 15748 11196 15804
rect 11196 15748 11252 15804
rect 11252 15748 11256 15804
rect 11192 15744 11256 15748
rect 20952 15804 21016 15808
rect 20952 15748 20956 15804
rect 20956 15748 21012 15804
rect 21012 15748 21016 15804
rect 20952 15744 21016 15748
rect 21032 15804 21096 15808
rect 21032 15748 21036 15804
rect 21036 15748 21092 15804
rect 21092 15748 21096 15804
rect 21032 15744 21096 15748
rect 21112 15804 21176 15808
rect 21112 15748 21116 15804
rect 21116 15748 21172 15804
rect 21172 15748 21176 15804
rect 21112 15744 21176 15748
rect 21192 15804 21256 15808
rect 21192 15748 21196 15804
rect 21196 15748 21252 15804
rect 21252 15748 21256 15804
rect 21192 15744 21256 15748
rect 5952 15260 6016 15264
rect 5952 15204 5956 15260
rect 5956 15204 6012 15260
rect 6012 15204 6016 15260
rect 5952 15200 6016 15204
rect 6032 15260 6096 15264
rect 6032 15204 6036 15260
rect 6036 15204 6092 15260
rect 6092 15204 6096 15260
rect 6032 15200 6096 15204
rect 6112 15260 6176 15264
rect 6112 15204 6116 15260
rect 6116 15204 6172 15260
rect 6172 15204 6176 15260
rect 6112 15200 6176 15204
rect 6192 15260 6256 15264
rect 6192 15204 6196 15260
rect 6196 15204 6252 15260
rect 6252 15204 6256 15260
rect 6192 15200 6256 15204
rect 15952 15260 16016 15264
rect 15952 15204 15956 15260
rect 15956 15204 16012 15260
rect 16012 15204 16016 15260
rect 15952 15200 16016 15204
rect 16032 15260 16096 15264
rect 16032 15204 16036 15260
rect 16036 15204 16092 15260
rect 16092 15204 16096 15260
rect 16032 15200 16096 15204
rect 16112 15260 16176 15264
rect 16112 15204 16116 15260
rect 16116 15204 16172 15260
rect 16172 15204 16176 15260
rect 16112 15200 16176 15204
rect 16192 15260 16256 15264
rect 16192 15204 16196 15260
rect 16196 15204 16252 15260
rect 16252 15204 16256 15260
rect 16192 15200 16256 15204
rect 25952 15260 26016 15264
rect 25952 15204 25956 15260
rect 25956 15204 26012 15260
rect 26012 15204 26016 15260
rect 25952 15200 26016 15204
rect 26032 15260 26096 15264
rect 26032 15204 26036 15260
rect 26036 15204 26092 15260
rect 26092 15204 26096 15260
rect 26032 15200 26096 15204
rect 26112 15260 26176 15264
rect 26112 15204 26116 15260
rect 26116 15204 26172 15260
rect 26172 15204 26176 15260
rect 26112 15200 26176 15204
rect 26192 15260 26256 15264
rect 26192 15204 26196 15260
rect 26196 15204 26252 15260
rect 26252 15204 26256 15260
rect 26192 15200 26256 15204
rect 10952 14716 11016 14720
rect 10952 14660 10956 14716
rect 10956 14660 11012 14716
rect 11012 14660 11016 14716
rect 10952 14656 11016 14660
rect 11032 14716 11096 14720
rect 11032 14660 11036 14716
rect 11036 14660 11092 14716
rect 11092 14660 11096 14716
rect 11032 14656 11096 14660
rect 11112 14716 11176 14720
rect 11112 14660 11116 14716
rect 11116 14660 11172 14716
rect 11172 14660 11176 14716
rect 11112 14656 11176 14660
rect 11192 14716 11256 14720
rect 11192 14660 11196 14716
rect 11196 14660 11252 14716
rect 11252 14660 11256 14716
rect 11192 14656 11256 14660
rect 20952 14716 21016 14720
rect 20952 14660 20956 14716
rect 20956 14660 21012 14716
rect 21012 14660 21016 14716
rect 20952 14656 21016 14660
rect 21032 14716 21096 14720
rect 21032 14660 21036 14716
rect 21036 14660 21092 14716
rect 21092 14660 21096 14716
rect 21032 14656 21096 14660
rect 21112 14716 21176 14720
rect 21112 14660 21116 14716
rect 21116 14660 21172 14716
rect 21172 14660 21176 14716
rect 21112 14656 21176 14660
rect 21192 14716 21256 14720
rect 21192 14660 21196 14716
rect 21196 14660 21252 14716
rect 21252 14660 21256 14716
rect 21192 14656 21256 14660
rect 5952 14172 6016 14176
rect 5952 14116 5956 14172
rect 5956 14116 6012 14172
rect 6012 14116 6016 14172
rect 5952 14112 6016 14116
rect 6032 14172 6096 14176
rect 6032 14116 6036 14172
rect 6036 14116 6092 14172
rect 6092 14116 6096 14172
rect 6032 14112 6096 14116
rect 6112 14172 6176 14176
rect 6112 14116 6116 14172
rect 6116 14116 6172 14172
rect 6172 14116 6176 14172
rect 6112 14112 6176 14116
rect 6192 14172 6256 14176
rect 6192 14116 6196 14172
rect 6196 14116 6252 14172
rect 6252 14116 6256 14172
rect 6192 14112 6256 14116
rect 15952 14172 16016 14176
rect 15952 14116 15956 14172
rect 15956 14116 16012 14172
rect 16012 14116 16016 14172
rect 15952 14112 16016 14116
rect 16032 14172 16096 14176
rect 16032 14116 16036 14172
rect 16036 14116 16092 14172
rect 16092 14116 16096 14172
rect 16032 14112 16096 14116
rect 16112 14172 16176 14176
rect 16112 14116 16116 14172
rect 16116 14116 16172 14172
rect 16172 14116 16176 14172
rect 16112 14112 16176 14116
rect 16192 14172 16256 14176
rect 16192 14116 16196 14172
rect 16196 14116 16252 14172
rect 16252 14116 16256 14172
rect 16192 14112 16256 14116
rect 25952 14172 26016 14176
rect 25952 14116 25956 14172
rect 25956 14116 26012 14172
rect 26012 14116 26016 14172
rect 25952 14112 26016 14116
rect 26032 14172 26096 14176
rect 26032 14116 26036 14172
rect 26036 14116 26092 14172
rect 26092 14116 26096 14172
rect 26032 14112 26096 14116
rect 26112 14172 26176 14176
rect 26112 14116 26116 14172
rect 26116 14116 26172 14172
rect 26172 14116 26176 14172
rect 26112 14112 26176 14116
rect 26192 14172 26256 14176
rect 26192 14116 26196 14172
rect 26196 14116 26252 14172
rect 26252 14116 26256 14172
rect 26192 14112 26256 14116
rect 10952 13628 11016 13632
rect 10952 13572 10956 13628
rect 10956 13572 11012 13628
rect 11012 13572 11016 13628
rect 10952 13568 11016 13572
rect 11032 13628 11096 13632
rect 11032 13572 11036 13628
rect 11036 13572 11092 13628
rect 11092 13572 11096 13628
rect 11032 13568 11096 13572
rect 11112 13628 11176 13632
rect 11112 13572 11116 13628
rect 11116 13572 11172 13628
rect 11172 13572 11176 13628
rect 11112 13568 11176 13572
rect 11192 13628 11256 13632
rect 11192 13572 11196 13628
rect 11196 13572 11252 13628
rect 11252 13572 11256 13628
rect 11192 13568 11256 13572
rect 20952 13628 21016 13632
rect 20952 13572 20956 13628
rect 20956 13572 21012 13628
rect 21012 13572 21016 13628
rect 20952 13568 21016 13572
rect 21032 13628 21096 13632
rect 21032 13572 21036 13628
rect 21036 13572 21092 13628
rect 21092 13572 21096 13628
rect 21032 13568 21096 13572
rect 21112 13628 21176 13632
rect 21112 13572 21116 13628
rect 21116 13572 21172 13628
rect 21172 13572 21176 13628
rect 21112 13568 21176 13572
rect 21192 13628 21256 13632
rect 21192 13572 21196 13628
rect 21196 13572 21252 13628
rect 21252 13572 21256 13628
rect 21192 13568 21256 13572
rect 9628 13228 9692 13292
rect 5952 13084 6016 13088
rect 5952 13028 5956 13084
rect 5956 13028 6012 13084
rect 6012 13028 6016 13084
rect 5952 13024 6016 13028
rect 6032 13084 6096 13088
rect 6032 13028 6036 13084
rect 6036 13028 6092 13084
rect 6092 13028 6096 13084
rect 6032 13024 6096 13028
rect 6112 13084 6176 13088
rect 6112 13028 6116 13084
rect 6116 13028 6172 13084
rect 6172 13028 6176 13084
rect 6112 13024 6176 13028
rect 6192 13084 6256 13088
rect 6192 13028 6196 13084
rect 6196 13028 6252 13084
rect 6252 13028 6256 13084
rect 6192 13024 6256 13028
rect 15952 13084 16016 13088
rect 15952 13028 15956 13084
rect 15956 13028 16012 13084
rect 16012 13028 16016 13084
rect 15952 13024 16016 13028
rect 16032 13084 16096 13088
rect 16032 13028 16036 13084
rect 16036 13028 16092 13084
rect 16092 13028 16096 13084
rect 16032 13024 16096 13028
rect 16112 13084 16176 13088
rect 16112 13028 16116 13084
rect 16116 13028 16172 13084
rect 16172 13028 16176 13084
rect 16112 13024 16176 13028
rect 16192 13084 16256 13088
rect 16192 13028 16196 13084
rect 16196 13028 16252 13084
rect 16252 13028 16256 13084
rect 16192 13024 16256 13028
rect 25952 13084 26016 13088
rect 25952 13028 25956 13084
rect 25956 13028 26012 13084
rect 26012 13028 26016 13084
rect 25952 13024 26016 13028
rect 26032 13084 26096 13088
rect 26032 13028 26036 13084
rect 26036 13028 26092 13084
rect 26092 13028 26096 13084
rect 26032 13024 26096 13028
rect 26112 13084 26176 13088
rect 26112 13028 26116 13084
rect 26116 13028 26172 13084
rect 26172 13028 26176 13084
rect 26112 13024 26176 13028
rect 26192 13084 26256 13088
rect 26192 13028 26196 13084
rect 26196 13028 26252 13084
rect 26252 13028 26256 13084
rect 26192 13024 26256 13028
rect 9628 12880 9692 12884
rect 9628 12824 9642 12880
rect 9642 12824 9692 12880
rect 9628 12820 9692 12824
rect 10952 12540 11016 12544
rect 10952 12484 10956 12540
rect 10956 12484 11012 12540
rect 11012 12484 11016 12540
rect 10952 12480 11016 12484
rect 11032 12540 11096 12544
rect 11032 12484 11036 12540
rect 11036 12484 11092 12540
rect 11092 12484 11096 12540
rect 11032 12480 11096 12484
rect 11112 12540 11176 12544
rect 11112 12484 11116 12540
rect 11116 12484 11172 12540
rect 11172 12484 11176 12540
rect 11112 12480 11176 12484
rect 11192 12540 11256 12544
rect 11192 12484 11196 12540
rect 11196 12484 11252 12540
rect 11252 12484 11256 12540
rect 11192 12480 11256 12484
rect 20952 12540 21016 12544
rect 20952 12484 20956 12540
rect 20956 12484 21012 12540
rect 21012 12484 21016 12540
rect 20952 12480 21016 12484
rect 21032 12540 21096 12544
rect 21032 12484 21036 12540
rect 21036 12484 21092 12540
rect 21092 12484 21096 12540
rect 21032 12480 21096 12484
rect 21112 12540 21176 12544
rect 21112 12484 21116 12540
rect 21116 12484 21172 12540
rect 21172 12484 21176 12540
rect 21112 12480 21176 12484
rect 21192 12540 21256 12544
rect 21192 12484 21196 12540
rect 21196 12484 21252 12540
rect 21252 12484 21256 12540
rect 21192 12480 21256 12484
rect 25452 12472 25516 12476
rect 25452 12416 25502 12472
rect 25502 12416 25516 12472
rect 25452 12412 25516 12416
rect 5952 11996 6016 12000
rect 5952 11940 5956 11996
rect 5956 11940 6012 11996
rect 6012 11940 6016 11996
rect 5952 11936 6016 11940
rect 6032 11996 6096 12000
rect 6032 11940 6036 11996
rect 6036 11940 6092 11996
rect 6092 11940 6096 11996
rect 6032 11936 6096 11940
rect 6112 11996 6176 12000
rect 6112 11940 6116 11996
rect 6116 11940 6172 11996
rect 6172 11940 6176 11996
rect 6112 11936 6176 11940
rect 6192 11996 6256 12000
rect 6192 11940 6196 11996
rect 6196 11940 6252 11996
rect 6252 11940 6256 11996
rect 6192 11936 6256 11940
rect 15952 11996 16016 12000
rect 15952 11940 15956 11996
rect 15956 11940 16012 11996
rect 16012 11940 16016 11996
rect 15952 11936 16016 11940
rect 16032 11996 16096 12000
rect 16032 11940 16036 11996
rect 16036 11940 16092 11996
rect 16092 11940 16096 11996
rect 16032 11936 16096 11940
rect 16112 11996 16176 12000
rect 16112 11940 16116 11996
rect 16116 11940 16172 11996
rect 16172 11940 16176 11996
rect 16112 11936 16176 11940
rect 16192 11996 16256 12000
rect 16192 11940 16196 11996
rect 16196 11940 16252 11996
rect 16252 11940 16256 11996
rect 16192 11936 16256 11940
rect 25952 11996 26016 12000
rect 25952 11940 25956 11996
rect 25956 11940 26012 11996
rect 26012 11940 26016 11996
rect 25952 11936 26016 11940
rect 26032 11996 26096 12000
rect 26032 11940 26036 11996
rect 26036 11940 26092 11996
rect 26092 11940 26096 11996
rect 26032 11936 26096 11940
rect 26112 11996 26176 12000
rect 26112 11940 26116 11996
rect 26116 11940 26172 11996
rect 26172 11940 26176 11996
rect 26112 11936 26176 11940
rect 26192 11996 26256 12000
rect 26192 11940 26196 11996
rect 26196 11940 26252 11996
rect 26252 11940 26256 11996
rect 26192 11936 26256 11940
rect 10952 11452 11016 11456
rect 10952 11396 10956 11452
rect 10956 11396 11012 11452
rect 11012 11396 11016 11452
rect 10952 11392 11016 11396
rect 11032 11452 11096 11456
rect 11032 11396 11036 11452
rect 11036 11396 11092 11452
rect 11092 11396 11096 11452
rect 11032 11392 11096 11396
rect 11112 11452 11176 11456
rect 11112 11396 11116 11452
rect 11116 11396 11172 11452
rect 11172 11396 11176 11452
rect 11112 11392 11176 11396
rect 11192 11452 11256 11456
rect 11192 11396 11196 11452
rect 11196 11396 11252 11452
rect 11252 11396 11256 11452
rect 11192 11392 11256 11396
rect 20952 11452 21016 11456
rect 20952 11396 20956 11452
rect 20956 11396 21012 11452
rect 21012 11396 21016 11452
rect 20952 11392 21016 11396
rect 21032 11452 21096 11456
rect 21032 11396 21036 11452
rect 21036 11396 21092 11452
rect 21092 11396 21096 11452
rect 21032 11392 21096 11396
rect 21112 11452 21176 11456
rect 21112 11396 21116 11452
rect 21116 11396 21172 11452
rect 21172 11396 21176 11452
rect 21112 11392 21176 11396
rect 21192 11452 21256 11456
rect 21192 11396 21196 11452
rect 21196 11396 21252 11452
rect 21252 11396 21256 11452
rect 21192 11392 21256 11396
rect 5952 10908 6016 10912
rect 5952 10852 5956 10908
rect 5956 10852 6012 10908
rect 6012 10852 6016 10908
rect 5952 10848 6016 10852
rect 6032 10908 6096 10912
rect 6032 10852 6036 10908
rect 6036 10852 6092 10908
rect 6092 10852 6096 10908
rect 6032 10848 6096 10852
rect 6112 10908 6176 10912
rect 6112 10852 6116 10908
rect 6116 10852 6172 10908
rect 6172 10852 6176 10908
rect 6112 10848 6176 10852
rect 6192 10908 6256 10912
rect 6192 10852 6196 10908
rect 6196 10852 6252 10908
rect 6252 10852 6256 10908
rect 6192 10848 6256 10852
rect 15952 10908 16016 10912
rect 15952 10852 15956 10908
rect 15956 10852 16012 10908
rect 16012 10852 16016 10908
rect 15952 10848 16016 10852
rect 16032 10908 16096 10912
rect 16032 10852 16036 10908
rect 16036 10852 16092 10908
rect 16092 10852 16096 10908
rect 16032 10848 16096 10852
rect 16112 10908 16176 10912
rect 16112 10852 16116 10908
rect 16116 10852 16172 10908
rect 16172 10852 16176 10908
rect 16112 10848 16176 10852
rect 16192 10908 16256 10912
rect 16192 10852 16196 10908
rect 16196 10852 16252 10908
rect 16252 10852 16256 10908
rect 16192 10848 16256 10852
rect 25952 10908 26016 10912
rect 25952 10852 25956 10908
rect 25956 10852 26012 10908
rect 26012 10852 26016 10908
rect 25952 10848 26016 10852
rect 26032 10908 26096 10912
rect 26032 10852 26036 10908
rect 26036 10852 26092 10908
rect 26092 10852 26096 10908
rect 26032 10848 26096 10852
rect 26112 10908 26176 10912
rect 26112 10852 26116 10908
rect 26116 10852 26172 10908
rect 26172 10852 26176 10908
rect 26112 10848 26176 10852
rect 26192 10908 26256 10912
rect 26192 10852 26196 10908
rect 26196 10852 26252 10908
rect 26252 10852 26256 10908
rect 26192 10848 26256 10852
rect 10952 10364 11016 10368
rect 10952 10308 10956 10364
rect 10956 10308 11012 10364
rect 11012 10308 11016 10364
rect 10952 10304 11016 10308
rect 11032 10364 11096 10368
rect 11032 10308 11036 10364
rect 11036 10308 11092 10364
rect 11092 10308 11096 10364
rect 11032 10304 11096 10308
rect 11112 10364 11176 10368
rect 11112 10308 11116 10364
rect 11116 10308 11172 10364
rect 11172 10308 11176 10364
rect 11112 10304 11176 10308
rect 11192 10364 11256 10368
rect 11192 10308 11196 10364
rect 11196 10308 11252 10364
rect 11252 10308 11256 10364
rect 11192 10304 11256 10308
rect 20952 10364 21016 10368
rect 20952 10308 20956 10364
rect 20956 10308 21012 10364
rect 21012 10308 21016 10364
rect 20952 10304 21016 10308
rect 21032 10364 21096 10368
rect 21032 10308 21036 10364
rect 21036 10308 21092 10364
rect 21092 10308 21096 10364
rect 21032 10304 21096 10308
rect 21112 10364 21176 10368
rect 21112 10308 21116 10364
rect 21116 10308 21172 10364
rect 21172 10308 21176 10364
rect 21112 10304 21176 10308
rect 21192 10364 21256 10368
rect 21192 10308 21196 10364
rect 21196 10308 21252 10364
rect 21252 10308 21256 10364
rect 21192 10304 21256 10308
rect 5952 9820 6016 9824
rect 5952 9764 5956 9820
rect 5956 9764 6012 9820
rect 6012 9764 6016 9820
rect 5952 9760 6016 9764
rect 6032 9820 6096 9824
rect 6032 9764 6036 9820
rect 6036 9764 6092 9820
rect 6092 9764 6096 9820
rect 6032 9760 6096 9764
rect 6112 9820 6176 9824
rect 6112 9764 6116 9820
rect 6116 9764 6172 9820
rect 6172 9764 6176 9820
rect 6112 9760 6176 9764
rect 6192 9820 6256 9824
rect 6192 9764 6196 9820
rect 6196 9764 6252 9820
rect 6252 9764 6256 9820
rect 6192 9760 6256 9764
rect 15952 9820 16016 9824
rect 15952 9764 15956 9820
rect 15956 9764 16012 9820
rect 16012 9764 16016 9820
rect 15952 9760 16016 9764
rect 16032 9820 16096 9824
rect 16032 9764 16036 9820
rect 16036 9764 16092 9820
rect 16092 9764 16096 9820
rect 16032 9760 16096 9764
rect 16112 9820 16176 9824
rect 16112 9764 16116 9820
rect 16116 9764 16172 9820
rect 16172 9764 16176 9820
rect 16112 9760 16176 9764
rect 16192 9820 16256 9824
rect 16192 9764 16196 9820
rect 16196 9764 16252 9820
rect 16252 9764 16256 9820
rect 16192 9760 16256 9764
rect 25952 9820 26016 9824
rect 25952 9764 25956 9820
rect 25956 9764 26012 9820
rect 26012 9764 26016 9820
rect 25952 9760 26016 9764
rect 26032 9820 26096 9824
rect 26032 9764 26036 9820
rect 26036 9764 26092 9820
rect 26092 9764 26096 9820
rect 26032 9760 26096 9764
rect 26112 9820 26176 9824
rect 26112 9764 26116 9820
rect 26116 9764 26172 9820
rect 26172 9764 26176 9820
rect 26112 9760 26176 9764
rect 26192 9820 26256 9824
rect 26192 9764 26196 9820
rect 26196 9764 26252 9820
rect 26252 9764 26256 9820
rect 26192 9760 26256 9764
rect 10952 9276 11016 9280
rect 10952 9220 10956 9276
rect 10956 9220 11012 9276
rect 11012 9220 11016 9276
rect 10952 9216 11016 9220
rect 11032 9276 11096 9280
rect 11032 9220 11036 9276
rect 11036 9220 11092 9276
rect 11092 9220 11096 9276
rect 11032 9216 11096 9220
rect 11112 9276 11176 9280
rect 11112 9220 11116 9276
rect 11116 9220 11172 9276
rect 11172 9220 11176 9276
rect 11112 9216 11176 9220
rect 11192 9276 11256 9280
rect 11192 9220 11196 9276
rect 11196 9220 11252 9276
rect 11252 9220 11256 9276
rect 11192 9216 11256 9220
rect 20952 9276 21016 9280
rect 20952 9220 20956 9276
rect 20956 9220 21012 9276
rect 21012 9220 21016 9276
rect 20952 9216 21016 9220
rect 21032 9276 21096 9280
rect 21032 9220 21036 9276
rect 21036 9220 21092 9276
rect 21092 9220 21096 9276
rect 21032 9216 21096 9220
rect 21112 9276 21176 9280
rect 21112 9220 21116 9276
rect 21116 9220 21172 9276
rect 21172 9220 21176 9276
rect 21112 9216 21176 9220
rect 21192 9276 21256 9280
rect 21192 9220 21196 9276
rect 21196 9220 21252 9276
rect 21252 9220 21256 9276
rect 21192 9216 21256 9220
rect 5952 8732 6016 8736
rect 5952 8676 5956 8732
rect 5956 8676 6012 8732
rect 6012 8676 6016 8732
rect 5952 8672 6016 8676
rect 6032 8732 6096 8736
rect 6032 8676 6036 8732
rect 6036 8676 6092 8732
rect 6092 8676 6096 8732
rect 6032 8672 6096 8676
rect 6112 8732 6176 8736
rect 6112 8676 6116 8732
rect 6116 8676 6172 8732
rect 6172 8676 6176 8732
rect 6112 8672 6176 8676
rect 6192 8732 6256 8736
rect 6192 8676 6196 8732
rect 6196 8676 6252 8732
rect 6252 8676 6256 8732
rect 6192 8672 6256 8676
rect 15952 8732 16016 8736
rect 15952 8676 15956 8732
rect 15956 8676 16012 8732
rect 16012 8676 16016 8732
rect 15952 8672 16016 8676
rect 16032 8732 16096 8736
rect 16032 8676 16036 8732
rect 16036 8676 16092 8732
rect 16092 8676 16096 8732
rect 16032 8672 16096 8676
rect 16112 8732 16176 8736
rect 16112 8676 16116 8732
rect 16116 8676 16172 8732
rect 16172 8676 16176 8732
rect 16112 8672 16176 8676
rect 16192 8732 16256 8736
rect 16192 8676 16196 8732
rect 16196 8676 16252 8732
rect 16252 8676 16256 8732
rect 16192 8672 16256 8676
rect 25952 8732 26016 8736
rect 25952 8676 25956 8732
rect 25956 8676 26012 8732
rect 26012 8676 26016 8732
rect 25952 8672 26016 8676
rect 26032 8732 26096 8736
rect 26032 8676 26036 8732
rect 26036 8676 26092 8732
rect 26092 8676 26096 8732
rect 26032 8672 26096 8676
rect 26112 8732 26176 8736
rect 26112 8676 26116 8732
rect 26116 8676 26172 8732
rect 26172 8676 26176 8732
rect 26112 8672 26176 8676
rect 26192 8732 26256 8736
rect 26192 8676 26196 8732
rect 26196 8676 26252 8732
rect 26252 8676 26256 8732
rect 26192 8672 26256 8676
rect 10952 8188 11016 8192
rect 10952 8132 10956 8188
rect 10956 8132 11012 8188
rect 11012 8132 11016 8188
rect 10952 8128 11016 8132
rect 11032 8188 11096 8192
rect 11032 8132 11036 8188
rect 11036 8132 11092 8188
rect 11092 8132 11096 8188
rect 11032 8128 11096 8132
rect 11112 8188 11176 8192
rect 11112 8132 11116 8188
rect 11116 8132 11172 8188
rect 11172 8132 11176 8188
rect 11112 8128 11176 8132
rect 11192 8188 11256 8192
rect 11192 8132 11196 8188
rect 11196 8132 11252 8188
rect 11252 8132 11256 8188
rect 11192 8128 11256 8132
rect 20952 8188 21016 8192
rect 20952 8132 20956 8188
rect 20956 8132 21012 8188
rect 21012 8132 21016 8188
rect 20952 8128 21016 8132
rect 21032 8188 21096 8192
rect 21032 8132 21036 8188
rect 21036 8132 21092 8188
rect 21092 8132 21096 8188
rect 21032 8128 21096 8132
rect 21112 8188 21176 8192
rect 21112 8132 21116 8188
rect 21116 8132 21172 8188
rect 21172 8132 21176 8188
rect 21112 8128 21176 8132
rect 21192 8188 21256 8192
rect 21192 8132 21196 8188
rect 21196 8132 21252 8188
rect 21252 8132 21256 8188
rect 21192 8128 21256 8132
rect 5952 7644 6016 7648
rect 5952 7588 5956 7644
rect 5956 7588 6012 7644
rect 6012 7588 6016 7644
rect 5952 7584 6016 7588
rect 6032 7644 6096 7648
rect 6032 7588 6036 7644
rect 6036 7588 6092 7644
rect 6092 7588 6096 7644
rect 6032 7584 6096 7588
rect 6112 7644 6176 7648
rect 6112 7588 6116 7644
rect 6116 7588 6172 7644
rect 6172 7588 6176 7644
rect 6112 7584 6176 7588
rect 6192 7644 6256 7648
rect 6192 7588 6196 7644
rect 6196 7588 6252 7644
rect 6252 7588 6256 7644
rect 6192 7584 6256 7588
rect 15952 7644 16016 7648
rect 15952 7588 15956 7644
rect 15956 7588 16012 7644
rect 16012 7588 16016 7644
rect 15952 7584 16016 7588
rect 16032 7644 16096 7648
rect 16032 7588 16036 7644
rect 16036 7588 16092 7644
rect 16092 7588 16096 7644
rect 16032 7584 16096 7588
rect 16112 7644 16176 7648
rect 16112 7588 16116 7644
rect 16116 7588 16172 7644
rect 16172 7588 16176 7644
rect 16112 7584 16176 7588
rect 16192 7644 16256 7648
rect 16192 7588 16196 7644
rect 16196 7588 16252 7644
rect 16252 7588 16256 7644
rect 16192 7584 16256 7588
rect 25952 7644 26016 7648
rect 25952 7588 25956 7644
rect 25956 7588 26012 7644
rect 26012 7588 26016 7644
rect 25952 7584 26016 7588
rect 26032 7644 26096 7648
rect 26032 7588 26036 7644
rect 26036 7588 26092 7644
rect 26092 7588 26096 7644
rect 26032 7584 26096 7588
rect 26112 7644 26176 7648
rect 26112 7588 26116 7644
rect 26116 7588 26172 7644
rect 26172 7588 26176 7644
rect 26112 7584 26176 7588
rect 26192 7644 26256 7648
rect 26192 7588 26196 7644
rect 26196 7588 26252 7644
rect 26252 7588 26256 7644
rect 26192 7584 26256 7588
rect 10952 7100 11016 7104
rect 10952 7044 10956 7100
rect 10956 7044 11012 7100
rect 11012 7044 11016 7100
rect 10952 7040 11016 7044
rect 11032 7100 11096 7104
rect 11032 7044 11036 7100
rect 11036 7044 11092 7100
rect 11092 7044 11096 7100
rect 11032 7040 11096 7044
rect 11112 7100 11176 7104
rect 11112 7044 11116 7100
rect 11116 7044 11172 7100
rect 11172 7044 11176 7100
rect 11112 7040 11176 7044
rect 11192 7100 11256 7104
rect 11192 7044 11196 7100
rect 11196 7044 11252 7100
rect 11252 7044 11256 7100
rect 11192 7040 11256 7044
rect 20952 7100 21016 7104
rect 20952 7044 20956 7100
rect 20956 7044 21012 7100
rect 21012 7044 21016 7100
rect 20952 7040 21016 7044
rect 21032 7100 21096 7104
rect 21032 7044 21036 7100
rect 21036 7044 21092 7100
rect 21092 7044 21096 7100
rect 21032 7040 21096 7044
rect 21112 7100 21176 7104
rect 21112 7044 21116 7100
rect 21116 7044 21172 7100
rect 21172 7044 21176 7100
rect 21112 7040 21176 7044
rect 21192 7100 21256 7104
rect 21192 7044 21196 7100
rect 21196 7044 21252 7100
rect 21252 7044 21256 7100
rect 21192 7040 21256 7044
rect 5952 6556 6016 6560
rect 5952 6500 5956 6556
rect 5956 6500 6012 6556
rect 6012 6500 6016 6556
rect 5952 6496 6016 6500
rect 6032 6556 6096 6560
rect 6032 6500 6036 6556
rect 6036 6500 6092 6556
rect 6092 6500 6096 6556
rect 6032 6496 6096 6500
rect 6112 6556 6176 6560
rect 6112 6500 6116 6556
rect 6116 6500 6172 6556
rect 6172 6500 6176 6556
rect 6112 6496 6176 6500
rect 6192 6556 6256 6560
rect 6192 6500 6196 6556
rect 6196 6500 6252 6556
rect 6252 6500 6256 6556
rect 6192 6496 6256 6500
rect 15952 6556 16016 6560
rect 15952 6500 15956 6556
rect 15956 6500 16012 6556
rect 16012 6500 16016 6556
rect 15952 6496 16016 6500
rect 16032 6556 16096 6560
rect 16032 6500 16036 6556
rect 16036 6500 16092 6556
rect 16092 6500 16096 6556
rect 16032 6496 16096 6500
rect 16112 6556 16176 6560
rect 16112 6500 16116 6556
rect 16116 6500 16172 6556
rect 16172 6500 16176 6556
rect 16112 6496 16176 6500
rect 16192 6556 16256 6560
rect 16192 6500 16196 6556
rect 16196 6500 16252 6556
rect 16252 6500 16256 6556
rect 16192 6496 16256 6500
rect 25952 6556 26016 6560
rect 25952 6500 25956 6556
rect 25956 6500 26012 6556
rect 26012 6500 26016 6556
rect 25952 6496 26016 6500
rect 26032 6556 26096 6560
rect 26032 6500 26036 6556
rect 26036 6500 26092 6556
rect 26092 6500 26096 6556
rect 26032 6496 26096 6500
rect 26112 6556 26176 6560
rect 26112 6500 26116 6556
rect 26116 6500 26172 6556
rect 26172 6500 26176 6556
rect 26112 6496 26176 6500
rect 26192 6556 26256 6560
rect 26192 6500 26196 6556
rect 26196 6500 26252 6556
rect 26252 6500 26256 6556
rect 26192 6496 26256 6500
rect 10952 6012 11016 6016
rect 10952 5956 10956 6012
rect 10956 5956 11012 6012
rect 11012 5956 11016 6012
rect 10952 5952 11016 5956
rect 11032 6012 11096 6016
rect 11032 5956 11036 6012
rect 11036 5956 11092 6012
rect 11092 5956 11096 6012
rect 11032 5952 11096 5956
rect 11112 6012 11176 6016
rect 11112 5956 11116 6012
rect 11116 5956 11172 6012
rect 11172 5956 11176 6012
rect 11112 5952 11176 5956
rect 11192 6012 11256 6016
rect 11192 5956 11196 6012
rect 11196 5956 11252 6012
rect 11252 5956 11256 6012
rect 11192 5952 11256 5956
rect 20952 6012 21016 6016
rect 20952 5956 20956 6012
rect 20956 5956 21012 6012
rect 21012 5956 21016 6012
rect 20952 5952 21016 5956
rect 21032 6012 21096 6016
rect 21032 5956 21036 6012
rect 21036 5956 21092 6012
rect 21092 5956 21096 6012
rect 21032 5952 21096 5956
rect 21112 6012 21176 6016
rect 21112 5956 21116 6012
rect 21116 5956 21172 6012
rect 21172 5956 21176 6012
rect 21112 5952 21176 5956
rect 21192 6012 21256 6016
rect 21192 5956 21196 6012
rect 21196 5956 21252 6012
rect 21252 5956 21256 6012
rect 21192 5952 21256 5956
rect 5952 5468 6016 5472
rect 5952 5412 5956 5468
rect 5956 5412 6012 5468
rect 6012 5412 6016 5468
rect 5952 5408 6016 5412
rect 6032 5468 6096 5472
rect 6032 5412 6036 5468
rect 6036 5412 6092 5468
rect 6092 5412 6096 5468
rect 6032 5408 6096 5412
rect 6112 5468 6176 5472
rect 6112 5412 6116 5468
rect 6116 5412 6172 5468
rect 6172 5412 6176 5468
rect 6112 5408 6176 5412
rect 6192 5468 6256 5472
rect 6192 5412 6196 5468
rect 6196 5412 6252 5468
rect 6252 5412 6256 5468
rect 6192 5408 6256 5412
rect 15952 5468 16016 5472
rect 15952 5412 15956 5468
rect 15956 5412 16012 5468
rect 16012 5412 16016 5468
rect 15952 5408 16016 5412
rect 16032 5468 16096 5472
rect 16032 5412 16036 5468
rect 16036 5412 16092 5468
rect 16092 5412 16096 5468
rect 16032 5408 16096 5412
rect 16112 5468 16176 5472
rect 16112 5412 16116 5468
rect 16116 5412 16172 5468
rect 16172 5412 16176 5468
rect 16112 5408 16176 5412
rect 16192 5468 16256 5472
rect 16192 5412 16196 5468
rect 16196 5412 16252 5468
rect 16252 5412 16256 5468
rect 16192 5408 16256 5412
rect 25952 5468 26016 5472
rect 25952 5412 25956 5468
rect 25956 5412 26012 5468
rect 26012 5412 26016 5468
rect 25952 5408 26016 5412
rect 26032 5468 26096 5472
rect 26032 5412 26036 5468
rect 26036 5412 26092 5468
rect 26092 5412 26096 5468
rect 26032 5408 26096 5412
rect 26112 5468 26176 5472
rect 26112 5412 26116 5468
rect 26116 5412 26172 5468
rect 26172 5412 26176 5468
rect 26112 5408 26176 5412
rect 26192 5468 26256 5472
rect 26192 5412 26196 5468
rect 26196 5412 26252 5468
rect 26252 5412 26256 5468
rect 26192 5408 26256 5412
rect 10952 4924 11016 4928
rect 10952 4868 10956 4924
rect 10956 4868 11012 4924
rect 11012 4868 11016 4924
rect 10952 4864 11016 4868
rect 11032 4924 11096 4928
rect 11032 4868 11036 4924
rect 11036 4868 11092 4924
rect 11092 4868 11096 4924
rect 11032 4864 11096 4868
rect 11112 4924 11176 4928
rect 11112 4868 11116 4924
rect 11116 4868 11172 4924
rect 11172 4868 11176 4924
rect 11112 4864 11176 4868
rect 11192 4924 11256 4928
rect 11192 4868 11196 4924
rect 11196 4868 11252 4924
rect 11252 4868 11256 4924
rect 11192 4864 11256 4868
rect 20952 4924 21016 4928
rect 20952 4868 20956 4924
rect 20956 4868 21012 4924
rect 21012 4868 21016 4924
rect 20952 4864 21016 4868
rect 21032 4924 21096 4928
rect 21032 4868 21036 4924
rect 21036 4868 21092 4924
rect 21092 4868 21096 4924
rect 21032 4864 21096 4868
rect 21112 4924 21176 4928
rect 21112 4868 21116 4924
rect 21116 4868 21172 4924
rect 21172 4868 21176 4924
rect 21112 4864 21176 4868
rect 21192 4924 21256 4928
rect 21192 4868 21196 4924
rect 21196 4868 21252 4924
rect 21252 4868 21256 4924
rect 21192 4864 21256 4868
rect 5952 4380 6016 4384
rect 5952 4324 5956 4380
rect 5956 4324 6012 4380
rect 6012 4324 6016 4380
rect 5952 4320 6016 4324
rect 6032 4380 6096 4384
rect 6032 4324 6036 4380
rect 6036 4324 6092 4380
rect 6092 4324 6096 4380
rect 6032 4320 6096 4324
rect 6112 4380 6176 4384
rect 6112 4324 6116 4380
rect 6116 4324 6172 4380
rect 6172 4324 6176 4380
rect 6112 4320 6176 4324
rect 6192 4380 6256 4384
rect 6192 4324 6196 4380
rect 6196 4324 6252 4380
rect 6252 4324 6256 4380
rect 6192 4320 6256 4324
rect 15952 4380 16016 4384
rect 15952 4324 15956 4380
rect 15956 4324 16012 4380
rect 16012 4324 16016 4380
rect 15952 4320 16016 4324
rect 16032 4380 16096 4384
rect 16032 4324 16036 4380
rect 16036 4324 16092 4380
rect 16092 4324 16096 4380
rect 16032 4320 16096 4324
rect 16112 4380 16176 4384
rect 16112 4324 16116 4380
rect 16116 4324 16172 4380
rect 16172 4324 16176 4380
rect 16112 4320 16176 4324
rect 16192 4380 16256 4384
rect 16192 4324 16196 4380
rect 16196 4324 16252 4380
rect 16252 4324 16256 4380
rect 16192 4320 16256 4324
rect 25952 4380 26016 4384
rect 25952 4324 25956 4380
rect 25956 4324 26012 4380
rect 26012 4324 26016 4380
rect 25952 4320 26016 4324
rect 26032 4380 26096 4384
rect 26032 4324 26036 4380
rect 26036 4324 26092 4380
rect 26092 4324 26096 4380
rect 26032 4320 26096 4324
rect 26112 4380 26176 4384
rect 26112 4324 26116 4380
rect 26116 4324 26172 4380
rect 26172 4324 26176 4380
rect 26112 4320 26176 4324
rect 26192 4380 26256 4384
rect 26192 4324 26196 4380
rect 26196 4324 26252 4380
rect 26252 4324 26256 4380
rect 26192 4320 26256 4324
rect 10952 3836 11016 3840
rect 10952 3780 10956 3836
rect 10956 3780 11012 3836
rect 11012 3780 11016 3836
rect 10952 3776 11016 3780
rect 11032 3836 11096 3840
rect 11032 3780 11036 3836
rect 11036 3780 11092 3836
rect 11092 3780 11096 3836
rect 11032 3776 11096 3780
rect 11112 3836 11176 3840
rect 11112 3780 11116 3836
rect 11116 3780 11172 3836
rect 11172 3780 11176 3836
rect 11112 3776 11176 3780
rect 11192 3836 11256 3840
rect 11192 3780 11196 3836
rect 11196 3780 11252 3836
rect 11252 3780 11256 3836
rect 11192 3776 11256 3780
rect 20952 3836 21016 3840
rect 20952 3780 20956 3836
rect 20956 3780 21012 3836
rect 21012 3780 21016 3836
rect 20952 3776 21016 3780
rect 21032 3836 21096 3840
rect 21032 3780 21036 3836
rect 21036 3780 21092 3836
rect 21092 3780 21096 3836
rect 21032 3776 21096 3780
rect 21112 3836 21176 3840
rect 21112 3780 21116 3836
rect 21116 3780 21172 3836
rect 21172 3780 21176 3836
rect 21112 3776 21176 3780
rect 21192 3836 21256 3840
rect 21192 3780 21196 3836
rect 21196 3780 21252 3836
rect 21252 3780 21256 3836
rect 21192 3776 21256 3780
rect 5952 3292 6016 3296
rect 5952 3236 5956 3292
rect 5956 3236 6012 3292
rect 6012 3236 6016 3292
rect 5952 3232 6016 3236
rect 6032 3292 6096 3296
rect 6032 3236 6036 3292
rect 6036 3236 6092 3292
rect 6092 3236 6096 3292
rect 6032 3232 6096 3236
rect 6112 3292 6176 3296
rect 6112 3236 6116 3292
rect 6116 3236 6172 3292
rect 6172 3236 6176 3292
rect 6112 3232 6176 3236
rect 6192 3292 6256 3296
rect 6192 3236 6196 3292
rect 6196 3236 6252 3292
rect 6252 3236 6256 3292
rect 6192 3232 6256 3236
rect 15952 3292 16016 3296
rect 15952 3236 15956 3292
rect 15956 3236 16012 3292
rect 16012 3236 16016 3292
rect 15952 3232 16016 3236
rect 16032 3292 16096 3296
rect 16032 3236 16036 3292
rect 16036 3236 16092 3292
rect 16092 3236 16096 3292
rect 16032 3232 16096 3236
rect 16112 3292 16176 3296
rect 16112 3236 16116 3292
rect 16116 3236 16172 3292
rect 16172 3236 16176 3292
rect 16112 3232 16176 3236
rect 16192 3292 16256 3296
rect 16192 3236 16196 3292
rect 16196 3236 16252 3292
rect 16252 3236 16256 3292
rect 16192 3232 16256 3236
rect 25952 3292 26016 3296
rect 25952 3236 25956 3292
rect 25956 3236 26012 3292
rect 26012 3236 26016 3292
rect 25952 3232 26016 3236
rect 26032 3292 26096 3296
rect 26032 3236 26036 3292
rect 26036 3236 26092 3292
rect 26092 3236 26096 3292
rect 26032 3232 26096 3236
rect 26112 3292 26176 3296
rect 26112 3236 26116 3292
rect 26116 3236 26172 3292
rect 26172 3236 26176 3292
rect 26112 3232 26176 3236
rect 26192 3292 26256 3296
rect 26192 3236 26196 3292
rect 26196 3236 26252 3292
rect 26252 3236 26256 3292
rect 26192 3232 26256 3236
rect 10952 2748 11016 2752
rect 10952 2692 10956 2748
rect 10956 2692 11012 2748
rect 11012 2692 11016 2748
rect 10952 2688 11016 2692
rect 11032 2748 11096 2752
rect 11032 2692 11036 2748
rect 11036 2692 11092 2748
rect 11092 2692 11096 2748
rect 11032 2688 11096 2692
rect 11112 2748 11176 2752
rect 11112 2692 11116 2748
rect 11116 2692 11172 2748
rect 11172 2692 11176 2748
rect 11112 2688 11176 2692
rect 11192 2748 11256 2752
rect 11192 2692 11196 2748
rect 11196 2692 11252 2748
rect 11252 2692 11256 2748
rect 11192 2688 11256 2692
rect 20952 2748 21016 2752
rect 20952 2692 20956 2748
rect 20956 2692 21012 2748
rect 21012 2692 21016 2748
rect 20952 2688 21016 2692
rect 21032 2748 21096 2752
rect 21032 2692 21036 2748
rect 21036 2692 21092 2748
rect 21092 2692 21096 2748
rect 21032 2688 21096 2692
rect 21112 2748 21176 2752
rect 21112 2692 21116 2748
rect 21116 2692 21172 2748
rect 21172 2692 21176 2748
rect 21112 2688 21176 2692
rect 21192 2748 21256 2752
rect 21192 2692 21196 2748
rect 21196 2692 21252 2748
rect 21252 2692 21256 2748
rect 21192 2688 21256 2692
rect 5952 2204 6016 2208
rect 5952 2148 5956 2204
rect 5956 2148 6012 2204
rect 6012 2148 6016 2204
rect 5952 2144 6016 2148
rect 6032 2204 6096 2208
rect 6032 2148 6036 2204
rect 6036 2148 6092 2204
rect 6092 2148 6096 2204
rect 6032 2144 6096 2148
rect 6112 2204 6176 2208
rect 6112 2148 6116 2204
rect 6116 2148 6172 2204
rect 6172 2148 6176 2204
rect 6112 2144 6176 2148
rect 6192 2204 6256 2208
rect 6192 2148 6196 2204
rect 6196 2148 6252 2204
rect 6252 2148 6256 2204
rect 6192 2144 6256 2148
rect 15952 2204 16016 2208
rect 15952 2148 15956 2204
rect 15956 2148 16012 2204
rect 16012 2148 16016 2204
rect 15952 2144 16016 2148
rect 16032 2204 16096 2208
rect 16032 2148 16036 2204
rect 16036 2148 16092 2204
rect 16092 2148 16096 2204
rect 16032 2144 16096 2148
rect 16112 2204 16176 2208
rect 16112 2148 16116 2204
rect 16116 2148 16172 2204
rect 16172 2148 16176 2204
rect 16112 2144 16176 2148
rect 16192 2204 16256 2208
rect 16192 2148 16196 2204
rect 16196 2148 16252 2204
rect 16252 2148 16256 2204
rect 16192 2144 16256 2148
rect 25952 2204 26016 2208
rect 25952 2148 25956 2204
rect 25956 2148 26012 2204
rect 26012 2148 26016 2204
rect 25952 2144 26016 2148
rect 26032 2204 26096 2208
rect 26032 2148 26036 2204
rect 26036 2148 26092 2204
rect 26092 2148 26096 2204
rect 26032 2144 26096 2148
rect 26112 2204 26176 2208
rect 26112 2148 26116 2204
rect 26116 2148 26172 2204
rect 26172 2148 26176 2204
rect 26112 2144 26176 2148
rect 26192 2204 26256 2208
rect 26192 2148 26196 2204
rect 26196 2148 26252 2204
rect 26252 2148 26256 2204
rect 26192 2144 26256 2148
<< metal4 >>
rect 5944 21792 6264 21808
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 20704 6264 21728
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 19616 6264 20640
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 18528 6264 19552
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 17440 6264 18464
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 16352 6264 17376
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 15264 6264 16288
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 14176 6264 15200
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 13088 6264 14112
rect 10944 21248 11264 21808
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 20160 11264 21184
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 19072 11264 20096
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 17984 11264 19008
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 16896 11264 17920
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 15808 11264 16832
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 14720 11264 15744
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 13632 11264 14656
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 9627 13292 9693 13293
rect 9627 13228 9628 13292
rect 9692 13228 9693 13292
rect 9627 13227 9693 13228
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 12000 6264 13024
rect 9630 12885 9690 13227
rect 9627 12884 9693 12885
rect 9627 12820 9628 12884
rect 9692 12820 9693 12884
rect 9627 12819 9693 12820
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 10912 6264 11936
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 9824 6264 10848
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 8736 6264 9760
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 7648 6264 8672
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 6560 6264 7584
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 5472 6264 6496
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 4384 6264 5408
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 3296 6264 4320
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 2208 6264 3232
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2128 6264 2144
rect 10944 12544 11264 13568
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 11456 11264 12480
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 10368 11264 11392
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 9280 11264 10304
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 8192 11264 9216
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 7104 11264 8128
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 6016 11264 7040
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 4928 11264 5952
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 3840 11264 4864
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 2752 11264 3776
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2128 11264 2688
rect 15944 21792 16264 21808
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 20704 16264 21728
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 19616 16264 20640
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 18528 16264 19552
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 17440 16264 18464
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 16352 16264 17376
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 15264 16264 16288
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 14176 16264 15200
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 13088 16264 14112
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 12000 16264 13024
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 10912 16264 11936
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 9824 16264 10848
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 8736 16264 9760
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 7648 16264 8672
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 6560 16264 7584
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 5472 16264 6496
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 4384 16264 5408
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 3296 16264 4320
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 2208 16264 3232
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2128 16264 2144
rect 20944 21248 21264 21808
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 20944 20160 21264 21184
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 19072 21264 20096
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 17984 21264 19008
rect 25944 21792 26264 21808
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 20704 26264 21728
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 19616 26264 20640
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 18528 26264 19552
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25451 18324 25517 18325
rect 25451 18260 25452 18324
rect 25516 18260 25517 18324
rect 25451 18259 25517 18260
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 16896 21264 17920
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 15808 21264 16832
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 20944 14720 21264 15744
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 13632 21264 14656
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 12544 21264 13568
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 11456 21264 12480
rect 25454 12477 25514 18259
rect 25944 17440 26264 18464
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 16352 26264 17376
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 15264 26264 16288
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 25944 14176 26264 15200
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 13088 26264 14112
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25451 12476 25517 12477
rect 25451 12412 25452 12476
rect 25516 12412 25517 12476
rect 25451 12411 25517 12412
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 10368 21264 11392
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 20944 9280 21264 10304
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 20944 8192 21264 9216
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 7104 21264 8128
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 6016 21264 7040
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 4928 21264 5952
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 3840 21264 4864
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 20944 2752 21264 3776
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2128 21264 2688
rect 25944 12000 26264 13024
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 10912 26264 11936
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 9824 26264 10848
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 25944 8736 26264 9760
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 7648 26264 8672
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 6560 26264 7584
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 5472 26264 6496
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 4384 26264 5408
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 25944 3296 26264 4320
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 25944 2208 26264 3232
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2128 26264 2144
use sky130_fd_sc_hd__decap_4  FILLER_0_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1564 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_13 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2300 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_9
timestamp 1604681595
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17
timestamp 1604681595
transform 1 0 2668 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1604681595
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 2116 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 2852 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_21 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26
timestamp 1604681595
transform 1 0 3496 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21
timestamp 1604681595
transform 1 0 3036 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3312 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3128 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3312 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_37
timestamp 1604681595
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_33
timestamp 1604681595
transform 1 0 4140 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 4692 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1604681595
transform 1 0 4324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 4324 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41
timestamp 1604681595
transform 1 0 4876 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4876 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_45
timestamp 1604681595
transform 1 0 5244 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48
timestamp 1604681595
transform 1 0 5520 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45
timestamp 1604681595
transform 1 0 5244 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 5336 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1604681595
transform 1 0 5428 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_53
timestamp 1604681595
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_49
timestamp 1604681595
transform 1 0 5612 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53
timestamp 1604681595
transform 1 0 5980 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 5796 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1604681595
transform 1 0 6164 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604681595
transform 1 0 5612 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1604681595
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1604681595
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1604681595
transform 1 0 6348 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_72
timestamp 1604681595
transform 1 0 7728 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_68
timestamp 1604681595
transform 1 0 7360 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69
timestamp 1604681595
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 7636 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7544 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_83
timestamp 1604681595
transform 1 0 8740 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73
timestamp 1604681595
transform 1 0 7820 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 7912 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8188 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_76 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8096 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10488 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100
timestamp 1604681595
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_104
timestamp 1604681595
transform 1 0 10672 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_88
timestamp 1604681595
transform 1 0 9200 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_100
timestamp 1604681595
transform 1 0 10304 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_1_112
timestamp 1604681595
transform 1 0 11408 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1604681595
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_123
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_134
timestamp 1604681595
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_127
timestamp 1604681595
transform 1 0 12788 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_131
timestamp 1604681595
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13340 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 12880 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_144
timestamp 1604681595
transform 1 0 14352 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_138
timestamp 1604681595
transform 1 0 13800 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14444 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_135
timestamp 1604681595
transform 1 0 13524 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15640 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15180 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_147
timestamp 1604681595
transform 1 0 14628 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_151
timestamp 1604681595
transform 1 0 14996 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_155
timestamp 1604681595
transform 1 0 15364 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_160
timestamp 1604681595
transform 1 0 15824 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1604681595
transform 1 0 16928 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_168
timestamp 1604681595
transform 1 0 16560 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16744 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16928 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_182
timestamp 1604681595
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_178
timestamp 1604681595
transform 1 0 17480 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1604681595
transform 1 0 17848 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_178
timestamp 1604681595
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17296 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 17664 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_187
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19136 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 18768 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 19872 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1604681595
transform 1 0 19044 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_202
timestamp 1604681595
transform 1 0 19688 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_206
timestamp 1604681595
transform 1 0 20056 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_190
timestamp 1604681595
transform 1 0 18584 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_194
timestamp 1604681595
transform 1 0 18952 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_206
timestamp 1604681595
transform 1 0 20056 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_217
timestamp 1604681595
transform 1 0 21068 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_214
timestamp 1604681595
transform 1 0 20792 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_214
timestamp 1604681595
transform 1 0 20792 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1604681595
transform 1 0 21436 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_224
timestamp 1604681595
transform 1 0 21712 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 21620 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 21252 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 21804 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_225
timestamp 1604681595
transform 1 0 21804 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_237
timestamp 1604681595
transform 1 0 22908 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_231
timestamp 1604681595
transform 1 0 22356 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 22540 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_249
timestamp 1604681595
transform 1 0 24012 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_243
timestamp 1604681595
transform 1 0 23460 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_247
timestamp 1604681595
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_235
timestamp 1604681595
transform 1 0 22724 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_253
timestamp 1604681595
transform 1 0 24380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_255
timestamp 1604681595
transform 1 0 24564 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24748 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1604681595
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1604681595
transform 1 0 24748 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_265
timestamp 1604681595
transform 1 0 25484 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_261
timestamp 1604681595
transform 1 0 25116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_259
timestamp 1604681595
transform 1 0 24932 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1604681595
transform 1 0 25300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 25668 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_279
timestamp 1604681595
transform 1 0 26772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_273
timestamp 1604681595
transform 1 0 26220 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_275
timestamp 1604681595
transform 1 0 26404 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_271
timestamp 1604681595
transform 1 0 26036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1604681595
transform 1 0 26220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1604681595
transform 1 0 26956 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604681595
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604681595
transform 1 0 26404 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1604681595
transform 1 0 26864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_291
timestamp 1604681595
transform 1 0 27876 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_283
timestamp 1604681595
transform 1 0 27140 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1604681595
transform 1 0 27324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 27508 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_284
timestamp 1604681595
transform 1 0 27232 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 28888 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 28888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1604681595
transform 1 0 28060 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_296
timestamp 1604681595
transform 1 0 28336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_295
timestamp 1604681595
transform 1 0 28244 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1604681595
transform 1 0 1932 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2760 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1604681595
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_7
timestamp 1604681595
transform 1 0 1748 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1604681595
transform 1 0 2300 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_17
timestamp 1604681595
transform 1 0 2668 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_20
timestamp 1604681595
transform 1 0 2944 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3312 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_26
timestamp 1604681595
transform 1 0 3496 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_30
timestamp 1604681595
transform 1 0 3864 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_36
timestamp 1604681595
transform 1 0 4416 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 5336 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_44
timestamp 1604681595
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_55
timestamp 1604681595
transform 1 0 6164 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6900 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_2_72
timestamp 1604681595
transform 1 0 7728 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9844 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_84
timestamp 1604681595
transform 1 0 8832 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_97
timestamp 1604681595
transform 1 0 10028 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 11316 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_109
timestamp 1604681595
transform 1 0 11132 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_113
timestamp 1604681595
transform 1 0 11500 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_125
timestamp 1604681595
transform 1 0 12604 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_137
timestamp 1604681595
transform 1 0 13708 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15640 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1604681595
transform 1 0 14812 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_164
timestamp 1604681595
transform 1 0 16192 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 17664 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_176
timestamp 1604681595
transform 1 0 17296 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 19228 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_189
timestamp 1604681595
transform 1 0 18492 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_199
timestamp 1604681595
transform 1 0 19412 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_203
timestamp 1604681595
transform 1 0 19780 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_207
timestamp 1604681595
transform 1 0 20148 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 22172 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_210
timestamp 1604681595
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_224
timestamp 1604681595
transform 1 0 21712 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_228
timestamp 1604681595
transform 1 0 22080 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_231
timestamp 1604681595
transform 1 0 22356 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_243
timestamp 1604681595
transform 1 0 23460 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_255
timestamp 1604681595
transform 1 0 24564 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_267
timestamp 1604681595
transform 1 0 25668 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_280
timestamp 1604681595
transform 1 0 26864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 28888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_292
timestamp 1604681595
transform 1 0 27968 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_298
timestamp 1604681595
transform 1 0 28520 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2760 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1604681595
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_7
timestamp 1604681595
transform 1 0 1748 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_11
timestamp 1604681595
transform 1 0 2116 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_14
timestamp 1604681595
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604681595
transform 1 0 4324 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1604681595
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1604681595
transform 1 0 4876 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1604681595
transform 1 0 3588 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_31
timestamp 1604681595
transform 1 0 3956 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_34
timestamp 1604681595
transform 1 0 4232 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_39
timestamp 1604681595
transform 1 0 4692 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5612 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_43
timestamp 1604681595
transform 1 0 5060 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_51
timestamp 1604681595
transform 1 0 5796 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_55
timestamp 1604681595
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_62
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 7636 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 7452 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 7084 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_67
timestamp 1604681595
transform 1 0 7268 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9844 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_87
timestamp 1604681595
transform 1 0 9108 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11500 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11868 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_111
timestamp 1604681595
transform 1 0 11316 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_115
timestamp 1604681595
transform 1 0 11684 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp 1604681595
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12880 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_127
timestamp 1604681595
transform 1 0 12788 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_130
timestamp 1604681595
transform 1 0 13064 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_134
timestamp 1604681595
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_138
timestamp 1604681595
transform 1 0 13800 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 16376 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_150
timestamp 1604681595
transform 1 0 14904 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_164
timestamp 1604681595
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_168
timestamp 1604681595
transform 1 0 16560 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_180
timestamp 1604681595
transform 1 0 17664 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20240 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20056 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 19688 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_200
timestamp 1604681595
transform 1 0 19504 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_204
timestamp 1604681595
transform 1 0 19872 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1604681595
transform 1 0 21804 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 21620 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_217
timestamp 1604681595
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1604681595
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_234
timestamp 1604681595
transform 1 0 22632 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_238
timestamp 1604681595
transform 1 0 23000 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1604681595
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_269
timestamp 1604681595
transform 1 0 25852 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 27508 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 26404 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1604681595
transform 1 0 26956 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604681595
transform 1 0 27324 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_279
timestamp 1604681595
transform 1 0 26772 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_283
timestamp 1604681595
transform 1 0 27140 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_291
timestamp 1604681595
transform 1 0 27876 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 28888 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 28060 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_295
timestamp 1604681595
transform 1 0 28244 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1604681595
transform 1 0 1932 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 2300 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_7
timestamp 1604681595
transform 1 0 1748 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_11
timestamp 1604681595
transform 1 0 2116 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_19
timestamp 1604681595
transform 1 0 2852 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3036 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_23
timestamp 1604681595
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604681595
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_36
timestamp 1604681595
transform 1 0 4416 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 5980 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_48
timestamp 1604681595
transform 1 0 5520 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_52
timestamp 1604681595
transform 1 0 5888 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_62
timestamp 1604681595
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_66
timestamp 1604681595
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_70
timestamp 1604681595
transform 1 0 7544 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_82
timestamp 1604681595
transform 1 0 8648 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10672 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1604681595
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_101
timestamp 1604681595
transform 1 0 10396 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11316 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 12328 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11040 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_106
timestamp 1604681595
transform 1 0 10856 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_110
timestamp 1604681595
transform 1 0 11224 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_120
timestamp 1604681595
transform 1 0 12144 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_124
timestamp 1604681595
transform 1 0 12512 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12880 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 12696 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_137
timestamp 1604681595
transform 1 0 13708 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 16008 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 15456 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1604681595
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_158
timestamp 1604681595
transform 1 0 15640 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_178
timestamp 1604681595
transform 1 0 17480 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_186
timestamp 1604681595
transform 1 0 18216 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_194
timestamp 1604681595
transform 1 0 18952 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_206
timestamp 1604681595
transform 1 0 20056 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 22172 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 21804 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 21068 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 20424 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1604681595
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_215
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_219
timestamp 1604681595
transform 1 0 21252 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_227
timestamp 1604681595
transform 1 0 21988 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_245
timestamp 1604681595
transform 1 0 23644 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_257
timestamp 1604681595
transform 1 0 24748 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_269
timestamp 1604681595
transform 1 0 25852 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_280
timestamp 1604681595
transform 1 0 26864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 28888 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_292
timestamp 1604681595
transform 1 0 27968 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_298
timestamp 1604681595
transform 1 0 28520 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 2944 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1604681595
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 2300 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_7
timestamp 1604681595
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_11
timestamp 1604681595
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_36
timestamp 1604681595
transform 1 0 4416 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 5152 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_42
timestamp 1604681595
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_46
timestamp 1604681595
transform 1 0 5336 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_54
timestamp 1604681595
transform 1 0 6072 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1604681595
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_71
timestamp 1604681595
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_75
timestamp 1604681595
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_79
timestamp 1604681595
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10672 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_91
timestamp 1604681595
transform 1 0 9476 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_95
timestamp 1604681595
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_99
timestamp 1604681595
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_103
timestamp 1604681595
transform 1 0 10580 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12604 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_113
timestamp 1604681595
transform 1 0 11500 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_117
timestamp 1604681595
transform 1 0 11868 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_141
timestamp 1604681595
transform 1 0 14076 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 14812 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 14628 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_165
timestamp 1604681595
transform 1 0 16284 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 16468 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1604681595
transform 1 0 16652 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp 1604681595
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_179
timestamp 1604681595
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 19872 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_196
timestamp 1604681595
transform 1 0 19136 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_206
timestamp 1604681595
transform 1 0 20056 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1604681595
transform 1 0 20424 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_219
timestamp 1604681595
transform 1 0 21252 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_223
timestamp 1604681595
transform 1 0 21620 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_235
timestamp 1604681595
transform 1 0 22724 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_241
timestamp 1604681595
transform 1 0 23276 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1604681595
transform 1 0 25116 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 26404 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604681595
transform 1 0 26956 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 26220 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_279
timestamp 1604681595
transform 1 0 26772 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_283
timestamp 1604681595
transform 1 0 27140 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 28888 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_295
timestamp 1604681595
transform 1 0 28244 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7
timestamp 1604681595
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1604681595
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_19
timestamp 1604681595
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_15
timestamp 1604681595
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_11
timestamp 1604681595
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 2668 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 1748 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 4784 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_23
timestamp 1604681595
transform 1 0 3220 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_23
timestamp 1604681595
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_35
timestamp 1604681595
transform 1 0 4324 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_48
timestamp 1604681595
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_43
timestamp 1604681595
transform 1 0 5060 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 5336 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_56
timestamp 1604681595
transform 1 0 6256 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_52
timestamp 1604681595
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_56
timestamp 1604681595
transform 1 0 6256 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 6992 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 8740 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 7820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_73
timestamp 1604681595
transform 1 0 7820 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_81
timestamp 1604681595
transform 1 0 8556 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_71
timestamp 1604681595
transform 1 0 7636 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_75
timestamp 1604681595
transform 1 0 8004 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_92
timestamp 1604681595
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1604681595
transform 1 0 9476 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85
timestamp 1604681595
transform 1 0 8924 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_96
timestamp 1604681595
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9752 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10304 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10396 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_7_109
timestamp 1604681595
transform 1 0 11132 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_114
timestamp 1604681595
transform 1 0 11592 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_110
timestamp 1604681595
transform 1 0 11224 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11408 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_118
timestamp 1604681595
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_115
timestamp 1604681595
transform 1 0 11684 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 11960 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 12604 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_135
timestamp 1604681595
transform 1 0 13524 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_127
timestamp 1604681595
transform 1 0 12788 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_131
timestamp 1604681595
transform 1 0 13156 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_127
timestamp 1604681595
transform 1 0 12788 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 13340 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12972 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 13340 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_139
timestamp 1604681595
transform 1 0 13892 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 14076 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 13708 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_143
timestamp 1604681595
transform 1 0 14260 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_135
timestamp 1604681595
transform 1 0 13524 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_155
timestamp 1604681595
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_154
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_147
timestamp 1604681595
transform 1 0 14628 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_159
timestamp 1604681595
transform 1 0 15732 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_165
timestamp 1604681595
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 15916 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1604681595
transform 1 0 15456 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16100 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_176
timestamp 1604681595
transform 1 0 17296 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_172
timestamp 1604681595
transform 1 0 16928 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_169
timestamp 1604681595
transform 1 0 16652 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 16836 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 16468 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 17020 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_187
timestamp 1604681595
transform 1 0 18308 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_180
timestamp 1604681595
transform 1 0 17664 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _20_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_182
timestamp 1604681595
transform 1 0 17848 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_195
timestamp 1604681595
transform 1 0 19044 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_191
timestamp 1604681595
transform 1 0 18676 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_194
timestamp 1604681595
transform 1 0 18952 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 18492 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_199
timestamp 1604681595
transform 1 0 19412 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_204
timestamp 1604681595
transform 1 0 19872 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 19688 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 19504 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 19688 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_7_218
timestamp 1604681595
transform 1 0 21160 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1604681595
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 20424 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_229
timestamp 1604681595
transform 1 0 22172 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1604681595
transform 1 0 21528 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 21712 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 21344 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1604681595
transform 1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_224
timestamp 1604681595
transform 1 0 21712 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_233
timestamp 1604681595
transform 1 0 22540 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_236
timestamp 1604681595
transform 1 0 22816 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 22356 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_249
timestamp 1604681595
transform 1 0 24012 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_245
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_241
timestamp 1604681595
transform 1 0 23276 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_244
timestamp 1604681595
transform 1 0 23552 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23644 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 23828 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_247
timestamp 1604681595
transform 1 0 23828 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 24196 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_259
timestamp 1604681595
transform 1 0 24932 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_253
timestamp 1604681595
transform 1 0 24380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_265
timestamp 1604681595
transform 1 0 25484 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 26404 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604681595
transform 1 0 26956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 26220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_271
timestamp 1604681595
transform 1 0 26036 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_280
timestamp 1604681595
transform 1 0 26864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_279
timestamp 1604681595
transform 1 0 26772 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_283
timestamp 1604681595
transform 1 0 27140 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 28888 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 28888 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_292
timestamp 1604681595
transform 1 0 27968 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_298
timestamp 1604681595
transform 1 0 28520 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_295
timestamp 1604681595
transform 1 0 28244 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 2300 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 1564 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_7
timestamp 1604681595
transform 1 0 1748 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 4232 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_22
timestamp 1604681595
transform 1 0 3128 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_26
timestamp 1604681595
transform 1 0 3496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1604681595
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_36
timestamp 1604681595
transform 1 0 4416 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 5336 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_55
timestamp 1604681595
transform 1 0 6164 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1604681595
transform 1 0 6900 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 8280 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_66
timestamp 1604681595
transform 1 0 7176 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_80
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 10304 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_85
timestamp 1604681595
transform 1 0 8924 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1604681595
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_93
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_99
timestamp 1604681595
transform 1 0 10212 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_102
timestamp 1604681595
transform 1 0 10488 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 11776 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_114
timestamp 1604681595
transform 1 0 11592 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_125
timestamp 1604681595
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 13340 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_129
timestamp 1604681595
transform 1 0 12972 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_142
timestamp 1604681595
transform 1 0 14168 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_146
timestamp 1604681595
transform 1 0 14536 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1604681595
transform 1 0 14812 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_162
timestamp 1604681595
transform 1 0 16008 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_165
timestamp 1604681595
transform 1 0 16284 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1604681595
transform 1 0 18032 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1604681595
transform 1 0 16468 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_176
timestamp 1604681595
transform 1 0 17296 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_193
timestamp 1604681595
transform 1 0 18860 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_205
timestamp 1604681595
transform 1 0 19964 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 21988 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1604681595
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_224
timestamp 1604681595
transform 1 0 21712 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_229
timestamp 1604681595
transform 1 0 22172 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1604681595
transform 1 0 23460 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 22356 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 22724 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_233
timestamp 1604681595
transform 1 0 22540 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_237
timestamp 1604681595
transform 1 0 22908 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24472 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 25300 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_252
timestamp 1604681595
transform 1 0 24288 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_256
timestamp 1604681595
transform 1 0 24656 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_262
timestamp 1604681595
transform 1 0 25208 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_265
timestamp 1604681595
transform 1 0 25484 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_273
timestamp 1604681595
transform 1 0 26220 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_280
timestamp 1604681595
transform 1 0 26864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 28888 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_292
timestamp 1604681595
transform 1 0 27968 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_298
timestamp 1604681595
transform 1 0 28520 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_19
timestamp 1604681595
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 3588 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_23
timestamp 1604681595
transform 1 0 3220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_36
timestamp 1604681595
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_40
timestamp 1604681595
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_53
timestamp 1604681595
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1604681595
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 8280 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_65
timestamp 1604681595
transform 1 0 7084 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_73
timestamp 1604681595
transform 1 0 7820 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_94
timestamp 1604681595
transform 1 0 9752 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_102
timestamp 1604681595
transform 1 0 10488 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_111
timestamp 1604681595
transform 1 0 11316 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_107
timestamp 1604681595
transform 1 0 10948 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 10764 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1604681595
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_115
timestamp 1604681595
transform 1 0 11684 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 14444 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_132
timestamp 1604681595
transform 1 0 13248 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_144
timestamp 1604681595
transform 1 0 14352 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 14628 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 1604681595
transform 1 0 16100 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_174
timestamp 1604681595
transform 1 0 17112 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_170
timestamp 1604681595
transform 1 0 16744 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1604681595
transform 1 0 16468 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16560 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17296 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_178
timestamp 1604681595
transform 1 0 17480 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1604681595
transform 1 0 18860 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1604681595
transform 1 0 19964 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 21068 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_219
timestamp 1604681595
transform 1 0 21252 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_223
timestamp 1604681595
transform 1 0 21620 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_236
timestamp 1604681595
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_240
timestamp 1604681595
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 25300 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_254
timestamp 1604681595
transform 1 0 24472 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_258
timestamp 1604681595
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_262
timestamp 1604681595
transform 1 0 25208 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 26956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_279
timestamp 1604681595
transform 1 0 26772 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_283
timestamp 1604681595
transform 1 0 27140 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 28888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_295
timestamp 1604681595
transform 1 0 28244 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 1564 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_3
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_7
timestamp 1604681595
transform 1 0 1748 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_11
timestamp 1604681595
transform 1 0 2116 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 4784 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_23
timestamp 1604681595
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1604681595
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 5152 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_42
timestamp 1604681595
transform 1 0 4968 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_60
timestamp 1604681595
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_64
timestamp 1604681595
transform 1 0 6992 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_76
timestamp 1604681595
transform 1 0 8096 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_84
timestamp 1604681595
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_88
timestamp 1604681595
transform 1 0 9200 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 11132 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_105
timestamp 1604681595
transform 1 0 10764 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_125
timestamp 1604681595
transform 1 0 12604 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604681595
transform 1 0 13340 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_136
timestamp 1604681595
transform 1 0 13616 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16376 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_148
timestamp 1604681595
transform 1 0 14720 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1604681595
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16928 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_168
timestamp 1604681595
transform 1 0 16560 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_181
timestamp 1604681595
transform 1 0 17756 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_186
timestamp 1604681595
transform 1 0 18216 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 18400 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 19964 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1604681595
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_202
timestamp 1604681595
transform 1 0 19688 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_207
timestamp 1604681595
transform 1 0 20148 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1604681595
transform 1 0 21988 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 21068 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 21436 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 20516 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1604681595
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_219
timestamp 1604681595
transform 1 0 21252 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_223
timestamp 1604681595
transform 1 0 21620 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1604681595
transform 1 0 23552 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 23368 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_236
timestamp 1604681595
transform 1 0 22816 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 25300 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_253
timestamp 1604681595
transform 1 0 24380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_261
timestamp 1604681595
transform 1 0 25116 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_265
timestamp 1604681595
transform 1 0 25484 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_273
timestamp 1604681595
transform 1 0 26220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_280
timestamp 1604681595
transform 1 0 26864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 28888 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_292
timestamp 1604681595
transform 1 0 27968 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_298
timestamp 1604681595
transform 1 0 28520 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1604681595
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_7
timestamp 1604681595
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_11
timestamp 1604681595
transform 1 0 2116 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_16
timestamp 1604681595
transform 1 0 2576 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 3128 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4784 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_31
timestamp 1604681595
transform 1 0 3956 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_35
timestamp 1604681595
transform 1 0 4324 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_49
timestamp 1604681595
transform 1 0 5612 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1604681595
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604681595
transform 1 0 6900 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 7360 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_66
timestamp 1604681595
transform 1 0 7176 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_70
timestamp 1604681595
transform 1 0 7544 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_78
timestamp 1604681595
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_82
timestamp 1604681595
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 9016 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 8832 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 10672 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_102
timestamp 1604681595
transform 1 0 10488 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_106
timestamp 1604681595
transform 1 0 10856 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_110
timestamp 1604681595
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1604681595
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_159
timestamp 1604681595
transform 1 0 15732 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_163
timestamp 1604681595
transform 1 0 16100 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_175
timestamp 1604681595
transform 1 0 17204 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_179
timestamp 1604681595
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 19964 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 19780 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 19320 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_196
timestamp 1604681595
transform 1 0 19136 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_200
timestamp 1604681595
transform 1 0 19504 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 21620 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1604681595
transform 1 0 21436 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_225
timestamp 1604681595
transform 1 0 21804 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 22448 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_231
timestamp 1604681595
transform 1 0 22356 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_234
timestamp 1604681595
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_238
timestamp 1604681595
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_242
timestamp 1604681595
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_245
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 24196 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 24564 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 24932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_253
timestamp 1604681595
transform 1 0 24380 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_257
timestamp 1604681595
transform 1 0 24748 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1604681595
transform 1 0 25116 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 26404 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604681595
transform 1 0 26956 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_273
timestamp 1604681595
transform 1 0 26220 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_279
timestamp 1604681595
transform 1 0 26772 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_283
timestamp 1604681595
transform 1 0 27140 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 28888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_295
timestamp 1604681595
transform 1 0 28244 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1604681595
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_7
timestamp 1604681595
transform 1 0 1748 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_11
timestamp 1604681595
transform 1 0 2116 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 4784 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_23
timestamp 1604681595
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1604681595
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 6808 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 5980 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_42
timestamp 1604681595
transform 1 0 4968 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_50
timestamp 1604681595
transform 1 0 5704 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_55
timestamp 1604681595
transform 1 0 6164 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_59
timestamp 1604681595
transform 1 0 6532 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_71
timestamp 1604681595
transform 1 0 7636 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_83
timestamp 1604681595
transform 1 0 8740 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 10212 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8924 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1604681595
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_93
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_115
timestamp 1604681595
transform 1 0 11684 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 13616 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_129
timestamp 1604681595
transform 1 0 12972 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_135
timestamp 1604681595
transform 1 0 13524 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1604681595
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_142
timestamp 1604681595
transform 1 0 14168 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 16376 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_150
timestamp 1604681595
transform 1 0 14904 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 17112 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_12_168
timestamp 1604681595
transform 1 0 16560 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1604681595
transform 1 0 19320 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_190
timestamp 1604681595
transform 1 0 18584 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_12_201
timestamp 1604681595
transform 1 0 19596 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_209
timestamp 1604681595
transform 1 0 20332 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_224
timestamp 1604681595
transform 1 0 21712 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1604681595
transform 1 0 22448 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 23644 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_241
timestamp 1604681595
transform 1 0 23276 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_247
timestamp 1604681595
transform 1 0 23828 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1604681595
transform 1 0 24196 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 25852 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 25208 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_260
timestamp 1604681595
transform 1 0 25024 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_264
timestamp 1604681595
transform 1 0 25392 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_268
timestamp 1604681595
transform 1 0 25760 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_271
timestamp 1604681595
transform 1 0 26036 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_276
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_288
timestamp 1604681595
transform 1 0 27600 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 28888 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_296
timestamp 1604681595
transform 1 0 28336 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_7
timestamp 1604681595
transform 1 0 1748 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1604681595
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_17
timestamp 1604681595
transform 1 0 2668 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_11
timestamp 1604681595
transform 1 0 2116 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1604681595
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1604681595
transform 1 0 2484 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_19
timestamp 1604681595
transform 1 0 2852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 3496 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 3036 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 3312 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 3496 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_23
timestamp 1604681595
transform 1 0 3220 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_23
timestamp 1604681595
transform 1 0 3220 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_28
timestamp 1604681595
transform 1 0 3680 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_49
timestamp 1604681595
transform 1 0 5612 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_46
timestamp 1604681595
transform 1 0 5336 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_42
timestamp 1604681595
transform 1 0 4968 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 5428 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_56
timestamp 1604681595
transform 1 0 6256 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_56
timestamp 1604681595
transform 1 0 6256 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 5980 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 6348 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1604681595
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_70
timestamp 1604681595
transform 1 0 7544 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_66
timestamp 1604681595
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_71
timestamp 1604681595
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 7728 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1604681595
transform 1 0 8648 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_77
timestamp 1604681595
transform 1 0 8188 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_75
timestamp 1604681595
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8464 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 7912 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_79
timestamp 1604681595
transform 1 0 8372 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_86
timestamp 1604681595
transform 1 0 9016 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_91
timestamp 1604681595
transform 1 0 9476 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 9660 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_99
timestamp 1604681595
transform 1 0 10212 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_99
timestamp 1604681595
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_95
timestamp 1604681595
transform 1 0 9844 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10028 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10396 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10580 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10580 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_112
timestamp 1604681595
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_124
timestamp 1604681595
transform 1 0 12512 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1604681595
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_116
timestamp 1604681595
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 12604 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_112
timestamp 1604681595
transform 1 0 11408 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 12788 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 14444 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_143
timestamp 1604681595
transform 1 0 14260 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_129
timestamp 1604681595
transform 1 0 12972 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_135
timestamp 1604681595
transform 1 0 13524 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_145
timestamp 1604681595
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_149
timestamp 1604681595
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_147
timestamp 1604681595
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 15456 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 14812 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_158
timestamp 1604681595
transform 1 0 15640 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 14996 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_167
timestamp 1604681595
transform 1 0 16468 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_179
timestamp 1604681595
transform 1 0 17572 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_170
timestamp 1604681595
transform 1 0 16744 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_182
timestamp 1604681595
transform 1 0 17848 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_190
timestamp 1604681595
transform 1 0 18584 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_196
timestamp 1604681595
transform 1 0 19136 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_192
timestamp 1604681595
transform 1 0 18768 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 18584 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 18952 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 18676 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18952 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_14_203
timestamp 1604681595
transform 1 0 19780 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_204
timestamp 1604681595
transform 1 0 19872 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_200
timestamp 1604681595
transform 1 0 19504 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19688 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 19320 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 20976 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 20792 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 20424 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_212
timestamp 1604681595
transform 1 0 20608 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_211
timestamp 1604681595
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1604681595
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_232
timestamp 1604681595
transform 1 0 22448 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_240
timestamp 1604681595
transform 1 0 23184 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1604681595
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_255
timestamp 1604681595
transform 1 0 24564 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_251
timestamp 1604681595
transform 1 0 24196 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 24656 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1604681595
transform 1 0 24840 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_267
timestamp 1604681595
transform 1 0 25668 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_265
timestamp 1604681595
transform 1 0 25484 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_261
timestamp 1604681595
transform 1 0 25116 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 25852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 25300 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 25668 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1604681595
transform 1 0 25852 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604681595
transform 1 0 26864 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1604681595
transform 1 0 26680 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_282
timestamp 1604681595
transform 1 0 27048 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_271
timestamp 1604681595
transform 1 0 26036 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_280
timestamp 1604681595
transform 1 0 26864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 28888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 28888 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_294
timestamp 1604681595
transform 1 0 28152 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_298
timestamp 1604681595
transform 1 0 28520 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_292
timestamp 1604681595
transform 1 0 27968 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_298
timestamp 1604681595
transform 1 0 28520 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 2392 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1604681595
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1604681595
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_7
timestamp 1604681595
transform 1 0 1748 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_11
timestamp 1604681595
transform 1 0 2116 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_30
timestamp 1604681595
transform 1 0 3864 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_50
timestamp 1604681595
transform 1 0 5704 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_46
timestamp 1604681595
transform 1 0 5336 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_42
timestamp 1604681595
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 5152 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1604681595
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_54
timestamp 1604681595
transform 1 0 6072 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8464 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_71
timestamp 1604681595
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_75
timestamp 1604681595
transform 1 0 8004 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10028 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 9476 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_89
timestamp 1604681595
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_93
timestamp 1604681595
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11408 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_106
timestamp 1604681595
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1604681595
transform 1 0 11224 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_114
timestamp 1604681595
transform 1 0 11592 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1604681595
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 12788 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 13616 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_129
timestamp 1604681595
transform 1 0 12972 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_134
timestamp 1604681595
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_138
timestamp 1604681595
transform 1 0 13800 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_142
timestamp 1604681595
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1604681595
transform 1 0 16100 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1604681595
transform 1 0 14536 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 15548 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_155
timestamp 1604681595
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_159
timestamp 1604681595
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_166
timestamp 1604681595
transform 1 0 16376 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_178
timestamp 1604681595
transform 1 0 17480 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1604681595
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18952 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18768 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 19964 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_190
timestamp 1604681595
transform 1 0 18584 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_203
timestamp 1604681595
transform 1 0 19780 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_207
timestamp 1604681595
transform 1 0 20148 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 20332 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 20700 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 21896 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_211
timestamp 1604681595
transform 1 0 20516 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_215
timestamp 1604681595
transform 1 0 20884 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_223
timestamp 1604681595
transform 1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_228
timestamp 1604681595
transform 1 0 22080 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 22264 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_232
timestamp 1604681595
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1604681595
transform 1 0 25208 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_257
timestamp 1604681595
transform 1 0 24748 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_261
timestamp 1604681595
transform 1 0 25116 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_265
timestamp 1604681595
transform 1 0 25484 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 26404 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 27508 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604681595
transform 1 0 26956 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1604681595
transform 1 0 27324 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_273
timestamp 1604681595
transform 1 0 26220 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_279
timestamp 1604681595
transform 1 0 26772 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_283
timestamp 1604681595
transform 1 0 27140 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_291
timestamp 1604681595
transform 1 0 27876 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 28888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604681595
transform 1 0 28060 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_295
timestamp 1604681595
transform 1 0 28244 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1604681595
transform 1 0 2484 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 1932 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 2300 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_7
timestamp 1604681595
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_11
timestamp 1604681595
transform 1 0 2116 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_19
timestamp 1604681595
transform 1 0 2852 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 3036 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_23
timestamp 1604681595
transform 1 0 3220 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 5152 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_60
timestamp 1604681595
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_64
timestamp 1604681595
transform 1 0 6992 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10028 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_84
timestamp 1604681595
transform 1 0 8832 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_106
timestamp 1604681595
transform 1 0 10856 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_118
timestamp 1604681595
transform 1 0 11960 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_122
timestamp 1604681595
transform 1 0 12328 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_125
timestamp 1604681595
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 12788 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_143
timestamp 1604681595
transform 1 0 14260 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1604681595
transform 1 0 15364 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 16376 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_147
timestamp 1604681595
transform 1 0 14628 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_164
timestamp 1604681595
transform 1 0 16192 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 16928 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_168
timestamp 1604681595
transform 1 0 16560 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_174
timestamp 1604681595
transform 1 0 17112 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_186
timestamp 1604681595
transform 1 0 18216 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18952 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18768 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18400 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_190
timestamp 1604681595
transform 1 0 18584 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_203
timestamp 1604681595
transform 1 0 19780 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 21896 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 21436 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_211
timestamp 1604681595
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_16_223
timestamp 1604681595
transform 1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_242
timestamp 1604681595
transform 1 0 23368 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1604681595
transform 1 0 25392 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 24472 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 24840 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_256
timestamp 1604681595
transform 1 0 24656 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_260
timestamp 1604681595
transform 1 0 25024 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_267
timestamp 1604681595
transform 1 0 25668 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 27048 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 27416 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_280
timestamp 1604681595
transform 1 0 26864 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_284
timestamp 1604681595
transform 1 0 27232 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_288
timestamp 1604681595
transform 1 0 27600 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 28888 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_296
timestamp 1604681595
transform 1 0 28336 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1604681595
transform 1 0 1932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 2668 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1604681595
transform 1 0 1748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_11
timestamp 1604681595
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_15
timestamp 1604681595
transform 1 0 2484 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_19
timestamp 1604681595
transform 1 0 2852 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_31
timestamp 1604681595
transform 1 0 3956 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 5612 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_43
timestamp 1604681595
transform 1 0 5060 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_51
timestamp 1604681595
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_55
timestamp 1604681595
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1604681595
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_74
timestamp 1604681595
transform 1 0 7912 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_82
timestamp 1604681595
transform 1 0 8648 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10120 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_87
timestamp 1604681595
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_91
timestamp 1604681595
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_95
timestamp 1604681595
transform 1 0 9844 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1604681595
transform 1 0 10948 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1604681595
transform 1 0 11316 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 11408 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 1604681595
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_114
timestamp 1604681595
transform 1 0 11592 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12604 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13984 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 12972 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 13800 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 13432 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_127
timestamp 1604681595
transform 1 0 12788 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_131
timestamp 1604681595
transform 1 0 13156 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_136
timestamp 1604681595
transform 1 0 13616 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1604681595
transform 1 0 15548 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_149
timestamp 1604681595
transform 1 0 14812 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_153
timestamp 1604681595
transform 1 0 15180 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_156
timestamp 1604681595
transform 1 0 15456 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1604681595
transform 1 0 16376 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_170
timestamp 1604681595
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 16560 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_174
timestamp 1604681595
transform 1 0 17112 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_178
timestamp 1604681595
transform 1 0 17480 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 17296 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 18308 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18492 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19504 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19872 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_198
timestamp 1604681595
transform 1 0 19320 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_202
timestamp 1604681595
transform 1 0 19688 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_206
timestamp 1604681595
transform 1 0 20056 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1604681595
transform 1 0 21436 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_210
timestamp 1604681595
transform 1 0 20424 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_213
timestamp 1604681595
transform 1 0 20700 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_217
timestamp 1604681595
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 22448 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 24012 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_230
timestamp 1604681595
transform 1 0 22264 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_234
timestamp 1604681595
transform 1 0 22632 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_238
timestamp 1604681595
transform 1 0 23000 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1604681595
transform 1 0 25300 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 25116 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 24748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 24380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_251
timestamp 1604681595
transform 1 0 24196 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_255
timestamp 1604681595
transform 1 0 24564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_259
timestamp 1604681595
transform 1 0 24932 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1604681595
transform 1 0 26864 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604681595
transform 1 0 26496 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 27876 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_272
timestamp 1604681595
transform 1 0 26128 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_278
timestamp 1604681595
transform 1 0 26680 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_289
timestamp 1604681595
transform 1 0 27692 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 28888 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_293
timestamp 1604681595
transform 1 0 28060 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 1564 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 4508 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_21
timestamp 1604681595
transform 1 0 3036 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_36
timestamp 1604681595
transform 1 0 4416 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_39
timestamp 1604681595
transform 1 0 4692 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 5612 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_43
timestamp 1604681595
transform 1 0 5060 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_46
timestamp 1604681595
transform 1 0 5336 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_58
timestamp 1604681595
transform 1 0 6440 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_70
timestamp 1604681595
transform 1 0 7544 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_78
timestamp 1604681595
transform 1 0 8280 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_83
timestamp 1604681595
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 10672 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8924 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_87
timestamp 1604681595
transform 1 0 9108 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1604681595
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1604681595
transform 1 0 10488 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12420 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1604681595
transform 1 0 11408 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_106
timestamp 1604681595
transform 1 0 10856 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_110
timestamp 1604681595
transform 1 0 11224 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_121
timestamp 1604681595
transform 1 0 12236 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 14260 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 13616 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_132
timestamp 1604681595
transform 1 0 13248 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1604681595
transform 1 0 13800 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_142
timestamp 1604681595
transform 1 0 14168 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1604681595
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_163
timestamp 1604681595
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1604681595
transform 1 0 16928 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 18308 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 16652 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 17940 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_167
timestamp 1604681595
transform 1 0 16468 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_171
timestamp 1604681595
transform 1 0 16836 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_181
timestamp 1604681595
transform 1 0 17756 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_185
timestamp 1604681595
transform 1 0 18124 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18492 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_18_198
timestamp 1604681595
transform 1 0 19320 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_206
timestamp 1604681595
transform 1 0 20056 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1604681595
transform 1 0 21436 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 21068 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 20332 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_211
timestamp 1604681595
transform 1 0 20516 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_215
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_219
timestamp 1604681595
transform 1 0 21252 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1604681595
transform 1 0 23000 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 23920 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 23460 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_230
timestamp 1604681595
transform 1 0 22264 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_241
timestamp 1604681595
transform 1 0 23276 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_245
timestamp 1604681595
transform 1 0 23644 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1604681595
transform 1 0 24104 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1604681595
transform 1 0 24472 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 25484 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 25852 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 24288 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_263
timestamp 1604681595
transform 1 0 25300 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_267
timestamp 1604681595
transform 1 0 25668 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 27048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_271
timestamp 1604681595
transform 1 0 26036 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_280
timestamp 1604681595
transform 1 0 26864 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_284
timestamp 1604681595
transform 1 0 27232 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 28888 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_296
timestamp 1604681595
transform 1 0 28336 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 1564 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 1748 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 1840 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_17
timestamp 1604681595
transform 1 0 2668 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_16
timestamp 1604681595
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_20
timestamp 1604681595
transform 1 0 2944 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_21
timestamp 1604681595
transform 1 0 3036 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_24
timestamp 1604681595
transform 1 0 3312 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 3128 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 3404 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_39
timestamp 1604681595
transform 1 0 4692 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_34
timestamp 1604681595
transform 1 0 4232 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4324 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4508 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_50
timestamp 1604681595
transform 1 0 5704 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_46
timestamp 1604681595
transform 1 0 5336 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 5520 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_57
timestamp 1604681595
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_53
timestamp 1604681595
transform 1 0 5980 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 6164 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 6072 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_70
timestamp 1604681595
transform 1 0 7544 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_66
timestamp 1604681595
transform 1 0 7176 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 6992 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_77
timestamp 1604681595
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_73
timestamp 1604681595
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8556 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_20_63
timestamp 1604681595
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_93
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_88
timestamp 1604681595
transform 1 0 9200 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1604681595
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_90
timestamp 1604681595
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_100
timestamp 1604681595
transform 1 0 10304 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_97
timestamp 1604681595
transform 1 0 10028 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_94
timestamp 1604681595
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 10120 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1604681595
transform 1 0 10120 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_111
timestamp 1604681595
transform 1 0 11316 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_107
timestamp 1604681595
transform 1 0 10948 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 11500 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 11132 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1604681595
transform 1 0 10856 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_115
timestamp 1604681595
transform 1 0 11684 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1604681595
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_115
timestamp 1604681595
transform 1 0 11684 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1604681595
transform 1 0 12420 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13524 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 13340 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 12972 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_131
timestamp 1604681595
transform 1 0 13156 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_126
timestamp 1604681595
transform 1 0 12696 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_134
timestamp 1604681595
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_145
timestamp 1604681595
transform 1 0 14444 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_155
timestamp 1604681595
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_163
timestamp 1604681595
transform 1 0 16100 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_159
timestamp 1604681595
transform 1 0 15732 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 16284 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_163
timestamp 1604681595
transform 1 0 16100 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_175
timestamp 1604681595
transform 1 0 17204 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_175
timestamp 1604681595
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_167
timestamp 1604681595
transform 1 0 16468 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_179
timestamp 1604681595
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18124 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 17756 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 20148 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19136 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 19504 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_194
timestamp 1604681595
transform 1 0 18952 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_198
timestamp 1604681595
transform 1 0 19320 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_202
timestamp 1604681595
transform 1 0 19688 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_206
timestamp 1604681595
transform 1 0 20056 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1604681595
transform 1 0 19228 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 20332 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 21988 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1604681595
transform 1 0 21804 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_229
timestamp 1604681595
transform 1 0 22172 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_209
timestamp 1604681595
transform 1 0 20332 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1604681595
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_224
timestamp 1604681595
transform 1 0 21712 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_236
timestamp 1604681595
transform 1 0 22816 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_238
timestamp 1604681595
transform 1 0 23000 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_233
timestamp 1604681595
transform 1 0 22540 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 22816 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 22356 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_245
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_242
timestamp 1604681595
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 23184 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1604681595
transform 1 0 23184 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1604681595
transform 1 0 23920 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_249
timestamp 1604681595
transform 1 0 24012 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_253
timestamp 1604681595
transform 1 0 24380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_257
timestamp 1604681595
transform 1 0 24748 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 24196 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24656 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24932 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24840 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_20_267
timestamp 1604681595
transform 1 0 25668 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_261
timestamp 1604681595
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 25300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 25484 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1604681595
transform 1 0 26680 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_274
timestamp 1604681595
transform 1 0 26312 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 26496 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 26864 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_291
timestamp 1604681595
transform 1 0 27876 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 27048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1604681595
transform 1 0 27048 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_20_284
timestamp 1604681595
transform 1 0 27232 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 28888 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 28888 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_296
timestamp 1604681595
transform 1 0 28336 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 1564 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 2944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_14
timestamp 1604681595
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_18
timestamp 1604681595
transform 1 0 2760 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 3312 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_22
timestamp 1604681595
transform 1 0 3128 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_26
timestamp 1604681595
transform 1 0 3496 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_34
timestamp 1604681595
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_38
timestamp 1604681595
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4968 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_51
timestamp 1604681595
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_55
timestamp 1604681595
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1604681595
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8556 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8372 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_70
timestamp 1604681595
transform 1 0 7544 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_73
timestamp 1604681595
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_77
timestamp 1604681595
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_90
timestamp 1604681595
transform 1 0 9384 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_102
timestamp 1604681595
transform 1 0 10488 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 10948 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_105
timestamp 1604681595
transform 1 0 10764 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_109
timestamp 1604681595
transform 1 0 11132 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1604681595
transform 1 0 12236 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_135
timestamp 1604681595
transform 1 0 13524 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_143
timestamp 1604681595
transform 1 0 14260 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 15272 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15088 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 14720 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_146
timestamp 1604681595
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_150
timestamp 1604681595
transform 1 0 14904 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 16928 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_170
timestamp 1604681595
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_174
timestamp 1604681595
transform 1 0 17112 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1604681595
transform 1 0 17848 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 19504 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 19964 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 18768 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_190
timestamp 1604681595
transform 1 0 18584 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_194
timestamp 1604681595
transform 1 0 18952 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_203
timestamp 1604681595
transform 1 0 19780 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_207
timestamp 1604681595
transform 1 0 20148 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_219
timestamp 1604681595
transform 1 0 21252 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_227
timestamp 1604681595
transform 1 0 21988 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 22264 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 22632 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_232
timestamp 1604681595
transform 1 0 22448 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_236
timestamp 1604681595
transform 1 0 22816 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_245
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 25484 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 25300 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_257
timestamp 1604681595
transform 1 0 24748 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1604681595
transform 1 0 26956 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 28888 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_293
timestamp 1604681595
transform 1 0 28060 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 1840 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 1564 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1604681595
transform 1 0 1748 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_17
timestamp 1604681595
transform 1 0 2668 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1604681595
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_40
timestamp 1604681595
transform 1 0 4784 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 5520 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 4968 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_44
timestamp 1604681595
transform 1 0 5152 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 8096 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8556 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_64
timestamp 1604681595
transform 1 0 6992 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_79
timestamp 1604681595
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_83
timestamp 1604681595
transform 1 0 8740 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 10580 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1604681595
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_101
timestamp 1604681595
transform 1 0 10396 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_119
timestamp 1604681595
transform 1 0 12052 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 13524 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_131
timestamp 1604681595
transform 1 0 13156 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_137
timestamp 1604681595
transform 1 0 13708 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_149
timestamp 1604681595
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_163
timestamp 1604681595
transform 1 0 16100 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_175
timestamp 1604681595
transform 1 0 17204 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_187
timestamp 1604681595
transform 1 0 18308 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 18400 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_204
timestamp 1604681595
transform 1 0 19872 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_208
timestamp 1604681595
transform 1 0 20240 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_227
timestamp 1604681595
transform 1 0 21988 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 22264 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_22_246
timestamp 1604681595
transform 1 0 23736 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 25484 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_258
timestamp 1604681595
transform 1 0 24840 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_264
timestamp 1604681595
transform 1 0 25392 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_267
timestamp 1604681595
transform 1 0 25668 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_288
timestamp 1604681595
transform 1 0 27600 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 28888 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_296
timestamp 1604681595
transform 1 0 28336 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2300 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 2116 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 1564 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_7
timestamp 1604681595
transform 1 0 1748 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4048 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_29
timestamp 1604681595
transform 1 0 3772 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_34
timestamp 1604681595
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_38
timestamp 1604681595
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_51
timestamp 1604681595
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_48
timestamp 1604681595
transform 1 0 5520 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_42
timestamp 1604681595
transform 1 0 4968 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 5612 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_55
timestamp 1604681595
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 8372 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 8188 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_74
timestamp 1604681595
transform 1 0 7912 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_95
timestamp 1604681595
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_99
timestamp 1604681595
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_103
timestamp 1604681595
transform 1 0 10580 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 11868 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12604 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_115
timestamp 1604681595
transform 1 0 11684 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_119
timestamp 1604681595
transform 1 0 12052 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_123
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 13524 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_127
timestamp 1604681595
transform 1 0 12788 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15548 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 15916 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 16284 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_151
timestamp 1604681595
transform 1 0 14996 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_159
timestamp 1604681595
transform 1 0 15732 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_163
timestamp 1604681595
transform 1 0 16100 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_167
timestamp 1604681595
transform 1 0 16468 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1604681595
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 19320 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19136 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18768 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18400 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_190
timestamp 1604681595
transform 1 0 18584 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_194
timestamp 1604681595
transform 1 0 18952 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 21620 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 20976 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_214
timestamp 1604681595
transform 1 0 20792 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_218
timestamp 1604681595
transform 1 0 21160 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_222
timestamp 1604681595
transform 1 0 21528 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_225
timestamp 1604681595
transform 1 0 21804 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 22632 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_233
timestamp 1604681595
transform 1 0 22540 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_236
timestamp 1604681595
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_240
timestamp 1604681595
transform 1 0 23184 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 25668 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 25484 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 25116 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_257
timestamp 1604681595
transform 1 0 24748 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_263
timestamp 1604681595
transform 1 0 25300 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 27324 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_283
timestamp 1604681595
transform 1 0 27140 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_287
timestamp 1604681595
transform 1 0 27508 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 28888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1604681595
transform 1 0 1840 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 2300 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1604681595
transform 1 0 1748 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_11
timestamp 1604681595
transform 1 0 2116 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1604681595
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1604681595
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_41
timestamp 1604681595
transform 1 0 4876 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5980 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 5704 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_49
timestamp 1604681595
transform 1 0 5612 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 8372 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_69
timestamp 1604681595
transform 1 0 7452 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_77
timestamp 1604681595
transform 1 0 8188 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_81
timestamp 1604681595
transform 1 0 8556 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_89
timestamp 1604681595
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 11868 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_109
timestamp 1604681595
transform 1 0 11132 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 13524 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 13892 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14260 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_133
timestamp 1604681595
transform 1 0 13340 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_137
timestamp 1604681595
transform 1 0 13708 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1604681595
transform 1 0 14076 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_145
timestamp 1604681595
transform 1 0 14444 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15548 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_154
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1604681595
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 17848 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_178
timestamp 1604681595
transform 1 0 17480 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_185
timestamp 1604681595
transform 1 0 18124 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 18676 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_193
timestamp 1604681595
transform 1 0 18860 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_206
timestamp 1604681595
transform 1 0 20056 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 21068 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_219
timestamp 1604681595
transform 1 0 21252 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_226
timestamp 1604681595
transform 1 0 21896 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 22632 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_24_250
timestamp 1604681595
transform 1 0 24104 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 25852 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 24840 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 25208 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_260
timestamp 1604681595
transform 1 0 25024 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_264
timestamp 1604681595
transform 1 0 25392 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_268
timestamp 1604681595
transform 1 0 25760 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_271
timestamp 1604681595
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_280
timestamp 1604681595
transform 1 0 26864 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 28888 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_292
timestamp 1604681595
transform 1 0 27968 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_298
timestamp 1604681595
transform 1 0 28520 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_19
timestamp 1604681595
transform 1 0 2852 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 3588 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_36
timestamp 1604681595
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_40
timestamp 1604681595
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_44
timestamp 1604681595
transform 1 0 5152 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5336 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_48
timestamp 1604681595
transform 1 0 5520 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_55
timestamp 1604681595
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_52
timestamp 1604681595
transform 1 0 5888 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_62
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 6992 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_66
timestamp 1604681595
transform 1 0 7176 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_78
timestamp 1604681595
transform 1 0 8280 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 9384 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10488 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 9200 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_86
timestamp 1604681595
transform 1 0 9016 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_93
timestamp 1604681595
transform 1 0 9660 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_97
timestamp 1604681595
transform 1 0 10028 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_100
timestamp 1604681595
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_104
timestamp 1604681595
transform 1 0 10672 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 10856 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_108
timestamp 1604681595
transform 1 0 11040 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_120
timestamp 1604681595
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_123
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1604681595
transform 1 0 13340 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 13156 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 12788 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 14352 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_129
timestamp 1604681595
transform 1 0 12972 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_142
timestamp 1604681595
transform 1 0 14168 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 14996 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 16100 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14812 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_146
timestamp 1604681595
transform 1 0 14536 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_160
timestamp 1604681595
transform 1 0 15824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_165
timestamp 1604681595
transform 1 0 16284 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 16468 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1604681595
transform 1 0 16652 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_181
timestamp 1604681595
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1604681595
transform 1 0 19412 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 18492 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_188
timestamp 1604681595
transform 1 0 18400 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_191
timestamp 1604681595
transform 1 0 18676 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_195
timestamp 1604681595
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_208
timestamp 1604681595
transform 1 0 20240 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 20976 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 20792 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 20424 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_212
timestamp 1604681595
transform 1 0 20608 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1604681595
transform 1 0 21804 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_237
timestamp 1604681595
transform 1 0 22908 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_240
timestamp 1604681595
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 25852 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 25668 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 25300 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_261
timestamp 1604681595
transform 1 0 25116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_265
timestamp 1604681595
transform 1 0 25484 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1604681595
transform 1 0 26864 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1604681595
transform 1 0 26680 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_282
timestamp 1604681595
transform 1 0 27048 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 28888 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_294
timestamp 1604681595
transform 1 0 28152 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_298
timestamp 1604681595
transform 1 0 28520 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_7
timestamp 1604681595
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_7
timestamp 1604681595
transform 1 0 1748 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 1932 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1604681595
transform 1 0 1564 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1604681595
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_19
timestamp 1604681595
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_11
timestamp 1604681595
transform 1 0 2116 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_11
timestamp 1604681595
transform 1 0 2116 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1604681595
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_25
timestamp 1604681595
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3036 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 3220 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_40
timestamp 1604681595
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_36
timestamp 1604681595
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_32
timestamp 1604681595
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1604681595
transform 1 0 4876 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_44
timestamp 1604681595
transform 1 0 5152 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_60
timestamp 1604681595
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_56
timestamp 1604681595
transform 1 0 6256 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_52
timestamp 1604681595
transform 1 0 5888 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_53
timestamp 1604681595
transform 1 0 5980 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 6440 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 6072 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 6348 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 7176 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 6992 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 7360 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_66
timestamp 1604681595
transform 1 0 7176 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_70
timestamp 1604681595
transform 1 0 7544 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_82
timestamp 1604681595
transform 1 0 8648 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_82
timestamp 1604681595
transform 1 0 8648 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_93
timestamp 1604681595
transform 1 0 9660 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_89
timestamp 1604681595
transform 1 0 9292 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_86
timestamp 1604681595
transform 1 0 9016 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_93
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1604681595
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9108 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_97
timestamp 1604681595
transform 1 0 10028 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 9844 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 10028 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 10120 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_27_114
timestamp 1604681595
transform 1 0 11592 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1604681595
transform 1 0 11224 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_106
timestamp 1604681595
transform 1 0 10856 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 11040 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_119
timestamp 1604681595
transform 1 0 12052 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_107
timestamp 1604681595
transform 1 0 10948 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_130
timestamp 1604681595
transform 1 0 13064 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_127
timestamp 1604681595
transform 1 0 12788 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_130
timestamp 1604681595
transform 1 0 13064 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_127
timestamp 1604681595
transform 1 0 12788 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 12880 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 12880 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 13340 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 13432 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_142
timestamp 1604681595
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_143
timestamp 1604681595
transform 1 0 14260 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_154
timestamp 1604681595
transform 1 0 15272 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_150
timestamp 1604681595
transform 1 0 14904 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_146
timestamp 1604681595
transform 1 0 14536 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14720 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15364 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1604681595
transform 1 0 16376 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_159
timestamp 1604681595
transform 1 0 15732 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15548 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15548 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 16100 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_27_174
timestamp 1604681595
transform 1 0 17112 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_170
timestamp 1604681595
transform 1 0 16744 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 17296 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 16928 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 16560 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_182
timestamp 1604681595
transform 1 0 17848 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_178
timestamp 1604681595
transform 1 0 17480 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 18216 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_179
timestamp 1604681595
transform 1 0 17572 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_192
timestamp 1604681595
transform 1 0 18768 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_188
timestamp 1604681595
transform 1 0 18400 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_191
timestamp 1604681595
transform 1 0 18676 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 18952 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 18584 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 18952 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1604681595
transform 1 0 19136 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1604681595
transform 1 0 19136 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_205
timestamp 1604681595
transform 1 0 19964 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_205
timestamp 1604681595
transform 1 0 19964 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 20148 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_217
timestamp 1604681595
transform 1 0 21068 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_213
timestamp 1604681595
transform 1 0 20700 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_209
timestamp 1604681595
transform 1 0 20332 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_213
timestamp 1604681595
transform 1 0 20700 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 20516 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 21160 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1604681595
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 21344 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_222
timestamp 1604681595
transform 1 0 21528 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 21344 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_27_236
timestamp 1604681595
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_234
timestamp 1604681595
transform 1 0 22632 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 23000 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_240
timestamp 1604681595
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_247
timestamp 1604681595
transform 1 0 23828 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_244
timestamp 1604681595
transform 1 0 23552 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_240
timestamp 1604681595
transform 1 0 23184 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 23644 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 24012 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_260
timestamp 1604681595
transform 1 0 25024 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_254
timestamp 1604681595
transform 1 0 24472 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_255
timestamp 1604681595
transform 1 0 24564 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_251
timestamp 1604681595
transform 1 0 24196 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 24656 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24840 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1604681595
transform 1 0 24840 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_264
timestamp 1604681595
transform 1 0 25392 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_267
timestamp 1604681595
transform 1 0 25668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 25484 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 25852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 25668 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_271
timestamp 1604681595
transform 1 0 26036 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_280
timestamp 1604681595
transform 1 0 26864 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_283
timestamp 1604681595
transform 1 0 27140 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 28888 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 28888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_292
timestamp 1604681595
transform 1 0 27968 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_298
timestamp 1604681595
transform 1 0 28520 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_295
timestamp 1604681595
transform 1 0 28244 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1604681595
transform 1 0 2944 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 2116 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_7
timestamp 1604681595
transform 1 0 1748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_13
timestamp 1604681595
transform 1 0 2300 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_19
timestamp 1604681595
transform 1 0 2852 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_23
timestamp 1604681595
transform 1 0 3220 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_41
timestamp 1604681595
transform 1 0 4876 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 6072 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 5060 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_45
timestamp 1604681595
transform 1 0 5244 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_53
timestamp 1604681595
transform 1 0 5980 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8096 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_70
timestamp 1604681595
transform 1 0 7544 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_78
timestamp 1604681595
transform 1 0 8280 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 10212 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 10028 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_93
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_108
timestamp 1604681595
transform 1 0 11040 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_120
timestamp 1604681595
transform 1 0 12144 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1604681595
transform 1 0 12880 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 13892 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_137
timestamp 1604681595
transform 1 0 13708 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1604681595
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1604681595
transform 1 0 16192 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 15548 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 15916 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_154
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_159
timestamp 1604681595
transform 1 0 15732 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_163
timestamp 1604681595
transform 1 0 16100 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_173
timestamp 1604681595
transform 1 0 17020 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_185
timestamp 1604681595
transform 1 0 18124 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1604681595
transform 1 0 19228 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 19044 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_193
timestamp 1604681595
transform 1 0 18860 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_206
timestamp 1604681595
transform 1 0 20056 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 21068 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_215
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_219
timestamp 1604681595
transform 1 0 21252 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23000 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 22816 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_231
timestamp 1604681595
transform 1 0 22356 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_235
timestamp 1604681595
transform 1 0 22724 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_247
timestamp 1604681595
transform 1 0 23828 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24840 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 24656 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 25852 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_255
timestamp 1604681595
transform 1 0 24564 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_267
timestamp 1604681595
transform 1 0 25668 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_271
timestamp 1604681595
transform 1 0 26036 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_276
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_288
timestamp 1604681595
transform 1 0 27600 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 28888 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_296
timestamp 1604681595
transform 1 0 28336 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 2116 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 1932 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4324 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_27
timestamp 1604681595
transform 1 0 3588 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_31
timestamp 1604681595
transform 1 0 3956 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_34
timestamp 1604681595
transform 1 0 4232 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 5336 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 5704 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_44
timestamp 1604681595
transform 1 0 5152 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_48
timestamp 1604681595
transform 1 0 5520 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_52
timestamp 1604681595
transform 1 0 5888 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_60
timestamp 1604681595
transform 1 0 6624 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 8096 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7912 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 9660 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 9476 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 9108 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10672 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_85
timestamp 1604681595
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_89
timestamp 1604681595
transform 1 0 9292 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_102
timestamp 1604681595
transform 1 0 10488 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 12604 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11040 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_106
timestamp 1604681595
transform 1 0 10856 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1604681595
transform 1 0 11224 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_114
timestamp 1604681595
transform 1 0 11592 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_123
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 12788 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 14444 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_143
timestamp 1604681595
transform 1 0 14260 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1604681595
transform 1 0 15364 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 15180 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 14812 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 16376 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_147
timestamp 1604681595
transform 1 0 14628 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_151
timestamp 1604681595
transform 1 0 14996 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_164
timestamp 1604681595
transform 1 0 16192 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1604681595
transform 1 0 16928 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_168
timestamp 1604681595
transform 1 0 16560 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_175
timestamp 1604681595
transform 1 0 17204 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1604681595
transform 1 0 19412 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 18492 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_188
timestamp 1604681595
transform 1 0 18400 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_191
timestamp 1604681595
transform 1 0 18676 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_195
timestamp 1604681595
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_208
timestamp 1604681595
transform 1 0 20240 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1604681595
transform 1 0 20976 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 20792 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 20424 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_212
timestamp 1604681595
transform 1 0 20608 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1604681595
transform 1 0 21804 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 23828 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_237
timestamp 1604681595
transform 1 0 22908 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_240
timestamp 1604681595
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_245
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_249
timestamp 1604681595
transform 1 0 24012 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_261
timestamp 1604681595
transform 1 0 25116 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_273
timestamp 1604681595
transform 1 0 26220 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_285
timestamp 1604681595
transform 1 0 27324 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 28888 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_297
timestamp 1604681595
transform 1 0 28428 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604681595
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_41
timestamp 1604681595
transform 1 0 4876 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 5060 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 6808 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_45
timestamp 1604681595
transform 1 0 5244 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_57
timestamp 1604681595
transform 1 0 6348 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_61
timestamp 1604681595
transform 1 0 6716 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8096 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 8464 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_64
timestamp 1604681595
transform 1 0 6992 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_78
timestamp 1604681595
transform 1 0 8280 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_82
timestamp 1604681595
transform 1 0 8648 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1604681595
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_102
timestamp 1604681595
transform 1 0 10488 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_106
timestamp 1604681595
transform 1 0 10856 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_118
timestamp 1604681595
transform 1 0 11960 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 12788 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_126
timestamp 1604681595
transform 1 0 12696 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1604681595
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1604681595
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_170
timestamp 1604681595
transform 1 0 16744 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_182
timestamp 1604681595
transform 1 0 17848 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1604681595
transform 1 0 19412 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_194
timestamp 1604681595
transform 1 0 18952 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_198
timestamp 1604681595
transform 1 0 19320 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1604681595
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 21988 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_229
timestamp 1604681595
transform 1 0 22172 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23000 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 24012 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 22816 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_235
timestamp 1604681595
transform 1 0 22724 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_247
timestamp 1604681595
transform 1 0 23828 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 25484 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 24380 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_251
timestamp 1604681595
transform 1 0 24196 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_255
timestamp 1604681595
transform 1 0 24564 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_263
timestamp 1604681595
transform 1 0 25300 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_267
timestamp 1604681595
transform 1 0 25668 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 27048 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_279
timestamp 1604681595
transform 1 0 26772 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_284
timestamp 1604681595
transform 1 0 27232 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 28888 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_296
timestamp 1604681595
transform 1 0 28336 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_39
timestamp 1604681595
transform 1 0 4692 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 5612 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_47
timestamp 1604681595
transform 1 0 5428 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_51
timestamp 1604681595
transform 1 0 5796 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_55
timestamp 1604681595
transform 1 0 6164 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 8464 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_78
timestamp 1604681595
transform 1 0 8280 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_82
timestamp 1604681595
transform 1 0 8648 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 10120 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 9936 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 9568 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 9200 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 8832 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_86
timestamp 1604681595
transform 1 0 9016 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_90
timestamp 1604681595
transform 1 0 9384 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_94
timestamp 1604681595
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 11132 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_107
timestamp 1604681595
transform 1 0 10948 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_111
timestamp 1604681595
transform 1 0 11316 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_119
timestamp 1604681595
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1604681595
transform 1 0 12788 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1604681595
transform 1 0 13156 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_129
timestamp 1604681595
transform 1 0 12972 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_133
timestamp 1604681595
transform 1 0 13340 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_145
timestamp 1604681595
transform 1 0 14444 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1604681595
transform 1 0 16100 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 15548 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_159
timestamp 1604681595
transform 1 0 15732 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_172
timestamp 1604681595
transform 1 0 16928 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_180
timestamp 1604681595
transform 1 0 17664 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 19596 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_196
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1604681595
transform 1 0 21252 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 21804 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_217
timestamp 1604681595
transform 1 0 21068 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_221
timestamp 1604681595
transform 1 0 21436 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1604681595
transform 1 0 23920 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 23000 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_236
timestamp 1604681595
transform 1 0 22816 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_240
timestamp 1604681595
transform 1 0 23184 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_245
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1604681595
transform 1 0 25484 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 25300 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_257
timestamp 1604681595
transform 1 0 24748 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1604681595
transform 1 0 27048 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 26864 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_274
timestamp 1604681595
transform 1 0 26312 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_291
timestamp 1604681595
transform 1 0 27876 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 28888 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1604681595
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 5612 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_32_44
timestamp 1604681595
transform 1 0 5152 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_48
timestamp 1604681595
transform 1 0 5520 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_65
timestamp 1604681595
transform 1 0 7084 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_73
timestamp 1604681595
transform 1 0 7820 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 10488 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 10120 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_84
timestamp 1604681595
transform 1 0 8832 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_97
timestamp 1604681595
transform 1 0 10028 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_100
timestamp 1604681595
transform 1 0 10304 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_111
timestamp 1604681595
transform 1 0 11316 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_125
timestamp 1604681595
transform 1 0 12604 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1604681595
transform 1 0 12788 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_32_143
timestamp 1604681595
transform 1 0 14260 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 16100 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_151
timestamp 1604681595
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_162
timestamp 1604681595
transform 1 0 16008 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_165
timestamp 1604681595
transform 1 0 16284 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_177
timestamp 1604681595
transform 1 0 17388 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 19596 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_189
timestamp 1604681595
transform 1 0 18492 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_203
timestamp 1604681595
transform 1 0 19780 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 21988 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_211
timestamp 1604681595
transform 1 0 20516 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_219
timestamp 1604681595
transform 1 0 21252 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_229
timestamp 1604681595
transform 1 0 22172 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 22816 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_32_235
timestamp 1604681595
transform 1 0 22724 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 25484 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_252
timestamp 1604681595
transform 1 0 24288 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_264
timestamp 1604681595
transform 1 0 25392 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_267
timestamp 1604681595
transform 1 0 25668 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 27048 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_276
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_284
timestamp 1604681595
transform 1 0 27232 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 28888 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_296
timestamp 1604681595
transform 1 0 28336 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1604681595
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1604681595
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1604681595
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_62
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604681595
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1604681595
transform 1 0 6900 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1604681595
transform 1 0 8740 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1604681595
transform 1 0 8556 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1604681595
transform 1 0 8740 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_67
timestamp 1604681595
transform 1 0 7268 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_79
timestamp 1604681595
transform 1 0 8372 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1604681595
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_80
timestamp 1604681595
transform 1 0 8464 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 10396 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_99
timestamp 1604681595
transform 1 0 10212 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_103
timestamp 1604681595
transform 1 0 10580 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_85
timestamp 1604681595
transform 1 0 8924 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1604681595
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_102
timestamp 1604681595
transform 1 0 10488 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1604681595
transform 1 0 10948 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 10764 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1604681595
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_114
timestamp 1604681595
transform 1 0 11592 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_114
timestamp 1604681595
transform 1 0 11592 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_139
timestamp 1604681595
transform 1 0 13892 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_126
timestamp 1604681595
transform 1 0 12696 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_138
timestamp 1604681595
transform 1 0 13800 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 15824 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_151
timestamp 1604681595
transform 1 0 14996 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_159
timestamp 1604681595
transform 1 0 15732 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1604681595
transform 1 0 16376 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_150
timestamp 1604681595
transform 1 0 14904 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1604681595
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 16560 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_170
timestamp 1604681595
transform 1 0 16744 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_182
timestamp 1604681595
transform 1 0 17848 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1604681595
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1604681595
transform 1 0 19688 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1604681595
transform 1 0 19504 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_io_mode_io__0.ltile_io_physical__iopad_0.EMBEDDED_IO_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1604681595
transform 1 0 19688 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_196
timestamp 1604681595
transform 1 0 19136 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1604681595
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_204
timestamp 1604681595
transform 1 0 19872 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_218
timestamp 1604681595
transform 1 0 21160 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_212
timestamp 1604681595
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_227
timestamp 1604681595
transform 1 0 21988 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1604681595
transform 1 0 22264 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1604681595
transform 1 0 22264 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1604681595
transform 1 0 22632 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_232
timestamp 1604681595
transform 1 0 22448 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_236
timestamp 1604681595
transform 1 0 22816 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_246
timestamp 1604681595
transform 1 0 23736 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1604681595
transform 1 0 25852 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1604681595
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_258
timestamp 1604681595
transform 1 0 24840 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_270
timestamp 1604681595
transform 1 0 25944 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_274
timestamp 1604681595
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_277
timestamp 1604681595
transform 1 0 26588 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_273
timestamp 1604681595
transform 1 0 26220 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1604681595
transform 1 0 26404 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1604681595
transform 1 0 26956 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_288
timestamp 1604681595
transform 1 0 27600 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_289
timestamp 1604681595
transform 1 0 27692 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_285
timestamp 1604681595
transform 1 0 27324 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A
timestamp 1604681595
transform 1 0 27508 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 28888 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 28888 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_297
timestamp 1604681595
transform 1 0 28428 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_296
timestamp 1604681595
transform 1 0 28336 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_32
timestamp 1604681595
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_44
timestamp 1604681595
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_56
timestamp 1604681595
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_63
timestamp 1604681595
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_75
timestamp 1604681595
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_87
timestamp 1604681595
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1604681595
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_106
timestamp 1604681595
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_118
timestamp 1604681595
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1604681595
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1604681595
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_149
timestamp 1604681595
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_156
timestamp 1604681595
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_168
timestamp 1604681595
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_180
timestamp 1604681595
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_187
timestamp 1604681595
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_199
timestamp 1604681595
transform 1 0 19412 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_211
timestamp 1604681595
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_218
timestamp 1604681595
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23920 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_230
timestamp 1604681595
transform 1 0 22264 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_242
timestamp 1604681595
transform 1 0 23368 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1604681595
transform 1 0 24012 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1604681595
transform 1 0 25116 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 26772 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1604681595
transform 1 0 26220 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_280
timestamp 1604681595
transform 1 0 26864 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 28888 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_292
timestamp 1604681595
transform 1 0 27968 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_298
timestamp 1604681595
transform 1 0 28520 0 1 21216
box -38 -48 130 592
<< labels >>
rlabel metal2 s 27710 0 27766 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 4986 23520 5042 24000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 29182 0 29238 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 8298 23520 8354 24000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 2042 0 2098 480 6 bottom_grid_pin_0_
port 4 nsew default tristate
rlabel metal2 s 16302 0 16358 480 6 bottom_grid_pin_10_
port 5 nsew default tristate
rlabel metal2 s 17774 0 17830 480 6 bottom_grid_pin_11_
port 6 nsew default tristate
rlabel metal2 s 19154 0 19210 480 6 bottom_grid_pin_12_
port 7 nsew default tristate
rlabel metal2 s 20626 0 20682 480 6 bottom_grid_pin_13_
port 8 nsew default tristate
rlabel metal2 s 22006 0 22062 480 6 bottom_grid_pin_14_
port 9 nsew default tristate
rlabel metal2 s 23478 0 23534 480 6 bottom_grid_pin_15_
port 10 nsew default tristate
rlabel metal2 s 3514 0 3570 480 6 bottom_grid_pin_1_
port 11 nsew default tristate
rlabel metal2 s 4894 0 4950 480 6 bottom_grid_pin_2_
port 12 nsew default tristate
rlabel metal2 s 6366 0 6422 480 6 bottom_grid_pin_3_
port 13 nsew default tristate
rlabel metal2 s 7746 0 7802 480 6 bottom_grid_pin_4_
port 14 nsew default tristate
rlabel metal2 s 9218 0 9274 480 6 bottom_grid_pin_5_
port 15 nsew default tristate
rlabel metal2 s 10598 0 10654 480 6 bottom_grid_pin_6_
port 16 nsew default tristate
rlabel metal2 s 12070 0 12126 480 6 bottom_grid_pin_7_
port 17 nsew default tristate
rlabel metal2 s 13450 0 13506 480 6 bottom_grid_pin_8_
port 18 nsew default tristate
rlabel metal2 s 14922 0 14978 480 6 bottom_grid_pin_9_
port 19 nsew default tristate
rlabel metal2 s 24858 0 24914 480 6 bottom_width_0_height_0__pin_0_
port 20 nsew default input
rlabel metal2 s 26330 0 26386 480 6 bottom_width_0_height_0__pin_1_lower
port 21 nsew default tristate
rlabel metal2 s 662 0 718 480 6 bottom_width_0_height_0__pin_1_upper
port 22 nsew default tristate
rlabel metal2 s 11610 23520 11666 24000 6 ccff_head
port 23 nsew default input
rlabel metal2 s 14922 23520 14978 24000 6 ccff_tail
port 24 nsew default tristate
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[0]
port 25 nsew default input
rlabel metal3 s 0 18232 480 18352 6 chanx_left_in[10]
port 26 nsew default input
rlabel metal3 s 0 18776 480 18896 6 chanx_left_in[11]
port 27 nsew default input
rlabel metal3 s 0 19320 480 19440 6 chanx_left_in[12]
port 28 nsew default input
rlabel metal3 s 0 20000 480 20120 6 chanx_left_in[13]
port 29 nsew default input
rlabel metal3 s 0 20544 480 20664 6 chanx_left_in[14]
port 30 nsew default input
rlabel metal3 s 0 21224 480 21344 6 chanx_left_in[15]
port 31 nsew default input
rlabel metal3 s 0 21768 480 21888 6 chanx_left_in[16]
port 32 nsew default input
rlabel metal3 s 0 22312 480 22432 6 chanx_left_in[17]
port 33 nsew default input
rlabel metal3 s 0 22992 480 23112 6 chanx_left_in[18]
port 34 nsew default input
rlabel metal3 s 0 23536 480 23656 6 chanx_left_in[19]
port 35 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[1]
port 36 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_left_in[2]
port 37 nsew default input
rlabel metal3 s 0 14016 480 14136 6 chanx_left_in[3]
port 38 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[4]
port 39 nsew default input
rlabel metal3 s 0 15240 480 15360 6 chanx_left_in[5]
port 40 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[6]
port 41 nsew default input
rlabel metal3 s 0 16328 480 16448 6 chanx_left_in[7]
port 42 nsew default input
rlabel metal3 s 0 17008 480 17128 6 chanx_left_in[8]
port 43 nsew default input
rlabel metal3 s 0 17552 480 17672 6 chanx_left_in[9]
port 44 nsew default input
rlabel metal3 s 0 280 480 400 6 chanx_left_out[0]
port 45 nsew default tristate
rlabel metal3 s 0 6264 480 6384 6 chanx_left_out[10]
port 46 nsew default tristate
rlabel metal3 s 0 6808 480 6928 6 chanx_left_out[11]
port 47 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 chanx_left_out[12]
port 48 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 chanx_left_out[13]
port 49 nsew default tristate
rlabel metal3 s 0 8576 480 8696 6 chanx_left_out[14]
port 50 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[15]
port 51 nsew default tristate
rlabel metal3 s 0 9800 480 9920 6 chanx_left_out[16]
port 52 nsew default tristate
rlabel metal3 s 0 10344 480 10464 6 chanx_left_out[17]
port 53 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 chanx_left_out[18]
port 54 nsew default tristate
rlabel metal3 s 0 11568 480 11688 6 chanx_left_out[19]
port 55 nsew default tristate
rlabel metal3 s 0 824 480 944 6 chanx_left_out[1]
port 56 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[2]
port 57 nsew default tristate
rlabel metal3 s 0 2048 480 2168 6 chanx_left_out[3]
port 58 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 chanx_left_out[4]
port 59 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 chanx_left_out[5]
port 60 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_out[6]
port 61 nsew default tristate
rlabel metal3 s 0 4360 480 4480 6 chanx_left_out[7]
port 62 nsew default tristate
rlabel metal3 s 0 5040 480 5160 6 chanx_left_out[8]
port 63 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 chanx_left_out[9]
port 64 nsew default tristate
rlabel metal3 s 29520 12248 30000 12368 6 chanx_right_in[0]
port 65 nsew default input
rlabel metal3 s 29520 18232 30000 18352 6 chanx_right_in[10]
port 66 nsew default input
rlabel metal3 s 29520 18776 30000 18896 6 chanx_right_in[11]
port 67 nsew default input
rlabel metal3 s 29520 19320 30000 19440 6 chanx_right_in[12]
port 68 nsew default input
rlabel metal3 s 29520 20000 30000 20120 6 chanx_right_in[13]
port 69 nsew default input
rlabel metal3 s 29520 20544 30000 20664 6 chanx_right_in[14]
port 70 nsew default input
rlabel metal3 s 29520 21224 30000 21344 6 chanx_right_in[15]
port 71 nsew default input
rlabel metal3 s 29520 21768 30000 21888 6 chanx_right_in[16]
port 72 nsew default input
rlabel metal3 s 29520 22312 30000 22432 6 chanx_right_in[17]
port 73 nsew default input
rlabel metal3 s 29520 22992 30000 23112 6 chanx_right_in[18]
port 74 nsew default input
rlabel metal3 s 29520 23536 30000 23656 6 chanx_right_in[19]
port 75 nsew default input
rlabel metal3 s 29520 12792 30000 12912 6 chanx_right_in[1]
port 76 nsew default input
rlabel metal3 s 29520 13336 30000 13456 6 chanx_right_in[2]
port 77 nsew default input
rlabel metal3 s 29520 14016 30000 14136 6 chanx_right_in[3]
port 78 nsew default input
rlabel metal3 s 29520 14560 30000 14680 6 chanx_right_in[4]
port 79 nsew default input
rlabel metal3 s 29520 15240 30000 15360 6 chanx_right_in[5]
port 80 nsew default input
rlabel metal3 s 29520 15784 30000 15904 6 chanx_right_in[6]
port 81 nsew default input
rlabel metal3 s 29520 16328 30000 16448 6 chanx_right_in[7]
port 82 nsew default input
rlabel metal3 s 29520 17008 30000 17128 6 chanx_right_in[8]
port 83 nsew default input
rlabel metal3 s 29520 17552 30000 17672 6 chanx_right_in[9]
port 84 nsew default input
rlabel metal3 s 29520 280 30000 400 6 chanx_right_out[0]
port 85 nsew default tristate
rlabel metal3 s 29520 6264 30000 6384 6 chanx_right_out[10]
port 86 nsew default tristate
rlabel metal3 s 29520 6808 30000 6928 6 chanx_right_out[11]
port 87 nsew default tristate
rlabel metal3 s 29520 7352 30000 7472 6 chanx_right_out[12]
port 88 nsew default tristate
rlabel metal3 s 29520 8032 30000 8152 6 chanx_right_out[13]
port 89 nsew default tristate
rlabel metal3 s 29520 8576 30000 8696 6 chanx_right_out[14]
port 90 nsew default tristate
rlabel metal3 s 29520 9256 30000 9376 6 chanx_right_out[15]
port 91 nsew default tristate
rlabel metal3 s 29520 9800 30000 9920 6 chanx_right_out[16]
port 92 nsew default tristate
rlabel metal3 s 29520 10344 30000 10464 6 chanx_right_out[17]
port 93 nsew default tristate
rlabel metal3 s 29520 11024 30000 11144 6 chanx_right_out[18]
port 94 nsew default tristate
rlabel metal3 s 29520 11568 30000 11688 6 chanx_right_out[19]
port 95 nsew default tristate
rlabel metal3 s 29520 824 30000 944 6 chanx_right_out[1]
port 96 nsew default tristate
rlabel metal3 s 29520 1368 30000 1488 6 chanx_right_out[2]
port 97 nsew default tristate
rlabel metal3 s 29520 2048 30000 2168 6 chanx_right_out[3]
port 98 nsew default tristate
rlabel metal3 s 29520 2592 30000 2712 6 chanx_right_out[4]
port 99 nsew default tristate
rlabel metal3 s 29520 3272 30000 3392 6 chanx_right_out[5]
port 100 nsew default tristate
rlabel metal3 s 29520 3816 30000 3936 6 chanx_right_out[6]
port 101 nsew default tristate
rlabel metal3 s 29520 4360 30000 4480 6 chanx_right_out[7]
port 102 nsew default tristate
rlabel metal3 s 29520 5040 30000 5160 6 chanx_right_out[8]
port 103 nsew default tristate
rlabel metal3 s 29520 5584 30000 5704 6 chanx_right_out[9]
port 104 nsew default tristate
rlabel metal2 s 21638 23520 21694 24000 6 gfpga_pad_EMBEDDED_IO_SOC_DIR
port 105 nsew default tristate
rlabel metal2 s 24950 23520 25006 24000 6 gfpga_pad_EMBEDDED_IO_SOC_IN
port 106 nsew default input
rlabel metal2 s 28262 23520 28318 24000 6 gfpga_pad_EMBEDDED_IO_SOC_OUT
port 107 nsew default tristate
rlabel metal2 s 1674 23520 1730 24000 6 prog_clk
port 108 nsew default input
rlabel metal2 s 18326 23520 18382 24000 6 top_grid_pin_0_
port 109 nsew default tristate
rlabel metal4 s 5944 2128 6264 21808 6 VPWR
port 110 nsew default input
rlabel metal4 s 10944 2128 11264 21808 6 VGND
port 111 nsew default input
<< properties >>
string FIXED_BBOX 0 0 30000 24000
<< end >>
