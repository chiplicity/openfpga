magic
tech sky130A
magscale 1 2
timestamp 1606930436
<< locali >>
rect 16773 18207 16807 18377
rect 14289 17595 14323 17697
rect 13829 17051 13863 17289
rect 9781 16439 9815 16745
rect 16681 14943 16715 15045
rect 12173 14399 12207 14569
rect 15301 14467 15335 14569
rect 7297 13243 7331 13481
rect 16129 13311 16163 13481
rect 8033 12699 8067 12869
rect 20269 11543 20303 11781
rect 19257 10999 19291 11305
rect 4905 10523 4939 10761
rect 8401 10591 8435 10761
rect 7849 10047 7883 10217
rect 5457 8959 5491 9129
rect 15025 8959 15059 9129
rect 19625 8959 19659 9129
rect 4169 8279 4203 8381
rect 7573 8347 7607 8449
rect 5641 7871 5675 8041
rect 7757 7871 7791 8041
rect 15025 2839 15059 3009
<< viali >>
rect 1961 20009 1995 20043
rect 8677 20009 8711 20043
rect 10333 20009 10367 20043
rect 14473 20009 14507 20043
rect 16037 20009 16071 20043
rect 18521 20009 18555 20043
rect 19625 20009 19659 20043
rect 20177 20009 20211 20043
rect 20729 20009 20763 20043
rect 1777 19873 1811 19907
rect 2329 19873 2363 19907
rect 2881 19873 2915 19907
rect 7665 19873 7699 19907
rect 8585 19873 8619 19907
rect 9229 19873 9263 19907
rect 10241 19873 10275 19907
rect 11345 19873 11379 19907
rect 11437 19873 11471 19907
rect 11989 19873 12023 19907
rect 13277 19873 13311 19907
rect 14289 19873 14323 19907
rect 14841 19873 14875 19907
rect 15853 19873 15887 19907
rect 17233 19873 17267 19907
rect 18337 19873 18371 19907
rect 18889 19873 18923 19907
rect 19441 19873 19475 19907
rect 19993 19873 20027 19907
rect 20545 19873 20579 19907
rect 8769 19805 8803 19839
rect 10425 19805 10459 19839
rect 11529 19805 11563 19839
rect 13369 19805 13403 19839
rect 13553 19805 13587 19839
rect 17325 19805 17359 19839
rect 17417 19805 17451 19839
rect 2513 19737 2547 19771
rect 7849 19737 7883 19771
rect 15025 19737 15059 19771
rect 19073 19737 19107 19771
rect 3065 19669 3099 19703
rect 8217 19669 8251 19703
rect 9873 19669 9907 19703
rect 10977 19669 11011 19703
rect 12173 19669 12207 19703
rect 12909 19669 12943 19703
rect 16865 19669 16899 19703
rect 1961 19465 1995 19499
rect 3433 19465 3467 19499
rect 8493 19465 8527 19499
rect 9413 19329 9447 19363
rect 14289 19329 14323 19363
rect 15485 19329 15519 19363
rect 17417 19329 17451 19363
rect 17601 19329 17635 19363
rect 1777 19261 1811 19295
rect 2329 19261 2363 19295
rect 3249 19261 3283 19295
rect 3985 19261 4019 19295
rect 5917 19261 5951 19295
rect 7113 19261 7147 19295
rect 9229 19261 9263 19295
rect 10333 19261 10367 19295
rect 10600 19261 10634 19295
rect 12449 19261 12483 19295
rect 14105 19261 14139 19295
rect 15853 19261 15887 19295
rect 18061 19261 18095 19295
rect 18889 19261 18923 19295
rect 19993 19261 20027 19295
rect 20545 19261 20579 19295
rect 4629 19193 4663 19227
rect 7380 19193 7414 19227
rect 12716 19193 12750 19227
rect 16129 19193 16163 19227
rect 18337 19193 18371 19227
rect 19165 19193 19199 19227
rect 2513 19125 2547 19159
rect 6101 19125 6135 19159
rect 8769 19125 8803 19159
rect 9137 19125 9171 19159
rect 11713 19125 11747 19159
rect 13829 19125 13863 19159
rect 14841 19125 14875 19159
rect 15209 19125 15243 19159
rect 15301 19125 15335 19159
rect 16957 19125 16991 19159
rect 17325 19125 17359 19159
rect 20177 19125 20211 19159
rect 20729 19125 20763 19159
rect 2053 18921 2087 18955
rect 2605 18921 2639 18955
rect 5549 18921 5583 18955
rect 9137 18921 9171 18955
rect 12173 18921 12207 18955
rect 16865 18921 16899 18955
rect 18521 18921 18555 18955
rect 6561 18853 6595 18887
rect 7297 18853 7331 18887
rect 8024 18853 8058 18887
rect 9934 18853 9968 18887
rect 11713 18853 11747 18887
rect 12633 18853 12667 18887
rect 13452 18853 13486 18887
rect 15730 18853 15764 18887
rect 17408 18853 17442 18887
rect 19042 18853 19076 18887
rect 1869 18785 1903 18819
rect 2421 18785 2455 18819
rect 2973 18785 3007 18819
rect 5365 18785 5399 18819
rect 6285 18785 6319 18819
rect 7021 18785 7055 18819
rect 7757 18785 7791 18819
rect 11437 18785 11471 18819
rect 12541 18785 12575 18819
rect 9689 18717 9723 18751
rect 12725 18717 12759 18751
rect 13185 18717 13219 18751
rect 15485 18717 15519 18751
rect 17141 18717 17175 18751
rect 18797 18717 18831 18751
rect 3157 18649 3191 18683
rect 11069 18649 11103 18683
rect 14565 18581 14599 18615
rect 20177 18581 20211 18615
rect 1961 18377 1995 18411
rect 8217 18377 8251 18411
rect 11437 18377 11471 18411
rect 12909 18377 12943 18411
rect 15669 18377 15703 18411
rect 15945 18377 15979 18411
rect 16773 18377 16807 18411
rect 16957 18377 16991 18411
rect 20729 18377 20763 18411
rect 3801 18309 3835 18343
rect 2513 18241 2547 18275
rect 4813 18241 4847 18275
rect 7481 18241 7515 18275
rect 8769 18241 8803 18275
rect 13461 18241 13495 18275
rect 14289 18241 14323 18275
rect 16497 18241 16531 18275
rect 18521 18309 18555 18343
rect 17509 18241 17543 18275
rect 19165 18241 19199 18275
rect 20177 18241 20211 18275
rect 1777 18173 1811 18207
rect 2318 18173 2352 18207
rect 3065 18173 3099 18207
rect 3617 18173 3651 18207
rect 4537 18173 4571 18207
rect 8585 18173 8619 18207
rect 9229 18173 9263 18207
rect 10057 18173 10091 18207
rect 12449 18173 12483 18207
rect 14556 18173 14590 18207
rect 16773 18173 16807 18207
rect 20545 18173 20579 18207
rect 7297 18105 7331 18139
rect 7389 18105 7423 18139
rect 9505 18105 9539 18139
rect 10302 18105 10336 18139
rect 11897 18105 11931 18139
rect 13277 18105 13311 18139
rect 13369 18105 13403 18139
rect 16313 18105 16347 18139
rect 17325 18105 17359 18139
rect 18061 18105 18095 18139
rect 18889 18105 18923 18139
rect 19901 18105 19935 18139
rect 3249 18037 3283 18071
rect 6929 18037 6963 18071
rect 8677 18037 8711 18071
rect 16405 18037 16439 18071
rect 17417 18037 17451 18071
rect 18981 18037 19015 18071
rect 19533 18037 19567 18071
rect 19993 18037 20027 18071
rect 1961 17833 1995 17867
rect 2513 17833 2547 17867
rect 7205 17833 7239 17867
rect 9045 17833 9079 17867
rect 11069 17833 11103 17867
rect 11345 17833 11379 17867
rect 13185 17833 13219 17867
rect 15301 17833 15335 17867
rect 16589 17833 16623 17867
rect 17877 17833 17911 17867
rect 18613 17833 18647 17867
rect 20913 17833 20947 17867
rect 9956 17765 9990 17799
rect 11805 17765 11839 17799
rect 15669 17765 15703 17799
rect 19248 17765 19282 17799
rect 1777 17697 1811 17731
rect 2329 17697 2363 17731
rect 2881 17697 2915 17731
rect 4445 17697 4479 17731
rect 4537 17697 4571 17731
rect 5816 17697 5850 17731
rect 7573 17697 7607 17731
rect 8953 17697 8987 17731
rect 11713 17697 11747 17731
rect 12357 17697 12391 17731
rect 13921 17697 13955 17731
rect 14289 17697 14323 17731
rect 14473 17697 14507 17731
rect 14749 17697 14783 17731
rect 15761 17697 15795 17731
rect 16405 17697 16439 17731
rect 16957 17697 16991 17731
rect 17693 17697 17727 17731
rect 18429 17697 18463 17731
rect 4721 17629 4755 17663
rect 5549 17629 5583 17663
rect 7665 17629 7699 17663
rect 7757 17629 7791 17663
rect 9229 17629 9263 17663
rect 9689 17629 9723 17663
rect 11897 17629 11931 17663
rect 13277 17629 13311 17663
rect 13461 17629 13495 17663
rect 15853 17629 15887 17663
rect 17141 17629 17175 17663
rect 18981 17629 19015 17663
rect 14289 17561 14323 17595
rect 3065 17493 3099 17527
rect 4077 17493 4111 17527
rect 6929 17493 6963 17527
rect 8585 17493 8619 17527
rect 12817 17493 12851 17527
rect 14105 17493 14139 17527
rect 20361 17493 20395 17527
rect 2513 17289 2547 17323
rect 6837 17289 6871 17323
rect 11161 17289 11195 17323
rect 12909 17289 12943 17323
rect 13829 17289 13863 17323
rect 14105 17289 14139 17323
rect 15393 17289 15427 17323
rect 15945 17289 15979 17323
rect 18061 17289 18095 17323
rect 19257 17289 19291 17323
rect 3525 17221 3559 17255
rect 5917 17221 5951 17255
rect 3985 17153 4019 17187
rect 4169 17153 4203 17187
rect 7297 17153 7331 17187
rect 7389 17153 7423 17187
rect 8401 17153 8435 17187
rect 9413 17153 9447 17187
rect 9597 17153 9631 17187
rect 10517 17153 10551 17187
rect 11805 17153 11839 17187
rect 13553 17153 13587 17187
rect 1777 17085 1811 17119
rect 2329 17085 2363 17119
rect 2881 17085 2915 17119
rect 4537 17085 4571 17119
rect 13277 17085 13311 17119
rect 13369 17085 13403 17119
rect 20729 17221 20763 17255
rect 18705 17153 18739 17187
rect 19809 17153 19843 17187
rect 13921 17085 13955 17119
rect 14473 17085 14507 17119
rect 14749 17085 14783 17119
rect 15209 17085 15243 17119
rect 15761 17085 15795 17119
rect 16313 17085 16347 17119
rect 16580 17085 16614 17119
rect 19625 17085 19659 17119
rect 20545 17085 20579 17119
rect 4804 17017 4838 17051
rect 7205 17017 7239 17051
rect 8309 17017 8343 17051
rect 10333 17017 10367 17051
rect 10425 17017 10459 17051
rect 11529 17017 11563 17051
rect 13829 17017 13863 17051
rect 1961 16949 1995 16983
rect 3065 16949 3099 16983
rect 3893 16949 3927 16983
rect 7849 16949 7883 16983
rect 8217 16949 8251 16983
rect 8953 16949 8987 16983
rect 9321 16949 9355 16983
rect 9965 16949 9999 16983
rect 11621 16949 11655 16983
rect 12449 16949 12483 16983
rect 17693 16949 17727 16983
rect 18429 16949 18463 16983
rect 18521 16949 18555 16983
rect 19717 16949 19751 16983
rect 3709 16745 3743 16779
rect 5457 16745 5491 16779
rect 7481 16745 7515 16779
rect 9781 16745 9815 16779
rect 9873 16745 9907 16779
rect 10517 16745 10551 16779
rect 11897 16745 11931 16779
rect 11989 16745 12023 16779
rect 12541 16745 12575 16779
rect 14105 16745 14139 16779
rect 14565 16745 14599 16779
rect 19625 16745 19659 16779
rect 4344 16677 4378 16711
rect 6368 16677 6402 16711
rect 8002 16677 8036 16711
rect 1777 16609 1811 16643
rect 2596 16609 2630 16643
rect 4077 16609 4111 16643
rect 6101 16609 6135 16643
rect 2329 16541 2363 16575
rect 7757 16541 7791 16575
rect 1961 16473 1995 16507
rect 9137 16473 9171 16507
rect 13645 16677 13679 16711
rect 15669 16677 15703 16711
rect 20177 16677 20211 16711
rect 10057 16609 10091 16643
rect 10885 16609 10919 16643
rect 12909 16609 12943 16643
rect 13001 16609 13035 16643
rect 14473 16609 14507 16643
rect 15761 16609 15795 16643
rect 16865 16609 16899 16643
rect 17509 16609 17543 16643
rect 18512 16609 18546 16643
rect 19901 16609 19935 16643
rect 20913 16609 20947 16643
rect 10977 16541 11011 16575
rect 11161 16541 11195 16575
rect 12173 16541 12207 16575
rect 13185 16541 13219 16575
rect 14749 16541 14783 16575
rect 15853 16541 15887 16575
rect 16957 16541 16991 16575
rect 17141 16541 17175 16575
rect 18245 16541 18279 16575
rect 11529 16473 11563 16507
rect 9781 16405 9815 16439
rect 15301 16405 15335 16439
rect 16497 16405 16531 16439
rect 17693 16405 17727 16439
rect 4353 16201 4387 16235
rect 6837 16201 6871 16235
rect 8953 16201 8987 16235
rect 11345 16201 11379 16235
rect 13829 16201 13863 16235
rect 15485 16201 15519 16235
rect 17601 16201 17635 16235
rect 20361 16201 20395 16235
rect 2605 16133 2639 16167
rect 3157 16065 3191 16099
rect 4905 16065 4939 16099
rect 7389 16065 7423 16099
rect 8401 16065 8435 16099
rect 9505 16065 9539 16099
rect 9965 16065 9999 16099
rect 11897 16065 11931 16099
rect 18245 16065 18279 16099
rect 1777 15997 1811 16031
rect 2973 15997 3007 16031
rect 8309 15997 8343 16031
rect 9321 15997 9355 16031
rect 9413 15997 9447 16031
rect 10221 15997 10255 16031
rect 11621 15997 11655 16031
rect 12449 15997 12483 16031
rect 14105 15997 14139 16031
rect 14361 15997 14395 16031
rect 15761 15997 15795 16031
rect 16017 15997 16051 16031
rect 17417 15997 17451 16031
rect 18061 15997 18095 16031
rect 18981 15997 19015 16031
rect 20637 15997 20671 16031
rect 4721 15929 4755 15963
rect 7205 15929 7239 15963
rect 12716 15929 12750 15963
rect 19248 15929 19282 15963
rect 20913 15929 20947 15963
rect 1961 15861 1995 15895
rect 3065 15861 3099 15895
rect 4813 15861 4847 15895
rect 7297 15861 7331 15895
rect 7849 15861 7883 15895
rect 8217 15861 8251 15895
rect 17141 15861 17175 15895
rect 1961 15657 1995 15691
rect 2513 15657 2547 15691
rect 4077 15657 4111 15691
rect 4445 15657 4479 15691
rect 5089 15657 5123 15691
rect 6101 15657 6135 15691
rect 7389 15657 7423 15691
rect 7757 15657 7791 15691
rect 8585 15657 8619 15691
rect 8953 15657 8987 15691
rect 10333 15657 10367 15691
rect 13461 15657 13495 15691
rect 14105 15657 14139 15691
rect 14473 15657 14507 15691
rect 15669 15657 15703 15691
rect 18153 15657 18187 15691
rect 18705 15657 18739 15691
rect 19073 15657 19107 15691
rect 2881 15589 2915 15623
rect 2973 15589 3007 15623
rect 6929 15589 6963 15623
rect 13369 15589 13403 15623
rect 16304 15589 16338 15623
rect 1777 15521 1811 15555
rect 3525 15521 3559 15555
rect 5457 15521 5491 15555
rect 6285 15521 6319 15555
rect 10701 15521 10735 15555
rect 10793 15521 10827 15555
rect 11345 15521 11379 15555
rect 11601 15521 11635 15555
rect 15485 15521 15519 15555
rect 18061 15521 18095 15555
rect 20085 15521 20119 15555
rect 3157 15453 3191 15487
rect 4537 15453 4571 15487
rect 4721 15453 4755 15487
rect 5549 15453 5583 15487
rect 5641 15453 5675 15487
rect 7849 15453 7883 15487
rect 7941 15453 7975 15487
rect 9045 15453 9079 15487
rect 9229 15453 9263 15487
rect 10885 15453 10919 15487
rect 13553 15453 13587 15487
rect 14565 15453 14599 15487
rect 14657 15453 14691 15487
rect 16037 15453 16071 15487
rect 18245 15453 18279 15487
rect 19165 15453 19199 15487
rect 19257 15453 19291 15487
rect 20177 15453 20211 15487
rect 20269 15453 20303 15487
rect 12725 15385 12759 15419
rect 13001 15385 13035 15419
rect 17417 15385 17451 15419
rect 19717 15385 19751 15419
rect 17693 15317 17727 15351
rect 4537 15113 4571 15147
rect 7849 15113 7883 15147
rect 10149 15113 10183 15147
rect 10609 15113 10643 15147
rect 13645 15113 13679 15147
rect 14289 15113 14323 15147
rect 14657 15113 14691 15147
rect 16773 15113 16807 15147
rect 19441 15113 19475 15147
rect 19717 15113 19751 15147
rect 20913 15113 20947 15147
rect 16681 15045 16715 15079
rect 1869 14977 1903 15011
rect 5181 14977 5215 15011
rect 7297 14977 7331 15011
rect 7481 14977 7515 15011
rect 8769 14977 8803 15011
rect 11253 14977 11287 15011
rect 13277 14977 13311 15011
rect 15209 14977 15243 15011
rect 17417 14977 17451 15011
rect 20269 14977 20303 15011
rect 1593 14909 1627 14943
rect 2329 14909 2363 14943
rect 8033 14909 8067 14943
rect 9036 14909 9070 14943
rect 11805 14909 11839 14943
rect 13829 14909 13863 14943
rect 14105 14909 14139 14943
rect 15669 14909 15703 14943
rect 16221 14909 16255 14943
rect 16681 14909 16715 14943
rect 17233 14909 17267 14943
rect 18061 14909 18095 14943
rect 18317 14909 18351 14943
rect 20177 14909 20211 14943
rect 20729 14909 20763 14943
rect 2596 14841 2630 14875
rect 4905 14841 4939 14875
rect 7205 14841 7239 14875
rect 11069 14841 11103 14875
rect 13093 14841 13127 14875
rect 15025 14841 15059 14875
rect 3709 14773 3743 14807
rect 4997 14773 5031 14807
rect 6837 14773 6871 14807
rect 10977 14773 11011 14807
rect 11989 14773 12023 14807
rect 12633 14773 12667 14807
rect 13001 14773 13035 14807
rect 15117 14773 15151 14807
rect 15853 14773 15887 14807
rect 16405 14773 16439 14807
rect 17141 14773 17175 14807
rect 20085 14773 20119 14807
rect 1961 14569 1995 14603
rect 2697 14569 2731 14603
rect 5825 14569 5859 14603
rect 8125 14569 8159 14603
rect 10057 14569 10091 14603
rect 10793 14569 10827 14603
rect 11253 14569 11287 14603
rect 11621 14569 11655 14603
rect 12173 14569 12207 14603
rect 14657 14569 14691 14603
rect 15301 14569 15335 14603
rect 16313 14569 16347 14603
rect 18337 14569 18371 14603
rect 18613 14569 18647 14603
rect 6346 14501 6380 14535
rect 8217 14501 8251 14535
rect 1777 14433 1811 14467
rect 3065 14433 3099 14467
rect 4445 14433 4479 14467
rect 4712 14433 4746 14467
rect 10149 14433 10183 14467
rect 17224 14501 17258 14535
rect 18981 14501 19015 14535
rect 20913 14501 20947 14535
rect 12532 14433 12566 14467
rect 14105 14433 14139 14467
rect 14565 14433 14599 14467
rect 15301 14433 15335 14467
rect 15393 14433 15427 14467
rect 16405 14433 16439 14467
rect 19993 14433 20027 14467
rect 3157 14365 3191 14399
rect 3249 14365 3283 14399
rect 6101 14365 6135 14399
rect 8309 14365 8343 14399
rect 10333 14365 10367 14399
rect 11713 14365 11747 14399
rect 11897 14365 11931 14399
rect 12173 14365 12207 14399
rect 12265 14365 12299 14399
rect 14749 14365 14783 14399
rect 16497 14365 16531 14399
rect 16957 14365 16991 14399
rect 19073 14365 19107 14399
rect 19165 14365 19199 14399
rect 20085 14365 20119 14399
rect 20177 14365 20211 14399
rect 13921 14297 13955 14331
rect 15577 14297 15611 14331
rect 7481 14229 7515 14263
rect 7757 14229 7791 14263
rect 9689 14229 9723 14263
rect 13645 14229 13679 14263
rect 14197 14229 14231 14263
rect 15945 14229 15979 14263
rect 19625 14229 19659 14263
rect 5089 14025 5123 14059
rect 5365 14025 5399 14059
rect 8769 14025 8803 14059
rect 11345 14025 11379 14059
rect 15025 14025 15059 14059
rect 8861 13957 8895 13991
rect 10517 13957 10551 13991
rect 1685 13889 1719 13923
rect 3709 13889 3743 13923
rect 5917 13889 5951 13923
rect 9321 13889 9355 13923
rect 9413 13889 9447 13923
rect 10333 13889 10367 13923
rect 10977 13889 11011 13923
rect 11069 13889 11103 13923
rect 11805 13889 11839 13923
rect 11989 13889 12023 13923
rect 13369 13889 13403 13923
rect 15577 13889 15611 13923
rect 16589 13889 16623 13923
rect 17509 13889 17543 13923
rect 20821 13889 20855 13923
rect 1409 13821 1443 13855
rect 2145 13821 2179 13855
rect 3976 13821 4010 13855
rect 5825 13821 5859 13855
rect 7389 13821 7423 13855
rect 10149 13821 10183 13855
rect 13636 13821 13670 13855
rect 16497 13821 16531 13855
rect 17233 13821 17267 13855
rect 18061 13821 18095 13855
rect 18613 13821 18647 13855
rect 18880 13821 18914 13855
rect 20729 13821 20763 13855
rect 2421 13753 2455 13787
rect 7656 13753 7690 13787
rect 10057 13753 10091 13787
rect 11713 13753 11747 13787
rect 5733 13685 5767 13719
rect 9229 13685 9263 13719
rect 9689 13685 9723 13719
rect 10885 13685 10919 13719
rect 12909 13685 12943 13719
rect 14749 13685 14783 13719
rect 15393 13685 15427 13719
rect 15485 13685 15519 13719
rect 16037 13685 16071 13719
rect 16405 13685 16439 13719
rect 18245 13685 18279 13719
rect 19993 13685 20027 13719
rect 20269 13685 20303 13719
rect 20637 13685 20671 13719
rect 1777 13481 1811 13515
rect 4445 13481 4479 13515
rect 5825 13481 5859 13515
rect 6929 13481 6963 13515
rect 7297 13481 7331 13515
rect 8861 13481 8895 13515
rect 11437 13481 11471 13515
rect 13001 13481 13035 13515
rect 13461 13481 13495 13515
rect 14841 13481 14875 13515
rect 15301 13481 15335 13515
rect 16129 13481 16163 13515
rect 17693 13481 17727 13515
rect 19625 13481 19659 13515
rect 2237 13413 2271 13447
rect 2789 13413 2823 13447
rect 1593 13345 1627 13379
rect 2697 13345 2731 13379
rect 4813 13345 4847 13379
rect 6837 13345 6871 13379
rect 2973 13277 3007 13311
rect 4905 13277 4939 13311
rect 5089 13277 5123 13311
rect 5917 13277 5951 13311
rect 6009 13277 6043 13311
rect 7113 13277 7147 13311
rect 7748 13413 7782 13447
rect 10324 13413 10358 13447
rect 11774 13413 11808 13447
rect 15669 13413 15703 13447
rect 15761 13413 15795 13447
rect 11529 13345 11563 13379
rect 13369 13345 13403 13379
rect 14197 13345 14231 13379
rect 14657 13345 14691 13379
rect 16580 13413 16614 13447
rect 18236 13345 18270 13379
rect 19993 13345 20027 13379
rect 7481 13277 7515 13311
rect 10057 13277 10091 13311
rect 13645 13277 13679 13311
rect 14289 13277 14323 13311
rect 14473 13277 14507 13311
rect 15945 13277 15979 13311
rect 16129 13277 16163 13311
rect 16313 13277 16347 13311
rect 17969 13277 18003 13311
rect 20085 13277 20119 13311
rect 20177 13277 20211 13311
rect 5457 13209 5491 13243
rect 7297 13209 7331 13243
rect 12909 13209 12943 13243
rect 2329 13141 2363 13175
rect 6469 13141 6503 13175
rect 13829 13141 13863 13175
rect 19349 13141 19383 13175
rect 1961 12937 1995 12971
rect 4721 12937 4755 12971
rect 7205 12937 7239 12971
rect 18981 12937 19015 12971
rect 3893 12869 3927 12903
rect 5733 12869 5767 12903
rect 8033 12869 8067 12903
rect 8217 12869 8251 12903
rect 9689 12869 9723 12903
rect 16957 12869 16991 12903
rect 4261 12801 4295 12835
rect 5273 12801 5307 12835
rect 6285 12801 6319 12835
rect 7665 12801 7699 12835
rect 7849 12801 7883 12835
rect 1777 12733 1811 12767
rect 2513 12733 2547 12767
rect 5181 12733 5215 12767
rect 8861 12801 8895 12835
rect 13737 12801 13771 12835
rect 13829 12801 13863 12835
rect 14105 12801 14139 12835
rect 15853 12801 15887 12835
rect 16497 12801 16531 12835
rect 17509 12801 17543 12835
rect 18429 12801 18463 12835
rect 19625 12801 19659 12835
rect 20545 12801 20579 12835
rect 8677 12733 8711 12767
rect 9873 12733 9907 12767
rect 11989 12733 12023 12767
rect 13001 12733 13035 12767
rect 14372 12733 14406 12767
rect 18245 12733 18279 12767
rect 19349 12733 19383 12767
rect 2780 12665 2814 12699
rect 6193 12665 6227 12699
rect 7573 12665 7607 12699
rect 8033 12665 8067 12699
rect 8585 12665 8619 12699
rect 9229 12665 9263 12699
rect 10425 12665 10459 12699
rect 16313 12665 16347 12699
rect 17325 12665 17359 12699
rect 17417 12665 17451 12699
rect 19441 12665 19475 12699
rect 20361 12665 20395 12699
rect 5089 12597 5123 12631
rect 6101 12597 6135 12631
rect 12817 12597 12851 12631
rect 13277 12597 13311 12631
rect 13645 12597 13679 12631
rect 15485 12597 15519 12631
rect 15945 12597 15979 12631
rect 16405 12597 16439 12631
rect 19993 12597 20027 12631
rect 20453 12597 20487 12631
rect 2973 12393 3007 12427
rect 12633 12393 12667 12427
rect 14289 12393 14323 12427
rect 15301 12393 15335 12427
rect 15669 12393 15703 12427
rect 17877 12393 17911 12427
rect 19625 12393 19659 12427
rect 19993 12393 20027 12427
rect 20913 12393 20947 12427
rect 4804 12325 4838 12359
rect 10609 12325 10643 12359
rect 13176 12325 13210 12359
rect 14749 12325 14783 12359
rect 1593 12257 1627 12291
rect 1860 12257 1894 12291
rect 6449 12257 6483 12291
rect 8116 12257 8150 12291
rect 11520 12257 11554 12291
rect 12909 12257 12943 12291
rect 15761 12257 15795 12291
rect 16497 12257 16531 12291
rect 16764 12257 16798 12291
rect 18981 12257 19015 12291
rect 19073 12257 19107 12291
rect 4537 12189 4571 12223
rect 6193 12189 6227 12223
rect 7849 12189 7883 12223
rect 10701 12189 10735 12223
rect 10885 12189 10919 12223
rect 11253 12189 11287 12223
rect 15945 12189 15979 12223
rect 19257 12189 19291 12223
rect 20085 12189 20119 12223
rect 20177 12189 20211 12223
rect 7573 12121 7607 12155
rect 18613 12121 18647 12155
rect 5917 12053 5951 12087
rect 9229 12053 9263 12087
rect 10241 12053 10275 12087
rect 1777 11849 1811 11883
rect 3801 11849 3835 11883
rect 10149 11849 10183 11883
rect 15761 11849 15795 11883
rect 17509 11849 17543 11883
rect 18153 11849 18187 11883
rect 20269 11781 20303 11815
rect 2421 11713 2455 11747
rect 3341 11713 3375 11747
rect 4445 11713 4479 11747
rect 5457 11713 5491 11747
rect 7941 11713 7975 11747
rect 10793 11713 10827 11747
rect 11713 11713 11747 11747
rect 15301 11713 15335 11747
rect 18797 11713 18831 11747
rect 19993 11713 20027 11747
rect 3157 11645 3191 11679
rect 7205 11645 7239 11679
rect 8309 11645 8343 11679
rect 8576 11645 8610 11679
rect 10517 11645 10551 11679
rect 11529 11645 11563 11679
rect 13093 11645 13127 11679
rect 13360 11645 13394 11679
rect 15117 11645 15151 11679
rect 15945 11645 15979 11679
rect 16129 11645 16163 11679
rect 3249 11577 3283 11611
rect 7757 11577 7791 11611
rect 11621 11577 11655 11611
rect 15209 11577 15243 11611
rect 16396 11577 16430 11611
rect 18521 11577 18555 11611
rect 19809 11577 19843 11611
rect 20729 11713 20763 11747
rect 20453 11645 20487 11679
rect 2145 11509 2179 11543
rect 2237 11509 2271 11543
rect 2789 11509 2823 11543
rect 4169 11509 4203 11543
rect 4261 11509 4295 11543
rect 4813 11509 4847 11543
rect 5181 11509 5215 11543
rect 5273 11509 5307 11543
rect 7021 11509 7055 11543
rect 7297 11509 7331 11543
rect 7665 11509 7699 11543
rect 9689 11509 9723 11543
rect 10609 11509 10643 11543
rect 11161 11509 11195 11543
rect 14473 11509 14507 11543
rect 14749 11509 14783 11543
rect 18613 11509 18647 11543
rect 19441 11509 19475 11543
rect 19901 11509 19935 11543
rect 20269 11509 20303 11543
rect 2881 11305 2915 11339
rect 5733 11305 5767 11339
rect 6193 11305 6227 11339
rect 6745 11305 6779 11339
rect 8585 11305 8619 11339
rect 8953 11305 8987 11339
rect 10425 11305 10459 11339
rect 12725 11305 12759 11339
rect 13369 11305 13403 11339
rect 13737 11305 13771 11339
rect 17417 11305 17451 11339
rect 18429 11305 18463 11339
rect 18797 11305 18831 11339
rect 18889 11305 18923 11339
rect 19257 11305 19291 11339
rect 19901 11305 19935 11339
rect 7205 11237 7239 11271
rect 12817 11237 12851 11271
rect 1501 11169 1535 11203
rect 1768 11169 1802 11203
rect 4077 11169 4111 11203
rect 4344 11169 4378 11203
rect 6101 11169 6135 11203
rect 7113 11169 7147 11203
rect 9045 11169 9079 11203
rect 10793 11169 10827 11203
rect 12265 11169 12299 11203
rect 14565 11169 14599 11203
rect 15301 11169 15335 11203
rect 15557 11169 15591 11203
rect 17325 11169 17359 11203
rect 3157 11101 3191 11135
rect 6377 11101 6411 11135
rect 7297 11101 7331 11135
rect 9229 11101 9263 11135
rect 10885 11101 10919 11135
rect 10977 11101 11011 11135
rect 13001 11101 13035 11135
rect 13829 11101 13863 11135
rect 13921 11101 13955 11135
rect 17509 11101 17543 11135
rect 17969 11101 18003 11135
rect 18981 11101 19015 11135
rect 5457 11033 5491 11067
rect 12357 11033 12391 11067
rect 14381 11033 14415 11067
rect 16681 11033 16715 11067
rect 19809 11237 19843 11271
rect 19993 11101 20027 11135
rect 19441 11033 19475 11067
rect 12081 10965 12115 10999
rect 16957 10965 16991 10999
rect 19257 10965 19291 10999
rect 1777 10761 1811 10795
rect 3985 10761 4019 10795
rect 4905 10761 4939 10795
rect 2329 10625 2363 10659
rect 3341 10625 3375 10659
rect 4629 10625 4663 10659
rect 3157 10557 3191 10591
rect 8401 10761 8435 10795
rect 12449 10761 12483 10795
rect 14933 10761 14967 10795
rect 16129 10761 16163 10795
rect 18521 10761 18555 10795
rect 19533 10761 19567 10795
rect 5641 10625 5675 10659
rect 7941 10625 7975 10659
rect 8125 10625 8159 10659
rect 9229 10625 9263 10659
rect 9321 10625 9355 10659
rect 12909 10625 12943 10659
rect 13001 10625 13035 10659
rect 14013 10625 14047 10659
rect 15485 10625 15519 10659
rect 16589 10625 16623 10659
rect 16681 10625 16715 10659
rect 19073 10625 19107 10659
rect 20085 10625 20119 10659
rect 8401 10557 8435 10591
rect 8677 10557 8711 10591
rect 10701 10557 10735 10591
rect 10968 10557 11002 10591
rect 16497 10557 16531 10591
rect 20545 10557 20579 10591
rect 2145 10489 2179 10523
rect 4445 10489 4479 10523
rect 4905 10489 4939 10523
rect 5457 10489 5491 10523
rect 12817 10489 12851 10523
rect 15301 10489 15335 10523
rect 18981 10489 19015 10523
rect 19901 10489 19935 10523
rect 20821 10489 20855 10523
rect 2237 10421 2271 10455
rect 2789 10421 2823 10455
rect 3249 10421 3283 10455
rect 4353 10421 4387 10455
rect 4997 10421 5031 10455
rect 5365 10421 5399 10455
rect 6009 10421 6043 10455
rect 7481 10421 7515 10455
rect 7849 10421 7883 10455
rect 8493 10421 8527 10455
rect 8769 10421 8803 10455
rect 9137 10421 9171 10455
rect 12081 10421 12115 10455
rect 13461 10421 13495 10455
rect 13829 10421 13863 10455
rect 13921 10421 13955 10455
rect 15393 10421 15427 10455
rect 18889 10421 18923 10455
rect 19993 10421 20027 10455
rect 1961 10217 1995 10251
rect 3433 10217 3467 10251
rect 4169 10217 4203 10251
rect 4537 10217 4571 10251
rect 6929 10217 6963 10251
rect 7849 10217 7883 10251
rect 9689 10217 9723 10251
rect 10057 10217 10091 10251
rect 13093 10217 13127 10251
rect 13645 10217 13679 10251
rect 14013 10217 14047 10251
rect 17693 10217 17727 10251
rect 18705 10217 18739 10251
rect 19165 10217 19199 10251
rect 4629 10149 4663 10183
rect 1409 10081 1443 10115
rect 2329 10081 2363 10115
rect 2421 10081 2455 10115
rect 3341 10081 3375 10115
rect 5365 10081 5399 10115
rect 5549 10081 5583 10115
rect 5816 10081 5850 10115
rect 11612 10149 11646 10183
rect 18245 10149 18279 10183
rect 8197 10081 8231 10115
rect 10149 10081 10183 10115
rect 14105 10081 14139 10115
rect 15117 10081 15151 10115
rect 15669 10081 15703 10115
rect 16569 10081 16603 10115
rect 17969 10081 18003 10115
rect 19073 10081 19107 10115
rect 20085 10081 20119 10115
rect 2605 10013 2639 10047
rect 3617 10013 3651 10047
rect 4813 10013 4847 10047
rect 7849 10013 7883 10047
rect 7941 10013 7975 10047
rect 10241 10013 10275 10047
rect 11345 10013 11379 10047
rect 14197 10013 14231 10047
rect 15761 10013 15795 10047
rect 15945 10013 15979 10047
rect 16313 10013 16347 10047
rect 19257 10013 19291 10047
rect 20177 10013 20211 10047
rect 20361 10013 20395 10047
rect 1593 9945 1627 9979
rect 2973 9945 3007 9979
rect 14933 9945 14967 9979
rect 5181 9877 5215 9911
rect 9321 9877 9355 9911
rect 12725 9877 12759 9911
rect 15301 9877 15335 9911
rect 19717 9877 19751 9911
rect 4445 9673 4479 9707
rect 16221 9673 16255 9707
rect 4169 9605 4203 9639
rect 18245 9605 18279 9639
rect 19533 9605 19567 9639
rect 1961 9537 1995 9571
rect 5089 9537 5123 9571
rect 6101 9537 6135 9571
rect 7297 9537 7331 9571
rect 7757 9537 7791 9571
rect 12909 9537 12943 9571
rect 13093 9537 13127 9571
rect 17049 9537 17083 9571
rect 18705 9537 18739 9571
rect 18889 9537 18923 9571
rect 20453 9537 20487 9571
rect 1777 9469 1811 9503
rect 2789 9469 2823 9503
rect 4813 9469 4847 9503
rect 5917 9469 5951 9503
rect 9873 9469 9907 9503
rect 10140 9469 10174 9503
rect 14841 9469 14875 9503
rect 18613 9469 18647 9503
rect 19349 9469 19383 9503
rect 3034 9401 3068 9435
rect 8024 9401 8058 9435
rect 12817 9401 12851 9435
rect 15086 9401 15120 9435
rect 16865 9401 16899 9435
rect 20361 9401 20395 9435
rect 4905 9333 4939 9367
rect 5457 9333 5491 9367
rect 5825 9333 5859 9367
rect 9137 9333 9171 9367
rect 11253 9333 11287 9367
rect 12449 9333 12483 9367
rect 14381 9333 14415 9367
rect 16497 9333 16531 9367
rect 16957 9333 16991 9367
rect 19901 9333 19935 9367
rect 20269 9333 20303 9367
rect 2237 9129 2271 9163
rect 4537 9129 4571 9163
rect 5457 9129 5491 9163
rect 5549 9129 5583 9163
rect 7297 9129 7331 9163
rect 7757 9129 7791 9163
rect 8309 9129 8343 9163
rect 8677 9129 8711 9163
rect 8769 9129 8803 9163
rect 10885 9129 10919 9163
rect 14933 9129 14967 9163
rect 15025 9129 15059 9163
rect 15301 9129 15335 9163
rect 15761 9129 15795 9163
rect 16313 9129 16347 9163
rect 16681 9129 16715 9163
rect 19625 9129 19659 9163
rect 19809 9129 19843 9163
rect 20913 9129 20947 9163
rect 1501 8993 1535 9027
rect 2605 8993 2639 9027
rect 4905 8993 4939 9027
rect 7665 9061 7699 9095
rect 10057 9061 10091 9095
rect 10149 9061 10183 9095
rect 11253 9061 11287 9095
rect 5917 8993 5951 9027
rect 12153 8993 12187 9027
rect 13820 8993 13854 9027
rect 15669 9061 15703 9095
rect 16773 8993 16807 9027
rect 18420 8993 18454 9027
rect 20177 8993 20211 9027
rect 1685 8925 1719 8959
rect 2697 8925 2731 8959
rect 2881 8925 2915 8959
rect 4997 8925 5031 8959
rect 5089 8925 5123 8959
rect 5457 8925 5491 8959
rect 6009 8925 6043 8959
rect 6193 8925 6227 8959
rect 7849 8925 7883 8959
rect 8953 8925 8987 8959
rect 10241 8925 10275 8959
rect 11345 8925 11379 8959
rect 11529 8925 11563 8959
rect 11897 8925 11931 8959
rect 13553 8925 13587 8959
rect 15025 8925 15059 8959
rect 15853 8925 15887 8959
rect 16957 8925 16991 8959
rect 18153 8925 18187 8959
rect 19625 8925 19659 8959
rect 20269 8925 20303 8959
rect 20361 8925 20395 8959
rect 9689 8857 9723 8891
rect 13277 8857 13311 8891
rect 19533 8789 19567 8823
rect 2973 8585 3007 8619
rect 3249 8585 3283 8619
rect 14841 8585 14875 8619
rect 16957 8585 16991 8619
rect 19441 8585 19475 8619
rect 19717 8585 19751 8619
rect 20913 8585 20947 8619
rect 7665 8517 7699 8551
rect 10057 8517 10091 8551
rect 11345 8517 11379 8551
rect 3709 8449 3743 8483
rect 3893 8449 3927 8483
rect 4721 8449 4755 8483
rect 4905 8449 4939 8483
rect 5917 8449 5951 8483
rect 7573 8449 7607 8483
rect 8217 8449 8251 8483
rect 10793 8449 10827 8483
rect 10885 8449 10919 8483
rect 11897 8449 11931 8483
rect 12449 8449 12483 8483
rect 15393 8449 15427 8483
rect 16497 8449 16531 8483
rect 17601 8449 17635 8483
rect 20177 8449 20211 8483
rect 20269 8449 20303 8483
rect 1593 8381 1627 8415
rect 4169 8381 4203 8415
rect 1860 8313 1894 8347
rect 8677 8381 8711 8415
rect 11713 8381 11747 8415
rect 15301 8381 15335 8415
rect 16221 8381 16255 8415
rect 18068 8381 18102 8415
rect 20085 8381 20119 8415
rect 20729 8381 20763 8415
rect 4629 8313 4663 8347
rect 5641 8313 5675 8347
rect 5733 8313 5767 8347
rect 7573 8313 7607 8347
rect 8033 8313 8067 8347
rect 8125 8313 8159 8347
rect 8922 8313 8956 8347
rect 11805 8313 11839 8347
rect 12716 8313 12750 8347
rect 15209 8313 15243 8347
rect 16313 8313 16347 8347
rect 17325 8313 17359 8347
rect 18328 8313 18362 8347
rect 3617 8245 3651 8279
rect 4169 8245 4203 8279
rect 4261 8245 4295 8279
rect 5273 8245 5307 8279
rect 10333 8245 10367 8279
rect 10701 8245 10735 8279
rect 13829 8245 13863 8279
rect 15853 8245 15887 8279
rect 17417 8245 17451 8279
rect 4077 8041 4111 8075
rect 4537 8041 4571 8075
rect 5641 8041 5675 8075
rect 7113 8041 7147 8075
rect 7757 8041 7791 8075
rect 9229 8041 9263 8075
rect 10425 8041 10459 8075
rect 10885 8041 10919 8075
rect 12357 8041 12391 8075
rect 12725 8041 12759 8075
rect 18429 8041 18463 8075
rect 19441 8041 19475 8075
rect 19809 8041 19843 8075
rect 2596 7905 2630 7939
rect 4445 7905 4479 7939
rect 6000 7905 6034 7939
rect 12817 7973 12851 8007
rect 8116 7905 8150 7939
rect 10793 7905 10827 7939
rect 17040 7905 17074 7939
rect 18797 7905 18831 7939
rect 18889 7905 18923 7939
rect 2329 7837 2363 7871
rect 4721 7837 4755 7871
rect 5641 7837 5675 7871
rect 5733 7837 5767 7871
rect 7757 7837 7791 7871
rect 7849 7837 7883 7871
rect 10977 7837 11011 7871
rect 12909 7837 12943 7871
rect 16773 7837 16807 7871
rect 18981 7837 19015 7871
rect 19901 7837 19935 7871
rect 19993 7837 20027 7871
rect 3709 7769 3743 7803
rect 18153 7769 18187 7803
rect 2513 7497 2547 7531
rect 6377 7497 6411 7531
rect 8309 7497 8343 7531
rect 8585 7497 8619 7531
rect 16313 7497 16347 7531
rect 19809 7497 19843 7531
rect 3157 7361 3191 7395
rect 4169 7361 4203 7395
rect 4997 7361 5031 7395
rect 6929 7361 6963 7395
rect 9137 7361 9171 7395
rect 16957 7361 16991 7395
rect 20361 7361 20395 7395
rect 5264 7293 5298 7327
rect 16773 7293 16807 7327
rect 19073 7293 19107 7327
rect 20177 7293 20211 7327
rect 2881 7225 2915 7259
rect 3985 7225 4019 7259
rect 7174 7225 7208 7259
rect 8953 7225 8987 7259
rect 19349 7225 19383 7259
rect 2973 7157 3007 7191
rect 3525 7157 3559 7191
rect 3893 7157 3927 7191
rect 4537 7157 4571 7191
rect 9045 7157 9079 7191
rect 16681 7157 16715 7191
rect 20269 7157 20303 7191
rect 3341 6953 3375 6987
rect 6561 6953 6595 6987
rect 17969 6953 18003 6987
rect 7573 6885 7607 6919
rect 1593 6817 1627 6851
rect 1860 6817 1894 6851
rect 4537 6817 4571 6851
rect 5549 6817 5583 6851
rect 6653 6817 6687 6851
rect 7665 6817 7699 6851
rect 16856 6817 16890 6851
rect 19340 6817 19374 6851
rect 4629 6749 4663 6783
rect 4813 6749 4847 6783
rect 5641 6749 5675 6783
rect 5825 6749 5859 6783
rect 6745 6749 6779 6783
rect 7849 6749 7883 6783
rect 16589 6749 16623 6783
rect 19073 6749 19107 6783
rect 20913 6749 20947 6783
rect 2973 6681 3007 6715
rect 4169 6681 4203 6715
rect 6193 6681 6227 6715
rect 5181 6613 5215 6647
rect 7205 6613 7239 6647
rect 20453 6613 20487 6647
rect 2973 6409 3007 6443
rect 4997 6409 5031 6443
rect 20637 6409 20671 6443
rect 3617 6273 3651 6307
rect 5549 6273 5583 6307
rect 19257 6273 19291 6307
rect 5365 6205 5399 6239
rect 19524 6205 19558 6239
rect 3433 6137 3467 6171
rect 3341 6069 3375 6103
rect 5457 6069 5491 6103
rect 19809 5865 19843 5899
rect 20177 5865 20211 5899
rect 20269 5661 20303 5695
rect 20361 5661 20395 5695
rect 20085 5321 20119 5355
rect 20637 5185 20671 5219
rect 19901 4981 19935 5015
rect 20453 4981 20487 5015
rect 20545 4981 20579 5015
rect 15025 3009 15059 3043
rect 15301 3009 15335 3043
rect 4629 2941 4663 2975
rect 4905 2941 4939 2975
rect 5549 2941 5583 2975
rect 5825 2873 5859 2907
rect 15117 2941 15151 2975
rect 15025 2805 15059 2839
<< metal1 >>
rect 3878 20952 3884 21004
rect 3936 20992 3942 21004
rect 5534 20992 5540 21004
rect 3936 20964 5540 20992
rect 3936 20952 3942 20964
rect 5534 20952 5540 20964
rect 5592 20952 5598 21004
rect 2222 20612 2228 20664
rect 2280 20652 2286 20664
rect 8662 20652 8668 20664
rect 2280 20624 8668 20652
rect 2280 20612 2286 20624
rect 8662 20612 8668 20624
rect 8720 20612 8726 20664
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 1949 20043 2007 20049
rect 1949 20009 1961 20043
rect 1995 20040 2007 20043
rect 2774 20040 2780 20052
rect 1995 20012 2780 20040
rect 1995 20009 2007 20012
rect 1949 20003 2007 20009
rect 2774 20000 2780 20012
rect 2832 20000 2838 20052
rect 8662 20040 8668 20052
rect 8623 20012 8668 20040
rect 8662 20000 8668 20012
rect 8720 20000 8726 20052
rect 10226 20000 10232 20052
rect 10284 20040 10290 20052
rect 10321 20043 10379 20049
rect 10321 20040 10333 20043
rect 10284 20012 10333 20040
rect 10284 20000 10290 20012
rect 10321 20009 10333 20012
rect 10367 20009 10379 20043
rect 10321 20003 10379 20009
rect 11606 20000 11612 20052
rect 11664 20040 11670 20052
rect 12250 20040 12256 20052
rect 11664 20012 12256 20040
rect 11664 20000 11670 20012
rect 12250 20000 12256 20012
rect 12308 20000 12314 20052
rect 14461 20043 14519 20049
rect 14461 20009 14473 20043
rect 14507 20009 14519 20043
rect 14461 20003 14519 20009
rect 16025 20043 16083 20049
rect 16025 20009 16037 20043
rect 16071 20040 16083 20043
rect 16666 20040 16672 20052
rect 16071 20012 16672 20040
rect 16071 20009 16083 20012
rect 16025 20003 16083 20009
rect 14476 19972 14504 20003
rect 16666 20000 16672 20012
rect 16724 20000 16730 20052
rect 17494 20000 17500 20052
rect 17552 20040 17558 20052
rect 18509 20043 18567 20049
rect 18509 20040 18521 20043
rect 17552 20012 18521 20040
rect 17552 20000 17558 20012
rect 18509 20009 18521 20012
rect 18555 20009 18567 20043
rect 19610 20040 19616 20052
rect 19571 20012 19616 20040
rect 18509 20003 18567 20009
rect 19610 20000 19616 20012
rect 19668 20000 19674 20052
rect 20162 20040 20168 20052
rect 20123 20012 20168 20040
rect 20162 20000 20168 20012
rect 20220 20000 20226 20052
rect 20622 20000 20628 20052
rect 20680 20040 20686 20052
rect 20717 20043 20775 20049
rect 20717 20040 20729 20043
rect 20680 20012 20729 20040
rect 20680 20000 20686 20012
rect 20717 20009 20729 20012
rect 20763 20009 20775 20043
rect 20717 20003 20775 20009
rect 17862 19972 17868 19984
rect 14476 19944 17868 19972
rect 17862 19932 17868 19944
rect 17920 19932 17926 19984
rect 1765 19907 1823 19913
rect 1765 19873 1777 19907
rect 1811 19873 1823 19907
rect 2314 19904 2320 19916
rect 2275 19876 2320 19904
rect 1765 19867 1823 19873
rect 1780 19768 1808 19867
rect 2314 19864 2320 19876
rect 2372 19864 2378 19916
rect 2866 19904 2872 19916
rect 2827 19876 2872 19904
rect 2866 19864 2872 19876
rect 2924 19864 2930 19916
rect 7282 19864 7288 19916
rect 7340 19904 7346 19916
rect 7653 19907 7711 19913
rect 7653 19904 7665 19907
rect 7340 19876 7665 19904
rect 7340 19864 7346 19876
rect 7653 19873 7665 19876
rect 7699 19873 7711 19907
rect 7653 19867 7711 19873
rect 8478 19864 8484 19916
rect 8536 19904 8542 19916
rect 8573 19907 8631 19913
rect 8573 19904 8585 19907
rect 8536 19876 8585 19904
rect 8536 19864 8542 19876
rect 8573 19873 8585 19876
rect 8619 19873 8631 19907
rect 8573 19867 8631 19873
rect 8662 19864 8668 19916
rect 8720 19904 8726 19916
rect 9217 19907 9275 19913
rect 9217 19904 9229 19907
rect 8720 19876 9229 19904
rect 8720 19864 8726 19876
rect 9217 19873 9229 19876
rect 9263 19873 9275 19907
rect 9217 19867 9275 19873
rect 10134 19864 10140 19916
rect 10192 19904 10198 19916
rect 10229 19907 10287 19913
rect 10229 19904 10241 19907
rect 10192 19876 10241 19904
rect 10192 19864 10198 19876
rect 10229 19873 10241 19876
rect 10275 19873 10287 19907
rect 10229 19867 10287 19873
rect 11146 19864 11152 19916
rect 11204 19904 11210 19916
rect 11333 19907 11391 19913
rect 11333 19904 11345 19907
rect 11204 19876 11345 19904
rect 11204 19864 11210 19876
rect 11333 19873 11345 19876
rect 11379 19873 11391 19907
rect 11333 19867 11391 19873
rect 11425 19907 11483 19913
rect 11425 19873 11437 19907
rect 11471 19904 11483 19907
rect 11606 19904 11612 19916
rect 11471 19876 11612 19904
rect 11471 19873 11483 19876
rect 11425 19867 11483 19873
rect 11606 19864 11612 19876
rect 11664 19864 11670 19916
rect 11977 19907 12035 19913
rect 11977 19873 11989 19907
rect 12023 19904 12035 19907
rect 12066 19904 12072 19916
rect 12023 19876 12072 19904
rect 12023 19873 12035 19876
rect 11977 19867 12035 19873
rect 12066 19864 12072 19876
rect 12124 19864 12130 19916
rect 13262 19904 13268 19916
rect 13223 19876 13268 19904
rect 13262 19864 13268 19876
rect 13320 19864 13326 19916
rect 14274 19904 14280 19916
rect 14235 19876 14280 19904
rect 14274 19864 14280 19876
rect 14332 19864 14338 19916
rect 14829 19907 14887 19913
rect 14829 19873 14841 19907
rect 14875 19873 14887 19907
rect 14829 19867 14887 19873
rect 3050 19796 3056 19848
rect 3108 19796 3114 19848
rect 8754 19796 8760 19848
rect 8812 19836 8818 19848
rect 10410 19836 10416 19848
rect 8812 19808 8857 19836
rect 10371 19808 10416 19836
rect 8812 19796 8818 19808
rect 10410 19796 10416 19808
rect 10468 19796 10474 19848
rect 11517 19839 11575 19845
rect 11517 19805 11529 19839
rect 11563 19836 11575 19839
rect 11882 19836 11888 19848
rect 11563 19808 11888 19836
rect 11563 19805 11575 19808
rect 11517 19799 11575 19805
rect 11882 19796 11888 19808
rect 11940 19796 11946 19848
rect 13354 19836 13360 19848
rect 13315 19808 13360 19836
rect 13354 19796 13360 19808
rect 13412 19796 13418 19848
rect 13538 19836 13544 19848
rect 13499 19808 13544 19836
rect 13538 19796 13544 19808
rect 13596 19796 13602 19848
rect 2406 19768 2412 19780
rect 1780 19740 2412 19768
rect 2406 19728 2412 19740
rect 2464 19728 2470 19780
rect 2501 19771 2559 19777
rect 2501 19737 2513 19771
rect 2547 19768 2559 19771
rect 3068 19768 3096 19796
rect 2547 19740 3096 19768
rect 7837 19771 7895 19777
rect 2547 19737 2559 19740
rect 2501 19731 2559 19737
rect 7837 19737 7849 19771
rect 7883 19768 7895 19771
rect 11790 19768 11796 19780
rect 7883 19740 11796 19768
rect 7883 19737 7895 19740
rect 7837 19731 7895 19737
rect 11790 19728 11796 19740
rect 11848 19728 11854 19780
rect 13170 19728 13176 19780
rect 13228 19768 13234 19780
rect 14844 19768 14872 19867
rect 15286 19864 15292 19916
rect 15344 19904 15350 19916
rect 15841 19907 15899 19913
rect 15841 19904 15853 19907
rect 15344 19876 15853 19904
rect 15344 19864 15350 19876
rect 15841 19873 15853 19876
rect 15887 19873 15899 19907
rect 17218 19904 17224 19916
rect 17179 19876 17224 19904
rect 15841 19867 15899 19873
rect 17218 19864 17224 19876
rect 17276 19864 17282 19916
rect 18325 19907 18383 19913
rect 18325 19873 18337 19907
rect 18371 19904 18383 19907
rect 18598 19904 18604 19916
rect 18371 19876 18604 19904
rect 18371 19873 18383 19876
rect 18325 19867 18383 19873
rect 18598 19864 18604 19876
rect 18656 19864 18662 19916
rect 18690 19864 18696 19916
rect 18748 19904 18754 19916
rect 18877 19907 18935 19913
rect 18877 19904 18889 19907
rect 18748 19876 18889 19904
rect 18748 19864 18754 19876
rect 18877 19873 18889 19876
rect 18923 19873 18935 19907
rect 19426 19904 19432 19916
rect 19387 19876 19432 19904
rect 18877 19867 18935 19873
rect 19426 19864 19432 19876
rect 19484 19864 19490 19916
rect 19610 19864 19616 19916
rect 19668 19904 19674 19916
rect 19981 19907 20039 19913
rect 19981 19904 19993 19907
rect 19668 19876 19993 19904
rect 19668 19864 19674 19876
rect 19981 19873 19993 19876
rect 20027 19873 20039 19907
rect 19981 19867 20039 19873
rect 20533 19907 20591 19913
rect 20533 19873 20545 19907
rect 20579 19873 20591 19907
rect 20533 19867 20591 19873
rect 17313 19839 17371 19845
rect 17313 19836 17325 19839
rect 13228 19740 14872 19768
rect 14936 19808 17325 19836
rect 13228 19728 13234 19740
rect 3050 19700 3056 19712
rect 3011 19672 3056 19700
rect 3050 19660 3056 19672
rect 3108 19660 3114 19712
rect 8205 19703 8263 19709
rect 8205 19669 8217 19703
rect 8251 19700 8263 19703
rect 8938 19700 8944 19712
rect 8251 19672 8944 19700
rect 8251 19669 8263 19672
rect 8205 19663 8263 19669
rect 8938 19660 8944 19672
rect 8996 19660 9002 19712
rect 9398 19660 9404 19712
rect 9456 19700 9462 19712
rect 9861 19703 9919 19709
rect 9861 19700 9873 19703
rect 9456 19672 9873 19700
rect 9456 19660 9462 19672
rect 9861 19669 9873 19672
rect 9907 19669 9919 19703
rect 9861 19663 9919 19669
rect 10965 19703 11023 19709
rect 10965 19669 10977 19703
rect 11011 19700 11023 19703
rect 11054 19700 11060 19712
rect 11011 19672 11060 19700
rect 11011 19669 11023 19672
rect 10965 19663 11023 19669
rect 11054 19660 11060 19672
rect 11112 19660 11118 19712
rect 12158 19700 12164 19712
rect 12119 19672 12164 19700
rect 12158 19660 12164 19672
rect 12216 19660 12222 19712
rect 12897 19703 12955 19709
rect 12897 19669 12909 19703
rect 12943 19700 12955 19703
rect 14090 19700 14096 19712
rect 12943 19672 14096 19700
rect 12943 19669 12955 19672
rect 12897 19663 12955 19669
rect 14090 19660 14096 19672
rect 14148 19660 14154 19712
rect 14182 19660 14188 19712
rect 14240 19700 14246 19712
rect 14936 19700 14964 19808
rect 17313 19805 17325 19808
rect 17359 19805 17371 19839
rect 17313 19799 17371 19805
rect 17402 19796 17408 19848
rect 17460 19836 17466 19848
rect 17460 19808 17505 19836
rect 17460 19796 17466 19808
rect 19334 19796 19340 19848
rect 19392 19836 19398 19848
rect 20548 19836 20576 19867
rect 19392 19808 20576 19836
rect 19392 19796 19398 19808
rect 15013 19771 15071 19777
rect 15013 19737 15025 19771
rect 15059 19768 15071 19771
rect 17034 19768 17040 19780
rect 15059 19740 17040 19768
rect 15059 19737 15071 19740
rect 15013 19731 15071 19737
rect 17034 19728 17040 19740
rect 17092 19728 17098 19780
rect 19058 19768 19064 19780
rect 19019 19740 19064 19768
rect 19058 19728 19064 19740
rect 19116 19728 19122 19780
rect 16850 19700 16856 19712
rect 14240 19672 14964 19700
rect 16811 19672 16856 19700
rect 14240 19660 14246 19672
rect 16850 19660 16856 19672
rect 16908 19660 16914 19712
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 1946 19496 1952 19508
rect 1907 19468 1952 19496
rect 1946 19456 1952 19468
rect 2004 19456 2010 19508
rect 3418 19496 3424 19508
rect 3379 19468 3424 19496
rect 3418 19456 3424 19468
rect 3476 19456 3482 19508
rect 8481 19499 8539 19505
rect 5368 19468 8432 19496
rect 5368 19440 5396 19468
rect 2314 19388 2320 19440
rect 2372 19428 2378 19440
rect 5350 19428 5356 19440
rect 2372 19400 5356 19428
rect 2372 19388 2378 19400
rect 5350 19388 5356 19400
rect 5408 19388 5414 19440
rect 8404 19360 8432 19468
rect 8481 19465 8493 19499
rect 8527 19496 8539 19499
rect 8754 19496 8760 19508
rect 8527 19468 8760 19496
rect 8527 19465 8539 19468
rect 8481 19459 8539 19465
rect 8754 19456 8760 19468
rect 8812 19456 8818 19508
rect 8846 19456 8852 19508
rect 8904 19496 8910 19508
rect 12710 19496 12716 19508
rect 8904 19468 12716 19496
rect 8904 19456 8910 19468
rect 12710 19456 12716 19468
rect 12768 19456 12774 19508
rect 8570 19388 8576 19440
rect 8628 19428 8634 19440
rect 9582 19428 9588 19440
rect 8628 19400 9588 19428
rect 8628 19388 8634 19400
rect 9582 19388 9588 19400
rect 9640 19388 9646 19440
rect 17218 19388 17224 19440
rect 17276 19428 17282 19440
rect 18046 19428 18052 19440
rect 17276 19400 18052 19428
rect 17276 19388 17282 19400
rect 18046 19388 18052 19400
rect 18104 19388 18110 19440
rect 8846 19360 8852 19372
rect 8404 19332 8852 19360
rect 8846 19320 8852 19332
rect 8904 19320 8910 19372
rect 8938 19320 8944 19372
rect 8996 19360 9002 19372
rect 9401 19363 9459 19369
rect 9401 19360 9413 19363
rect 8996 19332 9260 19360
rect 8996 19320 9002 19332
rect 1762 19292 1768 19304
rect 1723 19264 1768 19292
rect 1762 19252 1768 19264
rect 1820 19252 1826 19304
rect 2317 19295 2375 19301
rect 2317 19261 2329 19295
rect 2363 19292 2375 19295
rect 2498 19292 2504 19304
rect 2363 19264 2504 19292
rect 2363 19261 2375 19264
rect 2317 19255 2375 19261
rect 2498 19252 2504 19264
rect 2556 19252 2562 19304
rect 3237 19295 3295 19301
rect 3237 19261 3249 19295
rect 3283 19292 3295 19295
rect 3418 19292 3424 19304
rect 3283 19264 3424 19292
rect 3283 19261 3295 19264
rect 3237 19255 3295 19261
rect 3418 19252 3424 19264
rect 3476 19292 3482 19304
rect 3786 19292 3792 19304
rect 3476 19264 3792 19292
rect 3476 19252 3482 19264
rect 3786 19252 3792 19264
rect 3844 19252 3850 19304
rect 3970 19292 3976 19304
rect 3931 19264 3976 19292
rect 3970 19252 3976 19264
rect 4028 19252 4034 19304
rect 5902 19292 5908 19304
rect 5863 19264 5908 19292
rect 5902 19252 5908 19264
rect 5960 19252 5966 19304
rect 7098 19292 7104 19304
rect 7059 19264 7104 19292
rect 7098 19252 7104 19264
rect 7156 19252 7162 19304
rect 7742 19252 7748 19304
rect 7800 19292 7806 19304
rect 9122 19292 9128 19304
rect 7800 19264 9128 19292
rect 7800 19252 7806 19264
rect 9122 19252 9128 19264
rect 9180 19252 9186 19304
rect 9232 19301 9260 19332
rect 9324 19332 9413 19360
rect 9324 19304 9352 19332
rect 9401 19329 9413 19332
rect 9447 19329 9459 19363
rect 14274 19360 14280 19372
rect 14235 19332 14280 19360
rect 9401 19323 9459 19329
rect 14274 19320 14280 19332
rect 14332 19320 14338 19372
rect 15470 19360 15476 19372
rect 15431 19332 15476 19360
rect 15470 19320 15476 19332
rect 15528 19320 15534 19372
rect 16850 19320 16856 19372
rect 16908 19360 16914 19372
rect 17405 19363 17463 19369
rect 17405 19360 17417 19363
rect 16908 19332 17417 19360
rect 16908 19320 16914 19332
rect 17405 19329 17417 19332
rect 17451 19329 17463 19363
rect 17405 19323 17463 19329
rect 17589 19363 17647 19369
rect 17589 19329 17601 19363
rect 17635 19360 17647 19363
rect 18506 19360 18512 19372
rect 17635 19332 18512 19360
rect 17635 19329 17647 19332
rect 17589 19323 17647 19329
rect 18506 19320 18512 19332
rect 18564 19320 18570 19372
rect 19058 19320 19064 19372
rect 19116 19360 19122 19372
rect 19116 19332 19288 19360
rect 19116 19320 19122 19332
rect 9217 19295 9275 19301
rect 9217 19261 9229 19295
rect 9263 19261 9275 19295
rect 9217 19255 9275 19261
rect 9306 19252 9312 19304
rect 9364 19252 9370 19304
rect 9582 19252 9588 19304
rect 9640 19292 9646 19304
rect 10321 19295 10379 19301
rect 10321 19292 10333 19295
rect 9640 19264 10333 19292
rect 9640 19252 9646 19264
rect 10321 19261 10333 19264
rect 10367 19261 10379 19295
rect 10321 19255 10379 19261
rect 10588 19295 10646 19301
rect 10588 19261 10600 19295
rect 10634 19292 10646 19295
rect 11698 19292 11704 19304
rect 10634 19264 11704 19292
rect 10634 19261 10646 19264
rect 10588 19255 10646 19261
rect 11698 19252 11704 19264
rect 11756 19252 11762 19304
rect 12437 19295 12495 19301
rect 12437 19261 12449 19295
rect 12483 19292 12495 19295
rect 14090 19292 14096 19304
rect 12483 19264 12848 19292
rect 14051 19264 14096 19292
rect 12483 19261 12495 19264
rect 12437 19255 12495 19261
rect 12820 19236 12848 19264
rect 14090 19252 14096 19264
rect 14148 19252 14154 19304
rect 15841 19295 15899 19301
rect 15841 19292 15853 19295
rect 14844 19264 15853 19292
rect 198 19184 204 19236
rect 256 19224 262 19236
rect 2866 19224 2872 19236
rect 256 19196 2872 19224
rect 256 19184 262 19196
rect 2866 19184 2872 19196
rect 2924 19184 2930 19236
rect 4617 19227 4675 19233
rect 4617 19193 4629 19227
rect 4663 19224 4675 19227
rect 6546 19224 6552 19236
rect 4663 19196 6552 19224
rect 4663 19193 4675 19196
rect 4617 19187 4675 19193
rect 6546 19184 6552 19196
rect 6604 19184 6610 19236
rect 7368 19227 7426 19233
rect 7368 19193 7380 19227
rect 7414 19224 7426 19227
rect 11882 19224 11888 19236
rect 7414 19196 11888 19224
rect 7414 19193 7426 19196
rect 7368 19187 7426 19193
rect 2501 19159 2559 19165
rect 2501 19125 2513 19159
rect 2547 19156 2559 19159
rect 2958 19156 2964 19168
rect 2547 19128 2964 19156
rect 2547 19125 2559 19128
rect 2501 19119 2559 19125
rect 2958 19116 2964 19128
rect 3016 19116 3022 19168
rect 5534 19116 5540 19168
rect 5592 19156 5598 19168
rect 6089 19159 6147 19165
rect 6089 19156 6101 19159
rect 5592 19128 6101 19156
rect 5592 19116 5598 19128
rect 6089 19125 6101 19128
rect 6135 19125 6147 19159
rect 6089 19119 6147 19125
rect 6454 19116 6460 19168
rect 6512 19156 6518 19168
rect 8478 19156 8484 19168
rect 6512 19128 8484 19156
rect 6512 19116 6518 19128
rect 8478 19116 8484 19128
rect 8536 19116 8542 19168
rect 8757 19159 8815 19165
rect 8757 19125 8769 19159
rect 8803 19156 8815 19159
rect 8846 19156 8852 19168
rect 8803 19128 8852 19156
rect 8803 19125 8815 19128
rect 8757 19119 8815 19125
rect 8846 19116 8852 19128
rect 8904 19116 8910 19168
rect 9122 19156 9128 19168
rect 9083 19128 9128 19156
rect 9122 19116 9128 19128
rect 9180 19116 9186 19168
rect 9214 19116 9220 19168
rect 9272 19156 9278 19168
rect 10502 19156 10508 19168
rect 9272 19128 10508 19156
rect 9272 19116 9278 19128
rect 10502 19116 10508 19128
rect 10560 19116 10566 19168
rect 11716 19165 11744 19196
rect 11882 19184 11888 19196
rect 11940 19184 11946 19236
rect 12710 19233 12716 19236
rect 12704 19224 12716 19233
rect 12671 19196 12716 19224
rect 12704 19187 12716 19196
rect 12710 19184 12716 19187
rect 12768 19184 12774 19236
rect 12802 19184 12808 19236
rect 12860 19184 12866 19236
rect 14550 19224 14556 19236
rect 13464 19196 14556 19224
rect 11701 19159 11759 19165
rect 11701 19125 11713 19159
rect 11747 19125 11759 19159
rect 11701 19119 11759 19125
rect 11790 19116 11796 19168
rect 11848 19156 11854 19168
rect 13464 19156 13492 19196
rect 14550 19184 14556 19196
rect 14608 19184 14614 19236
rect 11848 19128 13492 19156
rect 11848 19116 11854 19128
rect 13538 19116 13544 19168
rect 13596 19156 13602 19168
rect 14844 19165 14872 19264
rect 15841 19261 15853 19264
rect 15887 19261 15899 19295
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 15841 19255 15899 19261
rect 16960 19264 18061 19292
rect 16117 19227 16175 19233
rect 16117 19193 16129 19227
rect 16163 19224 16175 19227
rect 16850 19224 16856 19236
rect 16163 19196 16856 19224
rect 16163 19193 16175 19196
rect 16117 19187 16175 19193
rect 16850 19184 16856 19196
rect 16908 19184 16914 19236
rect 13817 19159 13875 19165
rect 13817 19156 13829 19159
rect 13596 19128 13829 19156
rect 13596 19116 13602 19128
rect 13817 19125 13829 19128
rect 13863 19125 13875 19159
rect 13817 19119 13875 19125
rect 14829 19159 14887 19165
rect 14829 19125 14841 19159
rect 14875 19125 14887 19159
rect 15194 19156 15200 19168
rect 15155 19128 15200 19156
rect 14829 19119 14887 19125
rect 15194 19116 15200 19128
rect 15252 19116 15258 19168
rect 15289 19159 15347 19165
rect 15289 19125 15301 19159
rect 15335 19156 15347 19159
rect 15930 19156 15936 19168
rect 15335 19128 15936 19156
rect 15335 19125 15347 19128
rect 15289 19119 15347 19125
rect 15930 19116 15936 19128
rect 15988 19116 15994 19168
rect 16960 19165 16988 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18874 19292 18880 19304
rect 18835 19264 18880 19292
rect 18049 19255 18107 19261
rect 18874 19252 18880 19264
rect 18932 19252 18938 19304
rect 17494 19184 17500 19236
rect 17552 19224 17558 19236
rect 18325 19227 18383 19233
rect 18325 19224 18337 19227
rect 17552 19196 18337 19224
rect 17552 19184 17558 19196
rect 18325 19193 18337 19196
rect 18371 19193 18383 19227
rect 18325 19187 18383 19193
rect 19153 19227 19211 19233
rect 19153 19193 19165 19227
rect 19199 19193 19211 19227
rect 19260 19224 19288 19332
rect 19981 19295 20039 19301
rect 19981 19261 19993 19295
rect 20027 19292 20039 19295
rect 20346 19292 20352 19304
rect 20027 19264 20352 19292
rect 20027 19261 20039 19264
rect 19981 19255 20039 19261
rect 20346 19252 20352 19264
rect 20404 19252 20410 19304
rect 20530 19292 20536 19304
rect 20491 19264 20536 19292
rect 20530 19252 20536 19264
rect 20588 19252 20594 19304
rect 22094 19224 22100 19236
rect 19260 19196 22100 19224
rect 19153 19187 19211 19193
rect 16945 19159 17003 19165
rect 16945 19125 16957 19159
rect 16991 19125 17003 19159
rect 16945 19119 17003 19125
rect 17034 19116 17040 19168
rect 17092 19156 17098 19168
rect 17313 19159 17371 19165
rect 17313 19156 17325 19159
rect 17092 19128 17325 19156
rect 17092 19116 17098 19128
rect 17313 19125 17325 19128
rect 17359 19125 17371 19159
rect 17313 19119 17371 19125
rect 17770 19116 17776 19168
rect 17828 19156 17834 19168
rect 19168 19156 19196 19187
rect 22094 19184 22100 19196
rect 22152 19184 22158 19236
rect 17828 19128 19196 19156
rect 17828 19116 17834 19128
rect 19242 19116 19248 19168
rect 19300 19156 19306 19168
rect 20165 19159 20223 19165
rect 20165 19156 20177 19159
rect 19300 19128 20177 19156
rect 19300 19116 19306 19128
rect 20165 19125 20177 19128
rect 20211 19125 20223 19159
rect 20714 19156 20720 19168
rect 20675 19128 20720 19156
rect 20165 19119 20223 19125
rect 20714 19116 20720 19128
rect 20772 19116 20778 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 1578 18912 1584 18964
rect 1636 18952 1642 18964
rect 2041 18955 2099 18961
rect 2041 18952 2053 18955
rect 1636 18924 2053 18952
rect 1636 18912 1642 18924
rect 2041 18921 2053 18924
rect 2087 18921 2099 18955
rect 2041 18915 2099 18921
rect 2593 18955 2651 18961
rect 2593 18921 2605 18955
rect 2639 18952 2651 18955
rect 3234 18952 3240 18964
rect 2639 18924 3240 18952
rect 2639 18921 2651 18924
rect 2593 18915 2651 18921
rect 3234 18912 3240 18924
rect 3292 18912 3298 18964
rect 5537 18955 5595 18961
rect 5537 18921 5549 18955
rect 5583 18952 5595 18955
rect 9125 18955 9183 18961
rect 5583 18924 8984 18952
rect 5583 18921 5595 18924
rect 5537 18915 5595 18921
rect 1026 18844 1032 18896
rect 1084 18884 1090 18896
rect 5810 18884 5816 18896
rect 1084 18856 5816 18884
rect 1084 18844 1090 18856
rect 5810 18844 5816 18856
rect 5868 18844 5874 18896
rect 5902 18844 5908 18896
rect 5960 18884 5966 18896
rect 6549 18887 6607 18893
rect 6549 18884 6561 18887
rect 5960 18856 6561 18884
rect 5960 18844 5966 18856
rect 6549 18853 6561 18856
rect 6595 18853 6607 18887
rect 7282 18884 7288 18896
rect 7243 18856 7288 18884
rect 6549 18847 6607 18853
rect 7282 18844 7288 18856
rect 7340 18844 7346 18896
rect 8012 18887 8070 18893
rect 8012 18853 8024 18887
rect 8058 18884 8070 18887
rect 8754 18884 8760 18896
rect 8058 18856 8760 18884
rect 8058 18853 8070 18856
rect 8012 18847 8070 18853
rect 8754 18844 8760 18856
rect 8812 18844 8818 18896
rect 1857 18819 1915 18825
rect 1857 18785 1869 18819
rect 1903 18816 1915 18819
rect 2130 18816 2136 18828
rect 1903 18788 2136 18816
rect 1903 18785 1915 18788
rect 1857 18779 1915 18785
rect 2130 18776 2136 18788
rect 2188 18776 2194 18828
rect 2409 18819 2467 18825
rect 2409 18785 2421 18819
rect 2455 18785 2467 18819
rect 2409 18779 2467 18785
rect 2961 18819 3019 18825
rect 2961 18785 2973 18819
rect 3007 18816 3019 18819
rect 3694 18816 3700 18828
rect 3007 18788 3700 18816
rect 3007 18785 3019 18788
rect 2961 18779 3019 18785
rect 2424 18748 2452 18779
rect 3694 18776 3700 18788
rect 3752 18776 3758 18828
rect 4798 18776 4804 18828
rect 4856 18816 4862 18828
rect 5353 18819 5411 18825
rect 5353 18816 5365 18819
rect 4856 18788 5365 18816
rect 4856 18776 4862 18788
rect 5353 18785 5365 18788
rect 5399 18785 5411 18819
rect 6273 18819 6331 18825
rect 6273 18816 6285 18819
rect 5353 18779 5411 18785
rect 5920 18788 6285 18816
rect 5920 18760 5948 18788
rect 6273 18785 6285 18788
rect 6319 18785 6331 18819
rect 7006 18816 7012 18828
rect 6967 18788 7012 18816
rect 6273 18779 6331 18785
rect 7006 18776 7012 18788
rect 7064 18776 7070 18828
rect 7098 18776 7104 18828
rect 7156 18816 7162 18828
rect 7745 18819 7803 18825
rect 7745 18816 7757 18819
rect 7156 18788 7757 18816
rect 7156 18776 7162 18788
rect 7745 18785 7757 18788
rect 7791 18816 7803 18819
rect 8956 18816 8984 18924
rect 9125 18921 9137 18955
rect 9171 18952 9183 18955
rect 9306 18952 9312 18964
rect 9171 18924 9312 18952
rect 9171 18921 9183 18924
rect 9125 18915 9183 18921
rect 9306 18912 9312 18924
rect 9364 18912 9370 18964
rect 12161 18955 12219 18961
rect 12161 18921 12173 18955
rect 12207 18952 12219 18955
rect 13354 18952 13360 18964
rect 12207 18924 13360 18952
rect 12207 18921 12219 18924
rect 12161 18915 12219 18921
rect 13354 18912 13360 18924
rect 13412 18912 13418 18964
rect 16853 18955 16911 18961
rect 16853 18921 16865 18955
rect 16899 18921 16911 18955
rect 18506 18952 18512 18964
rect 18467 18924 18512 18952
rect 16853 18915 16911 18921
rect 9324 18884 9352 18912
rect 9922 18887 9980 18893
rect 9922 18884 9934 18887
rect 9324 18856 9934 18884
rect 9922 18853 9934 18856
rect 9968 18853 9980 18887
rect 9922 18847 9980 18853
rect 11701 18887 11759 18893
rect 11701 18853 11713 18887
rect 11747 18884 11759 18887
rect 12342 18884 12348 18896
rect 11747 18856 12348 18884
rect 11747 18853 11759 18856
rect 11701 18847 11759 18853
rect 12342 18844 12348 18856
rect 12400 18844 12406 18896
rect 12618 18884 12624 18896
rect 12579 18856 12624 18884
rect 12618 18844 12624 18856
rect 12676 18844 12682 18896
rect 13440 18887 13498 18893
rect 13440 18853 13452 18887
rect 13486 18884 13498 18887
rect 13538 18884 13544 18896
rect 13486 18856 13544 18884
rect 13486 18853 13498 18856
rect 13440 18847 13498 18853
rect 13538 18844 13544 18856
rect 13596 18844 13602 18896
rect 15470 18844 15476 18896
rect 15528 18884 15534 18896
rect 15718 18887 15776 18893
rect 15718 18884 15730 18887
rect 15528 18856 15730 18884
rect 15528 18844 15534 18856
rect 15718 18853 15730 18856
rect 15764 18853 15776 18887
rect 16868 18884 16896 18915
rect 18506 18912 18512 18924
rect 18564 18912 18570 18964
rect 17402 18893 17408 18896
rect 17396 18884 17408 18893
rect 16868 18856 17408 18884
rect 15718 18847 15776 18853
rect 17396 18847 17408 18856
rect 17402 18844 17408 18847
rect 17460 18844 17466 18896
rect 18524 18884 18552 18912
rect 19030 18887 19088 18893
rect 19030 18884 19042 18887
rect 18524 18856 19042 18884
rect 19030 18853 19042 18856
rect 19076 18853 19088 18887
rect 19030 18847 19088 18853
rect 10870 18816 10876 18828
rect 7791 18788 8800 18816
rect 8956 18788 10876 18816
rect 7791 18785 7803 18788
rect 7745 18779 7803 18785
rect 2424 18720 5856 18748
rect 3142 18680 3148 18692
rect 3103 18652 3148 18680
rect 3142 18640 3148 18652
rect 3200 18640 3206 18692
rect 3234 18640 3240 18692
rect 3292 18680 3298 18692
rect 4982 18680 4988 18692
rect 3292 18652 4988 18680
rect 3292 18640 3298 18652
rect 4982 18640 4988 18652
rect 5040 18640 5046 18692
rect 5828 18680 5856 18720
rect 5902 18708 5908 18760
rect 5960 18708 5966 18760
rect 8772 18748 8800 18788
rect 10870 18776 10876 18788
rect 10928 18776 10934 18828
rect 11054 18776 11060 18828
rect 11112 18816 11118 18828
rect 11425 18819 11483 18825
rect 11425 18816 11437 18819
rect 11112 18788 11437 18816
rect 11112 18776 11118 18788
rect 11425 18785 11437 18788
rect 11471 18785 11483 18819
rect 11425 18779 11483 18785
rect 12158 18776 12164 18828
rect 12216 18816 12222 18828
rect 12529 18819 12587 18825
rect 12529 18816 12541 18819
rect 12216 18788 12541 18816
rect 12216 18776 12222 18788
rect 12529 18785 12541 18788
rect 12575 18785 12587 18819
rect 18598 18816 18604 18828
rect 12529 18779 12587 18785
rect 14384 18788 18604 18816
rect 9306 18748 9312 18760
rect 8772 18720 9312 18748
rect 9306 18708 9312 18720
rect 9364 18748 9370 18760
rect 9674 18748 9680 18760
rect 9364 18720 9680 18748
rect 9364 18708 9370 18720
rect 9674 18708 9680 18720
rect 9732 18748 9738 18760
rect 12710 18748 12716 18760
rect 9732 18720 9825 18748
rect 12623 18720 12716 18748
rect 9732 18708 9738 18720
rect 12710 18708 12716 18720
rect 12768 18708 12774 18760
rect 13173 18751 13231 18757
rect 13173 18717 13185 18751
rect 13219 18717 13231 18751
rect 13173 18711 13231 18717
rect 6454 18680 6460 18692
rect 5828 18652 6460 18680
rect 6454 18640 6460 18652
rect 6512 18640 6518 18692
rect 11057 18683 11115 18689
rect 11057 18649 11069 18683
rect 11103 18680 11115 18683
rect 12728 18680 12756 18708
rect 11103 18652 12756 18680
rect 11103 18649 11115 18652
rect 11057 18643 11115 18649
rect 12802 18640 12808 18692
rect 12860 18680 12866 18692
rect 13188 18680 13216 18711
rect 12860 18652 13216 18680
rect 12860 18640 12866 18652
rect 1394 18572 1400 18624
rect 1452 18612 1458 18624
rect 2038 18612 2044 18624
rect 1452 18584 2044 18612
rect 1452 18572 1458 18584
rect 2038 18572 2044 18584
rect 2096 18572 2102 18624
rect 2222 18572 2228 18624
rect 2280 18612 2286 18624
rect 3326 18612 3332 18624
rect 2280 18584 3332 18612
rect 2280 18572 2286 18584
rect 3326 18572 3332 18584
rect 3384 18572 3390 18624
rect 3510 18572 3516 18624
rect 3568 18612 3574 18624
rect 8386 18612 8392 18624
rect 3568 18584 8392 18612
rect 3568 18572 3574 18584
rect 8386 18572 8392 18584
rect 8444 18572 8450 18624
rect 9674 18572 9680 18624
rect 9732 18612 9738 18624
rect 14384 18612 14412 18788
rect 18598 18776 18604 18788
rect 18656 18776 18662 18828
rect 15473 18751 15531 18757
rect 15473 18717 15485 18751
rect 15519 18717 15531 18751
rect 17129 18751 17187 18757
rect 17129 18748 17141 18751
rect 15473 18711 15531 18717
rect 16592 18720 17141 18748
rect 14550 18612 14556 18624
rect 9732 18584 14412 18612
rect 14511 18584 14556 18612
rect 9732 18572 9738 18584
rect 14550 18572 14556 18584
rect 14608 18572 14614 18624
rect 15488 18612 15516 18711
rect 16114 18612 16120 18624
rect 15488 18584 16120 18612
rect 16114 18572 16120 18584
rect 16172 18612 16178 18624
rect 16592 18612 16620 18720
rect 17129 18717 17141 18720
rect 17175 18717 17187 18751
rect 17129 18711 17187 18717
rect 18506 18708 18512 18760
rect 18564 18748 18570 18760
rect 18785 18751 18843 18757
rect 18785 18748 18797 18751
rect 18564 18720 18797 18748
rect 18564 18708 18570 18720
rect 18785 18717 18797 18720
rect 18831 18717 18843 18751
rect 18785 18711 18843 18717
rect 16172 18584 16620 18612
rect 16172 18572 16178 18584
rect 16666 18572 16672 18624
rect 16724 18612 16730 18624
rect 18966 18612 18972 18624
rect 16724 18584 18972 18612
rect 16724 18572 16730 18584
rect 18966 18572 18972 18584
rect 19024 18572 19030 18624
rect 20162 18612 20168 18624
rect 20123 18584 20168 18612
rect 20162 18572 20168 18584
rect 20220 18572 20226 18624
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 1946 18408 1952 18420
rect 1907 18380 1952 18408
rect 1946 18368 1952 18380
rect 2004 18368 2010 18420
rect 2038 18368 2044 18420
rect 2096 18408 2102 18420
rect 2866 18408 2872 18420
rect 2096 18380 2872 18408
rect 2096 18368 2102 18380
rect 2866 18368 2872 18380
rect 2924 18408 2930 18420
rect 3510 18408 3516 18420
rect 2924 18380 3516 18408
rect 2924 18368 2930 18380
rect 3510 18368 3516 18380
rect 3568 18368 3574 18420
rect 8205 18411 8263 18417
rect 8205 18377 8217 18411
rect 8251 18408 8263 18411
rect 9122 18408 9128 18420
rect 8251 18380 9128 18408
rect 8251 18377 8263 18380
rect 8205 18371 8263 18377
rect 9122 18368 9128 18380
rect 9180 18368 9186 18420
rect 9214 18368 9220 18420
rect 9272 18408 9278 18420
rect 9950 18408 9956 18420
rect 9272 18380 9956 18408
rect 9272 18368 9278 18380
rect 9950 18368 9956 18380
rect 10008 18368 10014 18420
rect 10778 18408 10784 18420
rect 10060 18380 10784 18408
rect 3786 18340 3792 18352
rect 3747 18312 3792 18340
rect 3786 18300 3792 18312
rect 3844 18300 3850 18352
rect 6822 18300 6828 18352
rect 6880 18340 6886 18352
rect 10060 18340 10088 18380
rect 10778 18368 10784 18380
rect 10836 18368 10842 18420
rect 11425 18411 11483 18417
rect 11425 18377 11437 18411
rect 11471 18408 11483 18411
rect 11698 18408 11704 18420
rect 11471 18380 11704 18408
rect 11471 18377 11483 18380
rect 11425 18371 11483 18377
rect 11698 18368 11704 18380
rect 11756 18368 11762 18420
rect 12897 18411 12955 18417
rect 12897 18377 12909 18411
rect 12943 18408 12955 18411
rect 13262 18408 13268 18420
rect 12943 18380 13268 18408
rect 12943 18377 12955 18380
rect 12897 18371 12955 18377
rect 13262 18368 13268 18380
rect 13320 18368 13326 18420
rect 15470 18368 15476 18420
rect 15528 18408 15534 18420
rect 15657 18411 15715 18417
rect 15657 18408 15669 18411
rect 15528 18380 15669 18408
rect 15528 18368 15534 18380
rect 15657 18377 15669 18380
rect 15703 18377 15715 18411
rect 15930 18408 15936 18420
rect 15891 18380 15936 18408
rect 15657 18371 15715 18377
rect 15930 18368 15936 18380
rect 15988 18368 15994 18420
rect 16022 18368 16028 18420
rect 16080 18408 16086 18420
rect 16761 18411 16819 18417
rect 16761 18408 16773 18411
rect 16080 18380 16773 18408
rect 16080 18368 16086 18380
rect 16761 18377 16773 18380
rect 16807 18377 16819 18411
rect 16761 18371 16819 18377
rect 16945 18411 17003 18417
rect 16945 18377 16957 18411
rect 16991 18408 17003 18411
rect 17034 18408 17040 18420
rect 16991 18380 17040 18408
rect 16991 18377 17003 18380
rect 16945 18371 17003 18377
rect 17034 18368 17040 18380
rect 17092 18368 17098 18420
rect 17126 18368 17132 18420
rect 17184 18408 17190 18420
rect 19610 18408 19616 18420
rect 17184 18380 19616 18408
rect 17184 18368 17190 18380
rect 19610 18368 19616 18380
rect 19668 18408 19674 18420
rect 20438 18408 20444 18420
rect 19668 18380 20444 18408
rect 19668 18368 19674 18380
rect 20438 18368 20444 18380
rect 20496 18368 20502 18420
rect 20714 18408 20720 18420
rect 20675 18380 20720 18408
rect 20714 18368 20720 18380
rect 20772 18368 20778 18420
rect 6880 18312 10088 18340
rect 6880 18300 6886 18312
rect 12802 18300 12808 18352
rect 12860 18340 12866 18352
rect 13078 18340 13084 18352
rect 12860 18312 13084 18340
rect 12860 18300 12866 18312
rect 13078 18300 13084 18312
rect 13136 18340 13142 18352
rect 13136 18312 14320 18340
rect 13136 18300 13142 18312
rect 2130 18232 2136 18284
rect 2188 18272 2194 18284
rect 2501 18275 2559 18281
rect 2501 18272 2513 18275
rect 2188 18244 2513 18272
rect 2188 18232 2194 18244
rect 2501 18241 2513 18244
rect 2547 18241 2559 18275
rect 4798 18272 4804 18284
rect 2501 18235 2559 18241
rect 3068 18244 3556 18272
rect 4759 18244 4804 18272
rect 1762 18204 1768 18216
rect 1723 18176 1768 18204
rect 1762 18164 1768 18176
rect 1820 18164 1826 18216
rect 2038 18164 2044 18216
rect 2096 18204 2102 18216
rect 3068 18213 3096 18244
rect 2306 18207 2364 18213
rect 2306 18204 2318 18207
rect 2096 18176 2318 18204
rect 2096 18164 2102 18176
rect 2306 18173 2318 18176
rect 2352 18173 2364 18207
rect 2306 18167 2364 18173
rect 3053 18207 3111 18213
rect 3053 18173 3065 18207
rect 3099 18173 3111 18207
rect 3053 18167 3111 18173
rect 3234 18164 3240 18216
rect 3292 18164 3298 18216
rect 566 18028 572 18080
rect 624 18068 630 18080
rect 2222 18068 2228 18080
rect 624 18040 2228 18068
rect 624 18028 630 18040
rect 2222 18028 2228 18040
rect 2280 18028 2286 18080
rect 3252 18077 3280 18164
rect 3528 18136 3556 18244
rect 4798 18232 4804 18244
rect 4856 18232 4862 18284
rect 7282 18232 7288 18284
rect 7340 18272 7346 18284
rect 7469 18275 7527 18281
rect 7469 18272 7481 18275
rect 7340 18244 7481 18272
rect 7340 18232 7346 18244
rect 7469 18241 7481 18244
rect 7515 18241 7527 18275
rect 8754 18272 8760 18284
rect 8715 18244 8760 18272
rect 7469 18235 7527 18241
rect 8754 18232 8760 18244
rect 8812 18232 8818 18284
rect 8938 18232 8944 18284
rect 8996 18272 9002 18284
rect 8996 18244 10180 18272
rect 8996 18232 9002 18244
rect 3605 18207 3663 18213
rect 3605 18173 3617 18207
rect 3651 18204 3663 18207
rect 3878 18204 3884 18216
rect 3651 18176 3884 18204
rect 3651 18173 3663 18176
rect 3605 18167 3663 18173
rect 3878 18164 3884 18176
rect 3936 18164 3942 18216
rect 4154 18164 4160 18216
rect 4212 18204 4218 18216
rect 4525 18207 4583 18213
rect 4525 18204 4537 18207
rect 4212 18176 4537 18204
rect 4212 18164 4218 18176
rect 4525 18173 4537 18176
rect 4571 18173 4583 18207
rect 4525 18167 4583 18173
rect 5810 18164 5816 18216
rect 5868 18204 5874 18216
rect 8573 18207 8631 18213
rect 5868 18176 7420 18204
rect 5868 18164 5874 18176
rect 3786 18136 3792 18148
rect 3528 18108 3792 18136
rect 3786 18096 3792 18108
rect 3844 18096 3850 18148
rect 6822 18096 6828 18148
rect 6880 18136 6886 18148
rect 7392 18145 7420 18176
rect 8573 18173 8585 18207
rect 8619 18204 8631 18207
rect 8662 18204 8668 18216
rect 8619 18176 8668 18204
rect 8619 18173 8631 18176
rect 8573 18167 8631 18173
rect 8662 18164 8668 18176
rect 8720 18164 8726 18216
rect 8846 18164 8852 18216
rect 8904 18204 8910 18216
rect 9217 18207 9275 18213
rect 9217 18204 9229 18207
rect 8904 18176 9229 18204
rect 8904 18164 8910 18176
rect 9217 18173 9229 18176
rect 9263 18173 9275 18207
rect 9217 18167 9275 18173
rect 9306 18164 9312 18216
rect 9364 18204 9370 18216
rect 10045 18207 10103 18213
rect 10045 18204 10057 18207
rect 9364 18176 10057 18204
rect 9364 18164 9370 18176
rect 10045 18173 10057 18176
rect 10091 18173 10103 18207
rect 10152 18204 10180 18244
rect 12710 18232 12716 18284
rect 12768 18272 12774 18284
rect 14292 18281 14320 18312
rect 15746 18300 15752 18352
rect 15804 18340 15810 18352
rect 17218 18340 17224 18352
rect 15804 18312 17224 18340
rect 15804 18300 15810 18312
rect 17218 18300 17224 18312
rect 17276 18300 17282 18352
rect 18509 18343 18567 18349
rect 18509 18309 18521 18343
rect 18555 18340 18567 18343
rect 20254 18340 20260 18352
rect 18555 18312 20260 18340
rect 18555 18309 18567 18312
rect 18509 18303 18567 18309
rect 20254 18300 20260 18312
rect 20312 18300 20318 18352
rect 13449 18275 13507 18281
rect 13449 18272 13461 18275
rect 12768 18244 13461 18272
rect 12768 18232 12774 18244
rect 13449 18241 13461 18244
rect 13495 18241 13507 18275
rect 13449 18235 13507 18241
rect 14277 18275 14335 18281
rect 14277 18241 14289 18275
rect 14323 18241 14335 18275
rect 14277 18235 14335 18241
rect 15838 18232 15844 18284
rect 15896 18272 15902 18284
rect 16485 18275 16543 18281
rect 16485 18272 16497 18275
rect 15896 18244 16497 18272
rect 15896 18232 15902 18244
rect 16485 18241 16497 18244
rect 16531 18241 16543 18275
rect 16485 18235 16543 18241
rect 17402 18232 17408 18284
rect 17460 18272 17466 18284
rect 17497 18275 17555 18281
rect 17497 18272 17509 18275
rect 17460 18244 17509 18272
rect 17460 18232 17466 18244
rect 17497 18241 17509 18244
rect 17543 18241 17555 18275
rect 17497 18235 17555 18241
rect 19153 18275 19211 18281
rect 19153 18241 19165 18275
rect 19199 18272 19211 18275
rect 19242 18272 19248 18284
rect 19199 18244 19248 18272
rect 19199 18241 19211 18244
rect 19153 18235 19211 18241
rect 19242 18232 19248 18244
rect 19300 18272 19306 18284
rect 20162 18272 20168 18284
rect 19300 18244 20168 18272
rect 19300 18232 19306 18244
rect 20162 18232 20168 18244
rect 20220 18232 20226 18284
rect 12437 18207 12495 18213
rect 10152 18176 11100 18204
rect 10045 18167 10103 18173
rect 7285 18139 7343 18145
rect 7285 18136 7297 18139
rect 6880 18108 7297 18136
rect 6880 18096 6886 18108
rect 7285 18105 7297 18108
rect 7331 18105 7343 18139
rect 7285 18099 7343 18105
rect 7377 18139 7435 18145
rect 7377 18105 7389 18139
rect 7423 18136 7435 18139
rect 9493 18139 9551 18145
rect 7423 18108 8800 18136
rect 7423 18105 7435 18108
rect 7377 18099 7435 18105
rect 3237 18071 3295 18077
rect 3237 18037 3249 18071
rect 3283 18037 3295 18071
rect 3237 18031 3295 18037
rect 5258 18028 5264 18080
rect 5316 18068 5322 18080
rect 5718 18068 5724 18080
rect 5316 18040 5724 18068
rect 5316 18028 5322 18040
rect 5718 18028 5724 18040
rect 5776 18028 5782 18080
rect 6914 18068 6920 18080
rect 6875 18040 6920 18068
rect 6914 18028 6920 18040
rect 6972 18028 6978 18080
rect 8662 18068 8668 18080
rect 8623 18040 8668 18068
rect 8662 18028 8668 18040
rect 8720 18028 8726 18080
rect 8772 18068 8800 18108
rect 9493 18105 9505 18139
rect 9539 18136 9551 18139
rect 9674 18136 9680 18148
rect 9539 18108 9680 18136
rect 9539 18105 9551 18108
rect 9493 18099 9551 18105
rect 9674 18096 9680 18108
rect 9732 18096 9738 18148
rect 9766 18096 9772 18148
rect 9824 18136 9830 18148
rect 10290 18139 10348 18145
rect 10290 18136 10302 18139
rect 9824 18108 10302 18136
rect 9824 18096 9830 18108
rect 10290 18105 10302 18108
rect 10336 18105 10348 18139
rect 10290 18099 10348 18105
rect 10962 18068 10968 18080
rect 8772 18040 10968 18068
rect 10962 18028 10968 18040
rect 11020 18028 11026 18080
rect 11072 18068 11100 18176
rect 12437 18173 12449 18207
rect 12483 18204 12495 18207
rect 14182 18204 14188 18216
rect 12483 18176 14188 18204
rect 12483 18173 12495 18176
rect 12437 18167 12495 18173
rect 14182 18164 14188 18176
rect 14240 18164 14246 18216
rect 14550 18213 14556 18216
rect 14544 18204 14556 18213
rect 14511 18176 14556 18204
rect 14544 18167 14556 18176
rect 14550 18164 14556 18167
rect 14608 18164 14614 18216
rect 16761 18207 16819 18213
rect 16761 18173 16773 18207
rect 16807 18204 16819 18207
rect 19426 18204 19432 18216
rect 16807 18176 19432 18204
rect 16807 18173 16819 18176
rect 16761 18167 16819 18173
rect 19426 18164 19432 18176
rect 19484 18164 19490 18216
rect 20070 18164 20076 18216
rect 20128 18204 20134 18216
rect 20533 18207 20591 18213
rect 20533 18204 20545 18207
rect 20128 18176 20545 18204
rect 20128 18164 20134 18176
rect 20533 18173 20545 18176
rect 20579 18173 20591 18207
rect 20533 18167 20591 18173
rect 11885 18139 11943 18145
rect 11885 18105 11897 18139
rect 11931 18136 11943 18139
rect 13265 18139 13323 18145
rect 13265 18136 13277 18139
rect 11931 18108 13277 18136
rect 11931 18105 11943 18108
rect 11885 18099 11943 18105
rect 13265 18105 13277 18108
rect 13311 18105 13323 18139
rect 13265 18099 13323 18105
rect 13354 18096 13360 18148
rect 13412 18136 13418 18148
rect 13412 18108 13457 18136
rect 13412 18096 13418 18108
rect 14366 18096 14372 18148
rect 14424 18136 14430 18148
rect 14424 18108 16160 18136
rect 14424 18096 14430 18108
rect 16022 18068 16028 18080
rect 11072 18040 16028 18068
rect 16022 18028 16028 18040
rect 16080 18028 16086 18080
rect 16132 18068 16160 18108
rect 16298 18096 16304 18148
rect 16356 18136 16362 18148
rect 17313 18139 17371 18145
rect 16356 18108 16401 18136
rect 16356 18096 16362 18108
rect 17313 18105 17325 18139
rect 17359 18136 17371 18139
rect 18049 18139 18107 18145
rect 18049 18136 18061 18139
rect 17359 18108 18061 18136
rect 17359 18105 17371 18108
rect 17313 18099 17371 18105
rect 18049 18105 18061 18108
rect 18095 18105 18107 18139
rect 18049 18099 18107 18105
rect 18877 18139 18935 18145
rect 18877 18105 18889 18139
rect 18923 18136 18935 18139
rect 19058 18136 19064 18148
rect 18923 18108 19064 18136
rect 18923 18105 18935 18108
rect 18877 18099 18935 18105
rect 19058 18096 19064 18108
rect 19116 18096 19122 18148
rect 19889 18139 19947 18145
rect 19889 18105 19901 18139
rect 19935 18136 19947 18139
rect 20898 18136 20904 18148
rect 19935 18108 20904 18136
rect 19935 18105 19947 18108
rect 19889 18099 19947 18105
rect 20898 18096 20904 18108
rect 20956 18096 20962 18148
rect 16393 18071 16451 18077
rect 16393 18068 16405 18071
rect 16132 18040 16405 18068
rect 16393 18037 16405 18040
rect 16439 18037 16451 18071
rect 17402 18068 17408 18080
rect 17363 18040 17408 18068
rect 16393 18031 16451 18037
rect 17402 18028 17408 18040
rect 17460 18028 17466 18080
rect 17586 18028 17592 18080
rect 17644 18068 17650 18080
rect 18782 18068 18788 18080
rect 17644 18040 18788 18068
rect 17644 18028 17650 18040
rect 18782 18028 18788 18040
rect 18840 18028 18846 18080
rect 18966 18068 18972 18080
rect 18927 18040 18972 18068
rect 18966 18028 18972 18040
rect 19024 18028 19030 18080
rect 19518 18068 19524 18080
rect 19479 18040 19524 18068
rect 19518 18028 19524 18040
rect 19576 18028 19582 18080
rect 19981 18071 20039 18077
rect 19981 18037 19993 18071
rect 20027 18068 20039 18071
rect 20530 18068 20536 18080
rect 20027 18040 20536 18068
rect 20027 18037 20039 18040
rect 19981 18031 20039 18037
rect 20530 18028 20536 18040
rect 20588 18028 20594 18080
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 1946 17864 1952 17876
rect 1907 17836 1952 17864
rect 1946 17824 1952 17836
rect 2004 17824 2010 17876
rect 2501 17867 2559 17873
rect 2501 17833 2513 17867
rect 2547 17864 2559 17867
rect 2774 17864 2780 17876
rect 2547 17836 2780 17864
rect 2547 17833 2559 17836
rect 2501 17827 2559 17833
rect 2774 17824 2780 17836
rect 2832 17824 2838 17876
rect 4062 17824 4068 17876
rect 4120 17864 4126 17876
rect 6638 17864 6644 17876
rect 4120 17836 6644 17864
rect 4120 17824 4126 17836
rect 6638 17824 6644 17836
rect 6696 17824 6702 17876
rect 7098 17824 7104 17876
rect 7156 17864 7162 17876
rect 7193 17867 7251 17873
rect 7193 17864 7205 17867
rect 7156 17836 7205 17864
rect 7156 17824 7162 17836
rect 7193 17833 7205 17836
rect 7239 17833 7251 17867
rect 9033 17867 9091 17873
rect 7193 17827 7251 17833
rect 7300 17836 8248 17864
rect 2332 17768 3464 17796
rect 2332 17737 2360 17768
rect 1765 17731 1823 17737
rect 1765 17697 1777 17731
rect 1811 17697 1823 17731
rect 1765 17691 1823 17697
rect 2317 17731 2375 17737
rect 2317 17697 2329 17731
rect 2363 17697 2375 17731
rect 2317 17691 2375 17697
rect 2869 17731 2927 17737
rect 2869 17697 2881 17731
rect 2915 17728 2927 17731
rect 3326 17728 3332 17740
rect 2915 17700 3332 17728
rect 2915 17697 2927 17700
rect 2869 17691 2927 17697
rect 1780 17660 1808 17691
rect 3326 17688 3332 17700
rect 3384 17688 3390 17740
rect 3436 17728 3464 17768
rect 3510 17756 3516 17808
rect 3568 17796 3574 17808
rect 7300 17796 7328 17836
rect 8110 17796 8116 17808
rect 3568 17768 7328 17796
rect 7392 17768 8116 17796
rect 3568 17756 3574 17768
rect 3436 17700 4200 17728
rect 4062 17660 4068 17672
rect 1780 17632 4068 17660
rect 4062 17620 4068 17632
rect 4120 17620 4126 17672
rect 4172 17660 4200 17700
rect 4246 17688 4252 17740
rect 4304 17728 4310 17740
rect 4433 17731 4491 17737
rect 4433 17728 4445 17731
rect 4304 17700 4445 17728
rect 4304 17688 4310 17700
rect 4433 17697 4445 17700
rect 4479 17697 4491 17731
rect 4433 17691 4491 17697
rect 4525 17731 4583 17737
rect 4525 17697 4537 17731
rect 4571 17728 4583 17731
rect 4798 17728 4804 17740
rect 4571 17700 4804 17728
rect 4571 17697 4583 17700
rect 4525 17691 4583 17697
rect 4798 17688 4804 17700
rect 4856 17688 4862 17740
rect 5810 17737 5816 17740
rect 5804 17691 5816 17737
rect 5868 17728 5874 17740
rect 7282 17728 7288 17740
rect 5868 17700 7288 17728
rect 5810 17688 5816 17691
rect 5868 17688 5874 17700
rect 7282 17688 7288 17700
rect 7340 17728 7346 17740
rect 7392 17728 7420 17768
rect 8110 17756 8116 17768
rect 8168 17756 8174 17808
rect 8220 17796 8248 17836
rect 9033 17833 9045 17867
rect 9079 17864 9091 17867
rect 9398 17864 9404 17876
rect 9079 17836 9404 17864
rect 9079 17833 9091 17836
rect 9033 17827 9091 17833
rect 9398 17824 9404 17836
rect 9456 17824 9462 17876
rect 9766 17824 9772 17876
rect 9824 17864 9830 17876
rect 11057 17867 11115 17873
rect 11057 17864 11069 17867
rect 9824 17836 11069 17864
rect 9824 17824 9830 17836
rect 11057 17833 11069 17836
rect 11103 17833 11115 17867
rect 11057 17827 11115 17833
rect 11146 17824 11152 17876
rect 11204 17864 11210 17876
rect 11333 17867 11391 17873
rect 11333 17864 11345 17867
rect 11204 17836 11345 17864
rect 11204 17824 11210 17836
rect 11333 17833 11345 17836
rect 11379 17833 11391 17867
rect 11333 17827 11391 17833
rect 12802 17824 12808 17876
rect 12860 17864 12866 17876
rect 13173 17867 13231 17873
rect 13173 17864 13185 17867
rect 12860 17836 13185 17864
rect 12860 17824 12866 17836
rect 13173 17833 13185 17836
rect 13219 17864 13231 17867
rect 13998 17864 14004 17876
rect 13219 17836 14004 17864
rect 13219 17833 13231 17836
rect 13173 17827 13231 17833
rect 13998 17824 14004 17836
rect 14056 17824 14062 17876
rect 15194 17824 15200 17876
rect 15252 17864 15258 17876
rect 15289 17867 15347 17873
rect 15289 17864 15301 17867
rect 15252 17836 15301 17864
rect 15252 17824 15258 17836
rect 15289 17833 15301 17836
rect 15335 17833 15347 17867
rect 16574 17864 16580 17876
rect 16535 17836 16580 17864
rect 15289 17827 15347 17833
rect 16574 17824 16580 17836
rect 16632 17824 16638 17876
rect 17865 17867 17923 17873
rect 17865 17833 17877 17867
rect 17911 17864 17923 17867
rect 17954 17864 17960 17876
rect 17911 17836 17960 17864
rect 17911 17833 17923 17836
rect 17865 17827 17923 17833
rect 17954 17824 17960 17836
rect 18012 17824 18018 17876
rect 18601 17867 18659 17873
rect 18601 17833 18613 17867
rect 18647 17864 18659 17867
rect 18782 17864 18788 17876
rect 18647 17836 18788 17864
rect 18647 17833 18659 17836
rect 18601 17827 18659 17833
rect 18782 17824 18788 17836
rect 18840 17824 18846 17876
rect 20898 17864 20904 17876
rect 20859 17836 20904 17864
rect 20898 17824 20904 17836
rect 20956 17824 20962 17876
rect 9944 17799 10002 17805
rect 8220 17768 9904 17796
rect 7558 17728 7564 17740
rect 7340 17700 7420 17728
rect 7519 17700 7564 17728
rect 7340 17688 7346 17700
rect 7558 17688 7564 17700
rect 7616 17688 7622 17740
rect 8941 17731 8999 17737
rect 8941 17697 8953 17731
rect 8987 17728 8999 17731
rect 9122 17728 9128 17740
rect 8987 17700 9128 17728
rect 8987 17697 8999 17700
rect 8941 17691 8999 17697
rect 9122 17688 9128 17700
rect 9180 17688 9186 17740
rect 9766 17728 9772 17740
rect 9232 17700 9772 17728
rect 4706 17660 4712 17672
rect 4172 17632 4568 17660
rect 4667 17632 4712 17660
rect 3234 17552 3240 17604
rect 3292 17592 3298 17604
rect 4540 17592 4568 17632
rect 4706 17620 4712 17632
rect 4764 17620 4770 17672
rect 5534 17660 5540 17672
rect 5495 17632 5540 17660
rect 5534 17620 5540 17632
rect 5592 17620 5598 17672
rect 6822 17620 6828 17672
rect 6880 17660 6886 17672
rect 7653 17663 7711 17669
rect 7653 17660 7665 17663
rect 6880 17632 7665 17660
rect 6880 17620 6886 17632
rect 7653 17629 7665 17632
rect 7699 17629 7711 17663
rect 7653 17623 7711 17629
rect 7742 17620 7748 17672
rect 7800 17660 7806 17672
rect 9232 17669 9260 17700
rect 9766 17688 9772 17700
rect 9824 17688 9830 17740
rect 9876 17728 9904 17768
rect 9944 17765 9956 17799
rect 9990 17796 10002 17799
rect 10410 17796 10416 17808
rect 9990 17768 10416 17796
rect 9990 17765 10002 17768
rect 9944 17759 10002 17765
rect 10410 17756 10416 17768
rect 10468 17756 10474 17808
rect 11790 17796 11796 17808
rect 11624 17768 11796 17796
rect 10226 17728 10232 17740
rect 9876 17700 10232 17728
rect 10226 17688 10232 17700
rect 10284 17688 10290 17740
rect 11146 17688 11152 17740
rect 11204 17728 11210 17740
rect 11624 17728 11652 17768
rect 11790 17756 11796 17768
rect 11848 17756 11854 17808
rect 14182 17756 14188 17808
rect 14240 17796 14246 17808
rect 15657 17799 15715 17805
rect 15657 17796 15669 17799
rect 14240 17768 15669 17796
rect 14240 17756 14246 17768
rect 15657 17765 15669 17768
rect 15703 17765 15715 17799
rect 15657 17759 15715 17765
rect 16850 17756 16856 17808
rect 16908 17796 16914 17808
rect 19242 17805 19248 17808
rect 19236 17796 19248 17805
rect 16908 17768 17724 17796
rect 19203 17768 19248 17796
rect 16908 17756 16914 17768
rect 11204 17700 11652 17728
rect 11701 17731 11759 17737
rect 11204 17688 11210 17700
rect 11701 17697 11713 17731
rect 11747 17728 11759 17731
rect 12345 17731 12403 17737
rect 12345 17728 12357 17731
rect 11747 17700 12357 17728
rect 11747 17697 11759 17700
rect 11701 17691 11759 17697
rect 12345 17697 12357 17700
rect 12391 17697 12403 17731
rect 12345 17691 12403 17697
rect 13909 17731 13967 17737
rect 13909 17697 13921 17731
rect 13955 17697 13967 17731
rect 13909 17691 13967 17697
rect 14277 17731 14335 17737
rect 14277 17697 14289 17731
rect 14323 17728 14335 17731
rect 14461 17731 14519 17737
rect 14461 17728 14473 17731
rect 14323 17700 14473 17728
rect 14323 17697 14335 17700
rect 14277 17691 14335 17697
rect 14461 17697 14473 17700
rect 14507 17697 14519 17731
rect 14461 17691 14519 17697
rect 14737 17731 14795 17737
rect 14737 17697 14749 17731
rect 14783 17728 14795 17731
rect 15286 17728 15292 17740
rect 14783 17700 15292 17728
rect 14783 17697 14795 17700
rect 14737 17691 14795 17697
rect 9217 17663 9275 17669
rect 7800 17632 7845 17660
rect 7800 17620 7806 17632
rect 9217 17629 9229 17663
rect 9263 17629 9275 17663
rect 9217 17623 9275 17629
rect 9306 17620 9312 17672
rect 9364 17660 9370 17672
rect 9490 17660 9496 17672
rect 9364 17632 9496 17660
rect 9364 17620 9370 17632
rect 9490 17620 9496 17632
rect 9548 17660 9554 17672
rect 9677 17663 9735 17669
rect 9677 17660 9689 17663
rect 9548 17632 9689 17660
rect 9548 17620 9554 17632
rect 9677 17629 9689 17632
rect 9723 17629 9735 17663
rect 9677 17623 9735 17629
rect 11790 17620 11796 17672
rect 11848 17660 11854 17672
rect 11885 17663 11943 17669
rect 11885 17660 11897 17663
rect 11848 17632 11897 17660
rect 11848 17620 11854 17632
rect 11885 17629 11897 17632
rect 11931 17629 11943 17663
rect 11885 17623 11943 17629
rect 12618 17620 12624 17672
rect 12676 17660 12682 17672
rect 13265 17663 13323 17669
rect 13265 17660 13277 17663
rect 12676 17632 13277 17660
rect 12676 17620 12682 17632
rect 13265 17629 13277 17632
rect 13311 17629 13323 17663
rect 13265 17623 13323 17629
rect 13449 17663 13507 17669
rect 13449 17629 13461 17663
rect 13495 17660 13507 17663
rect 13538 17660 13544 17672
rect 13495 17632 13544 17660
rect 13495 17629 13507 17632
rect 13449 17623 13507 17629
rect 13538 17620 13544 17632
rect 13596 17620 13602 17672
rect 13722 17620 13728 17672
rect 13780 17660 13786 17672
rect 13924 17660 13952 17691
rect 15286 17688 15292 17700
rect 15344 17688 15350 17740
rect 15746 17728 15752 17740
rect 15707 17700 15752 17728
rect 15746 17688 15752 17700
rect 15804 17688 15810 17740
rect 16393 17731 16451 17737
rect 16393 17697 16405 17731
rect 16439 17697 16451 17731
rect 16942 17728 16948 17740
rect 16903 17700 16948 17728
rect 16393 17691 16451 17697
rect 13780 17632 13952 17660
rect 13780 17620 13786 17632
rect 14550 17620 14556 17672
rect 14608 17660 14614 17672
rect 15838 17660 15844 17672
rect 14608 17632 15844 17660
rect 14608 17620 14614 17632
rect 15838 17620 15844 17632
rect 15896 17620 15902 17672
rect 16408 17660 16436 17691
rect 16942 17688 16948 17700
rect 17000 17688 17006 17740
rect 17696 17737 17724 17768
rect 19236 17759 19248 17768
rect 19242 17756 19248 17759
rect 19300 17756 19306 17808
rect 17681 17731 17739 17737
rect 17681 17697 17693 17731
rect 17727 17697 17739 17731
rect 18414 17728 18420 17740
rect 18375 17700 18420 17728
rect 17681 17691 17739 17697
rect 18414 17688 18420 17700
rect 18472 17688 18478 17740
rect 19610 17728 19616 17740
rect 18524 17700 19616 17728
rect 17129 17663 17187 17669
rect 17129 17660 17141 17663
rect 16408 17632 17141 17660
rect 17129 17629 17141 17632
rect 17175 17629 17187 17663
rect 17129 17623 17187 17629
rect 5442 17592 5448 17604
rect 3292 17564 4200 17592
rect 4540 17564 5448 17592
rect 3292 17552 3298 17564
rect 3050 17524 3056 17536
rect 3011 17496 3056 17524
rect 3050 17484 3056 17496
rect 3108 17484 3114 17536
rect 3970 17484 3976 17536
rect 4028 17524 4034 17536
rect 4065 17527 4123 17533
rect 4065 17524 4077 17527
rect 4028 17496 4077 17524
rect 4028 17484 4034 17496
rect 4065 17493 4077 17496
rect 4111 17493 4123 17527
rect 4172 17524 4200 17564
rect 5442 17552 5448 17564
rect 5500 17552 5506 17604
rect 9398 17592 9404 17604
rect 6472 17564 9404 17592
rect 6472 17524 6500 17564
rect 9398 17552 9404 17564
rect 9456 17552 9462 17604
rect 14277 17595 14335 17601
rect 14277 17592 14289 17595
rect 10612 17564 14289 17592
rect 4172 17496 6500 17524
rect 6917 17527 6975 17533
rect 4065 17487 4123 17493
rect 6917 17493 6929 17527
rect 6963 17524 6975 17527
rect 7374 17524 7380 17536
rect 6963 17496 7380 17524
rect 6963 17493 6975 17496
rect 6917 17487 6975 17493
rect 7374 17484 7380 17496
rect 7432 17484 7438 17536
rect 8573 17527 8631 17533
rect 8573 17493 8585 17527
rect 8619 17524 8631 17527
rect 10612 17524 10640 17564
rect 14277 17561 14289 17564
rect 14323 17561 14335 17595
rect 18524 17592 18552 17700
rect 19610 17688 19616 17700
rect 19668 17688 19674 17740
rect 18598 17620 18604 17672
rect 18656 17660 18662 17672
rect 18782 17660 18788 17672
rect 18656 17632 18788 17660
rect 18656 17620 18662 17632
rect 18782 17620 18788 17632
rect 18840 17660 18846 17672
rect 18969 17663 19027 17669
rect 18969 17660 18981 17663
rect 18840 17632 18981 17660
rect 18840 17620 18846 17632
rect 18969 17629 18981 17632
rect 19015 17629 19027 17663
rect 18969 17623 19027 17629
rect 14277 17555 14335 17561
rect 15856 17564 18552 17592
rect 8619 17496 10640 17524
rect 12805 17527 12863 17533
rect 8619 17493 8631 17496
rect 8573 17487 8631 17493
rect 12805 17493 12817 17527
rect 12851 17524 12863 17527
rect 13262 17524 13268 17536
rect 12851 17496 13268 17524
rect 12851 17493 12863 17496
rect 12805 17487 12863 17493
rect 13262 17484 13268 17496
rect 13320 17484 13326 17536
rect 14093 17527 14151 17533
rect 14093 17493 14105 17527
rect 14139 17524 14151 17527
rect 15856 17524 15884 17564
rect 14139 17496 15884 17524
rect 14139 17493 14151 17496
rect 14093 17487 14151 17493
rect 16758 17484 16764 17536
rect 16816 17524 16822 17536
rect 18966 17524 18972 17536
rect 16816 17496 18972 17524
rect 16816 17484 16822 17496
rect 18966 17484 18972 17496
rect 19024 17484 19030 17536
rect 19886 17484 19892 17536
rect 19944 17524 19950 17536
rect 20349 17527 20407 17533
rect 20349 17524 20361 17527
rect 19944 17496 20361 17524
rect 19944 17484 19950 17496
rect 20349 17493 20361 17496
rect 20395 17493 20407 17527
rect 20349 17487 20407 17493
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 2501 17323 2559 17329
rect 2501 17289 2513 17323
rect 2547 17320 2559 17323
rect 2774 17320 2780 17332
rect 2547 17292 2780 17320
rect 2547 17289 2559 17292
rect 2501 17283 2559 17289
rect 2774 17280 2780 17292
rect 2832 17280 2838 17332
rect 3050 17280 3056 17332
rect 3108 17320 3114 17332
rect 6822 17320 6828 17332
rect 3108 17292 6592 17320
rect 6783 17292 6828 17320
rect 3108 17280 3114 17292
rect 3513 17255 3571 17261
rect 3513 17221 3525 17255
rect 3559 17252 3571 17255
rect 4062 17252 4068 17264
rect 3559 17224 4068 17252
rect 3559 17221 3571 17224
rect 3513 17215 3571 17221
rect 4062 17212 4068 17224
rect 4120 17212 4126 17264
rect 5810 17212 5816 17264
rect 5868 17252 5874 17264
rect 5905 17255 5963 17261
rect 5905 17252 5917 17255
rect 5868 17224 5917 17252
rect 5868 17212 5874 17224
rect 5905 17221 5917 17224
rect 5951 17221 5963 17255
rect 6564 17252 6592 17292
rect 6822 17280 6828 17292
rect 6880 17280 6886 17332
rect 7098 17280 7104 17332
rect 7156 17320 7162 17332
rect 10870 17320 10876 17332
rect 7156 17292 10876 17320
rect 7156 17280 7162 17292
rect 10870 17280 10876 17292
rect 10928 17280 10934 17332
rect 11149 17323 11207 17329
rect 11149 17289 11161 17323
rect 11195 17320 11207 17323
rect 11606 17320 11612 17332
rect 11195 17292 11612 17320
rect 11195 17289 11207 17292
rect 11149 17283 11207 17289
rect 11606 17280 11612 17292
rect 11664 17280 11670 17332
rect 12897 17323 12955 17329
rect 12897 17289 12909 17323
rect 12943 17320 12955 17323
rect 13817 17323 13875 17329
rect 13817 17320 13829 17323
rect 12943 17292 13829 17320
rect 12943 17289 12955 17292
rect 12897 17283 12955 17289
rect 13817 17289 13829 17292
rect 13863 17289 13875 17323
rect 13817 17283 13875 17289
rect 14093 17323 14151 17329
rect 14093 17289 14105 17323
rect 14139 17320 14151 17323
rect 15102 17320 15108 17332
rect 14139 17292 15108 17320
rect 14139 17289 14151 17292
rect 14093 17283 14151 17289
rect 15102 17280 15108 17292
rect 15160 17280 15166 17332
rect 15378 17320 15384 17332
rect 15339 17292 15384 17320
rect 15378 17280 15384 17292
rect 15436 17280 15442 17332
rect 15933 17323 15991 17329
rect 15933 17289 15945 17323
rect 15979 17320 15991 17323
rect 16666 17320 16672 17332
rect 15979 17292 16672 17320
rect 15979 17289 15991 17292
rect 15933 17283 15991 17289
rect 16666 17280 16672 17292
rect 16724 17280 16730 17332
rect 16942 17280 16948 17332
rect 17000 17320 17006 17332
rect 18049 17323 18107 17329
rect 18049 17320 18061 17323
rect 17000 17292 18061 17320
rect 17000 17280 17006 17292
rect 18049 17289 18061 17292
rect 18095 17289 18107 17323
rect 18049 17283 18107 17289
rect 18874 17280 18880 17332
rect 18932 17320 18938 17332
rect 19245 17323 19303 17329
rect 19245 17320 19257 17323
rect 18932 17292 19257 17320
rect 18932 17280 18938 17292
rect 19245 17289 19257 17292
rect 19291 17289 19303 17323
rect 19245 17283 19303 17289
rect 19334 17280 19340 17332
rect 19392 17320 19398 17332
rect 21726 17320 21732 17332
rect 19392 17292 21732 17320
rect 19392 17280 19398 17292
rect 21726 17280 21732 17292
rect 21784 17280 21790 17332
rect 14182 17252 14188 17264
rect 6564 17224 14188 17252
rect 5905 17215 5963 17221
rect 14182 17212 14188 17224
rect 14240 17212 14246 17264
rect 17402 17212 17408 17264
rect 17460 17252 17466 17264
rect 17460 17224 19104 17252
rect 17460 17212 17466 17224
rect 3970 17184 3976 17196
rect 3931 17156 3976 17184
rect 3970 17144 3976 17156
rect 4028 17144 4034 17196
rect 4157 17187 4215 17193
rect 4157 17153 4169 17187
rect 4203 17184 4215 17187
rect 4203 17156 4660 17184
rect 4203 17153 4215 17156
rect 4157 17147 4215 17153
rect 1765 17119 1823 17125
rect 1765 17085 1777 17119
rect 1811 17085 1823 17119
rect 1765 17079 1823 17085
rect 1780 17048 1808 17079
rect 1854 17076 1860 17128
rect 1912 17116 1918 17128
rect 2317 17119 2375 17125
rect 2317 17116 2329 17119
rect 1912 17088 2329 17116
rect 1912 17076 1918 17088
rect 2317 17085 2329 17088
rect 2363 17085 2375 17119
rect 2317 17079 2375 17085
rect 2869 17119 2927 17125
rect 2869 17085 2881 17119
rect 2915 17116 2927 17119
rect 2958 17116 2964 17128
rect 2915 17088 2964 17116
rect 2915 17085 2927 17088
rect 2869 17079 2927 17085
rect 2958 17076 2964 17088
rect 3016 17076 3022 17128
rect 4522 17116 4528 17128
rect 4483 17088 4528 17116
rect 4522 17076 4528 17088
rect 4580 17076 4586 17128
rect 2130 17048 2136 17060
rect 1780 17020 2136 17048
rect 2130 17008 2136 17020
rect 2188 17008 2194 17060
rect 4632 17048 4660 17156
rect 6914 17144 6920 17196
rect 6972 17184 6978 17196
rect 7285 17187 7343 17193
rect 7285 17184 7297 17187
rect 6972 17156 7297 17184
rect 6972 17144 6978 17156
rect 7285 17153 7297 17156
rect 7331 17153 7343 17187
rect 7285 17147 7343 17153
rect 7374 17144 7380 17196
rect 7432 17184 7438 17196
rect 7432 17156 7477 17184
rect 7432 17144 7438 17156
rect 8110 17144 8116 17196
rect 8168 17184 8174 17196
rect 8389 17187 8447 17193
rect 8389 17184 8401 17187
rect 8168 17156 8401 17184
rect 8168 17144 8174 17156
rect 8389 17153 8401 17156
rect 8435 17153 8447 17187
rect 8389 17147 8447 17153
rect 9030 17144 9036 17196
rect 9088 17184 9094 17196
rect 9214 17184 9220 17196
rect 9088 17156 9220 17184
rect 9088 17144 9094 17156
rect 9214 17144 9220 17156
rect 9272 17144 9278 17196
rect 9398 17184 9404 17196
rect 9359 17156 9404 17184
rect 9398 17144 9404 17156
rect 9456 17144 9462 17196
rect 9585 17187 9643 17193
rect 9585 17153 9597 17187
rect 9631 17184 9643 17187
rect 9858 17184 9864 17196
rect 9631 17156 9864 17184
rect 9631 17153 9643 17156
rect 9585 17147 9643 17153
rect 9858 17144 9864 17156
rect 9916 17184 9922 17196
rect 10505 17187 10563 17193
rect 10505 17184 10517 17187
rect 9916 17156 10517 17184
rect 9916 17144 9922 17156
rect 10505 17153 10517 17156
rect 10551 17153 10563 17187
rect 10505 17147 10563 17153
rect 11793 17187 11851 17193
rect 11793 17153 11805 17187
rect 11839 17153 11851 17187
rect 11793 17147 11851 17153
rect 13541 17187 13599 17193
rect 13541 17153 13553 17187
rect 13587 17184 13599 17187
rect 13814 17184 13820 17196
rect 13587 17156 13820 17184
rect 13587 17153 13599 17156
rect 13541 17147 13599 17153
rect 6638 17076 6644 17128
rect 6696 17116 6702 17128
rect 6822 17116 6828 17128
rect 6696 17088 6828 17116
rect 6696 17076 6702 17088
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 7466 17076 7472 17128
rect 7524 17116 7530 17128
rect 10594 17116 10600 17128
rect 7524 17088 10600 17116
rect 7524 17076 7530 17088
rect 10594 17076 10600 17088
rect 10652 17076 10658 17128
rect 10870 17116 10876 17128
rect 10783 17088 10876 17116
rect 10870 17076 10876 17088
rect 10928 17116 10934 17128
rect 10928 17088 11652 17116
rect 10928 17076 10934 17088
rect 4792 17051 4850 17057
rect 4792 17048 4804 17051
rect 4632 17020 4804 17048
rect 4792 17017 4804 17020
rect 4838 17048 4850 17051
rect 5442 17048 5448 17060
rect 4838 17020 5448 17048
rect 4838 17017 4850 17020
rect 4792 17011 4850 17017
rect 5442 17008 5448 17020
rect 5500 17008 5506 17060
rect 7193 17051 7251 17057
rect 7193 17017 7205 17051
rect 7239 17048 7251 17051
rect 7239 17020 7880 17048
rect 7239 17017 7251 17020
rect 7193 17011 7251 17017
rect 1946 16980 1952 16992
rect 1907 16952 1952 16980
rect 1946 16940 1952 16952
rect 2004 16940 2010 16992
rect 3050 16980 3056 16992
rect 3011 16952 3056 16980
rect 3050 16940 3056 16952
rect 3108 16940 3114 16992
rect 3878 16980 3884 16992
rect 3839 16952 3884 16980
rect 3878 16940 3884 16952
rect 3936 16940 3942 16992
rect 7852 16989 7880 17020
rect 8018 17008 8024 17060
rect 8076 17048 8082 17060
rect 8297 17051 8355 17057
rect 8297 17048 8309 17051
rect 8076 17020 8309 17048
rect 8076 17008 8082 17020
rect 8297 17017 8309 17020
rect 8343 17048 8355 17051
rect 10042 17048 10048 17060
rect 8343 17020 10048 17048
rect 8343 17017 8355 17020
rect 8297 17011 8355 17017
rect 10042 17008 10048 17020
rect 10100 17008 10106 17060
rect 10226 17008 10232 17060
rect 10284 17048 10290 17060
rect 10321 17051 10379 17057
rect 10321 17048 10333 17051
rect 10284 17020 10333 17048
rect 10284 17008 10290 17020
rect 10321 17017 10333 17020
rect 10367 17017 10379 17051
rect 10321 17011 10379 17017
rect 10413 17051 10471 17057
rect 10413 17017 10425 17051
rect 10459 17048 10471 17051
rect 10888 17048 10916 17076
rect 10459 17020 10916 17048
rect 10459 17017 10471 17020
rect 10413 17011 10471 17017
rect 10962 17008 10968 17060
rect 11020 17048 11026 17060
rect 11514 17048 11520 17060
rect 11020 17020 11520 17048
rect 11020 17008 11026 17020
rect 11514 17008 11520 17020
rect 11572 17008 11578 17060
rect 11624 17048 11652 17088
rect 11698 17076 11704 17128
rect 11756 17116 11762 17128
rect 11808 17116 11836 17147
rect 13814 17144 13820 17156
rect 13872 17144 13878 17196
rect 18693 17187 18751 17193
rect 18693 17153 18705 17187
rect 18739 17153 18751 17187
rect 19076 17184 19104 17224
rect 19150 17212 19156 17264
rect 19208 17252 19214 17264
rect 20717 17255 20775 17261
rect 20717 17252 20729 17255
rect 19208 17224 20729 17252
rect 19208 17212 19214 17224
rect 20717 17221 20729 17224
rect 20763 17221 20775 17255
rect 20717 17215 20775 17221
rect 19076 17156 19748 17184
rect 18693 17147 18751 17153
rect 13262 17116 13268 17128
rect 11756 17088 11836 17116
rect 13223 17088 13268 17116
rect 11756 17076 11762 17088
rect 13262 17076 13268 17088
rect 13320 17076 13326 17128
rect 13354 17076 13360 17128
rect 13412 17116 13418 17128
rect 13909 17119 13967 17125
rect 13412 17088 13457 17116
rect 13412 17076 13418 17088
rect 13909 17085 13921 17119
rect 13955 17116 13967 17119
rect 13998 17116 14004 17128
rect 13955 17088 14004 17116
rect 13955 17085 13967 17088
rect 13909 17079 13967 17085
rect 13998 17076 14004 17088
rect 14056 17076 14062 17128
rect 14090 17076 14096 17128
rect 14148 17116 14154 17128
rect 14461 17119 14519 17125
rect 14461 17116 14473 17119
rect 14148 17088 14473 17116
rect 14148 17076 14154 17088
rect 14461 17085 14473 17088
rect 14507 17085 14519 17119
rect 14461 17079 14519 17085
rect 14737 17119 14795 17125
rect 14737 17085 14749 17119
rect 14783 17116 14795 17119
rect 15197 17119 15255 17125
rect 15197 17116 15209 17119
rect 14783 17088 15209 17116
rect 14783 17085 14795 17088
rect 14737 17079 14795 17085
rect 15197 17085 15209 17088
rect 15243 17085 15255 17119
rect 15197 17079 15255 17085
rect 15749 17119 15807 17125
rect 15749 17085 15761 17119
rect 15795 17085 15807 17119
rect 15749 17079 15807 17085
rect 13817 17051 13875 17057
rect 11624 17020 12848 17048
rect 7837 16983 7895 16989
rect 7837 16949 7849 16983
rect 7883 16949 7895 16983
rect 7837 16943 7895 16949
rect 8205 16983 8263 16989
rect 8205 16949 8217 16983
rect 8251 16980 8263 16983
rect 8386 16980 8392 16992
rect 8251 16952 8392 16980
rect 8251 16949 8263 16952
rect 8205 16943 8263 16949
rect 8386 16940 8392 16952
rect 8444 16940 8450 16992
rect 8938 16980 8944 16992
rect 8899 16952 8944 16980
rect 8938 16940 8944 16952
rect 8996 16940 9002 16992
rect 9030 16940 9036 16992
rect 9088 16980 9094 16992
rect 9309 16983 9367 16989
rect 9309 16980 9321 16983
rect 9088 16952 9321 16980
rect 9088 16940 9094 16952
rect 9309 16949 9321 16952
rect 9355 16949 9367 16983
rect 9309 16943 9367 16949
rect 9398 16940 9404 16992
rect 9456 16980 9462 16992
rect 9953 16983 10011 16989
rect 9953 16980 9965 16983
rect 9456 16952 9965 16980
rect 9456 16940 9462 16952
rect 9953 16949 9965 16952
rect 9999 16949 10011 16983
rect 9953 16943 10011 16949
rect 10778 16940 10784 16992
rect 10836 16980 10842 16992
rect 11609 16983 11667 16989
rect 11609 16980 11621 16983
rect 10836 16952 11621 16980
rect 10836 16940 10842 16952
rect 11609 16949 11621 16952
rect 11655 16980 11667 16983
rect 11698 16980 11704 16992
rect 11655 16952 11704 16980
rect 11655 16949 11667 16952
rect 11609 16943 11667 16949
rect 11698 16940 11704 16952
rect 11756 16940 11762 16992
rect 11882 16940 11888 16992
rect 11940 16980 11946 16992
rect 12437 16983 12495 16989
rect 12437 16980 12449 16983
rect 11940 16952 12449 16980
rect 11940 16940 11946 16952
rect 12437 16949 12449 16952
rect 12483 16949 12495 16983
rect 12820 16980 12848 17020
rect 13817 17017 13829 17051
rect 13863 17048 13875 17051
rect 14550 17048 14556 17060
rect 13863 17020 14556 17048
rect 13863 17017 13875 17020
rect 13817 17011 13875 17017
rect 14550 17008 14556 17020
rect 14608 17008 14614 17060
rect 15764 17048 15792 17079
rect 16022 17076 16028 17128
rect 16080 17116 16086 17128
rect 16301 17119 16359 17125
rect 16301 17116 16313 17119
rect 16080 17088 16313 17116
rect 16080 17076 16086 17088
rect 16301 17085 16313 17088
rect 16347 17085 16359 17119
rect 16301 17079 16359 17085
rect 16568 17119 16626 17125
rect 16568 17085 16580 17119
rect 16614 17116 16626 17119
rect 18046 17116 18052 17128
rect 16614 17088 18052 17116
rect 16614 17085 16626 17088
rect 16568 17079 16626 17085
rect 18046 17076 18052 17088
rect 18104 17076 18110 17128
rect 18708 17116 18736 17147
rect 19150 17116 19156 17128
rect 18708 17088 19156 17116
rect 19150 17076 19156 17088
rect 19208 17076 19214 17128
rect 19518 17076 19524 17128
rect 19576 17116 19582 17128
rect 19613 17119 19671 17125
rect 19613 17116 19625 17119
rect 19576 17088 19625 17116
rect 19576 17076 19582 17088
rect 19613 17085 19625 17088
rect 19659 17085 19671 17119
rect 19720 17116 19748 17156
rect 19794 17144 19800 17196
rect 19852 17184 19858 17196
rect 19852 17156 19897 17184
rect 19852 17144 19858 17156
rect 20533 17119 20591 17125
rect 20533 17116 20545 17119
rect 19720 17088 20545 17116
rect 19613 17079 19671 17085
rect 20533 17085 20545 17088
rect 20579 17085 20591 17119
rect 20533 17079 20591 17085
rect 17770 17048 17776 17060
rect 15764 17020 17776 17048
rect 17770 17008 17776 17020
rect 17828 17008 17834 17060
rect 17862 17008 17868 17060
rect 17920 17048 17926 17060
rect 20070 17048 20076 17060
rect 17920 17020 20076 17048
rect 17920 17008 17926 17020
rect 20070 17008 20076 17020
rect 20128 17008 20134 17060
rect 16758 16980 16764 16992
rect 12820 16952 16764 16980
rect 12437 16943 12495 16949
rect 16758 16940 16764 16952
rect 16816 16940 16822 16992
rect 17678 16980 17684 16992
rect 17639 16952 17684 16980
rect 17678 16940 17684 16952
rect 17736 16940 17742 16992
rect 18414 16980 18420 16992
rect 18375 16952 18420 16980
rect 18414 16940 18420 16952
rect 18472 16940 18478 16992
rect 18509 16983 18567 16989
rect 18509 16949 18521 16983
rect 18555 16980 18567 16983
rect 19610 16980 19616 16992
rect 18555 16952 19616 16980
rect 18555 16949 18567 16952
rect 18509 16943 18567 16949
rect 19610 16940 19616 16952
rect 19668 16940 19674 16992
rect 19705 16983 19763 16989
rect 19705 16949 19717 16983
rect 19751 16980 19763 16983
rect 20254 16980 20260 16992
rect 19751 16952 20260 16980
rect 19751 16949 19763 16952
rect 19705 16943 19763 16949
rect 20254 16940 20260 16952
rect 20312 16940 20318 16992
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 3697 16779 3755 16785
rect 3697 16745 3709 16779
rect 3743 16745 3755 16779
rect 3697 16739 3755 16745
rect 3712 16708 3740 16739
rect 4062 16736 4068 16788
rect 4120 16776 4126 16788
rect 5442 16776 5448 16788
rect 4120 16748 4844 16776
rect 5403 16748 5448 16776
rect 4120 16736 4126 16748
rect 4332 16711 4390 16717
rect 4332 16708 4344 16711
rect 3712 16680 4344 16708
rect 4332 16677 4344 16680
rect 4378 16708 4390 16711
rect 4706 16708 4712 16720
rect 4378 16680 4712 16708
rect 4378 16677 4390 16680
rect 4332 16671 4390 16677
rect 4706 16668 4712 16680
rect 4764 16668 4770 16720
rect 4816 16708 4844 16748
rect 5442 16736 5448 16748
rect 5500 16736 5506 16788
rect 7098 16776 7104 16788
rect 5552 16748 7104 16776
rect 5552 16708 5580 16748
rect 7098 16736 7104 16748
rect 7156 16736 7162 16788
rect 7469 16779 7527 16785
rect 7469 16745 7481 16779
rect 7515 16776 7527 16779
rect 7742 16776 7748 16788
rect 7515 16748 7748 16776
rect 7515 16745 7527 16748
rect 7469 16739 7527 16745
rect 7742 16736 7748 16748
rect 7800 16736 7806 16788
rect 9490 16736 9496 16788
rect 9548 16776 9554 16788
rect 9769 16779 9827 16785
rect 9769 16776 9781 16779
rect 9548 16748 9781 16776
rect 9548 16736 9554 16748
rect 9769 16745 9781 16748
rect 9815 16776 9827 16779
rect 9861 16779 9919 16785
rect 9861 16776 9873 16779
rect 9815 16748 9873 16776
rect 9815 16745 9827 16748
rect 9769 16739 9827 16745
rect 9861 16745 9873 16748
rect 9907 16745 9919 16779
rect 9861 16739 9919 16745
rect 10505 16779 10563 16785
rect 10505 16745 10517 16779
rect 10551 16776 10563 16779
rect 11606 16776 11612 16788
rect 10551 16748 11612 16776
rect 10551 16745 10563 16748
rect 10505 16739 10563 16745
rect 11606 16736 11612 16748
rect 11664 16736 11670 16788
rect 11882 16776 11888 16788
rect 11843 16748 11888 16776
rect 11882 16736 11888 16748
rect 11940 16736 11946 16788
rect 11977 16779 12035 16785
rect 11977 16745 11989 16779
rect 12023 16776 12035 16779
rect 12342 16776 12348 16788
rect 12023 16748 12348 16776
rect 12023 16745 12035 16748
rect 11977 16739 12035 16745
rect 12342 16736 12348 16748
rect 12400 16736 12406 16788
rect 12529 16779 12587 16785
rect 12529 16745 12541 16779
rect 12575 16776 12587 16779
rect 13354 16776 13360 16788
rect 12575 16748 13360 16776
rect 12575 16745 12587 16748
rect 12529 16739 12587 16745
rect 13354 16736 13360 16748
rect 13412 16736 13418 16788
rect 14090 16776 14096 16788
rect 14051 16748 14096 16776
rect 14090 16736 14096 16748
rect 14148 16736 14154 16788
rect 14550 16776 14556 16788
rect 14511 16748 14556 16776
rect 14550 16736 14556 16748
rect 14608 16736 14614 16788
rect 14844 16748 15792 16776
rect 4816 16680 5580 16708
rect 6356 16711 6414 16717
rect 6356 16677 6368 16711
rect 6402 16708 6414 16711
rect 7374 16708 7380 16720
rect 6402 16680 7380 16708
rect 6402 16677 6414 16680
rect 6356 16671 6414 16677
rect 7374 16668 7380 16680
rect 7432 16668 7438 16720
rect 7760 16708 7788 16736
rect 7990 16711 8048 16717
rect 7990 16708 8002 16711
rect 7760 16680 8002 16708
rect 7990 16677 8002 16680
rect 8036 16677 8048 16711
rect 7990 16671 8048 16677
rect 9122 16668 9128 16720
rect 9180 16708 9186 16720
rect 13633 16711 13691 16717
rect 9180 16680 11008 16708
rect 9180 16668 9186 16680
rect 1762 16640 1768 16652
rect 1723 16612 1768 16640
rect 1762 16600 1768 16612
rect 1820 16600 1826 16652
rect 2584 16643 2642 16649
rect 2584 16609 2596 16643
rect 2630 16640 2642 16643
rect 3142 16640 3148 16652
rect 2630 16612 3148 16640
rect 2630 16609 2642 16612
rect 2584 16603 2642 16609
rect 3142 16600 3148 16612
rect 3200 16600 3206 16652
rect 4065 16643 4123 16649
rect 4065 16609 4077 16643
rect 4111 16640 4123 16643
rect 4614 16640 4620 16652
rect 4111 16612 4620 16640
rect 4111 16609 4123 16612
rect 4065 16603 4123 16609
rect 4614 16600 4620 16612
rect 4672 16600 4678 16652
rect 6089 16643 6147 16649
rect 6089 16609 6101 16643
rect 6135 16640 6147 16643
rect 6135 16612 7512 16640
rect 6135 16609 6147 16612
rect 6089 16603 6147 16609
rect 7484 16584 7512 16612
rect 7650 16600 7656 16652
rect 7708 16640 7714 16652
rect 10045 16643 10103 16649
rect 10045 16640 10057 16643
rect 7708 16612 10057 16640
rect 7708 16600 7714 16612
rect 10045 16609 10057 16612
rect 10091 16609 10103 16643
rect 10870 16640 10876 16652
rect 10831 16612 10876 16640
rect 10045 16603 10103 16609
rect 10870 16600 10876 16612
rect 10928 16600 10934 16652
rect 10980 16640 11008 16680
rect 13633 16677 13645 16711
rect 13679 16708 13691 16711
rect 14734 16708 14740 16720
rect 13679 16680 14740 16708
rect 13679 16677 13691 16680
rect 13633 16671 13691 16677
rect 14734 16668 14740 16680
rect 14792 16668 14798 16720
rect 10980 16612 11560 16640
rect 2314 16572 2320 16584
rect 2275 16544 2320 16572
rect 2314 16532 2320 16544
rect 2372 16532 2378 16584
rect 7466 16532 7472 16584
rect 7524 16572 7530 16584
rect 7745 16575 7803 16581
rect 7745 16572 7757 16575
rect 7524 16544 7757 16572
rect 7524 16532 7530 16544
rect 7745 16541 7757 16544
rect 7791 16541 7803 16575
rect 7745 16535 7803 16541
rect 1946 16504 1952 16516
rect 1907 16476 1952 16504
rect 1946 16464 1952 16476
rect 2004 16464 2010 16516
rect 2222 16396 2228 16448
rect 2280 16436 2286 16448
rect 3418 16436 3424 16448
rect 2280 16408 3424 16436
rect 2280 16396 2286 16408
rect 3418 16396 3424 16408
rect 3476 16436 3482 16448
rect 4062 16436 4068 16448
rect 3476 16408 4068 16436
rect 3476 16396 3482 16408
rect 4062 16396 4068 16408
rect 4120 16396 4126 16448
rect 7760 16436 7788 16535
rect 9030 16532 9036 16584
rect 9088 16572 9094 16584
rect 10965 16575 11023 16581
rect 10965 16572 10977 16575
rect 9088 16544 10977 16572
rect 9088 16532 9094 16544
rect 10965 16541 10977 16544
rect 11011 16541 11023 16575
rect 11146 16572 11152 16584
rect 11107 16544 11152 16572
rect 10965 16535 11023 16541
rect 11146 16532 11152 16544
rect 11204 16532 11210 16584
rect 9125 16507 9183 16513
rect 9125 16473 9137 16507
rect 9171 16504 9183 16507
rect 9858 16504 9864 16516
rect 9171 16476 9864 16504
rect 9171 16473 9183 16476
rect 9125 16467 9183 16473
rect 9858 16464 9864 16476
rect 9916 16464 9922 16516
rect 11532 16513 11560 16612
rect 11698 16600 11704 16652
rect 11756 16640 11762 16652
rect 12897 16643 12955 16649
rect 12897 16640 12909 16643
rect 11756 16612 12909 16640
rect 11756 16600 11762 16612
rect 12897 16609 12909 16612
rect 12943 16609 12955 16643
rect 12897 16603 12955 16609
rect 12989 16643 13047 16649
rect 12989 16609 13001 16643
rect 13035 16640 13047 16643
rect 13722 16640 13728 16652
rect 13035 16612 13728 16640
rect 13035 16609 13047 16612
rect 12989 16603 13047 16609
rect 13722 16600 13728 16612
rect 13780 16640 13786 16652
rect 13780 16612 14044 16640
rect 13780 16600 13786 16612
rect 12161 16575 12219 16581
rect 12161 16541 12173 16575
rect 12207 16572 12219 16575
rect 12342 16572 12348 16584
rect 12207 16544 12348 16572
rect 12207 16541 12219 16544
rect 12161 16535 12219 16541
rect 12342 16532 12348 16544
rect 12400 16532 12406 16584
rect 13173 16575 13231 16581
rect 13173 16541 13185 16575
rect 13219 16541 13231 16575
rect 14016 16572 14044 16612
rect 14090 16600 14096 16652
rect 14148 16640 14154 16652
rect 14461 16643 14519 16649
rect 14461 16640 14473 16643
rect 14148 16612 14473 16640
rect 14148 16600 14154 16612
rect 14461 16609 14473 16612
rect 14507 16609 14519 16643
rect 14844 16640 14872 16748
rect 14918 16668 14924 16720
rect 14976 16708 14982 16720
rect 15657 16711 15715 16717
rect 15657 16708 15669 16711
rect 14976 16680 15669 16708
rect 14976 16668 14982 16680
rect 15657 16677 15669 16680
rect 15703 16677 15715 16711
rect 15764 16708 15792 16748
rect 18046 16736 18052 16788
rect 18104 16776 18110 16788
rect 19150 16776 19156 16788
rect 18104 16748 19156 16776
rect 18104 16736 18110 16748
rect 19150 16736 19156 16748
rect 19208 16776 19214 16788
rect 19613 16779 19671 16785
rect 19613 16776 19625 16779
rect 19208 16748 19625 16776
rect 19208 16736 19214 16748
rect 19613 16745 19625 16748
rect 19659 16745 19671 16779
rect 19613 16739 19671 16745
rect 16666 16708 16672 16720
rect 15764 16680 16672 16708
rect 15657 16671 15715 16677
rect 16666 16668 16672 16680
rect 16724 16668 16730 16720
rect 16942 16668 16948 16720
rect 17000 16708 17006 16720
rect 18966 16708 18972 16720
rect 17000 16680 18972 16708
rect 17000 16668 17006 16680
rect 18966 16668 18972 16680
rect 19024 16668 19030 16720
rect 19334 16668 19340 16720
rect 19392 16708 19398 16720
rect 20165 16711 20223 16717
rect 20165 16708 20177 16711
rect 19392 16680 20177 16708
rect 19392 16668 19398 16680
rect 20165 16677 20177 16680
rect 20211 16677 20223 16711
rect 20165 16671 20223 16677
rect 14461 16603 14519 16609
rect 14568 16612 14872 16640
rect 14568 16572 14596 16612
rect 15194 16600 15200 16652
rect 15252 16640 15258 16652
rect 15749 16643 15807 16649
rect 15749 16640 15761 16643
rect 15252 16612 15761 16640
rect 15252 16600 15258 16612
rect 15749 16609 15761 16612
rect 15795 16609 15807 16643
rect 15749 16603 15807 16609
rect 16853 16643 16911 16649
rect 16853 16609 16865 16643
rect 16899 16640 16911 16643
rect 17034 16640 17040 16652
rect 16899 16612 17040 16640
rect 16899 16609 16911 16612
rect 16853 16603 16911 16609
rect 17034 16600 17040 16612
rect 17092 16600 17098 16652
rect 17218 16600 17224 16652
rect 17276 16640 17282 16652
rect 17497 16643 17555 16649
rect 17276 16612 17448 16640
rect 17276 16600 17282 16612
rect 14016 16544 14596 16572
rect 14737 16575 14795 16581
rect 13173 16535 13231 16541
rect 14737 16541 14749 16575
rect 14783 16572 14795 16575
rect 15470 16572 15476 16584
rect 14783 16544 15476 16572
rect 14783 16541 14795 16544
rect 14737 16535 14795 16541
rect 11517 16507 11575 16513
rect 11517 16473 11529 16507
rect 11563 16473 11575 16507
rect 11517 16467 11575 16473
rect 12802 16464 12808 16516
rect 12860 16504 12866 16516
rect 13188 16504 13216 16535
rect 15470 16532 15476 16544
rect 15528 16532 15534 16584
rect 15841 16575 15899 16581
rect 15841 16541 15853 16575
rect 15887 16541 15899 16575
rect 15841 16535 15899 16541
rect 13538 16504 13544 16516
rect 12860 16476 13544 16504
rect 12860 16464 12866 16476
rect 13538 16464 13544 16476
rect 13596 16504 13602 16516
rect 15102 16504 15108 16516
rect 13596 16476 15108 16504
rect 13596 16464 13602 16476
rect 15102 16464 15108 16476
rect 15160 16504 15166 16516
rect 15856 16504 15884 16535
rect 16758 16532 16764 16584
rect 16816 16572 16822 16584
rect 16945 16575 17003 16581
rect 16945 16572 16957 16575
rect 16816 16544 16957 16572
rect 16816 16532 16822 16544
rect 16945 16541 16957 16544
rect 16991 16541 17003 16575
rect 17126 16572 17132 16584
rect 17087 16544 17132 16572
rect 16945 16535 17003 16541
rect 17126 16532 17132 16544
rect 17184 16532 17190 16584
rect 17420 16572 17448 16612
rect 17497 16609 17509 16643
rect 17543 16640 17555 16643
rect 17954 16640 17960 16652
rect 17543 16612 17960 16640
rect 17543 16609 17555 16612
rect 17497 16603 17555 16609
rect 17954 16600 17960 16612
rect 18012 16600 18018 16652
rect 18500 16643 18558 16649
rect 18500 16609 18512 16643
rect 18546 16640 18558 16643
rect 19242 16640 19248 16652
rect 18546 16612 19248 16640
rect 18546 16609 18558 16612
rect 18500 16603 18558 16609
rect 19242 16600 19248 16612
rect 19300 16600 19306 16652
rect 19889 16643 19947 16649
rect 19889 16640 19901 16643
rect 19352 16612 19901 16640
rect 18233 16575 18291 16581
rect 17420 16544 17724 16572
rect 15160 16476 15884 16504
rect 15160 16464 15166 16476
rect 9766 16436 9772 16448
rect 7760 16408 9772 16436
rect 9766 16396 9772 16408
rect 9824 16396 9830 16448
rect 12434 16396 12440 16448
rect 12492 16436 12498 16448
rect 13998 16436 14004 16448
rect 12492 16408 14004 16436
rect 12492 16396 12498 16408
rect 13998 16396 14004 16408
rect 14056 16396 14062 16448
rect 15286 16436 15292 16448
rect 15247 16408 15292 16436
rect 15286 16396 15292 16408
rect 15344 16396 15350 16448
rect 16485 16439 16543 16445
rect 16485 16405 16497 16439
rect 16531 16436 16543 16439
rect 17402 16436 17408 16448
rect 16531 16408 17408 16436
rect 16531 16405 16543 16408
rect 16485 16399 16543 16405
rect 17402 16396 17408 16408
rect 17460 16396 17466 16448
rect 17696 16445 17724 16544
rect 18233 16541 18245 16575
rect 18279 16541 18291 16575
rect 18233 16535 18291 16541
rect 17681 16439 17739 16445
rect 17681 16405 17693 16439
rect 17727 16405 17739 16439
rect 18248 16436 18276 16535
rect 18598 16436 18604 16448
rect 18248 16408 18604 16436
rect 17681 16399 17739 16405
rect 18598 16396 18604 16408
rect 18656 16436 18662 16448
rect 18874 16436 18880 16448
rect 18656 16408 18880 16436
rect 18656 16396 18662 16408
rect 18874 16396 18880 16408
rect 18932 16396 18938 16448
rect 19150 16396 19156 16448
rect 19208 16436 19214 16448
rect 19352 16436 19380 16612
rect 19889 16609 19901 16612
rect 19935 16609 19947 16643
rect 19889 16603 19947 16609
rect 19978 16600 19984 16652
rect 20036 16640 20042 16652
rect 20901 16643 20959 16649
rect 20901 16640 20913 16643
rect 20036 16612 20913 16640
rect 20036 16600 20042 16612
rect 20901 16609 20913 16612
rect 20947 16609 20959 16643
rect 20901 16603 20959 16609
rect 19208 16408 19380 16436
rect 19208 16396 19214 16408
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 4246 16192 4252 16244
rect 4304 16232 4310 16244
rect 4341 16235 4399 16241
rect 4341 16232 4353 16235
rect 4304 16204 4353 16232
rect 4304 16192 4310 16204
rect 4341 16201 4353 16204
rect 4387 16201 4399 16235
rect 4341 16195 4399 16201
rect 6825 16235 6883 16241
rect 6825 16201 6837 16235
rect 6871 16232 6883 16235
rect 7558 16232 7564 16244
rect 6871 16204 7564 16232
rect 6871 16201 6883 16204
rect 6825 16195 6883 16201
rect 7558 16192 7564 16204
rect 7616 16192 7622 16244
rect 8941 16235 8999 16241
rect 8941 16201 8953 16235
rect 8987 16232 8999 16235
rect 9030 16232 9036 16244
rect 8987 16204 9036 16232
rect 8987 16201 8999 16204
rect 8941 16195 8999 16201
rect 9030 16192 9036 16204
rect 9088 16192 9094 16244
rect 11146 16192 11152 16244
rect 11204 16232 11210 16244
rect 11333 16235 11391 16241
rect 11333 16232 11345 16235
rect 11204 16204 11345 16232
rect 11204 16192 11210 16204
rect 11333 16201 11345 16204
rect 11379 16201 11391 16235
rect 13814 16232 13820 16244
rect 13775 16204 13820 16232
rect 11333 16195 11391 16201
rect 13814 16192 13820 16204
rect 13872 16192 13878 16244
rect 15470 16232 15476 16244
rect 15431 16204 15476 16232
rect 15470 16192 15476 16204
rect 15528 16192 15534 16244
rect 16390 16192 16396 16244
rect 16448 16232 16454 16244
rect 17586 16232 17592 16244
rect 16448 16204 16712 16232
rect 17547 16204 17592 16232
rect 16448 16192 16454 16204
rect 2593 16167 2651 16173
rect 2593 16133 2605 16167
rect 2639 16164 2651 16167
rect 4798 16164 4804 16176
rect 2639 16136 4804 16164
rect 2639 16133 2651 16136
rect 2593 16127 2651 16133
rect 4798 16124 4804 16136
rect 4856 16124 4862 16176
rect 6914 16124 6920 16176
rect 6972 16164 6978 16176
rect 12434 16164 12440 16176
rect 6972 16136 8616 16164
rect 6972 16124 6978 16136
rect 3142 16096 3148 16108
rect 3103 16068 3148 16096
rect 3142 16056 3148 16068
rect 3200 16096 3206 16108
rect 4062 16096 4068 16108
rect 3200 16068 4068 16096
rect 3200 16056 3206 16068
rect 4062 16056 4068 16068
rect 4120 16096 4126 16108
rect 4893 16099 4951 16105
rect 4893 16096 4905 16099
rect 4120 16068 4905 16096
rect 4120 16056 4126 16068
rect 4893 16065 4905 16068
rect 4939 16065 4951 16099
rect 7374 16096 7380 16108
rect 7335 16068 7380 16096
rect 4893 16059 4951 16065
rect 7374 16056 7380 16068
rect 7432 16056 7438 16108
rect 7742 16056 7748 16108
rect 7800 16096 7806 16108
rect 8202 16096 8208 16108
rect 7800 16068 8208 16096
rect 7800 16056 7806 16068
rect 8202 16056 8208 16068
rect 8260 16096 8266 16108
rect 8389 16099 8447 16105
rect 8389 16096 8401 16099
rect 8260 16068 8401 16096
rect 8260 16056 8266 16068
rect 8389 16065 8401 16068
rect 8435 16065 8447 16099
rect 8389 16059 8447 16065
rect 1765 16031 1823 16037
rect 1765 15997 1777 16031
rect 1811 16028 1823 16031
rect 2222 16028 2228 16040
rect 1811 16000 2228 16028
rect 1811 15997 1823 16000
rect 1765 15991 1823 15997
rect 2222 15988 2228 16000
rect 2280 15988 2286 16040
rect 2961 16031 3019 16037
rect 2961 15997 2973 16031
rect 3007 16028 3019 16031
rect 3234 16028 3240 16040
rect 3007 16000 3240 16028
rect 3007 15997 3019 16000
rect 2961 15991 3019 15997
rect 3234 15988 3240 16000
rect 3292 15988 3298 16040
rect 7098 15988 7104 16040
rect 7156 16028 7162 16040
rect 8297 16031 8355 16037
rect 8297 16028 8309 16031
rect 7156 16000 8309 16028
rect 7156 15988 7162 16000
rect 8297 15997 8309 16000
rect 8343 15997 8355 16031
rect 8297 15991 8355 15997
rect 4709 15963 4767 15969
rect 4709 15929 4721 15963
rect 4755 15960 4767 15963
rect 6086 15960 6092 15972
rect 4755 15932 6092 15960
rect 4755 15929 4767 15932
rect 4709 15923 4767 15929
rect 6086 15920 6092 15932
rect 6144 15920 6150 15972
rect 7193 15963 7251 15969
rect 7193 15929 7205 15963
rect 7239 15960 7251 15963
rect 7239 15932 7880 15960
rect 7239 15929 7251 15932
rect 7193 15923 7251 15929
rect 1394 15852 1400 15904
rect 1452 15892 1458 15904
rect 1949 15895 2007 15901
rect 1949 15892 1961 15895
rect 1452 15864 1961 15892
rect 1452 15852 1458 15864
rect 1949 15861 1961 15864
rect 1995 15861 2007 15895
rect 1949 15855 2007 15861
rect 3050 15852 3056 15904
rect 3108 15892 3114 15904
rect 4801 15895 4859 15901
rect 3108 15864 3153 15892
rect 3108 15852 3114 15864
rect 4801 15861 4813 15895
rect 4847 15892 4859 15895
rect 4982 15892 4988 15904
rect 4847 15864 4988 15892
rect 4847 15861 4859 15864
rect 4801 15855 4859 15861
rect 4982 15852 4988 15864
rect 5040 15852 5046 15904
rect 7285 15895 7343 15901
rect 7285 15861 7297 15895
rect 7331 15892 7343 15895
rect 7374 15892 7380 15904
rect 7331 15864 7380 15892
rect 7331 15861 7343 15864
rect 7285 15855 7343 15861
rect 7374 15852 7380 15864
rect 7432 15852 7438 15904
rect 7852 15901 7880 15932
rect 7837 15895 7895 15901
rect 7837 15861 7849 15895
rect 7883 15861 7895 15895
rect 8202 15892 8208 15904
rect 8163 15864 8208 15892
rect 7837 15855 7895 15861
rect 8202 15852 8208 15864
rect 8260 15852 8266 15904
rect 8588 15892 8616 16136
rect 11900 16136 12440 16164
rect 9490 16096 9496 16108
rect 9451 16068 9496 16096
rect 9490 16056 9496 16068
rect 9548 16056 9554 16108
rect 9766 16056 9772 16108
rect 9824 16096 9830 16108
rect 11900 16105 11928 16136
rect 12434 16124 12440 16136
rect 12492 16124 12498 16176
rect 9953 16099 10011 16105
rect 9953 16096 9965 16099
rect 9824 16068 9965 16096
rect 9824 16056 9830 16068
rect 9953 16065 9965 16068
rect 9999 16065 10011 16099
rect 9953 16059 10011 16065
rect 11885 16099 11943 16105
rect 11885 16065 11897 16099
rect 11931 16065 11943 16099
rect 13832 16096 13860 16192
rect 15488 16096 15516 16192
rect 16684 16164 16712 16204
rect 17586 16192 17592 16204
rect 17644 16192 17650 16244
rect 19242 16192 19248 16244
rect 19300 16232 19306 16244
rect 20349 16235 20407 16241
rect 20349 16232 20361 16235
rect 19300 16204 20361 16232
rect 19300 16192 19306 16204
rect 20349 16201 20361 16204
rect 20395 16201 20407 16235
rect 20349 16195 20407 16201
rect 18966 16164 18972 16176
rect 16684 16136 18972 16164
rect 18966 16124 18972 16136
rect 19024 16124 19030 16176
rect 13832 16068 14228 16096
rect 15488 16068 15884 16096
rect 11885 16059 11943 16065
rect 8938 15988 8944 16040
rect 8996 16028 9002 16040
rect 9309 16031 9367 16037
rect 9309 16028 9321 16031
rect 8996 16000 9321 16028
rect 8996 15988 9002 16000
rect 9309 15997 9321 16000
rect 9355 15997 9367 16031
rect 9309 15991 9367 15997
rect 9398 15988 9404 16040
rect 9456 16028 9462 16040
rect 9456 16000 9501 16028
rect 9456 15988 9462 16000
rect 10042 15988 10048 16040
rect 10100 16028 10106 16040
rect 10209 16031 10267 16037
rect 10209 16028 10221 16031
rect 10100 16000 10221 16028
rect 10100 15988 10106 16000
rect 10209 15997 10221 16000
rect 10255 15997 10267 16031
rect 11606 16028 11612 16040
rect 11567 16000 11612 16028
rect 10209 15991 10267 15997
rect 11606 15988 11612 16000
rect 11664 15988 11670 16040
rect 12434 15988 12440 16040
rect 12492 16028 12498 16040
rect 13078 16028 13084 16040
rect 12492 16000 13084 16028
rect 12492 15988 12498 16000
rect 13078 15988 13084 16000
rect 13136 16028 13142 16040
rect 13538 16028 13544 16040
rect 13136 16000 13544 16028
rect 13136 15988 13142 16000
rect 13538 15988 13544 16000
rect 13596 16028 13602 16040
rect 14093 16031 14151 16037
rect 14093 16028 14105 16031
rect 13596 16000 14105 16028
rect 13596 15988 13602 16000
rect 14093 15997 14105 16000
rect 14139 15997 14151 16031
rect 14200 16028 14228 16068
rect 14366 16037 14372 16040
rect 14349 16031 14372 16037
rect 14349 16028 14361 16031
rect 14200 16000 14361 16028
rect 14093 15991 14151 15997
rect 14349 15997 14361 16000
rect 14424 16028 14430 16040
rect 15749 16031 15807 16037
rect 14424 16000 14497 16028
rect 14349 15991 14372 15997
rect 11974 15960 11980 15972
rect 11532 15932 11980 15960
rect 11532 15892 11560 15932
rect 11974 15920 11980 15932
rect 12032 15920 12038 15972
rect 12704 15963 12762 15969
rect 12704 15929 12716 15963
rect 12750 15960 12762 15963
rect 12802 15960 12808 15972
rect 12750 15932 12808 15960
rect 12750 15929 12762 15932
rect 12704 15923 12762 15929
rect 12802 15920 12808 15932
rect 12860 15920 12866 15972
rect 14108 15960 14136 15991
rect 14366 15988 14372 15991
rect 14424 15988 14430 16000
rect 15749 15997 15761 16031
rect 15795 15997 15807 16031
rect 15856 16028 15884 16068
rect 16850 16056 16856 16108
rect 16908 16096 16914 16108
rect 17678 16096 17684 16108
rect 16908 16068 17684 16096
rect 16908 16056 16914 16068
rect 17678 16056 17684 16068
rect 17736 16056 17742 16108
rect 17954 16056 17960 16108
rect 18012 16096 18018 16108
rect 18233 16099 18291 16105
rect 18233 16096 18245 16099
rect 18012 16068 18245 16096
rect 18012 16056 18018 16068
rect 18233 16065 18245 16068
rect 18279 16065 18291 16099
rect 18233 16059 18291 16065
rect 16005 16031 16063 16037
rect 16005 16028 16017 16031
rect 15856 16000 16017 16028
rect 15749 15991 15807 15997
rect 16005 15997 16017 16000
rect 16051 15997 16063 16031
rect 16005 15991 16063 15997
rect 17405 16031 17463 16037
rect 17405 15997 17417 16031
rect 17451 16028 17463 16031
rect 17494 16028 17500 16040
rect 17451 16000 17500 16028
rect 17451 15997 17463 16000
rect 17405 15991 17463 15997
rect 15764 15960 15792 15991
rect 17494 15988 17500 16000
rect 17552 15988 17558 16040
rect 18049 16031 18107 16037
rect 18049 15997 18061 16031
rect 18095 15997 18107 16031
rect 18049 15991 18107 15997
rect 14108 15932 15792 15960
rect 17954 15920 17960 15972
rect 18012 15960 18018 15972
rect 18064 15960 18092 15991
rect 18598 15988 18604 16040
rect 18656 16028 18662 16040
rect 18969 16031 19027 16037
rect 18969 16028 18981 16031
rect 18656 16000 18981 16028
rect 18656 15988 18662 16000
rect 18969 15997 18981 16000
rect 19015 15997 19027 16031
rect 18969 15991 19027 15997
rect 19610 15988 19616 16040
rect 19668 16028 19674 16040
rect 20625 16031 20683 16037
rect 20625 16028 20637 16031
rect 19668 16000 20637 16028
rect 19668 15988 19674 16000
rect 20625 15997 20637 16000
rect 20671 15997 20683 16031
rect 20625 15991 20683 15997
rect 18012 15932 18092 15960
rect 19236 15963 19294 15969
rect 18012 15920 18018 15932
rect 19236 15929 19248 15963
rect 19282 15960 19294 15963
rect 19426 15960 19432 15972
rect 19282 15932 19432 15960
rect 19282 15929 19294 15932
rect 19236 15923 19294 15929
rect 19426 15920 19432 15932
rect 19484 15920 19490 15972
rect 20901 15963 20959 15969
rect 20901 15929 20913 15963
rect 20947 15929 20959 15963
rect 20901 15923 20959 15929
rect 17126 15892 17132 15904
rect 8588 15864 11560 15892
rect 17087 15864 17132 15892
rect 17126 15852 17132 15864
rect 17184 15852 17190 15904
rect 17310 15852 17316 15904
rect 17368 15892 17374 15904
rect 20916 15892 20944 15923
rect 17368 15864 20944 15892
rect 17368 15852 17374 15864
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 1946 15688 1952 15700
rect 1907 15660 1952 15688
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 2501 15691 2559 15697
rect 2501 15657 2513 15691
rect 2547 15688 2559 15691
rect 3050 15688 3056 15700
rect 2547 15660 3056 15688
rect 2547 15657 2559 15660
rect 2501 15651 2559 15657
rect 3050 15648 3056 15660
rect 3108 15648 3114 15700
rect 3878 15648 3884 15700
rect 3936 15688 3942 15700
rect 4065 15691 4123 15697
rect 4065 15688 4077 15691
rect 3936 15660 4077 15688
rect 3936 15648 3942 15660
rect 4065 15657 4077 15660
rect 4111 15657 4123 15691
rect 4065 15651 4123 15657
rect 4433 15691 4491 15697
rect 4433 15657 4445 15691
rect 4479 15688 4491 15691
rect 5077 15691 5135 15697
rect 5077 15688 5089 15691
rect 4479 15660 5089 15688
rect 4479 15657 4491 15660
rect 4433 15651 4491 15657
rect 5077 15657 5089 15660
rect 5123 15657 5135 15691
rect 5077 15651 5135 15657
rect 5534 15648 5540 15700
rect 5592 15688 5598 15700
rect 6089 15691 6147 15697
rect 6089 15688 6101 15691
rect 5592 15660 6101 15688
rect 5592 15648 5598 15660
rect 6089 15657 6101 15660
rect 6135 15657 6147 15691
rect 7374 15688 7380 15700
rect 7335 15660 7380 15688
rect 6089 15651 6147 15657
rect 7374 15648 7380 15660
rect 7432 15648 7438 15700
rect 7558 15648 7564 15700
rect 7616 15688 7622 15700
rect 7745 15691 7803 15697
rect 7745 15688 7757 15691
rect 7616 15660 7757 15688
rect 7616 15648 7622 15660
rect 7745 15657 7757 15660
rect 7791 15657 7803 15691
rect 7745 15651 7803 15657
rect 8573 15691 8631 15697
rect 8573 15657 8585 15691
rect 8619 15657 8631 15691
rect 8573 15651 8631 15657
rect 8941 15691 8999 15697
rect 8941 15657 8953 15691
rect 8987 15688 8999 15691
rect 9582 15688 9588 15700
rect 8987 15660 9588 15688
rect 8987 15657 8999 15660
rect 8941 15651 8999 15657
rect 2866 15620 2872 15632
rect 2827 15592 2872 15620
rect 2866 15580 2872 15592
rect 2924 15580 2930 15632
rect 2961 15623 3019 15629
rect 2961 15589 2973 15623
rect 3007 15620 3019 15623
rect 3418 15620 3424 15632
rect 3007 15592 3424 15620
rect 3007 15589 3019 15592
rect 2961 15583 3019 15589
rect 3418 15580 3424 15592
rect 3476 15580 3482 15632
rect 6917 15623 6975 15629
rect 6917 15589 6929 15623
rect 6963 15620 6975 15623
rect 8202 15620 8208 15632
rect 6963 15592 8208 15620
rect 6963 15589 6975 15592
rect 6917 15583 6975 15589
rect 8202 15580 8208 15592
rect 8260 15580 8266 15632
rect 8588 15620 8616 15651
rect 9582 15648 9588 15660
rect 9640 15648 9646 15700
rect 10321 15691 10379 15697
rect 10321 15657 10333 15691
rect 10367 15688 10379 15691
rect 10870 15688 10876 15700
rect 10367 15660 10876 15688
rect 10367 15657 10379 15660
rect 10321 15651 10379 15657
rect 10870 15648 10876 15660
rect 10928 15648 10934 15700
rect 13449 15691 13507 15697
rect 13449 15688 13461 15691
rect 10980 15660 13461 15688
rect 10980 15620 11008 15660
rect 13449 15657 13461 15660
rect 13495 15657 13507 15691
rect 14090 15688 14096 15700
rect 14051 15660 14096 15688
rect 13449 15651 13507 15657
rect 14090 15648 14096 15660
rect 14148 15648 14154 15700
rect 14461 15691 14519 15697
rect 14461 15657 14473 15691
rect 14507 15688 14519 15691
rect 15286 15688 15292 15700
rect 14507 15660 15292 15688
rect 14507 15657 14519 15660
rect 14461 15651 14519 15657
rect 15286 15648 15292 15660
rect 15344 15648 15350 15700
rect 15657 15691 15715 15697
rect 15657 15657 15669 15691
rect 15703 15688 15715 15691
rect 15703 15660 17356 15688
rect 15703 15657 15715 15660
rect 15657 15651 15715 15657
rect 8588 15592 11008 15620
rect 11348 15592 11836 15620
rect 1765 15555 1823 15561
rect 1765 15521 1777 15555
rect 1811 15521 1823 15555
rect 1765 15515 1823 15521
rect 3513 15555 3571 15561
rect 3513 15521 3525 15555
rect 3559 15552 3571 15555
rect 5445 15555 5503 15561
rect 5445 15552 5457 15555
rect 3559 15524 5457 15552
rect 3559 15521 3571 15524
rect 3513 15515 3571 15521
rect 5445 15521 5457 15524
rect 5491 15521 5503 15555
rect 5445 15515 5503 15521
rect 6273 15555 6331 15561
rect 6273 15521 6285 15555
rect 6319 15552 6331 15555
rect 7650 15552 7656 15564
rect 6319 15524 7656 15552
rect 6319 15521 6331 15524
rect 6273 15515 6331 15521
rect 1780 15348 1808 15515
rect 7650 15512 7656 15524
rect 7708 15512 7714 15564
rect 7742 15512 7748 15564
rect 7800 15552 7806 15564
rect 10686 15552 10692 15564
rect 7800 15524 7972 15552
rect 10647 15524 10692 15552
rect 7800 15512 7806 15524
rect 3145 15487 3203 15493
rect 3145 15453 3157 15487
rect 3191 15484 3203 15487
rect 3234 15484 3240 15496
rect 3191 15456 3240 15484
rect 3191 15453 3203 15456
rect 3145 15447 3203 15453
rect 3234 15444 3240 15456
rect 3292 15444 3298 15496
rect 4154 15444 4160 15496
rect 4212 15484 4218 15496
rect 4525 15487 4583 15493
rect 4525 15484 4537 15487
rect 4212 15456 4537 15484
rect 4212 15444 4218 15456
rect 4525 15453 4537 15456
rect 4571 15453 4583 15487
rect 4706 15484 4712 15496
rect 4667 15456 4712 15484
rect 4525 15447 4583 15453
rect 4706 15444 4712 15456
rect 4764 15444 4770 15496
rect 5350 15444 5356 15496
rect 5408 15484 5414 15496
rect 5537 15487 5595 15493
rect 5537 15484 5549 15487
rect 5408 15456 5549 15484
rect 5408 15444 5414 15456
rect 5537 15453 5549 15456
rect 5583 15453 5595 15487
rect 5537 15447 5595 15453
rect 5629 15487 5687 15493
rect 5629 15453 5641 15487
rect 5675 15453 5687 15487
rect 5629 15447 5687 15453
rect 4062 15376 4068 15428
rect 4120 15416 4126 15428
rect 5644 15416 5672 15447
rect 7282 15444 7288 15496
rect 7340 15484 7346 15496
rect 7944 15493 7972 15524
rect 10686 15512 10692 15524
rect 10744 15512 10750 15564
rect 10781 15555 10839 15561
rect 10781 15521 10793 15555
rect 10827 15552 10839 15555
rect 11238 15552 11244 15564
rect 10827 15524 11244 15552
rect 10827 15521 10839 15524
rect 10781 15515 10839 15521
rect 11238 15512 11244 15524
rect 11296 15512 11302 15564
rect 11348 15561 11376 15592
rect 11333 15555 11391 15561
rect 11333 15521 11345 15555
rect 11379 15521 11391 15555
rect 11589 15555 11647 15561
rect 11589 15552 11601 15555
rect 11333 15515 11391 15521
rect 11440 15524 11601 15552
rect 7837 15487 7895 15493
rect 7837 15484 7849 15487
rect 7340 15456 7849 15484
rect 7340 15444 7346 15456
rect 7837 15453 7849 15456
rect 7883 15453 7895 15487
rect 7837 15447 7895 15453
rect 7929 15487 7987 15493
rect 7929 15453 7941 15487
rect 7975 15453 7987 15487
rect 7929 15447 7987 15453
rect 8478 15444 8484 15496
rect 8536 15484 8542 15496
rect 9030 15484 9036 15496
rect 8536 15456 9036 15484
rect 8536 15444 8542 15456
rect 9030 15444 9036 15456
rect 9088 15444 9094 15496
rect 9217 15487 9275 15493
rect 9217 15453 9229 15487
rect 9263 15453 9275 15487
rect 9217 15447 9275 15453
rect 4120 15388 5672 15416
rect 4120 15376 4126 15388
rect 6178 15376 6184 15428
rect 6236 15416 6242 15428
rect 9232 15416 9260 15447
rect 10042 15444 10048 15496
rect 10100 15484 10106 15496
rect 10873 15487 10931 15493
rect 10873 15484 10885 15487
rect 10100 15456 10885 15484
rect 10100 15444 10106 15456
rect 10873 15453 10885 15456
rect 10919 15453 10931 15487
rect 10873 15447 10931 15453
rect 11146 15444 11152 15496
rect 11204 15484 11210 15496
rect 11440 15484 11468 15524
rect 11589 15521 11601 15524
rect 11635 15521 11647 15555
rect 11808 15552 11836 15592
rect 12618 15580 12624 15632
rect 12676 15620 12682 15632
rect 13357 15623 13415 15629
rect 13357 15620 13369 15623
rect 12676 15592 13369 15620
rect 12676 15580 12682 15592
rect 13357 15589 13369 15592
rect 13403 15589 13415 15623
rect 13357 15583 13415 15589
rect 16292 15623 16350 15629
rect 16292 15589 16304 15623
rect 16338 15620 16350 15623
rect 17126 15620 17132 15632
rect 16338 15592 17132 15620
rect 16338 15589 16350 15592
rect 16292 15583 16350 15589
rect 17126 15580 17132 15592
rect 17184 15580 17190 15632
rect 17328 15620 17356 15660
rect 17402 15648 17408 15700
rect 17460 15688 17466 15700
rect 18141 15691 18199 15697
rect 18141 15688 18153 15691
rect 17460 15660 18153 15688
rect 17460 15648 17466 15660
rect 18141 15657 18153 15660
rect 18187 15657 18199 15691
rect 18690 15688 18696 15700
rect 18651 15660 18696 15688
rect 18141 15651 18199 15657
rect 18690 15648 18696 15660
rect 18748 15648 18754 15700
rect 19061 15691 19119 15697
rect 19061 15657 19073 15691
rect 19107 15688 19119 15691
rect 19978 15688 19984 15700
rect 19107 15660 19984 15688
rect 19107 15657 19119 15660
rect 19061 15651 19119 15657
rect 19978 15648 19984 15660
rect 20036 15648 20042 15700
rect 17862 15620 17868 15632
rect 17328 15592 17868 15620
rect 17862 15580 17868 15592
rect 17920 15580 17926 15632
rect 19518 15620 19524 15632
rect 17972 15592 19524 15620
rect 12434 15552 12440 15564
rect 11808 15524 12440 15552
rect 11589 15515 11647 15521
rect 12434 15512 12440 15524
rect 12492 15512 12498 15564
rect 14366 15512 14372 15564
rect 14424 15552 14430 15564
rect 14424 15524 14688 15552
rect 14424 15512 14430 15524
rect 11204 15456 11468 15484
rect 11204 15444 11210 15456
rect 13170 15444 13176 15496
rect 13228 15484 13234 15496
rect 13541 15487 13599 15493
rect 13541 15484 13553 15487
rect 13228 15456 13553 15484
rect 13228 15444 13234 15456
rect 13541 15453 13553 15456
rect 13587 15453 13599 15487
rect 14550 15484 14556 15496
rect 14511 15456 14556 15484
rect 13541 15447 13599 15453
rect 14550 15444 14556 15456
rect 14608 15444 14614 15496
rect 14660 15493 14688 15524
rect 15194 15512 15200 15564
rect 15252 15552 15258 15564
rect 15473 15555 15531 15561
rect 15473 15552 15485 15555
rect 15252 15524 15485 15552
rect 15252 15512 15258 15524
rect 15473 15521 15485 15524
rect 15519 15521 15531 15555
rect 17972 15552 18000 15592
rect 19518 15580 19524 15592
rect 19576 15580 19582 15632
rect 15473 15515 15531 15521
rect 15856 15524 18000 15552
rect 18049 15555 18107 15561
rect 14645 15487 14703 15493
rect 14645 15453 14657 15487
rect 14691 15453 14703 15487
rect 14645 15447 14703 15453
rect 10410 15416 10416 15428
rect 6236 15388 9168 15416
rect 9232 15388 10416 15416
rect 6236 15376 6242 15388
rect 7558 15348 7564 15360
rect 1780 15320 7564 15348
rect 7558 15308 7564 15320
rect 7616 15308 7622 15360
rect 9140 15348 9168 15388
rect 10410 15376 10416 15388
rect 10468 15376 10474 15428
rect 12713 15419 12771 15425
rect 12713 15385 12725 15419
rect 12759 15416 12771 15419
rect 12802 15416 12808 15428
rect 12759 15388 12808 15416
rect 12759 15385 12771 15388
rect 12713 15379 12771 15385
rect 12802 15376 12808 15388
rect 12860 15376 12866 15428
rect 12989 15419 13047 15425
rect 12989 15385 13001 15419
rect 13035 15416 13047 15419
rect 15856 15416 15884 15524
rect 18049 15521 18061 15555
rect 18095 15552 18107 15555
rect 18874 15552 18880 15564
rect 18095 15524 18880 15552
rect 18095 15521 18107 15524
rect 18049 15515 18107 15521
rect 18874 15512 18880 15524
rect 18932 15512 18938 15564
rect 20070 15552 20076 15564
rect 20031 15524 20076 15552
rect 20070 15512 20076 15524
rect 20128 15512 20134 15564
rect 16022 15484 16028 15496
rect 15983 15456 16028 15484
rect 16022 15444 16028 15456
rect 16080 15444 16086 15496
rect 17862 15484 17868 15496
rect 17420 15456 17868 15484
rect 17034 15416 17040 15428
rect 13035 15388 15884 15416
rect 16960 15388 17040 15416
rect 13035 15385 13047 15388
rect 12989 15379 13047 15385
rect 11698 15348 11704 15360
rect 9140 15320 11704 15348
rect 11698 15308 11704 15320
rect 11756 15308 11762 15360
rect 11974 15308 11980 15360
rect 12032 15348 12038 15360
rect 16960 15348 16988 15388
rect 17034 15376 17040 15388
rect 17092 15376 17098 15428
rect 17420 15425 17448 15456
rect 17862 15444 17868 15456
rect 17920 15484 17926 15496
rect 18233 15487 18291 15493
rect 18233 15484 18245 15487
rect 17920 15456 18245 15484
rect 17920 15444 17926 15456
rect 18233 15453 18245 15456
rect 18279 15453 18291 15487
rect 18233 15447 18291 15453
rect 18690 15444 18696 15496
rect 18748 15484 18754 15496
rect 19153 15487 19211 15493
rect 19153 15484 19165 15487
rect 18748 15456 19165 15484
rect 18748 15444 18754 15456
rect 19153 15453 19165 15456
rect 19199 15453 19211 15487
rect 19153 15447 19211 15453
rect 19242 15444 19248 15496
rect 19300 15484 19306 15496
rect 20162 15484 20168 15496
rect 19300 15456 20024 15484
rect 20123 15456 20168 15484
rect 19300 15444 19306 15456
rect 17405 15419 17463 15425
rect 17405 15385 17417 15419
rect 17451 15385 17463 15419
rect 17405 15379 17463 15385
rect 17770 15376 17776 15428
rect 17828 15416 17834 15428
rect 18598 15416 18604 15428
rect 17828 15388 18604 15416
rect 17828 15376 17834 15388
rect 18598 15376 18604 15388
rect 18656 15376 18662 15428
rect 19702 15416 19708 15428
rect 19663 15388 19708 15416
rect 19702 15376 19708 15388
rect 19760 15376 19766 15428
rect 19996 15416 20024 15456
rect 20162 15444 20168 15456
rect 20220 15444 20226 15496
rect 20257 15487 20315 15493
rect 20257 15453 20269 15487
rect 20303 15453 20315 15487
rect 20257 15447 20315 15453
rect 20272 15416 20300 15447
rect 19996 15388 20300 15416
rect 17678 15348 17684 15360
rect 12032 15320 16988 15348
rect 17639 15320 17684 15348
rect 12032 15308 12038 15320
rect 17678 15308 17684 15320
rect 17736 15308 17742 15360
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 4525 15147 4583 15153
rect 4525 15144 4537 15147
rect 1596 15116 4537 15144
rect 1596 14949 1624 15116
rect 4525 15113 4537 15116
rect 4571 15113 4583 15147
rect 4525 15107 4583 15113
rect 7650 15104 7656 15156
rect 7708 15144 7714 15156
rect 7837 15147 7895 15153
rect 7837 15144 7849 15147
rect 7708 15116 7849 15144
rect 7708 15104 7714 15116
rect 7837 15113 7849 15116
rect 7883 15113 7895 15147
rect 9766 15144 9772 15156
rect 7837 15107 7895 15113
rect 7944 15116 9772 15144
rect 3418 15036 3424 15088
rect 3476 15076 3482 15088
rect 7944 15076 7972 15116
rect 9766 15104 9772 15116
rect 9824 15104 9830 15156
rect 10042 15104 10048 15156
rect 10100 15144 10106 15156
rect 10137 15147 10195 15153
rect 10137 15144 10149 15147
rect 10100 15116 10149 15144
rect 10100 15104 10106 15116
rect 10137 15113 10149 15116
rect 10183 15113 10195 15147
rect 10137 15107 10195 15113
rect 10597 15147 10655 15153
rect 10597 15113 10609 15147
rect 10643 15144 10655 15147
rect 10686 15144 10692 15156
rect 10643 15116 10692 15144
rect 10643 15113 10655 15116
rect 10597 15107 10655 15113
rect 10686 15104 10692 15116
rect 10744 15104 10750 15156
rect 11698 15104 11704 15156
rect 11756 15144 11762 15156
rect 12158 15144 12164 15156
rect 11756 15116 12164 15144
rect 11756 15104 11762 15116
rect 12158 15104 12164 15116
rect 12216 15144 12222 15156
rect 13078 15144 13084 15156
rect 12216 15116 13084 15144
rect 12216 15104 12222 15116
rect 13078 15104 13084 15116
rect 13136 15104 13142 15156
rect 13538 15104 13544 15156
rect 13596 15144 13602 15156
rect 13633 15147 13691 15153
rect 13633 15144 13645 15147
rect 13596 15116 13645 15144
rect 13596 15104 13602 15116
rect 13633 15113 13645 15116
rect 13679 15113 13691 15147
rect 13633 15107 13691 15113
rect 14277 15147 14335 15153
rect 14277 15113 14289 15147
rect 14323 15144 14335 15147
rect 14458 15144 14464 15156
rect 14323 15116 14464 15144
rect 14323 15113 14335 15116
rect 14277 15107 14335 15113
rect 14458 15104 14464 15116
rect 14516 15104 14522 15156
rect 14550 15104 14556 15156
rect 14608 15144 14614 15156
rect 14645 15147 14703 15153
rect 14645 15144 14657 15147
rect 14608 15116 14657 15144
rect 14608 15104 14614 15116
rect 14645 15113 14657 15116
rect 14691 15113 14703 15147
rect 14645 15107 14703 15113
rect 16761 15147 16819 15153
rect 16761 15113 16773 15147
rect 16807 15144 16819 15147
rect 17954 15144 17960 15156
rect 16807 15116 17960 15144
rect 16807 15113 16819 15116
rect 16761 15107 16819 15113
rect 17954 15104 17960 15116
rect 18012 15104 18018 15156
rect 19242 15144 19248 15156
rect 18064 15116 19248 15144
rect 3476 15048 7972 15076
rect 3476 15036 3482 15048
rect 9950 15036 9956 15088
rect 10008 15076 10014 15088
rect 11514 15076 11520 15088
rect 10008 15048 11520 15076
rect 10008 15036 10014 15048
rect 11514 15036 11520 15048
rect 11572 15036 11578 15088
rect 11606 15036 11612 15088
rect 11664 15076 11670 15088
rect 12066 15076 12072 15088
rect 11664 15048 12072 15076
rect 11664 15036 11670 15048
rect 12066 15036 12072 15048
rect 12124 15036 12130 15088
rect 12710 15036 12716 15088
rect 12768 15076 12774 15088
rect 12986 15076 12992 15088
rect 12768 15048 12992 15076
rect 12768 15036 12774 15048
rect 12986 15036 12992 15048
rect 13044 15036 13050 15088
rect 16669 15079 16727 15085
rect 16669 15045 16681 15079
rect 16715 15076 16727 15079
rect 18064 15076 18092 15116
rect 19242 15104 19248 15116
rect 19300 15104 19306 15156
rect 19426 15144 19432 15156
rect 19387 15116 19432 15144
rect 19426 15104 19432 15116
rect 19484 15104 19490 15156
rect 19705 15147 19763 15153
rect 19705 15113 19717 15147
rect 19751 15144 19763 15147
rect 20162 15144 20168 15156
rect 19751 15116 20168 15144
rect 19751 15113 19763 15116
rect 19705 15107 19763 15113
rect 20162 15104 20168 15116
rect 20220 15104 20226 15156
rect 20622 15104 20628 15156
rect 20680 15144 20686 15156
rect 20901 15147 20959 15153
rect 20901 15144 20913 15147
rect 20680 15116 20913 15144
rect 20680 15104 20686 15116
rect 20901 15113 20913 15116
rect 20947 15113 20959 15147
rect 20901 15107 20959 15113
rect 16715 15048 18092 15076
rect 16715 15045 16727 15048
rect 16669 15039 16727 15045
rect 1854 15008 1860 15020
rect 1815 14980 1860 15008
rect 1854 14968 1860 14980
rect 1912 14968 1918 15020
rect 5169 15011 5227 15017
rect 5169 14977 5181 15011
rect 5215 15008 5227 15011
rect 5810 15008 5816 15020
rect 5215 14980 5816 15008
rect 5215 14977 5227 14980
rect 5169 14971 5227 14977
rect 5810 14968 5816 14980
rect 5868 14968 5874 15020
rect 7006 14968 7012 15020
rect 7064 15008 7070 15020
rect 7285 15011 7343 15017
rect 7285 15008 7297 15011
rect 7064 14980 7297 15008
rect 7064 14968 7070 14980
rect 7285 14977 7297 14980
rect 7331 14977 7343 15011
rect 7466 15008 7472 15020
rect 7427 14980 7472 15008
rect 7285 14971 7343 14977
rect 7466 14968 7472 14980
rect 7524 14968 7530 15020
rect 8757 15011 8815 15017
rect 8757 15008 8769 15011
rect 7944 14980 8769 15008
rect 1581 14943 1639 14949
rect 1581 14909 1593 14943
rect 1627 14909 1639 14943
rect 2314 14940 2320 14952
rect 2227 14912 2320 14940
rect 1581 14903 1639 14909
rect 2314 14900 2320 14912
rect 2372 14940 2378 14952
rect 3878 14940 3884 14952
rect 2372 14912 3884 14940
rect 2372 14900 2378 14912
rect 3878 14900 3884 14912
rect 3936 14900 3942 14952
rect 7374 14900 7380 14952
rect 7432 14940 7438 14952
rect 7944 14940 7972 14980
rect 8757 14977 8769 14980
rect 8803 14977 8815 15011
rect 11241 15011 11299 15017
rect 11241 15008 11253 15011
rect 8757 14971 8815 14977
rect 10244 14980 11253 15008
rect 7432 14912 7972 14940
rect 8021 14943 8079 14949
rect 7432 14900 7438 14912
rect 8021 14909 8033 14943
rect 8067 14940 8079 14943
rect 8202 14940 8208 14952
rect 8067 14912 8208 14940
rect 8067 14909 8079 14912
rect 8021 14903 8079 14909
rect 8202 14900 8208 14912
rect 8260 14900 8266 14952
rect 9024 14943 9082 14949
rect 9024 14909 9036 14943
rect 9070 14940 9082 14943
rect 9858 14940 9864 14952
rect 9070 14912 9864 14940
rect 9070 14909 9082 14912
rect 9024 14903 9082 14909
rect 9858 14900 9864 14912
rect 9916 14940 9922 14952
rect 10244 14940 10272 14980
rect 11241 14977 11253 14980
rect 11287 15008 11299 15011
rect 12158 15008 12164 15020
rect 11287 14980 12164 15008
rect 11287 14977 11299 14980
rect 11241 14971 11299 14977
rect 12158 14968 12164 14980
rect 12216 14968 12222 15020
rect 13265 15011 13323 15017
rect 13265 14977 13277 15011
rect 13311 15008 13323 15011
rect 13446 15008 13452 15020
rect 13311 14980 13452 15008
rect 13311 14977 13323 14980
rect 13265 14971 13323 14977
rect 13446 14968 13452 14980
rect 13504 14968 13510 15020
rect 15102 14968 15108 15020
rect 15160 15008 15166 15020
rect 15197 15011 15255 15017
rect 15197 15008 15209 15011
rect 15160 14980 15209 15008
rect 15160 14968 15166 14980
rect 15197 14977 15209 14980
rect 15243 14977 15255 15011
rect 17310 15008 17316 15020
rect 15197 14971 15255 14977
rect 15580 14980 17316 15008
rect 9916 14912 10272 14940
rect 9916 14900 9922 14912
rect 10318 14900 10324 14952
rect 10376 14940 10382 14952
rect 10594 14940 10600 14952
rect 10376 14912 10600 14940
rect 10376 14900 10382 14912
rect 10594 14900 10600 14912
rect 10652 14900 10658 14952
rect 10778 14900 10784 14952
rect 10836 14940 10842 14952
rect 11698 14940 11704 14952
rect 10836 14912 11704 14940
rect 10836 14900 10842 14912
rect 11698 14900 11704 14912
rect 11756 14940 11762 14952
rect 11793 14943 11851 14949
rect 11793 14940 11805 14943
rect 11756 14912 11805 14940
rect 11756 14900 11762 14912
rect 11793 14909 11805 14912
rect 11839 14909 11851 14943
rect 11793 14903 11851 14909
rect 11882 14900 11888 14952
rect 11940 14940 11946 14952
rect 12894 14940 12900 14952
rect 11940 14912 12900 14940
rect 11940 14900 11946 14912
rect 12894 14900 12900 14912
rect 12952 14900 12958 14952
rect 13814 14940 13820 14952
rect 13775 14912 13820 14940
rect 13814 14900 13820 14912
rect 13872 14900 13878 14952
rect 14093 14943 14151 14949
rect 14093 14909 14105 14943
rect 14139 14940 14151 14943
rect 15580 14940 15608 14980
rect 17310 14968 17316 14980
rect 17368 14968 17374 15020
rect 17405 15011 17463 15017
rect 17405 14977 17417 15011
rect 17451 15008 17463 15011
rect 19444 15008 19472 15104
rect 20257 15011 20315 15017
rect 20257 15008 20269 15011
rect 17451 14980 18184 15008
rect 19444 14980 20269 15008
rect 17451 14977 17463 14980
rect 17405 14971 17463 14977
rect 14139 14912 15608 14940
rect 14139 14909 14151 14912
rect 14093 14903 14151 14909
rect 15654 14900 15660 14952
rect 15712 14940 15718 14952
rect 16209 14943 16267 14949
rect 15712 14912 15757 14940
rect 15712 14900 15718 14912
rect 16209 14909 16221 14943
rect 16255 14940 16267 14943
rect 16669 14943 16727 14949
rect 16669 14940 16681 14943
rect 16255 14912 16681 14940
rect 16255 14909 16267 14912
rect 16209 14903 16267 14909
rect 16669 14909 16681 14912
rect 16715 14909 16727 14943
rect 16669 14903 16727 14909
rect 17221 14943 17279 14949
rect 17221 14909 17233 14943
rect 17267 14940 17279 14943
rect 17678 14940 17684 14952
rect 17267 14912 17684 14940
rect 17267 14909 17279 14912
rect 17221 14903 17279 14909
rect 17678 14900 17684 14912
rect 17736 14900 17742 14952
rect 17770 14900 17776 14952
rect 17828 14940 17834 14952
rect 18049 14943 18107 14949
rect 18049 14940 18061 14943
rect 17828 14912 18061 14940
rect 17828 14900 17834 14912
rect 18049 14909 18061 14912
rect 18095 14909 18107 14943
rect 18156 14940 18184 14980
rect 20257 14977 20269 14980
rect 20303 14977 20315 15011
rect 20257 14971 20315 14977
rect 18322 14949 18328 14952
rect 18305 14943 18328 14949
rect 18305 14940 18317 14943
rect 18156 14912 18317 14940
rect 18049 14903 18107 14909
rect 18305 14909 18317 14912
rect 18380 14940 18386 14952
rect 18380 14912 18453 14940
rect 18305 14903 18328 14909
rect 18322 14900 18328 14903
rect 18380 14900 18386 14912
rect 18598 14900 18604 14952
rect 18656 14940 18662 14952
rect 20165 14943 20223 14949
rect 20165 14940 20177 14943
rect 18656 14912 20177 14940
rect 18656 14900 18662 14912
rect 20165 14909 20177 14912
rect 20211 14909 20223 14943
rect 20165 14903 20223 14909
rect 20717 14943 20775 14949
rect 20717 14909 20729 14943
rect 20763 14909 20775 14943
rect 20717 14903 20775 14909
rect 2584 14875 2642 14881
rect 2584 14841 2596 14875
rect 2630 14872 2642 14875
rect 3234 14872 3240 14884
rect 2630 14844 3240 14872
rect 2630 14841 2642 14844
rect 2584 14835 2642 14841
rect 3234 14832 3240 14844
rect 3292 14832 3298 14884
rect 4893 14875 4951 14881
rect 4893 14841 4905 14875
rect 4939 14872 4951 14875
rect 5442 14872 5448 14884
rect 4939 14844 5448 14872
rect 4939 14841 4951 14844
rect 4893 14835 4951 14841
rect 5442 14832 5448 14844
rect 5500 14832 5506 14884
rect 7193 14875 7251 14881
rect 7193 14841 7205 14875
rect 7239 14872 7251 14875
rect 9950 14872 9956 14884
rect 7239 14844 9956 14872
rect 7239 14841 7251 14844
rect 7193 14835 7251 14841
rect 9950 14832 9956 14844
rect 10008 14832 10014 14884
rect 10870 14872 10876 14884
rect 10336 14844 10876 14872
rect 10336 14816 10364 14844
rect 10870 14832 10876 14844
rect 10928 14872 10934 14884
rect 11057 14875 11115 14881
rect 11057 14872 11069 14875
rect 10928 14844 11069 14872
rect 10928 14832 10934 14844
rect 11057 14841 11069 14844
rect 11103 14841 11115 14875
rect 11057 14835 11115 14841
rect 11238 14832 11244 14884
rect 11296 14872 11302 14884
rect 13081 14875 13139 14881
rect 13081 14872 13093 14875
rect 11296 14844 13093 14872
rect 11296 14832 11302 14844
rect 13081 14841 13093 14844
rect 13127 14841 13139 14875
rect 13081 14835 13139 14841
rect 15013 14875 15071 14881
rect 15013 14841 15025 14875
rect 15059 14872 15071 14875
rect 15930 14872 15936 14884
rect 15059 14844 15936 14872
rect 15059 14841 15071 14844
rect 15013 14835 15071 14841
rect 15930 14832 15936 14844
rect 15988 14832 15994 14884
rect 16850 14872 16856 14884
rect 16316 14844 16856 14872
rect 3142 14764 3148 14816
rect 3200 14804 3206 14816
rect 3697 14807 3755 14813
rect 3697 14804 3709 14807
rect 3200 14776 3709 14804
rect 3200 14764 3206 14776
rect 3697 14773 3709 14776
rect 3743 14773 3755 14807
rect 3697 14767 3755 14773
rect 4985 14807 5043 14813
rect 4985 14773 4997 14807
rect 5031 14804 5043 14807
rect 5350 14804 5356 14816
rect 5031 14776 5356 14804
rect 5031 14773 5043 14776
rect 4985 14767 5043 14773
rect 5350 14764 5356 14776
rect 5408 14764 5414 14816
rect 6822 14804 6828 14816
rect 6783 14776 6828 14804
rect 6822 14764 6828 14776
rect 6880 14764 6886 14816
rect 10318 14764 10324 14816
rect 10376 14764 10382 14816
rect 10778 14764 10784 14816
rect 10836 14804 10842 14816
rect 10965 14807 11023 14813
rect 10965 14804 10977 14807
rect 10836 14776 10977 14804
rect 10836 14764 10842 14776
rect 10965 14773 10977 14776
rect 11011 14773 11023 14807
rect 11974 14804 11980 14816
rect 11935 14776 11980 14804
rect 10965 14767 11023 14773
rect 11974 14764 11980 14776
rect 12032 14764 12038 14816
rect 12618 14804 12624 14816
rect 12579 14776 12624 14804
rect 12618 14764 12624 14776
rect 12676 14764 12682 14816
rect 12986 14804 12992 14816
rect 12947 14776 12992 14804
rect 12986 14764 12992 14776
rect 13044 14764 13050 14816
rect 15105 14807 15163 14813
rect 15105 14773 15117 14807
rect 15151 14804 15163 14807
rect 15470 14804 15476 14816
rect 15151 14776 15476 14804
rect 15151 14773 15163 14776
rect 15105 14767 15163 14773
rect 15470 14764 15476 14776
rect 15528 14764 15534 14816
rect 15841 14807 15899 14813
rect 15841 14773 15853 14807
rect 15887 14804 15899 14807
rect 16316 14804 16344 14844
rect 16850 14832 16856 14844
rect 16908 14832 16914 14884
rect 17494 14832 17500 14884
rect 17552 14872 17558 14884
rect 20732 14872 20760 14903
rect 17552 14844 20760 14872
rect 17552 14832 17558 14844
rect 15887 14776 16344 14804
rect 16393 14807 16451 14813
rect 15887 14773 15899 14776
rect 15841 14767 15899 14773
rect 16393 14773 16405 14807
rect 16439 14804 16451 14807
rect 16942 14804 16948 14816
rect 16439 14776 16948 14804
rect 16439 14773 16451 14776
rect 16393 14767 16451 14773
rect 16942 14764 16948 14776
rect 17000 14764 17006 14816
rect 17129 14807 17187 14813
rect 17129 14773 17141 14807
rect 17175 14804 17187 14807
rect 18598 14804 18604 14816
rect 17175 14776 18604 14804
rect 17175 14773 17187 14776
rect 17129 14767 17187 14773
rect 18598 14764 18604 14776
rect 18656 14764 18662 14816
rect 19334 14764 19340 14816
rect 19392 14804 19398 14816
rect 20073 14807 20131 14813
rect 20073 14804 20085 14807
rect 19392 14776 20085 14804
rect 19392 14764 19398 14776
rect 20073 14773 20085 14776
rect 20119 14773 20131 14807
rect 20073 14767 20131 14773
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 1946 14600 1952 14612
rect 1907 14572 1952 14600
rect 1946 14560 1952 14572
rect 2004 14560 2010 14612
rect 2685 14603 2743 14609
rect 2685 14569 2697 14603
rect 2731 14600 2743 14603
rect 4154 14600 4160 14612
rect 2731 14572 4160 14600
rect 2731 14569 2743 14572
rect 2685 14563 2743 14569
rect 4154 14560 4160 14572
rect 4212 14560 4218 14612
rect 4982 14560 4988 14612
rect 5040 14600 5046 14612
rect 5258 14600 5264 14612
rect 5040 14572 5264 14600
rect 5040 14560 5046 14572
rect 5258 14560 5264 14572
rect 5316 14560 5322 14612
rect 5810 14600 5816 14612
rect 5771 14572 5816 14600
rect 5810 14560 5816 14572
rect 5868 14560 5874 14612
rect 6914 14560 6920 14612
rect 6972 14600 6978 14612
rect 8113 14603 8171 14609
rect 8113 14600 8125 14603
rect 6972 14572 8125 14600
rect 6972 14560 6978 14572
rect 8113 14569 8125 14572
rect 8159 14569 8171 14603
rect 8113 14563 8171 14569
rect 9582 14560 9588 14612
rect 9640 14600 9646 14612
rect 10045 14603 10103 14609
rect 10045 14600 10057 14603
rect 9640 14572 10057 14600
rect 9640 14560 9646 14572
rect 10045 14569 10057 14572
rect 10091 14569 10103 14603
rect 10778 14600 10784 14612
rect 10739 14572 10784 14600
rect 10045 14563 10103 14569
rect 10778 14560 10784 14572
rect 10836 14560 10842 14612
rect 11238 14600 11244 14612
rect 11199 14572 11244 14600
rect 11238 14560 11244 14572
rect 11296 14560 11302 14612
rect 11514 14560 11520 14612
rect 11572 14600 11578 14612
rect 11609 14603 11667 14609
rect 11609 14600 11621 14603
rect 11572 14572 11621 14600
rect 11572 14560 11578 14572
rect 11609 14569 11621 14572
rect 11655 14569 11667 14603
rect 11609 14563 11667 14569
rect 12161 14603 12219 14609
rect 12161 14569 12173 14603
rect 12207 14600 12219 14603
rect 12434 14600 12440 14612
rect 12207 14572 12440 14600
rect 12207 14569 12219 14572
rect 12161 14563 12219 14569
rect 12434 14560 12440 14572
rect 12492 14560 12498 14612
rect 12526 14560 12532 14612
rect 12584 14560 12590 14612
rect 12618 14560 12624 14612
rect 12676 14600 12682 14612
rect 14645 14603 14703 14609
rect 14645 14600 14657 14603
rect 12676 14572 14657 14600
rect 12676 14560 12682 14572
rect 14645 14569 14657 14572
rect 14691 14569 14703 14603
rect 15289 14603 15347 14609
rect 15289 14600 15301 14603
rect 14645 14563 14703 14569
rect 14752 14572 15301 14600
rect 3142 14492 3148 14544
rect 3200 14492 3206 14544
rect 5534 14532 5540 14544
rect 4448 14504 5540 14532
rect 1670 14424 1676 14476
rect 1728 14464 1734 14476
rect 1765 14467 1823 14473
rect 1765 14464 1777 14467
rect 1728 14436 1777 14464
rect 1728 14424 1734 14436
rect 1765 14433 1777 14436
rect 1811 14433 1823 14467
rect 3050 14464 3056 14476
rect 3011 14436 3056 14464
rect 1765 14427 1823 14433
rect 3050 14424 3056 14436
rect 3108 14424 3114 14476
rect 3160 14464 3188 14492
rect 3160 14436 3280 14464
rect 2222 14356 2228 14408
rect 2280 14396 2286 14408
rect 3252 14405 3280 14436
rect 3878 14424 3884 14476
rect 3936 14464 3942 14476
rect 4448 14473 4476 14504
rect 5534 14492 5540 14504
rect 5592 14492 5598 14544
rect 5828 14532 5856 14560
rect 6334 14535 6392 14541
rect 6334 14532 6346 14535
rect 5828 14504 6346 14532
rect 6334 14501 6346 14504
rect 6380 14501 6392 14535
rect 6334 14495 6392 14501
rect 7006 14492 7012 14544
rect 7064 14532 7070 14544
rect 8205 14535 8263 14541
rect 7064 14504 8156 14532
rect 7064 14492 7070 14504
rect 4433 14467 4491 14473
rect 4433 14464 4445 14467
rect 3936 14436 4445 14464
rect 3936 14424 3942 14436
rect 4433 14433 4445 14436
rect 4479 14433 4491 14467
rect 4433 14427 4491 14433
rect 4700 14467 4758 14473
rect 4700 14433 4712 14467
rect 4746 14464 4758 14467
rect 5074 14464 5080 14476
rect 4746 14436 5080 14464
rect 4746 14433 4758 14436
rect 4700 14427 4758 14433
rect 5074 14424 5080 14436
rect 5132 14424 5138 14476
rect 5258 14424 5264 14476
rect 5316 14464 5322 14476
rect 8128 14464 8156 14504
rect 8205 14501 8217 14535
rect 8251 14532 8263 14535
rect 11882 14532 11888 14544
rect 8251 14504 11888 14532
rect 8251 14501 8263 14504
rect 8205 14495 8263 14501
rect 11882 14492 11888 14504
rect 11940 14492 11946 14544
rect 12066 14492 12072 14544
rect 12124 14532 12130 14544
rect 12544 14532 12572 14560
rect 14752 14532 14780 14572
rect 15289 14569 15301 14572
rect 15335 14569 15347 14603
rect 15289 14563 15347 14569
rect 16301 14603 16359 14609
rect 16301 14569 16313 14603
rect 16347 14600 16359 14603
rect 17402 14600 17408 14612
rect 16347 14572 17408 14600
rect 16347 14569 16359 14572
rect 16301 14563 16359 14569
rect 17402 14560 17408 14572
rect 17460 14560 17466 14612
rect 18322 14600 18328 14612
rect 18283 14572 18328 14600
rect 18322 14560 18328 14572
rect 18380 14560 18386 14612
rect 18598 14600 18604 14612
rect 18559 14572 18604 14600
rect 18598 14560 18604 14572
rect 18656 14560 18662 14612
rect 19150 14600 19156 14612
rect 18708 14572 19156 14600
rect 12124 14504 12572 14532
rect 13648 14504 14780 14532
rect 12124 14492 12130 14504
rect 5316 14436 7512 14464
rect 8128 14436 8708 14464
rect 5316 14424 5322 14436
rect 7484 14408 7512 14436
rect 3145 14399 3203 14405
rect 3145 14396 3157 14399
rect 2280 14368 3157 14396
rect 2280 14356 2286 14368
rect 3145 14365 3157 14368
rect 3191 14365 3203 14399
rect 3145 14359 3203 14365
rect 3237 14399 3295 14405
rect 3237 14365 3249 14399
rect 3283 14365 3295 14399
rect 3237 14359 3295 14365
rect 3160 14328 3188 14359
rect 5534 14356 5540 14408
rect 5592 14396 5598 14408
rect 6089 14399 6147 14405
rect 6089 14396 6101 14399
rect 5592 14368 6101 14396
rect 5592 14356 5598 14368
rect 6089 14365 6101 14368
rect 6135 14365 6147 14399
rect 6089 14359 6147 14365
rect 7466 14356 7472 14408
rect 7524 14396 7530 14408
rect 8297 14399 8355 14405
rect 8297 14396 8309 14399
rect 7524 14368 8309 14396
rect 7524 14356 7530 14368
rect 8297 14365 8309 14368
rect 8343 14365 8355 14399
rect 8680 14396 8708 14436
rect 9030 14424 9036 14476
rect 9088 14464 9094 14476
rect 10137 14467 10195 14473
rect 10137 14464 10149 14467
rect 9088 14436 10149 14464
rect 9088 14424 9094 14436
rect 10137 14433 10149 14436
rect 10183 14433 10195 14467
rect 12520 14467 12578 14473
rect 12520 14464 12532 14467
rect 10137 14427 10195 14433
rect 11900 14436 12532 14464
rect 10042 14396 10048 14408
rect 8680 14368 10048 14396
rect 8297 14359 8355 14365
rect 10042 14356 10048 14368
rect 10100 14356 10106 14408
rect 10321 14399 10379 14405
rect 10321 14365 10333 14399
rect 10367 14396 10379 14399
rect 10410 14396 10416 14408
rect 10367 14368 10416 14396
rect 10367 14365 10379 14368
rect 10321 14359 10379 14365
rect 10410 14356 10416 14368
rect 10468 14356 10474 14408
rect 10778 14356 10784 14408
rect 10836 14396 10842 14408
rect 11900 14405 11928 14436
rect 12520 14433 12532 14436
rect 12566 14464 12578 14467
rect 13538 14464 13544 14476
rect 12566 14436 13544 14464
rect 12566 14433 12578 14436
rect 12520 14427 12578 14433
rect 13538 14424 13544 14436
rect 13596 14424 13602 14476
rect 11701 14399 11759 14405
rect 11701 14396 11713 14399
rect 10836 14368 11713 14396
rect 10836 14356 10842 14368
rect 11701 14365 11713 14368
rect 11747 14365 11759 14399
rect 11701 14359 11759 14365
rect 11885 14399 11943 14405
rect 11885 14365 11897 14399
rect 11931 14365 11943 14399
rect 11885 14359 11943 14365
rect 12161 14399 12219 14405
rect 12161 14365 12173 14399
rect 12207 14396 12219 14399
rect 12253 14399 12311 14405
rect 12253 14396 12265 14399
rect 12207 14368 12265 14396
rect 12207 14365 12219 14368
rect 12161 14359 12219 14365
rect 12253 14365 12265 14368
rect 12299 14365 12311 14399
rect 12253 14359 12311 14365
rect 3418 14328 3424 14340
rect 3160 14300 3424 14328
rect 3418 14288 3424 14300
rect 3476 14288 3482 14340
rect 7098 14288 7104 14340
rect 7156 14328 7162 14340
rect 13648 14328 13676 14504
rect 14826 14492 14832 14544
rect 14884 14532 14890 14544
rect 17034 14532 17040 14544
rect 14884 14504 17040 14532
rect 14884 14492 14890 14504
rect 17034 14492 17040 14504
rect 17092 14492 17098 14544
rect 17212 14535 17270 14541
rect 17212 14501 17224 14535
rect 17258 14532 17270 14535
rect 17862 14532 17868 14544
rect 17258 14504 17868 14532
rect 17258 14501 17270 14504
rect 17212 14495 17270 14501
rect 17862 14492 17868 14504
rect 17920 14492 17926 14544
rect 17954 14492 17960 14544
rect 18012 14532 18018 14544
rect 18708 14532 18736 14572
rect 19150 14560 19156 14572
rect 19208 14560 19214 14612
rect 18012 14504 18736 14532
rect 18969 14535 19027 14541
rect 18012 14492 18018 14504
rect 18969 14501 18981 14535
rect 19015 14532 19027 14535
rect 20901 14535 20959 14541
rect 20901 14532 20913 14535
rect 19015 14504 20913 14532
rect 19015 14501 19027 14504
rect 18969 14495 19027 14501
rect 20901 14501 20913 14504
rect 20947 14501 20959 14535
rect 20901 14495 20959 14501
rect 14090 14464 14096 14476
rect 14051 14436 14096 14464
rect 14090 14424 14096 14436
rect 14148 14424 14154 14476
rect 14553 14467 14611 14473
rect 14553 14433 14565 14467
rect 14599 14464 14611 14467
rect 15010 14464 15016 14476
rect 14599 14436 15016 14464
rect 14599 14433 14611 14436
rect 14553 14427 14611 14433
rect 15010 14424 15016 14436
rect 15068 14424 15074 14476
rect 15289 14467 15347 14473
rect 15289 14433 15301 14467
rect 15335 14464 15347 14467
rect 15381 14467 15439 14473
rect 15381 14464 15393 14467
rect 15335 14436 15393 14464
rect 15335 14433 15347 14436
rect 15289 14427 15347 14433
rect 15381 14433 15393 14436
rect 15427 14464 15439 14467
rect 16206 14464 16212 14476
rect 15427 14436 16212 14464
rect 15427 14433 15439 14436
rect 15381 14427 15439 14433
rect 16206 14424 16212 14436
rect 16264 14424 16270 14476
rect 16393 14467 16451 14473
rect 16393 14433 16405 14467
rect 16439 14464 16451 14467
rect 17770 14464 17776 14476
rect 16439 14436 17776 14464
rect 16439 14433 16451 14436
rect 16393 14427 16451 14433
rect 17770 14424 17776 14436
rect 17828 14424 17834 14476
rect 17880 14464 17908 14492
rect 17880 14436 19196 14464
rect 14366 14356 14372 14408
rect 14424 14396 14430 14408
rect 14737 14399 14795 14405
rect 14737 14396 14749 14399
rect 14424 14368 14749 14396
rect 14424 14356 14430 14368
rect 14737 14365 14749 14368
rect 14783 14365 14795 14399
rect 16298 14396 16304 14408
rect 14737 14359 14795 14365
rect 15488 14368 16304 14396
rect 7156 14300 11100 14328
rect 7156 14288 7162 14300
rect 2038 14220 2044 14272
rect 2096 14260 2102 14272
rect 7006 14260 7012 14272
rect 2096 14232 7012 14260
rect 2096 14220 2102 14232
rect 7006 14220 7012 14232
rect 7064 14220 7070 14272
rect 7466 14260 7472 14272
rect 7427 14232 7472 14260
rect 7466 14220 7472 14232
rect 7524 14220 7530 14272
rect 7742 14260 7748 14272
rect 7703 14232 7748 14260
rect 7742 14220 7748 14232
rect 7800 14220 7806 14272
rect 8294 14220 8300 14272
rect 8352 14260 8358 14272
rect 9030 14260 9036 14272
rect 8352 14232 9036 14260
rect 8352 14220 8358 14232
rect 9030 14220 9036 14232
rect 9088 14220 9094 14272
rect 9677 14263 9735 14269
rect 9677 14229 9689 14263
rect 9723 14260 9735 14263
rect 10962 14260 10968 14272
rect 9723 14232 10968 14260
rect 9723 14229 9735 14232
rect 9677 14223 9735 14229
rect 10962 14220 10968 14232
rect 11020 14220 11026 14272
rect 11072 14260 11100 14300
rect 13372 14300 13676 14328
rect 13372 14260 13400 14300
rect 13814 14288 13820 14340
rect 13872 14328 13878 14340
rect 13909 14331 13967 14337
rect 13909 14328 13921 14331
rect 13872 14300 13921 14328
rect 13872 14288 13878 14300
rect 13909 14297 13921 14300
rect 13955 14328 13967 14331
rect 15378 14328 15384 14340
rect 13955 14300 15384 14328
rect 13955 14297 13967 14300
rect 13909 14291 13967 14297
rect 15378 14288 15384 14300
rect 15436 14288 15442 14340
rect 11072 14232 13400 14260
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 13633 14263 13691 14269
rect 13633 14260 13645 14263
rect 13504 14232 13645 14260
rect 13504 14220 13510 14232
rect 13633 14229 13645 14232
rect 13679 14229 13691 14263
rect 13633 14223 13691 14229
rect 14185 14263 14243 14269
rect 14185 14229 14197 14263
rect 14231 14260 14243 14263
rect 15488 14260 15516 14368
rect 16298 14356 16304 14368
rect 16356 14356 16362 14408
rect 16485 14399 16543 14405
rect 16485 14365 16497 14399
rect 16531 14396 16543 14399
rect 16574 14396 16580 14408
rect 16531 14368 16580 14396
rect 16531 14365 16543 14368
rect 16485 14359 16543 14365
rect 16574 14356 16580 14368
rect 16632 14356 16638 14408
rect 16850 14356 16856 14408
rect 16908 14396 16914 14408
rect 16945 14399 17003 14405
rect 16945 14396 16957 14399
rect 16908 14368 16957 14396
rect 16908 14356 16914 14368
rect 16945 14365 16957 14368
rect 16991 14365 17003 14399
rect 16945 14359 17003 14365
rect 18414 14356 18420 14408
rect 18472 14396 18478 14408
rect 18966 14396 18972 14408
rect 18472 14368 18972 14396
rect 18472 14356 18478 14368
rect 18966 14356 18972 14368
rect 19024 14396 19030 14408
rect 19168 14405 19196 14436
rect 19242 14424 19248 14476
rect 19300 14464 19306 14476
rect 19981 14467 20039 14473
rect 19981 14464 19993 14467
rect 19300 14436 19993 14464
rect 19300 14424 19306 14436
rect 19981 14433 19993 14436
rect 20027 14433 20039 14467
rect 19981 14427 20039 14433
rect 19061 14399 19119 14405
rect 19061 14396 19073 14399
rect 19024 14368 19073 14396
rect 19024 14356 19030 14368
rect 19061 14365 19073 14368
rect 19107 14365 19119 14399
rect 19061 14359 19119 14365
rect 19153 14399 19211 14405
rect 19153 14365 19165 14399
rect 19199 14365 19211 14399
rect 19153 14359 19211 14365
rect 19794 14356 19800 14408
rect 19852 14396 19858 14408
rect 20073 14399 20131 14405
rect 20073 14396 20085 14399
rect 19852 14368 20085 14396
rect 19852 14356 19858 14368
rect 20073 14365 20085 14368
rect 20119 14365 20131 14399
rect 20073 14359 20131 14365
rect 20162 14356 20168 14408
rect 20220 14396 20226 14408
rect 20220 14368 20265 14396
rect 20220 14356 20226 14368
rect 15565 14331 15623 14337
rect 15565 14297 15577 14331
rect 15611 14328 15623 14331
rect 16758 14328 16764 14340
rect 15611 14300 16764 14328
rect 15611 14297 15623 14300
rect 15565 14291 15623 14297
rect 16758 14288 16764 14300
rect 16816 14288 16822 14340
rect 14231 14232 15516 14260
rect 15933 14263 15991 14269
rect 14231 14229 14243 14232
rect 14185 14223 14243 14229
rect 15933 14229 15945 14263
rect 15979 14260 15991 14263
rect 17310 14260 17316 14272
rect 15979 14232 17316 14260
rect 15979 14229 15991 14232
rect 15933 14223 15991 14229
rect 17310 14220 17316 14232
rect 17368 14220 17374 14272
rect 17586 14220 17592 14272
rect 17644 14260 17650 14272
rect 19613 14263 19671 14269
rect 19613 14260 19625 14263
rect 17644 14232 19625 14260
rect 17644 14220 17650 14232
rect 19613 14229 19625 14232
rect 19659 14229 19671 14263
rect 19613 14223 19671 14229
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 3878 14056 3884 14068
rect 3712 14028 3884 14056
rect 1670 13920 1676 13932
rect 1631 13892 1676 13920
rect 1670 13880 1676 13892
rect 1728 13880 1734 13932
rect 3712 13929 3740 14028
rect 3878 14016 3884 14028
rect 3936 14016 3942 14068
rect 5074 14056 5080 14068
rect 5035 14028 5080 14056
rect 5074 14016 5080 14028
rect 5132 14016 5138 14068
rect 5350 14056 5356 14068
rect 5311 14028 5356 14056
rect 5350 14016 5356 14028
rect 5408 14016 5414 14068
rect 7006 14016 7012 14068
rect 7064 14056 7070 14068
rect 8754 14056 8760 14068
rect 7064 14028 8340 14056
rect 8667 14028 8760 14056
rect 7064 14016 7070 14028
rect 3697 13923 3755 13929
rect 3697 13889 3709 13923
rect 3743 13889 3755 13923
rect 5092 13920 5120 14016
rect 8312 13988 8340 14028
rect 8754 14016 8760 14028
rect 8812 14056 8818 14068
rect 8812 14028 11100 14056
rect 8812 14016 8818 14028
rect 8849 13991 8907 13997
rect 8849 13988 8861 13991
rect 8312 13960 8861 13988
rect 8849 13957 8861 13960
rect 8895 13957 8907 13991
rect 10505 13991 10563 13997
rect 10505 13988 10517 13991
rect 8849 13951 8907 13957
rect 9324 13960 10517 13988
rect 5905 13923 5963 13929
rect 5905 13920 5917 13923
rect 5092 13892 5917 13920
rect 3697 13883 3755 13889
rect 5905 13889 5917 13892
rect 5951 13920 5963 13923
rect 5994 13920 6000 13932
rect 5951 13892 6000 13920
rect 5951 13889 5963 13892
rect 5905 13883 5963 13889
rect 5994 13880 6000 13892
rect 6052 13880 6058 13932
rect 9324 13929 9352 13960
rect 10505 13957 10517 13960
rect 10551 13957 10563 13991
rect 10505 13951 10563 13957
rect 9309 13923 9367 13929
rect 9309 13889 9321 13923
rect 9355 13889 9367 13923
rect 9309 13883 9367 13889
rect 9398 13880 9404 13932
rect 9456 13920 9462 13932
rect 10321 13923 10379 13929
rect 10321 13920 10333 13923
rect 9456 13892 9501 13920
rect 9600 13892 10333 13920
rect 9456 13880 9462 13892
rect 1394 13852 1400 13864
rect 1355 13824 1400 13852
rect 1394 13812 1400 13824
rect 1452 13812 1458 13864
rect 2133 13855 2191 13861
rect 2133 13821 2145 13855
rect 2179 13852 2191 13855
rect 3602 13852 3608 13864
rect 2179 13824 3608 13852
rect 2179 13821 2191 13824
rect 2133 13815 2191 13821
rect 3602 13812 3608 13824
rect 3660 13812 3666 13864
rect 3964 13855 4022 13861
rect 3964 13821 3976 13855
rect 4010 13852 4022 13855
rect 5258 13852 5264 13864
rect 4010 13824 5264 13852
rect 4010 13821 4022 13824
rect 3964 13815 4022 13821
rect 5258 13812 5264 13824
rect 5316 13812 5322 13864
rect 5813 13855 5871 13861
rect 5813 13821 5825 13855
rect 5859 13852 5871 13855
rect 6822 13852 6828 13864
rect 5859 13824 6828 13852
rect 5859 13821 5871 13824
rect 5813 13815 5871 13821
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 7374 13852 7380 13864
rect 7335 13824 7380 13852
rect 7374 13812 7380 13824
rect 7432 13812 7438 13864
rect 1578 13744 1584 13796
rect 1636 13784 1642 13796
rect 2409 13787 2467 13793
rect 2409 13784 2421 13787
rect 1636 13756 2421 13784
rect 1636 13744 1642 13756
rect 2409 13753 2421 13756
rect 2455 13753 2467 13787
rect 2409 13747 2467 13753
rect 7466 13744 7472 13796
rect 7524 13784 7530 13796
rect 7644 13787 7702 13793
rect 7644 13784 7656 13787
rect 7524 13756 7656 13784
rect 7524 13744 7530 13756
rect 7644 13753 7656 13756
rect 7690 13784 7702 13787
rect 8938 13784 8944 13796
rect 7690 13756 8944 13784
rect 7690 13753 7702 13756
rect 7644 13747 7702 13753
rect 8938 13744 8944 13756
rect 8996 13784 9002 13796
rect 9600 13784 9628 13892
rect 10321 13889 10333 13892
rect 10367 13920 10379 13923
rect 10410 13920 10416 13932
rect 10367 13892 10416 13920
rect 10367 13889 10379 13892
rect 10321 13883 10379 13889
rect 10410 13880 10416 13892
rect 10468 13880 10474 13932
rect 10962 13920 10968 13932
rect 10923 13892 10968 13920
rect 10962 13880 10968 13892
rect 11020 13880 11026 13932
rect 11072 13929 11100 14028
rect 11146 14016 11152 14068
rect 11204 14056 11210 14068
rect 11333 14059 11391 14065
rect 11333 14056 11345 14059
rect 11204 14028 11345 14056
rect 11204 14016 11210 14028
rect 11333 14025 11345 14028
rect 11379 14025 11391 14059
rect 11333 14019 11391 14025
rect 11974 14016 11980 14068
rect 12032 14056 12038 14068
rect 14826 14056 14832 14068
rect 12032 14028 14832 14056
rect 12032 14016 12038 14028
rect 14826 14016 14832 14028
rect 14884 14016 14890 14068
rect 15010 14056 15016 14068
rect 14971 14028 15016 14056
rect 15010 14016 15016 14028
rect 15068 14016 15074 14068
rect 16574 14016 16580 14068
rect 16632 14056 16638 14068
rect 17034 14056 17040 14068
rect 16632 14028 17040 14056
rect 16632 14016 16638 14028
rect 17034 14016 17040 14028
rect 17092 14056 17098 14068
rect 20162 14056 20168 14068
rect 17092 14028 20168 14056
rect 17092 14016 17098 14028
rect 20162 14016 20168 14028
rect 20220 14016 20226 14068
rect 11514 13948 11520 14000
rect 11572 13988 11578 14000
rect 12434 13988 12440 14000
rect 11572 13960 12440 13988
rect 11572 13948 11578 13960
rect 12434 13948 12440 13960
rect 12492 13988 12498 14000
rect 12492 13960 13400 13988
rect 12492 13948 12498 13960
rect 11057 13923 11115 13929
rect 11057 13889 11069 13923
rect 11103 13889 11115 13923
rect 11057 13883 11115 13889
rect 11146 13880 11152 13932
rect 11204 13920 11210 13932
rect 11793 13923 11851 13929
rect 11793 13920 11805 13923
rect 11204 13892 11805 13920
rect 11204 13880 11210 13892
rect 11793 13889 11805 13892
rect 11839 13889 11851 13923
rect 11793 13883 11851 13889
rect 11977 13923 12035 13929
rect 11977 13889 11989 13923
rect 12023 13920 12035 13923
rect 12158 13920 12164 13932
rect 12023 13892 12164 13920
rect 12023 13889 12035 13892
rect 11977 13883 12035 13889
rect 12158 13880 12164 13892
rect 12216 13880 12222 13932
rect 13372 13929 13400 13960
rect 15102 13948 15108 14000
rect 15160 13988 15166 14000
rect 18506 13988 18512 14000
rect 15160 13960 18512 13988
rect 15160 13948 15166 13960
rect 18506 13948 18512 13960
rect 18564 13948 18570 14000
rect 13357 13923 13415 13929
rect 13357 13889 13369 13923
rect 13403 13889 13415 13923
rect 13357 13883 13415 13889
rect 15565 13923 15623 13929
rect 15565 13889 15577 13923
rect 15611 13889 15623 13923
rect 15565 13883 15623 13889
rect 10137 13855 10195 13861
rect 10137 13821 10149 13855
rect 10183 13852 10195 13855
rect 12066 13852 12072 13864
rect 10183 13824 12072 13852
rect 10183 13821 10195 13824
rect 10137 13815 10195 13821
rect 12066 13812 12072 13824
rect 12124 13812 12130 13864
rect 13446 13812 13452 13864
rect 13504 13852 13510 13864
rect 13624 13855 13682 13861
rect 13624 13852 13636 13855
rect 13504 13824 13636 13852
rect 13504 13812 13510 13824
rect 13624 13821 13636 13824
rect 13670 13852 13682 13855
rect 15580 13852 15608 13883
rect 16390 13880 16396 13932
rect 16448 13920 16454 13932
rect 16577 13923 16635 13929
rect 16577 13920 16589 13923
rect 16448 13892 16589 13920
rect 16448 13880 16454 13892
rect 16577 13889 16589 13892
rect 16623 13889 16635 13923
rect 17494 13920 17500 13932
rect 17455 13892 17500 13920
rect 16577 13883 16635 13889
rect 17494 13880 17500 13892
rect 17552 13880 17558 13932
rect 18064 13892 18736 13920
rect 16482 13852 16488 13864
rect 13670 13824 15608 13852
rect 16443 13824 16488 13852
rect 13670 13821 13682 13824
rect 13624 13815 13682 13821
rect 16482 13812 16488 13824
rect 16540 13812 16546 13864
rect 16666 13812 16672 13864
rect 16724 13852 16730 13864
rect 18064 13861 18092 13892
rect 18708 13864 18736 13892
rect 20162 13880 20168 13932
rect 20220 13920 20226 13932
rect 20809 13923 20867 13929
rect 20809 13920 20821 13923
rect 20220 13892 20821 13920
rect 20220 13880 20226 13892
rect 20809 13889 20821 13892
rect 20855 13889 20867 13923
rect 20809 13883 20867 13889
rect 17221 13855 17279 13861
rect 17221 13852 17233 13855
rect 16724 13824 17233 13852
rect 16724 13812 16730 13824
rect 17221 13821 17233 13824
rect 17267 13821 17279 13855
rect 18049 13855 18107 13861
rect 18049 13852 18061 13855
rect 17221 13815 17279 13821
rect 17788 13824 18061 13852
rect 10042 13784 10048 13796
rect 8996 13756 9628 13784
rect 10003 13756 10048 13784
rect 8996 13744 9002 13756
rect 10042 13744 10048 13756
rect 10100 13744 10106 13796
rect 11701 13787 11759 13793
rect 11701 13753 11713 13787
rect 11747 13784 11759 13787
rect 14550 13784 14556 13796
rect 11747 13756 14556 13784
rect 11747 13753 11759 13756
rect 11701 13747 11759 13753
rect 14550 13744 14556 13756
rect 14608 13744 14614 13796
rect 15010 13744 15016 13796
rect 15068 13784 15074 13796
rect 15068 13756 16160 13784
rect 15068 13744 15074 13756
rect 5721 13719 5779 13725
rect 5721 13685 5733 13719
rect 5767 13716 5779 13719
rect 7742 13716 7748 13728
rect 5767 13688 7748 13716
rect 5767 13685 5779 13688
rect 5721 13679 5779 13685
rect 7742 13676 7748 13688
rect 7800 13676 7806 13728
rect 9214 13716 9220 13728
rect 9175 13688 9220 13716
rect 9214 13676 9220 13688
rect 9272 13676 9278 13728
rect 9677 13719 9735 13725
rect 9677 13685 9689 13719
rect 9723 13716 9735 13719
rect 10873 13719 10931 13725
rect 10873 13716 10885 13719
rect 9723 13688 10885 13716
rect 9723 13685 9735 13688
rect 9677 13679 9735 13685
rect 10873 13685 10885 13688
rect 10919 13685 10931 13719
rect 10873 13679 10931 13685
rect 12897 13719 12955 13725
rect 12897 13685 12909 13719
rect 12943 13716 12955 13719
rect 13814 13716 13820 13728
rect 12943 13688 13820 13716
rect 12943 13685 12955 13688
rect 12897 13679 12955 13685
rect 13814 13676 13820 13688
rect 13872 13676 13878 13728
rect 14366 13676 14372 13728
rect 14424 13716 14430 13728
rect 14737 13719 14795 13725
rect 14737 13716 14749 13719
rect 14424 13688 14749 13716
rect 14424 13676 14430 13688
rect 14737 13685 14749 13688
rect 14783 13685 14795 13719
rect 14737 13679 14795 13685
rect 15286 13676 15292 13728
rect 15344 13716 15350 13728
rect 15381 13719 15439 13725
rect 15381 13716 15393 13719
rect 15344 13688 15393 13716
rect 15344 13676 15350 13688
rect 15381 13685 15393 13688
rect 15427 13685 15439 13719
rect 15381 13679 15439 13685
rect 15473 13719 15531 13725
rect 15473 13685 15485 13719
rect 15519 13716 15531 13719
rect 16025 13719 16083 13725
rect 16025 13716 16037 13719
rect 15519 13688 16037 13716
rect 15519 13685 15531 13688
rect 15473 13679 15531 13685
rect 16025 13685 16037 13688
rect 16071 13685 16083 13719
rect 16132 13716 16160 13756
rect 16206 13744 16212 13796
rect 16264 13784 16270 13796
rect 17788 13784 17816 13824
rect 18049 13821 18061 13824
rect 18095 13821 18107 13855
rect 18049 13815 18107 13821
rect 18138 13812 18144 13864
rect 18196 13852 18202 13864
rect 18601 13855 18659 13861
rect 18601 13852 18613 13855
rect 18196 13824 18613 13852
rect 18196 13812 18202 13824
rect 18601 13821 18613 13824
rect 18647 13821 18659 13855
rect 18601 13815 18659 13821
rect 18690 13812 18696 13864
rect 18748 13812 18754 13864
rect 18868 13855 18926 13861
rect 18868 13821 18880 13855
rect 18914 13852 18926 13855
rect 19426 13852 19432 13864
rect 18914 13824 19432 13852
rect 18914 13821 18926 13824
rect 18868 13815 18926 13821
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 20717 13855 20775 13861
rect 20717 13852 20729 13855
rect 19536 13824 20729 13852
rect 18966 13784 18972 13796
rect 16264 13756 17816 13784
rect 18156 13756 18972 13784
rect 16264 13744 16270 13756
rect 16393 13719 16451 13725
rect 16393 13716 16405 13719
rect 16132 13688 16405 13716
rect 16025 13679 16083 13685
rect 16393 13685 16405 13688
rect 16439 13716 16451 13719
rect 18156 13716 18184 13756
rect 18966 13744 18972 13756
rect 19024 13744 19030 13796
rect 19058 13744 19064 13796
rect 19116 13784 19122 13796
rect 19536 13784 19564 13824
rect 20717 13821 20729 13824
rect 20763 13821 20775 13855
rect 20717 13815 20775 13821
rect 19116 13756 19564 13784
rect 19116 13744 19122 13756
rect 16439 13688 18184 13716
rect 18233 13719 18291 13725
rect 16439 13685 16451 13688
rect 16393 13679 16451 13685
rect 18233 13685 18245 13719
rect 18279 13716 18291 13719
rect 18782 13716 18788 13728
rect 18279 13688 18788 13716
rect 18279 13685 18291 13688
rect 18233 13679 18291 13685
rect 18782 13676 18788 13688
rect 18840 13676 18846 13728
rect 19886 13676 19892 13728
rect 19944 13716 19950 13728
rect 19981 13719 20039 13725
rect 19981 13716 19993 13719
rect 19944 13688 19993 13716
rect 19944 13676 19950 13688
rect 19981 13685 19993 13688
rect 20027 13685 20039 13719
rect 20254 13716 20260 13728
rect 20215 13688 20260 13716
rect 19981 13679 20039 13685
rect 20254 13676 20260 13688
rect 20312 13676 20318 13728
rect 20438 13676 20444 13728
rect 20496 13716 20502 13728
rect 20625 13719 20683 13725
rect 20625 13716 20637 13719
rect 20496 13688 20637 13716
rect 20496 13676 20502 13688
rect 20625 13685 20637 13688
rect 20671 13685 20683 13719
rect 20625 13679 20683 13685
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 1762 13512 1768 13524
rect 1723 13484 1768 13512
rect 1762 13472 1768 13484
rect 1820 13472 1826 13524
rect 4433 13515 4491 13521
rect 4433 13481 4445 13515
rect 4479 13512 4491 13515
rect 5813 13515 5871 13521
rect 5813 13512 5825 13515
rect 4479 13484 5825 13512
rect 4479 13481 4491 13484
rect 4433 13475 4491 13481
rect 5813 13481 5825 13484
rect 5859 13481 5871 13515
rect 5813 13475 5871 13481
rect 6454 13472 6460 13524
rect 6512 13512 6518 13524
rect 6914 13512 6920 13524
rect 6512 13484 6920 13512
rect 6512 13472 6518 13484
rect 6914 13472 6920 13484
rect 6972 13472 6978 13524
rect 7285 13515 7343 13521
rect 7285 13481 7297 13515
rect 7331 13512 7343 13515
rect 7374 13512 7380 13524
rect 7331 13484 7380 13512
rect 7331 13481 7343 13484
rect 7285 13475 7343 13481
rect 7374 13472 7380 13484
rect 7432 13472 7438 13524
rect 8846 13512 8852 13524
rect 8759 13484 8852 13512
rect 8846 13472 8852 13484
rect 8904 13512 8910 13524
rect 9398 13512 9404 13524
rect 8904 13484 9404 13512
rect 8904 13472 8910 13484
rect 9398 13472 9404 13484
rect 9456 13472 9462 13524
rect 9858 13472 9864 13524
rect 9916 13512 9922 13524
rect 10226 13512 10232 13524
rect 9916 13484 10232 13512
rect 9916 13472 9922 13484
rect 10226 13472 10232 13484
rect 10284 13472 10290 13524
rect 10870 13472 10876 13524
rect 10928 13512 10934 13524
rect 11425 13515 11483 13521
rect 11425 13512 11437 13515
rect 10928 13484 11437 13512
rect 10928 13472 10934 13484
rect 11425 13481 11437 13484
rect 11471 13512 11483 13515
rect 11471 13484 11805 13512
rect 11471 13481 11483 13484
rect 11425 13475 11483 13481
rect 2130 13404 2136 13456
rect 2188 13444 2194 13456
rect 2225 13447 2283 13453
rect 2225 13444 2237 13447
rect 2188 13416 2237 13444
rect 2188 13404 2194 13416
rect 2225 13413 2237 13416
rect 2271 13444 2283 13447
rect 2777 13447 2835 13453
rect 2777 13444 2789 13447
rect 2271 13416 2789 13444
rect 2271 13413 2283 13416
rect 2225 13407 2283 13413
rect 2777 13413 2789 13416
rect 2823 13444 2835 13447
rect 3142 13444 3148 13456
rect 2823 13416 3148 13444
rect 2823 13413 2835 13416
rect 2777 13407 2835 13413
rect 3142 13404 3148 13416
rect 3200 13404 3206 13456
rect 4062 13404 4068 13456
rect 4120 13444 4126 13456
rect 7736 13447 7794 13453
rect 4120 13416 6960 13444
rect 4120 13404 4126 13416
rect 1578 13376 1584 13388
rect 1539 13348 1584 13376
rect 1578 13336 1584 13348
rect 1636 13336 1642 13388
rect 2406 13336 2412 13388
rect 2464 13376 2470 13388
rect 2685 13379 2743 13385
rect 2685 13376 2697 13379
rect 2464 13348 2697 13376
rect 2464 13336 2470 13348
rect 2685 13345 2697 13348
rect 2731 13345 2743 13379
rect 2685 13339 2743 13345
rect 4246 13336 4252 13388
rect 4304 13376 4310 13388
rect 4801 13379 4859 13385
rect 4801 13376 4813 13379
rect 4304 13348 4813 13376
rect 4304 13336 4310 13348
rect 4801 13345 4813 13348
rect 4847 13345 4859 13379
rect 4801 13339 4859 13345
rect 6638 13336 6644 13388
rect 6696 13376 6702 13388
rect 6825 13379 6883 13385
rect 6825 13376 6837 13379
rect 6696 13348 6837 13376
rect 6696 13336 6702 13348
rect 6825 13345 6837 13348
rect 6871 13345 6883 13379
rect 6932 13376 6960 13416
rect 7736 13413 7748 13447
rect 7782 13444 7794 13447
rect 7834 13444 7840 13456
rect 7782 13416 7840 13444
rect 7782 13413 7794 13416
rect 7736 13407 7794 13413
rect 7834 13404 7840 13416
rect 7892 13444 7898 13456
rect 8754 13444 8760 13456
rect 7892 13416 8760 13444
rect 7892 13404 7898 13416
rect 8754 13404 8760 13416
rect 8812 13404 8818 13456
rect 11777 13453 11805 13484
rect 11882 13472 11888 13524
rect 11940 13512 11946 13524
rect 12618 13512 12624 13524
rect 11940 13484 12624 13512
rect 11940 13472 11946 13484
rect 12618 13472 12624 13484
rect 12676 13472 12682 13524
rect 12986 13512 12992 13524
rect 12947 13484 12992 13512
rect 12986 13472 12992 13484
rect 13044 13472 13050 13524
rect 13449 13515 13507 13521
rect 13449 13481 13461 13515
rect 13495 13481 13507 13515
rect 13449 13475 13507 13481
rect 14829 13515 14887 13521
rect 14829 13481 14841 13515
rect 14875 13512 14887 13515
rect 15102 13512 15108 13524
rect 14875 13484 15108 13512
rect 14875 13481 14887 13484
rect 14829 13475 14887 13481
rect 10312 13447 10370 13453
rect 10312 13413 10324 13447
rect 10358 13444 10370 13447
rect 11762 13447 11820 13453
rect 10358 13416 11652 13444
rect 10358 13413 10370 13416
rect 10312 13407 10370 13413
rect 11514 13376 11520 13388
rect 6932 13348 11100 13376
rect 11475 13348 11520 13376
rect 6825 13339 6883 13345
rect 2961 13311 3019 13317
rect 2961 13277 2973 13311
rect 3007 13308 3019 13311
rect 3418 13308 3424 13320
rect 3007 13280 3424 13308
rect 3007 13277 3019 13280
rect 2961 13271 3019 13277
rect 3418 13268 3424 13280
rect 3476 13268 3482 13320
rect 4706 13268 4712 13320
rect 4764 13308 4770 13320
rect 4893 13311 4951 13317
rect 4893 13308 4905 13311
rect 4764 13280 4905 13308
rect 4764 13268 4770 13280
rect 4893 13277 4905 13280
rect 4939 13277 4951 13311
rect 4893 13271 4951 13277
rect 5077 13311 5135 13317
rect 5077 13277 5089 13311
rect 5123 13308 5135 13311
rect 5258 13308 5264 13320
rect 5123 13280 5264 13308
rect 5123 13277 5135 13280
rect 5077 13271 5135 13277
rect 5258 13268 5264 13280
rect 5316 13268 5322 13320
rect 5902 13308 5908 13320
rect 5863 13280 5908 13308
rect 5902 13268 5908 13280
rect 5960 13268 5966 13320
rect 5994 13268 6000 13320
rect 6052 13308 6058 13320
rect 7101 13311 7159 13317
rect 6052 13280 6097 13308
rect 6052 13268 6058 13280
rect 7101 13277 7113 13311
rect 7147 13308 7159 13311
rect 7374 13308 7380 13320
rect 7147 13280 7380 13308
rect 7147 13277 7159 13280
rect 7101 13271 7159 13277
rect 7374 13268 7380 13280
rect 7432 13268 7438 13320
rect 7469 13311 7527 13317
rect 7469 13277 7481 13311
rect 7515 13277 7527 13311
rect 7469 13271 7527 13277
rect 5442 13240 5448 13252
rect 5403 13212 5448 13240
rect 5442 13200 5448 13212
rect 5500 13200 5506 13252
rect 5626 13200 5632 13252
rect 5684 13240 5690 13252
rect 6822 13240 6828 13252
rect 5684 13212 6828 13240
rect 5684 13200 5690 13212
rect 6822 13200 6828 13212
rect 6880 13200 6886 13252
rect 7285 13243 7343 13249
rect 7285 13209 7297 13243
rect 7331 13240 7343 13243
rect 7484 13240 7512 13271
rect 8478 13268 8484 13320
rect 8536 13308 8542 13320
rect 10045 13311 10103 13317
rect 10045 13308 10057 13311
rect 8536 13280 10057 13308
rect 8536 13268 8542 13280
rect 10045 13277 10057 13280
rect 10091 13277 10103 13311
rect 10045 13271 10103 13277
rect 7331 13212 7512 13240
rect 7331 13209 7343 13212
rect 7285 13203 7343 13209
rect 2317 13175 2375 13181
rect 2317 13141 2329 13175
rect 2363 13172 2375 13175
rect 3142 13172 3148 13184
rect 2363 13144 3148 13172
rect 2363 13141 2375 13144
rect 2317 13135 2375 13141
rect 3142 13132 3148 13144
rect 3200 13132 3206 13184
rect 6457 13175 6515 13181
rect 6457 13141 6469 13175
rect 6503 13172 6515 13175
rect 7742 13172 7748 13184
rect 6503 13144 7748 13172
rect 6503 13141 6515 13144
rect 6457 13135 6515 13141
rect 7742 13132 7748 13144
rect 7800 13132 7806 13184
rect 11072 13172 11100 13348
rect 11514 13336 11520 13348
rect 11572 13336 11578 13388
rect 11624 13376 11652 13416
rect 11762 13413 11774 13447
rect 11808 13413 11820 13447
rect 11762 13407 11820 13413
rect 12894 13404 12900 13456
rect 12952 13444 12958 13456
rect 13464 13444 13492 13475
rect 15102 13472 15108 13484
rect 15160 13472 15166 13524
rect 15286 13512 15292 13524
rect 15247 13484 15292 13512
rect 15286 13472 15292 13484
rect 15344 13472 15350 13524
rect 15562 13472 15568 13524
rect 15620 13512 15626 13524
rect 16117 13515 16175 13521
rect 15620 13484 15792 13512
rect 15620 13472 15626 13484
rect 12952 13416 13492 13444
rect 12952 13404 12958 13416
rect 13814 13404 13820 13456
rect 13872 13444 13878 13456
rect 15764 13453 15792 13484
rect 16117 13481 16129 13515
rect 16163 13512 16175 13515
rect 16390 13512 16396 13524
rect 16163 13484 16396 13512
rect 16163 13481 16175 13484
rect 16117 13475 16175 13481
rect 16390 13472 16396 13484
rect 16448 13512 16454 13524
rect 17681 13515 17739 13521
rect 17681 13512 17693 13515
rect 16448 13484 17693 13512
rect 16448 13472 16454 13484
rect 17681 13481 17693 13484
rect 17727 13481 17739 13515
rect 19610 13512 19616 13524
rect 19571 13484 19616 13512
rect 17681 13475 17739 13481
rect 19610 13472 19616 13484
rect 19668 13472 19674 13524
rect 15657 13447 15715 13453
rect 15657 13444 15669 13447
rect 13872 13416 15669 13444
rect 13872 13404 13878 13416
rect 15657 13413 15669 13416
rect 15703 13413 15715 13447
rect 15657 13407 15715 13413
rect 15749 13447 15807 13453
rect 15749 13413 15761 13447
rect 15795 13444 15807 13447
rect 16298 13444 16304 13456
rect 15795 13416 16304 13444
rect 15795 13413 15807 13416
rect 15749 13407 15807 13413
rect 16298 13404 16304 13416
rect 16356 13404 16362 13456
rect 16568 13447 16626 13453
rect 16568 13413 16580 13447
rect 16614 13444 16626 13447
rect 19886 13444 19892 13456
rect 16614 13416 19892 13444
rect 16614 13413 16626 13416
rect 16568 13407 16626 13413
rect 19886 13404 19892 13416
rect 19944 13444 19950 13456
rect 19944 13416 20208 13444
rect 19944 13404 19950 13416
rect 11624 13348 12756 13376
rect 11882 13172 11888 13184
rect 11072 13144 11888 13172
rect 11882 13132 11888 13144
rect 11940 13132 11946 13184
rect 12728 13172 12756 13348
rect 12802 13336 12808 13388
rect 12860 13376 12866 13388
rect 13357 13379 13415 13385
rect 13357 13376 13369 13379
rect 12860 13348 13369 13376
rect 12860 13336 12866 13348
rect 13357 13345 13369 13348
rect 13403 13345 13415 13379
rect 13357 13339 13415 13345
rect 14185 13379 14243 13385
rect 14185 13345 14197 13379
rect 14231 13376 14243 13379
rect 14645 13379 14703 13385
rect 14231 13348 14596 13376
rect 14231 13345 14243 13348
rect 14185 13339 14243 13345
rect 13538 13268 13544 13320
rect 13596 13308 13602 13320
rect 13633 13311 13691 13317
rect 13633 13308 13645 13311
rect 13596 13280 13645 13308
rect 13596 13268 13602 13280
rect 13633 13277 13645 13280
rect 13679 13308 13691 13311
rect 14274 13308 14280 13320
rect 13679 13280 14136 13308
rect 14235 13280 14280 13308
rect 13679 13277 13691 13280
rect 13633 13271 13691 13277
rect 12897 13243 12955 13249
rect 12897 13209 12909 13243
rect 12943 13240 12955 13243
rect 13170 13240 13176 13252
rect 12943 13212 13176 13240
rect 12943 13209 12955 13212
rect 12897 13203 12955 13209
rect 13170 13200 13176 13212
rect 13228 13200 13234 13252
rect 14108 13240 14136 13280
rect 14274 13268 14280 13280
rect 14332 13268 14338 13320
rect 14458 13308 14464 13320
rect 14419 13280 14464 13308
rect 14458 13268 14464 13280
rect 14516 13268 14522 13320
rect 14568 13308 14596 13348
rect 14645 13345 14657 13379
rect 14691 13376 14703 13379
rect 17862 13376 17868 13388
rect 14691 13348 17868 13376
rect 14691 13345 14703 13348
rect 14645 13339 14703 13345
rect 17862 13336 17868 13348
rect 17920 13336 17926 13388
rect 18046 13376 18052 13388
rect 17972 13348 18052 13376
rect 15286 13308 15292 13320
rect 14568 13280 15292 13308
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 15933 13311 15991 13317
rect 15933 13277 15945 13311
rect 15979 13308 15991 13311
rect 16117 13311 16175 13317
rect 16117 13308 16129 13311
rect 15979 13280 16129 13308
rect 15979 13277 15991 13280
rect 15933 13271 15991 13277
rect 16117 13277 16129 13280
rect 16163 13277 16175 13311
rect 16298 13308 16304 13320
rect 16259 13280 16304 13308
rect 16117 13271 16175 13277
rect 15948 13240 15976 13271
rect 16298 13268 16304 13280
rect 16356 13268 16362 13320
rect 17770 13268 17776 13320
rect 17828 13308 17834 13320
rect 17972 13317 18000 13348
rect 18046 13336 18052 13348
rect 18104 13336 18110 13388
rect 18230 13385 18236 13388
rect 18224 13376 18236 13385
rect 18191 13348 18236 13376
rect 18224 13339 18236 13348
rect 18288 13376 18294 13388
rect 19150 13376 19156 13388
rect 18288 13348 19156 13376
rect 18230 13336 18236 13339
rect 18288 13336 18294 13348
rect 19150 13336 19156 13348
rect 19208 13336 19214 13388
rect 19610 13336 19616 13388
rect 19668 13376 19674 13388
rect 19981 13379 20039 13385
rect 19981 13376 19993 13379
rect 19668 13348 19993 13376
rect 19668 13336 19674 13348
rect 19981 13345 19993 13348
rect 20027 13345 20039 13379
rect 19981 13339 20039 13345
rect 17957 13311 18015 13317
rect 17957 13308 17969 13311
rect 17828 13280 17969 13308
rect 17828 13268 17834 13280
rect 17957 13277 17969 13280
rect 18003 13277 18015 13311
rect 17957 13271 18015 13277
rect 18966 13268 18972 13320
rect 19024 13308 19030 13320
rect 20180 13317 20208 13416
rect 20073 13311 20131 13317
rect 20073 13308 20085 13311
rect 19024 13280 20085 13308
rect 19024 13268 19030 13280
rect 20073 13277 20085 13280
rect 20119 13277 20131 13311
rect 20073 13271 20131 13277
rect 20165 13311 20223 13317
rect 20165 13277 20177 13311
rect 20211 13277 20223 13311
rect 20165 13271 20223 13277
rect 13648 13212 14044 13240
rect 14108 13212 15976 13240
rect 13648 13172 13676 13212
rect 12728 13144 13676 13172
rect 13722 13132 13728 13184
rect 13780 13172 13786 13184
rect 13817 13175 13875 13181
rect 13817 13172 13829 13175
rect 13780 13144 13829 13172
rect 13780 13132 13786 13144
rect 13817 13141 13829 13144
rect 13863 13141 13875 13175
rect 14016 13172 14044 13212
rect 17494 13172 17500 13184
rect 14016 13144 17500 13172
rect 13817 13135 13875 13141
rect 17494 13132 17500 13144
rect 17552 13132 17558 13184
rect 19337 13175 19395 13181
rect 19337 13141 19349 13175
rect 19383 13172 19395 13175
rect 19426 13172 19432 13184
rect 19383 13144 19432 13172
rect 19383 13141 19395 13144
rect 19337 13135 19395 13141
rect 19426 13132 19432 13144
rect 19484 13132 19490 13184
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 1949 12971 2007 12977
rect 1949 12937 1961 12971
rect 1995 12968 2007 12971
rect 2774 12968 2780 12980
rect 1995 12940 2780 12968
rect 1995 12937 2007 12940
rect 1949 12931 2007 12937
rect 2774 12928 2780 12940
rect 2832 12928 2838 12980
rect 4709 12971 4767 12977
rect 4709 12937 4721 12971
rect 4755 12968 4767 12971
rect 5902 12968 5908 12980
rect 4755 12940 5908 12968
rect 4755 12937 4767 12940
rect 4709 12931 4767 12937
rect 5902 12928 5908 12940
rect 5960 12928 5966 12980
rect 7193 12971 7251 12977
rect 7193 12937 7205 12971
rect 7239 12968 7251 12971
rect 9214 12968 9220 12980
rect 7239 12940 9220 12968
rect 7239 12937 7251 12940
rect 7193 12931 7251 12937
rect 9214 12928 9220 12940
rect 9272 12928 9278 12980
rect 11698 12928 11704 12980
rect 11756 12968 11762 12980
rect 12066 12968 12072 12980
rect 11756 12940 12072 12968
rect 11756 12928 11762 12940
rect 12066 12928 12072 12940
rect 12124 12928 12130 12980
rect 15746 12968 15752 12980
rect 14108 12940 15752 12968
rect 3881 12903 3939 12909
rect 3881 12869 3893 12903
rect 3927 12900 3939 12903
rect 5721 12903 5779 12909
rect 3927 12872 5304 12900
rect 3927 12869 3939 12872
rect 3881 12863 3939 12869
rect 5276 12844 5304 12872
rect 5721 12869 5733 12903
rect 5767 12900 5779 12903
rect 5994 12900 6000 12912
rect 5767 12872 6000 12900
rect 5767 12869 5779 12872
rect 5721 12863 5779 12869
rect 5994 12860 6000 12872
rect 6052 12860 6058 12912
rect 7098 12860 7104 12912
rect 7156 12900 7162 12912
rect 7466 12900 7472 12912
rect 7156 12872 7472 12900
rect 7156 12860 7162 12872
rect 7466 12860 7472 12872
rect 7524 12860 7530 12912
rect 8021 12903 8079 12909
rect 8021 12869 8033 12903
rect 8067 12900 8079 12903
rect 8205 12903 8263 12909
rect 8205 12900 8217 12903
rect 8067 12872 8217 12900
rect 8067 12869 8079 12872
rect 8021 12863 8079 12869
rect 8205 12869 8217 12872
rect 8251 12869 8263 12903
rect 8205 12863 8263 12869
rect 8294 12860 8300 12912
rect 8352 12900 8358 12912
rect 9677 12903 9735 12909
rect 9677 12900 9689 12903
rect 8352 12872 9689 12900
rect 8352 12860 8358 12872
rect 9677 12869 9689 12872
rect 9723 12869 9735 12903
rect 13538 12900 13544 12912
rect 9677 12863 9735 12869
rect 9784 12872 13544 12900
rect 4246 12832 4252 12844
rect 4207 12804 4252 12832
rect 4246 12792 4252 12804
rect 4304 12792 4310 12844
rect 5258 12832 5264 12844
rect 5219 12804 5264 12832
rect 5258 12792 5264 12804
rect 5316 12792 5322 12844
rect 6270 12832 6276 12844
rect 6231 12804 6276 12832
rect 6270 12792 6276 12804
rect 6328 12792 6334 12844
rect 7653 12835 7711 12841
rect 7653 12801 7665 12835
rect 7699 12832 7711 12835
rect 7742 12832 7748 12844
rect 7699 12804 7748 12832
rect 7699 12801 7711 12804
rect 7653 12795 7711 12801
rect 7742 12792 7748 12804
rect 7800 12792 7806 12844
rect 7834 12792 7840 12844
rect 7892 12832 7898 12844
rect 8849 12835 8907 12841
rect 7892 12804 7937 12832
rect 7892 12792 7898 12804
rect 8849 12801 8861 12835
rect 8895 12832 8907 12835
rect 8938 12832 8944 12844
rect 8895 12804 8944 12832
rect 8895 12801 8907 12804
rect 8849 12795 8907 12801
rect 8938 12792 8944 12804
rect 8996 12792 9002 12844
rect 1765 12767 1823 12773
rect 1765 12733 1777 12767
rect 1811 12764 1823 12767
rect 1854 12764 1860 12776
rect 1811 12736 1860 12764
rect 1811 12733 1823 12736
rect 1765 12727 1823 12733
rect 1854 12724 1860 12736
rect 1912 12724 1918 12776
rect 2501 12767 2559 12773
rect 2501 12733 2513 12767
rect 2547 12764 2559 12767
rect 2590 12764 2596 12776
rect 2547 12736 2596 12764
rect 2547 12733 2559 12736
rect 2501 12727 2559 12733
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 4982 12724 4988 12776
rect 5040 12764 5046 12776
rect 5169 12767 5227 12773
rect 5169 12764 5181 12767
rect 5040 12736 5181 12764
rect 5040 12724 5046 12736
rect 5169 12733 5181 12736
rect 5215 12733 5227 12767
rect 5169 12727 5227 12733
rect 5350 12724 5356 12776
rect 5408 12764 5414 12776
rect 8665 12767 8723 12773
rect 8665 12764 8677 12767
rect 5408 12736 8677 12764
rect 5408 12724 5414 12736
rect 8665 12733 8677 12736
rect 8711 12733 8723 12767
rect 8665 12727 8723 12733
rect 8754 12724 8760 12776
rect 8812 12764 8818 12776
rect 9784 12764 9812 12872
rect 13538 12860 13544 12872
rect 13596 12860 13602 12912
rect 13722 12832 13728 12844
rect 13683 12804 13728 12832
rect 13722 12792 13728 12804
rect 13780 12792 13786 12844
rect 14108 12841 14136 12940
rect 15746 12928 15752 12940
rect 15804 12968 15810 12980
rect 16022 12968 16028 12980
rect 15804 12940 16028 12968
rect 15804 12928 15810 12940
rect 16022 12928 16028 12940
rect 16080 12968 16086 12980
rect 16298 12968 16304 12980
rect 16080 12940 16304 12968
rect 16080 12928 16086 12940
rect 16298 12928 16304 12940
rect 16356 12968 16362 12980
rect 16758 12968 16764 12980
rect 16356 12940 16764 12968
rect 16356 12928 16362 12940
rect 16758 12928 16764 12940
rect 16816 12968 16822 12980
rect 17770 12968 17776 12980
rect 16816 12940 17776 12968
rect 16816 12928 16822 12940
rect 17770 12928 17776 12940
rect 17828 12928 17834 12980
rect 18966 12968 18972 12980
rect 18927 12940 18972 12968
rect 18966 12928 18972 12940
rect 19024 12928 19030 12980
rect 20162 12928 20168 12980
rect 20220 12928 20226 12980
rect 15470 12860 15476 12912
rect 15528 12900 15534 12912
rect 16850 12900 16856 12912
rect 15528 12872 16856 12900
rect 15528 12860 15534 12872
rect 16850 12860 16856 12872
rect 16908 12860 16914 12912
rect 16945 12903 17003 12909
rect 16945 12869 16957 12903
rect 16991 12869 17003 12903
rect 16945 12863 17003 12869
rect 13817 12835 13875 12841
rect 13817 12801 13829 12835
rect 13863 12801 13875 12835
rect 13817 12795 13875 12801
rect 14093 12835 14151 12841
rect 14093 12801 14105 12835
rect 14139 12801 14151 12835
rect 14093 12795 14151 12801
rect 15841 12835 15899 12841
rect 15841 12801 15853 12835
rect 15887 12832 15899 12835
rect 16114 12832 16120 12844
rect 15887 12804 16120 12832
rect 15887 12801 15899 12804
rect 15841 12795 15899 12801
rect 8812 12736 9812 12764
rect 9861 12767 9919 12773
rect 8812 12724 8818 12736
rect 9861 12733 9873 12767
rect 9907 12764 9919 12767
rect 11977 12767 12035 12773
rect 11977 12764 11989 12767
rect 9907 12736 11989 12764
rect 9907 12733 9919 12736
rect 9861 12727 9919 12733
rect 11977 12733 11989 12736
rect 12023 12764 12035 12767
rect 12989 12767 13047 12773
rect 12989 12764 13001 12767
rect 12023 12736 13001 12764
rect 12023 12733 12035 12736
rect 11977 12727 12035 12733
rect 12989 12733 13001 12736
rect 13035 12733 13047 12767
rect 12989 12727 13047 12733
rect 13630 12724 13636 12776
rect 13688 12764 13694 12776
rect 13832 12764 13860 12795
rect 16114 12792 16120 12804
rect 16172 12792 16178 12844
rect 16390 12792 16396 12844
rect 16448 12832 16454 12844
rect 16485 12835 16543 12841
rect 16485 12832 16497 12835
rect 16448 12804 16497 12832
rect 16448 12792 16454 12804
rect 16485 12801 16497 12804
rect 16531 12801 16543 12835
rect 16485 12795 16543 12801
rect 14366 12773 14372 12776
rect 13688 12736 13860 12764
rect 13688 12724 13694 12736
rect 14360 12727 14372 12773
rect 14424 12764 14430 12776
rect 16666 12764 16672 12776
rect 14424 12736 14460 12764
rect 15212 12736 16672 12764
rect 14366 12724 14372 12727
rect 14424 12724 14430 12736
rect 2768 12699 2826 12705
rect 2768 12665 2780 12699
rect 2814 12696 2826 12699
rect 2958 12696 2964 12708
rect 2814 12668 2964 12696
rect 2814 12665 2826 12668
rect 2768 12659 2826 12665
rect 2958 12656 2964 12668
rect 3016 12656 3022 12708
rect 6178 12696 6184 12708
rect 4908 12668 6184 12696
rect 2498 12588 2504 12640
rect 2556 12628 2562 12640
rect 4908 12628 4936 12668
rect 6178 12656 6184 12668
rect 6236 12656 6242 12708
rect 7561 12699 7619 12705
rect 7561 12665 7573 12699
rect 7607 12696 7619 12699
rect 8021 12699 8079 12705
rect 8021 12696 8033 12699
rect 7607 12668 8033 12696
rect 7607 12665 7619 12668
rect 7561 12659 7619 12665
rect 8021 12665 8033 12668
rect 8067 12665 8079 12699
rect 8021 12659 8079 12665
rect 8573 12699 8631 12705
rect 8573 12665 8585 12699
rect 8619 12696 8631 12699
rect 9217 12699 9275 12705
rect 9217 12696 9229 12699
rect 8619 12668 9229 12696
rect 8619 12665 8631 12668
rect 8573 12659 8631 12665
rect 9217 12665 9229 12668
rect 9263 12665 9275 12699
rect 9217 12659 9275 12665
rect 10413 12699 10471 12705
rect 10413 12665 10425 12699
rect 10459 12665 10471 12699
rect 15212 12696 15240 12736
rect 16666 12724 16672 12736
rect 16724 12724 16730 12776
rect 16960 12764 16988 12863
rect 19150 12860 19156 12912
rect 19208 12900 19214 12912
rect 19334 12900 19340 12912
rect 19208 12872 19340 12900
rect 19208 12860 19214 12872
rect 19334 12860 19340 12872
rect 19392 12900 19398 12912
rect 20180 12900 20208 12928
rect 19392 12872 20576 12900
rect 19392 12860 19398 12872
rect 17494 12832 17500 12844
rect 17455 12804 17500 12832
rect 17494 12792 17500 12804
rect 17552 12792 17558 12844
rect 17862 12792 17868 12844
rect 17920 12832 17926 12844
rect 18417 12835 18475 12841
rect 18417 12832 18429 12835
rect 17920 12804 18429 12832
rect 17920 12792 17926 12804
rect 18417 12801 18429 12804
rect 18463 12801 18475 12835
rect 18417 12795 18475 12801
rect 19426 12792 19432 12844
rect 19484 12832 19490 12844
rect 19613 12835 19671 12841
rect 19613 12832 19625 12835
rect 19484 12804 19625 12832
rect 19484 12792 19490 12804
rect 19613 12801 19625 12804
rect 19659 12832 19671 12835
rect 20162 12832 20168 12844
rect 19659 12804 20168 12832
rect 19659 12801 19671 12804
rect 19613 12795 19671 12801
rect 20162 12792 20168 12804
rect 20220 12792 20226 12844
rect 20548 12841 20576 12872
rect 20533 12835 20591 12841
rect 20533 12801 20545 12835
rect 20579 12801 20591 12835
rect 20533 12795 20591 12801
rect 18233 12767 18291 12773
rect 18233 12764 18245 12767
rect 16960 12736 18245 12764
rect 18233 12733 18245 12736
rect 18279 12733 18291 12767
rect 18233 12727 18291 12733
rect 19337 12767 19395 12773
rect 19337 12733 19349 12767
rect 19383 12764 19395 12767
rect 20254 12764 20260 12776
rect 19383 12736 20260 12764
rect 19383 12733 19395 12736
rect 19337 12727 19395 12733
rect 20254 12724 20260 12736
rect 20312 12724 20318 12776
rect 10413 12659 10471 12665
rect 13280 12668 15240 12696
rect 5074 12628 5080 12640
rect 2556 12600 4936 12628
rect 5035 12600 5080 12628
rect 2556 12588 2562 12600
rect 5074 12588 5080 12600
rect 5132 12588 5138 12640
rect 5810 12588 5816 12640
rect 5868 12628 5874 12640
rect 6089 12631 6147 12637
rect 6089 12628 6101 12631
rect 5868 12600 6101 12628
rect 5868 12588 5874 12600
rect 6089 12597 6101 12600
rect 6135 12597 6147 12631
rect 6089 12591 6147 12597
rect 6546 12588 6552 12640
rect 6604 12628 6610 12640
rect 10428 12628 10456 12659
rect 6604 12600 10456 12628
rect 12805 12631 12863 12637
rect 6604 12588 6610 12600
rect 12805 12597 12817 12631
rect 12851 12628 12863 12631
rect 12986 12628 12992 12640
rect 12851 12600 12992 12628
rect 12851 12597 12863 12600
rect 12805 12591 12863 12597
rect 12986 12588 12992 12600
rect 13044 12588 13050 12640
rect 13280 12637 13308 12668
rect 15562 12656 15568 12708
rect 15620 12696 15626 12708
rect 16301 12699 16359 12705
rect 16301 12696 16313 12699
rect 15620 12668 16313 12696
rect 15620 12656 15626 12668
rect 16301 12665 16313 12668
rect 16347 12665 16359 12699
rect 17310 12696 17316 12708
rect 17271 12668 17316 12696
rect 16301 12659 16359 12665
rect 17310 12656 17316 12668
rect 17368 12656 17374 12708
rect 17405 12699 17463 12705
rect 17405 12665 17417 12699
rect 17451 12696 17463 12699
rect 17586 12696 17592 12708
rect 17451 12668 17592 12696
rect 17451 12665 17463 12668
rect 17405 12659 17463 12665
rect 17586 12656 17592 12668
rect 17644 12656 17650 12708
rect 19429 12699 19487 12705
rect 19429 12665 19441 12699
rect 19475 12696 19487 12699
rect 19518 12696 19524 12708
rect 19475 12668 19524 12696
rect 19475 12665 19487 12668
rect 19429 12659 19487 12665
rect 19518 12656 19524 12668
rect 19576 12656 19582 12708
rect 20349 12699 20407 12705
rect 19628 12668 20116 12696
rect 13265 12631 13323 12637
rect 13265 12597 13277 12631
rect 13311 12597 13323 12631
rect 13265 12591 13323 12597
rect 13633 12631 13691 12637
rect 13633 12597 13645 12631
rect 13679 12628 13691 12631
rect 13998 12628 14004 12640
rect 13679 12600 14004 12628
rect 13679 12597 13691 12600
rect 13633 12591 13691 12597
rect 13998 12588 14004 12600
rect 14056 12588 14062 12640
rect 15470 12628 15476 12640
rect 15431 12600 15476 12628
rect 15470 12588 15476 12600
rect 15528 12588 15534 12640
rect 15838 12588 15844 12640
rect 15896 12628 15902 12640
rect 15933 12631 15991 12637
rect 15933 12628 15945 12631
rect 15896 12600 15945 12628
rect 15896 12588 15902 12600
rect 15933 12597 15945 12600
rect 15979 12597 15991 12631
rect 15933 12591 15991 12597
rect 16114 12588 16120 12640
rect 16172 12628 16178 12640
rect 16393 12631 16451 12637
rect 16393 12628 16405 12631
rect 16172 12600 16405 12628
rect 16172 12588 16178 12600
rect 16393 12597 16405 12600
rect 16439 12597 16451 12631
rect 16393 12591 16451 12597
rect 16666 12588 16672 12640
rect 16724 12628 16730 12640
rect 18966 12628 18972 12640
rect 16724 12600 18972 12628
rect 16724 12588 16730 12600
rect 18966 12588 18972 12600
rect 19024 12628 19030 12640
rect 19628 12628 19656 12668
rect 19978 12628 19984 12640
rect 19024 12600 19656 12628
rect 19939 12600 19984 12628
rect 19024 12588 19030 12600
rect 19978 12588 19984 12600
rect 20036 12588 20042 12640
rect 20088 12628 20116 12668
rect 20349 12665 20361 12699
rect 20395 12696 20407 12699
rect 20898 12696 20904 12708
rect 20395 12668 20904 12696
rect 20395 12665 20407 12668
rect 20349 12659 20407 12665
rect 20898 12656 20904 12668
rect 20956 12656 20962 12708
rect 20441 12631 20499 12637
rect 20441 12628 20453 12631
rect 20088 12600 20453 12628
rect 20441 12597 20453 12600
rect 20487 12597 20499 12631
rect 20441 12591 20499 12597
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 2958 12424 2964 12436
rect 2919 12396 2964 12424
rect 2958 12384 2964 12396
rect 3016 12384 3022 12436
rect 4062 12384 4068 12436
rect 4120 12424 4126 12436
rect 11882 12424 11888 12436
rect 4120 12396 11888 12424
rect 4120 12384 4126 12396
rect 11882 12384 11888 12396
rect 11940 12384 11946 12436
rect 12621 12427 12679 12433
rect 12621 12393 12633 12427
rect 12667 12424 12679 12427
rect 12667 12396 13207 12424
rect 12667 12393 12679 12396
rect 12621 12387 12679 12393
rect 2590 12356 2596 12368
rect 1596 12328 2596 12356
rect 1486 12248 1492 12300
rect 1544 12288 1550 12300
rect 1596 12297 1624 12328
rect 2590 12316 2596 12328
rect 2648 12316 2654 12368
rect 4792 12359 4850 12365
rect 4792 12325 4804 12359
rect 4838 12356 4850 12359
rect 5442 12356 5448 12368
rect 4838 12328 5448 12356
rect 4838 12325 4850 12328
rect 4792 12319 4850 12325
rect 5442 12316 5448 12328
rect 5500 12316 5506 12368
rect 10594 12356 10600 12368
rect 5552 12328 9444 12356
rect 10555 12328 10600 12356
rect 1581 12291 1639 12297
rect 1581 12288 1593 12291
rect 1544 12260 1593 12288
rect 1544 12248 1550 12260
rect 1581 12257 1593 12260
rect 1627 12257 1639 12291
rect 1581 12251 1639 12257
rect 1848 12291 1906 12297
rect 1848 12257 1860 12291
rect 1894 12288 1906 12291
rect 2314 12288 2320 12300
rect 1894 12260 2320 12288
rect 1894 12257 1906 12260
rect 1848 12251 1906 12257
rect 2314 12248 2320 12260
rect 2372 12248 2378 12300
rect 3970 12248 3976 12300
rect 4028 12288 4034 12300
rect 5552 12288 5580 12328
rect 6437 12291 6495 12297
rect 6437 12288 6449 12291
rect 4028 12260 5580 12288
rect 5920 12260 6449 12288
rect 4028 12248 4034 12260
rect 2590 12180 2596 12232
rect 2648 12220 2654 12232
rect 4062 12220 4068 12232
rect 2648 12192 4068 12220
rect 2648 12180 2654 12192
rect 4062 12180 4068 12192
rect 4120 12220 4126 12232
rect 4522 12220 4528 12232
rect 4120 12192 4528 12220
rect 4120 12180 4126 12192
rect 4522 12180 4528 12192
rect 4580 12180 4586 12232
rect 5258 12044 5264 12096
rect 5316 12084 5322 12096
rect 5920 12093 5948 12260
rect 6437 12257 6449 12260
rect 6483 12257 6495 12291
rect 8104 12291 8162 12297
rect 8104 12288 8116 12291
rect 6437 12251 6495 12257
rect 7576 12260 8116 12288
rect 6178 12220 6184 12232
rect 6139 12192 6184 12220
rect 6178 12180 6184 12192
rect 6236 12180 6242 12232
rect 7576 12161 7604 12260
rect 8104 12257 8116 12260
rect 8150 12288 8162 12291
rect 9306 12288 9312 12300
rect 8150 12260 9312 12288
rect 8150 12257 8162 12260
rect 8104 12251 8162 12257
rect 9306 12248 9312 12260
rect 9364 12248 9370 12300
rect 9416 12288 9444 12328
rect 10594 12316 10600 12328
rect 10652 12356 10658 12368
rect 10870 12356 10876 12368
rect 10652 12328 10876 12356
rect 10652 12316 10658 12328
rect 10870 12316 10876 12328
rect 10928 12316 10934 12368
rect 12342 12316 12348 12368
rect 12400 12356 12406 12368
rect 13179 12365 13207 12396
rect 13630 12384 13636 12436
rect 13688 12424 13694 12436
rect 14277 12427 14335 12433
rect 14277 12424 14289 12427
rect 13688 12396 14289 12424
rect 13688 12384 13694 12396
rect 14277 12393 14289 12396
rect 14323 12393 14335 12427
rect 15286 12424 15292 12436
rect 15247 12396 15292 12424
rect 14277 12387 14335 12393
rect 15286 12384 15292 12396
rect 15344 12384 15350 12436
rect 15657 12427 15715 12433
rect 15657 12393 15669 12427
rect 15703 12424 15715 12427
rect 15703 12396 17448 12424
rect 15703 12393 15715 12396
rect 15657 12387 15715 12393
rect 13164 12359 13222 12365
rect 12400 12328 12940 12356
rect 12400 12316 12406 12328
rect 10778 12288 10784 12300
rect 9416 12260 10784 12288
rect 10778 12248 10784 12260
rect 10836 12248 10842 12300
rect 11508 12291 11566 12297
rect 11508 12288 11520 12291
rect 11072 12260 11520 12288
rect 7834 12220 7840 12232
rect 7795 12192 7840 12220
rect 7834 12180 7840 12192
rect 7892 12180 7898 12232
rect 10689 12223 10747 12229
rect 10689 12220 10701 12223
rect 9140 12192 10701 12220
rect 7561 12155 7619 12161
rect 7561 12121 7573 12155
rect 7607 12121 7619 12155
rect 7561 12115 7619 12121
rect 5905 12087 5963 12093
rect 5905 12084 5917 12087
rect 5316 12056 5917 12084
rect 5316 12044 5322 12056
rect 5905 12053 5917 12056
rect 5951 12053 5963 12087
rect 5905 12047 5963 12053
rect 6086 12044 6092 12096
rect 6144 12084 6150 12096
rect 6454 12084 6460 12096
rect 6144 12056 6460 12084
rect 6144 12044 6150 12056
rect 6454 12044 6460 12056
rect 6512 12044 6518 12096
rect 7190 12044 7196 12096
rect 7248 12084 7254 12096
rect 9140 12084 9168 12192
rect 10689 12189 10701 12192
rect 10735 12189 10747 12223
rect 10689 12183 10747 12189
rect 10873 12223 10931 12229
rect 10873 12189 10885 12223
rect 10919 12220 10931 12223
rect 11072 12220 11100 12260
rect 11508 12257 11520 12260
rect 11554 12288 11566 12291
rect 12434 12288 12440 12300
rect 11554 12260 12440 12288
rect 11554 12257 11566 12260
rect 11508 12251 11566 12257
rect 12434 12248 12440 12260
rect 12492 12248 12498 12300
rect 12912 12297 12940 12328
rect 13164 12325 13176 12359
rect 13210 12356 13222 12359
rect 14458 12356 14464 12368
rect 13210 12328 14464 12356
rect 13210 12325 13222 12328
rect 13164 12319 13222 12325
rect 14458 12316 14464 12328
rect 14516 12316 14522 12368
rect 14737 12359 14795 12365
rect 14737 12325 14749 12359
rect 14783 12356 14795 12359
rect 15562 12356 15568 12368
rect 14783 12328 15568 12356
rect 14783 12325 14795 12328
rect 14737 12319 14795 12325
rect 15562 12316 15568 12328
rect 15620 12316 15626 12368
rect 17420 12356 17448 12396
rect 17494 12384 17500 12436
rect 17552 12424 17558 12436
rect 17865 12427 17923 12433
rect 17865 12424 17877 12427
rect 17552 12396 17877 12424
rect 17552 12384 17558 12396
rect 17865 12393 17877 12396
rect 17911 12393 17923 12427
rect 19610 12424 19616 12436
rect 19571 12396 19616 12424
rect 17865 12387 17923 12393
rect 19610 12384 19616 12396
rect 19668 12384 19674 12436
rect 19978 12424 19984 12436
rect 19939 12396 19984 12424
rect 19978 12384 19984 12396
rect 20036 12384 20042 12436
rect 20898 12424 20904 12436
rect 20859 12396 20904 12424
rect 20898 12384 20904 12396
rect 20956 12384 20962 12436
rect 18506 12356 18512 12368
rect 17420 12328 18512 12356
rect 18506 12316 18512 12328
rect 18564 12316 18570 12368
rect 12897 12291 12955 12297
rect 12897 12257 12909 12291
rect 12943 12257 12955 12291
rect 15749 12291 15807 12297
rect 15749 12288 15761 12291
rect 12897 12251 12955 12257
rect 13004 12260 15761 12288
rect 10919 12192 11100 12220
rect 10919 12189 10931 12192
rect 10873 12183 10931 12189
rect 10704 12152 10732 12183
rect 11146 12180 11152 12232
rect 11204 12220 11210 12232
rect 11241 12223 11299 12229
rect 11241 12220 11253 12223
rect 11204 12192 11253 12220
rect 11204 12180 11210 12192
rect 11241 12189 11253 12192
rect 11287 12189 11299 12223
rect 11241 12183 11299 12189
rect 12710 12180 12716 12232
rect 12768 12220 12774 12232
rect 13004 12220 13032 12260
rect 15749 12257 15761 12260
rect 15795 12257 15807 12291
rect 15749 12251 15807 12257
rect 16114 12248 16120 12300
rect 16172 12288 16178 12300
rect 16485 12291 16543 12297
rect 16485 12288 16497 12291
rect 16172 12260 16497 12288
rect 16172 12248 16178 12260
rect 16485 12257 16497 12260
rect 16531 12257 16543 12291
rect 16485 12251 16543 12257
rect 16752 12291 16810 12297
rect 16752 12257 16764 12291
rect 16798 12288 16810 12291
rect 17034 12288 17040 12300
rect 16798 12260 17040 12288
rect 16798 12257 16810 12260
rect 16752 12251 16810 12257
rect 17034 12248 17040 12260
rect 17092 12248 17098 12300
rect 18969 12291 19027 12297
rect 18969 12288 18981 12291
rect 17512 12260 18981 12288
rect 12768 12192 13032 12220
rect 15933 12223 15991 12229
rect 12768 12180 12774 12192
rect 15933 12189 15945 12223
rect 15979 12220 15991 12223
rect 16390 12220 16396 12232
rect 15979 12192 16396 12220
rect 15979 12189 15991 12192
rect 15933 12183 15991 12189
rect 10962 12152 10968 12164
rect 10704 12124 10968 12152
rect 10962 12112 10968 12124
rect 11020 12112 11026 12164
rect 7248 12056 9168 12084
rect 7248 12044 7254 12056
rect 9214 12044 9220 12096
rect 9272 12084 9278 12096
rect 10229 12087 10287 12093
rect 9272 12056 9317 12084
rect 9272 12044 9278 12056
rect 10229 12053 10241 12087
rect 10275 12084 10287 12087
rect 14274 12084 14280 12096
rect 10275 12056 14280 12084
rect 10275 12053 10287 12056
rect 10229 12047 10287 12053
rect 14274 12044 14280 12056
rect 14332 12044 14338 12096
rect 15470 12044 15476 12096
rect 15528 12084 15534 12096
rect 16132 12084 16160 12192
rect 16390 12180 16396 12192
rect 16448 12180 16454 12232
rect 15528 12056 16160 12084
rect 15528 12044 15534 12056
rect 16390 12044 16396 12096
rect 16448 12084 16454 12096
rect 17512 12084 17540 12260
rect 18969 12257 18981 12260
rect 19015 12257 19027 12291
rect 18969 12251 19027 12257
rect 19061 12291 19119 12297
rect 19061 12257 19073 12291
rect 19107 12288 19119 12291
rect 19610 12288 19616 12300
rect 19107 12260 19616 12288
rect 19107 12257 19119 12260
rect 19061 12251 19119 12257
rect 19610 12248 19616 12260
rect 19668 12248 19674 12300
rect 19245 12223 19303 12229
rect 19245 12189 19257 12223
rect 19291 12220 19303 12223
rect 19334 12220 19340 12232
rect 19291 12192 19340 12220
rect 19291 12189 19303 12192
rect 19245 12183 19303 12189
rect 19334 12180 19340 12192
rect 19392 12180 19398 12232
rect 20073 12223 20131 12229
rect 20073 12189 20085 12223
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 18601 12155 18659 12161
rect 18601 12121 18613 12155
rect 18647 12152 18659 12155
rect 20088 12152 20116 12183
rect 20162 12180 20168 12232
rect 20220 12220 20226 12232
rect 20220 12192 20265 12220
rect 20220 12180 20226 12192
rect 18647 12124 20116 12152
rect 18647 12121 18659 12124
rect 18601 12115 18659 12121
rect 16448 12056 17540 12084
rect 16448 12044 16454 12056
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 1394 11840 1400 11892
rect 1452 11880 1458 11892
rect 1765 11883 1823 11889
rect 1765 11880 1777 11883
rect 1452 11852 1777 11880
rect 1452 11840 1458 11852
rect 1765 11849 1777 11852
rect 1811 11849 1823 11883
rect 1765 11843 1823 11849
rect 3602 11840 3608 11892
rect 3660 11880 3666 11892
rect 3789 11883 3847 11889
rect 3789 11880 3801 11883
rect 3660 11852 3801 11880
rect 3660 11840 3666 11852
rect 3789 11849 3801 11852
rect 3835 11849 3847 11883
rect 9214 11880 9220 11892
rect 3789 11843 3847 11849
rect 8005 11852 9220 11880
rect 2314 11772 2320 11824
rect 2372 11812 2378 11824
rect 2372 11784 3372 11812
rect 2372 11772 2378 11784
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11744 2467 11747
rect 2958 11744 2964 11756
rect 2455 11716 2964 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 2958 11704 2964 11716
rect 3016 11704 3022 11756
rect 3344 11753 3372 11784
rect 3418 11772 3424 11824
rect 3476 11812 3482 11824
rect 8005 11812 8033 11852
rect 9214 11840 9220 11852
rect 9272 11840 9278 11892
rect 10137 11883 10195 11889
rect 10137 11849 10149 11883
rect 10183 11880 10195 11883
rect 11790 11880 11796 11892
rect 10183 11852 11796 11880
rect 10183 11849 10195 11852
rect 10137 11843 10195 11849
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 11882 11840 11888 11892
rect 11940 11880 11946 11892
rect 11940 11852 14044 11880
rect 11940 11840 11946 11852
rect 3476 11784 8033 11812
rect 3476 11772 3482 11784
rect 3329 11747 3387 11753
rect 3329 11713 3341 11747
rect 3375 11713 3387 11747
rect 3329 11707 3387 11713
rect 4433 11747 4491 11753
rect 4433 11713 4445 11747
rect 4479 11744 4491 11747
rect 5258 11744 5264 11756
rect 4479 11716 5264 11744
rect 4479 11713 4491 11716
rect 4433 11707 4491 11713
rect 5258 11704 5264 11716
rect 5316 11704 5322 11756
rect 5442 11744 5448 11756
rect 5403 11716 5448 11744
rect 5442 11704 5448 11716
rect 5500 11704 5506 11756
rect 7944 11753 7972 11784
rect 9306 11772 9312 11824
rect 9364 11812 9370 11824
rect 14016 11812 14044 11852
rect 15102 11840 15108 11892
rect 15160 11880 15166 11892
rect 15562 11880 15568 11892
rect 15160 11852 15568 11880
rect 15160 11840 15166 11852
rect 15562 11840 15568 11852
rect 15620 11840 15626 11892
rect 15746 11880 15752 11892
rect 15707 11852 15752 11880
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 16390 11880 16396 11892
rect 16132 11852 16396 11880
rect 15654 11812 15660 11824
rect 9364 11784 11744 11812
rect 14016 11784 15660 11812
rect 9364 11772 9370 11784
rect 7929 11747 7987 11753
rect 7929 11713 7941 11747
rect 7975 11713 7987 11747
rect 7929 11707 7987 11713
rect 9950 11704 9956 11756
rect 10008 11744 10014 11756
rect 10410 11744 10416 11756
rect 10008 11716 10416 11744
rect 10008 11704 10014 11716
rect 10410 11704 10416 11716
rect 10468 11704 10474 11756
rect 10778 11744 10784 11756
rect 10739 11716 10784 11744
rect 10778 11704 10784 11716
rect 10836 11704 10842 11756
rect 10870 11704 10876 11756
rect 10928 11744 10934 11756
rect 11716 11753 11744 11784
rect 15654 11772 15660 11784
rect 15712 11772 15718 11824
rect 11701 11747 11759 11753
rect 10928 11716 11560 11744
rect 10928 11704 10934 11716
rect 3142 11676 3148 11688
rect 3103 11648 3148 11676
rect 3142 11636 3148 11648
rect 3200 11636 3206 11688
rect 7193 11679 7251 11685
rect 7193 11645 7205 11679
rect 7239 11676 7251 11679
rect 8202 11676 8208 11688
rect 7239 11648 8208 11676
rect 7239 11645 7251 11648
rect 7193 11639 7251 11645
rect 8202 11636 8208 11648
rect 8260 11636 8266 11688
rect 8297 11679 8355 11685
rect 8297 11645 8309 11679
rect 8343 11676 8355 11679
rect 8386 11676 8392 11688
rect 8343 11648 8392 11676
rect 8343 11645 8355 11648
rect 8297 11639 8355 11645
rect 8386 11636 8392 11648
rect 8444 11636 8450 11688
rect 8564 11679 8622 11685
rect 8564 11645 8576 11679
rect 8610 11676 8622 11679
rect 8846 11676 8852 11688
rect 8610 11648 8852 11676
rect 8610 11645 8622 11648
rect 8564 11639 8622 11645
rect 8846 11636 8852 11648
rect 8904 11636 8910 11688
rect 9398 11636 9404 11688
rect 9456 11676 9462 11688
rect 10505 11679 10563 11685
rect 10505 11676 10517 11679
rect 9456 11648 10517 11676
rect 9456 11636 9462 11648
rect 10505 11645 10517 11648
rect 10551 11645 10563 11679
rect 10505 11639 10563 11645
rect 10962 11636 10968 11688
rect 11020 11676 11026 11688
rect 11532 11685 11560 11716
rect 11701 11713 11713 11747
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 14458 11704 14464 11756
rect 14516 11744 14522 11756
rect 15289 11747 15347 11753
rect 15289 11744 15301 11747
rect 14516 11716 15301 11744
rect 14516 11704 14522 11716
rect 15289 11713 15301 11716
rect 15335 11713 15347 11747
rect 15289 11707 15347 11713
rect 15562 11704 15568 11756
rect 15620 11744 15626 11756
rect 16132 11744 16160 11852
rect 16390 11840 16396 11852
rect 16448 11840 16454 11892
rect 17034 11840 17040 11892
rect 17092 11880 17098 11892
rect 17497 11883 17555 11889
rect 17497 11880 17509 11883
rect 17092 11852 17509 11880
rect 17092 11840 17098 11852
rect 17497 11849 17509 11852
rect 17543 11849 17555 11883
rect 17497 11843 17555 11849
rect 18141 11883 18199 11889
rect 18141 11849 18153 11883
rect 18187 11880 18199 11883
rect 19242 11880 19248 11892
rect 18187 11852 19248 11880
rect 18187 11849 18199 11852
rect 18141 11843 18199 11849
rect 19242 11840 19248 11852
rect 19300 11840 19306 11892
rect 17770 11772 17776 11824
rect 17828 11812 17834 11824
rect 20257 11815 20315 11821
rect 20257 11812 20269 11815
rect 17828 11784 20269 11812
rect 17828 11772 17834 11784
rect 20257 11781 20269 11784
rect 20303 11781 20315 11815
rect 20257 11775 20315 11781
rect 15620 11716 16160 11744
rect 18785 11747 18843 11753
rect 15620 11704 15626 11716
rect 18785 11713 18797 11747
rect 18831 11744 18843 11747
rect 18966 11744 18972 11756
rect 18831 11716 18972 11744
rect 18831 11713 18843 11716
rect 18785 11707 18843 11713
rect 18966 11704 18972 11716
rect 19024 11704 19030 11756
rect 19978 11744 19984 11756
rect 19939 11716 19984 11744
rect 19978 11704 19984 11716
rect 20036 11704 20042 11756
rect 20346 11704 20352 11756
rect 20404 11744 20410 11756
rect 20717 11747 20775 11753
rect 20717 11744 20729 11747
rect 20404 11716 20729 11744
rect 20404 11704 20410 11716
rect 20717 11713 20729 11716
rect 20763 11713 20775 11747
rect 20717 11707 20775 11713
rect 11517 11679 11575 11685
rect 11020 11648 11284 11676
rect 11020 11636 11026 11648
rect 3237 11611 3295 11617
rect 3237 11577 3249 11611
rect 3283 11608 3295 11611
rect 7745 11611 7803 11617
rect 3283 11580 7328 11608
rect 3283 11577 3295 11580
rect 3237 11571 3295 11577
rect 2130 11540 2136 11552
rect 2091 11512 2136 11540
rect 2130 11500 2136 11512
rect 2188 11500 2194 11552
rect 2225 11543 2283 11549
rect 2225 11509 2237 11543
rect 2271 11540 2283 11543
rect 2777 11543 2835 11549
rect 2777 11540 2789 11543
rect 2271 11512 2789 11540
rect 2271 11509 2283 11512
rect 2225 11503 2283 11509
rect 2777 11509 2789 11512
rect 2823 11509 2835 11543
rect 2777 11503 2835 11509
rect 3970 11500 3976 11552
rect 4028 11540 4034 11552
rect 4157 11543 4215 11549
rect 4157 11540 4169 11543
rect 4028 11512 4169 11540
rect 4028 11500 4034 11512
rect 4157 11509 4169 11512
rect 4203 11509 4215 11543
rect 4157 11503 4215 11509
rect 4249 11543 4307 11549
rect 4249 11509 4261 11543
rect 4295 11540 4307 11543
rect 4801 11543 4859 11549
rect 4801 11540 4813 11543
rect 4295 11512 4813 11540
rect 4295 11509 4307 11512
rect 4249 11503 4307 11509
rect 4801 11509 4813 11512
rect 4847 11509 4859 11543
rect 5166 11540 5172 11552
rect 5127 11512 5172 11540
rect 4801 11503 4859 11509
rect 5166 11500 5172 11512
rect 5224 11500 5230 11552
rect 5261 11543 5319 11549
rect 5261 11509 5273 11543
rect 5307 11540 5319 11543
rect 6730 11540 6736 11552
rect 5307 11512 6736 11540
rect 5307 11509 5319 11512
rect 5261 11503 5319 11509
rect 6730 11500 6736 11512
rect 6788 11500 6794 11552
rect 7006 11540 7012 11552
rect 6967 11512 7012 11540
rect 7006 11500 7012 11512
rect 7064 11500 7070 11552
rect 7300 11549 7328 11580
rect 7745 11577 7757 11611
rect 7791 11608 7803 11611
rect 11256 11608 11284 11648
rect 11517 11645 11529 11679
rect 11563 11645 11575 11679
rect 11517 11639 11575 11645
rect 13081 11679 13139 11685
rect 13081 11645 13093 11679
rect 13127 11645 13139 11679
rect 13081 11639 13139 11645
rect 13348 11679 13406 11685
rect 13348 11645 13360 11679
rect 13394 11676 13406 11679
rect 13630 11676 13636 11688
rect 13394 11648 13636 11676
rect 13394 11645 13406 11648
rect 13348 11639 13406 11645
rect 11609 11611 11667 11617
rect 11609 11608 11621 11611
rect 7791 11580 11192 11608
rect 11256 11580 11621 11608
rect 7791 11577 7803 11580
rect 7745 11571 7803 11577
rect 7285 11543 7343 11549
rect 7285 11509 7297 11543
rect 7331 11509 7343 11543
rect 7285 11503 7343 11509
rect 7653 11543 7711 11549
rect 7653 11509 7665 11543
rect 7699 11540 7711 11543
rect 9582 11540 9588 11552
rect 7699 11512 9588 11540
rect 7699 11509 7711 11512
rect 7653 11503 7711 11509
rect 9582 11500 9588 11512
rect 9640 11500 9646 11552
rect 9677 11543 9735 11549
rect 9677 11509 9689 11543
rect 9723 11540 9735 11543
rect 9766 11540 9772 11552
rect 9723 11512 9772 11540
rect 9723 11509 9735 11512
rect 9677 11503 9735 11509
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 9950 11500 9956 11552
rect 10008 11540 10014 11552
rect 11164 11549 11192 11580
rect 11609 11577 11621 11580
rect 11655 11577 11667 11611
rect 11609 11571 11667 11577
rect 11882 11568 11888 11620
rect 11940 11608 11946 11620
rect 12342 11608 12348 11620
rect 11940 11580 12348 11608
rect 11940 11568 11946 11580
rect 12342 11568 12348 11580
rect 12400 11608 12406 11620
rect 13096 11608 13124 11639
rect 13630 11636 13636 11648
rect 13688 11636 13694 11688
rect 13906 11636 13912 11688
rect 13964 11676 13970 11688
rect 15105 11679 15163 11685
rect 13964 11648 14228 11676
rect 13964 11636 13970 11648
rect 12400 11580 13124 11608
rect 14200 11608 14228 11648
rect 15105 11645 15117 11679
rect 15151 11676 15163 11679
rect 15151 11648 15332 11676
rect 15151 11645 15163 11648
rect 15105 11639 15163 11645
rect 14200 11580 14780 11608
rect 12400 11568 12406 11580
rect 10597 11543 10655 11549
rect 10597 11540 10609 11543
rect 10008 11512 10609 11540
rect 10008 11500 10014 11512
rect 10597 11509 10609 11512
rect 10643 11509 10655 11543
rect 10597 11503 10655 11509
rect 11149 11543 11207 11549
rect 11149 11509 11161 11543
rect 11195 11509 11207 11543
rect 11149 11503 11207 11509
rect 11698 11500 11704 11552
rect 11756 11540 11762 11552
rect 13906 11540 13912 11552
rect 11756 11512 13912 11540
rect 11756 11500 11762 11512
rect 13906 11500 13912 11512
rect 13964 11540 13970 11552
rect 14752 11549 14780 11580
rect 15010 11568 15016 11620
rect 15068 11608 15074 11620
rect 15197 11611 15255 11617
rect 15197 11608 15209 11611
rect 15068 11580 15209 11608
rect 15068 11568 15074 11580
rect 15197 11577 15209 11580
rect 15243 11577 15255 11611
rect 15304 11608 15332 11648
rect 15378 11636 15384 11688
rect 15436 11676 15442 11688
rect 15933 11679 15991 11685
rect 15933 11676 15945 11679
rect 15436 11648 15945 11676
rect 15436 11636 15442 11648
rect 15933 11645 15945 11648
rect 15979 11645 15991 11679
rect 16114 11676 16120 11688
rect 16075 11648 16120 11676
rect 15933 11639 15991 11645
rect 16114 11636 16120 11648
rect 16172 11636 16178 11688
rect 16758 11636 16764 11688
rect 16816 11676 16822 11688
rect 20441 11679 20499 11685
rect 20441 11676 20453 11679
rect 16816 11648 20453 11676
rect 16816 11636 16822 11648
rect 20441 11645 20453 11648
rect 20487 11645 20499 11679
rect 20441 11639 20499 11645
rect 15838 11608 15844 11620
rect 15304 11580 15844 11608
rect 15197 11571 15255 11577
rect 15838 11568 15844 11580
rect 15896 11568 15902 11620
rect 14461 11543 14519 11549
rect 14461 11540 14473 11543
rect 13964 11512 14473 11540
rect 13964 11500 13970 11512
rect 14461 11509 14473 11512
rect 14507 11509 14519 11543
rect 14461 11503 14519 11509
rect 14737 11543 14795 11549
rect 14737 11509 14749 11543
rect 14783 11509 14795 11543
rect 14737 11503 14795 11509
rect 15286 11500 15292 11552
rect 15344 11540 15350 11552
rect 16132 11540 16160 11636
rect 16384 11611 16442 11617
rect 16384 11577 16396 11611
rect 16430 11608 16442 11611
rect 16482 11608 16488 11620
rect 16430 11580 16488 11608
rect 16430 11577 16442 11580
rect 16384 11571 16442 11577
rect 16482 11568 16488 11580
rect 16540 11568 16546 11620
rect 18509 11611 18567 11617
rect 18509 11577 18521 11611
rect 18555 11608 18567 11611
rect 19518 11608 19524 11620
rect 18555 11580 19524 11608
rect 18555 11577 18567 11580
rect 18509 11571 18567 11577
rect 19518 11568 19524 11580
rect 19576 11568 19582 11620
rect 19610 11568 19616 11620
rect 19668 11608 19674 11620
rect 19797 11611 19855 11617
rect 19797 11608 19809 11611
rect 19668 11580 19809 11608
rect 19668 11568 19674 11580
rect 19797 11577 19809 11580
rect 19843 11608 19855 11611
rect 20162 11608 20168 11620
rect 19843 11580 20168 11608
rect 19843 11577 19855 11580
rect 19797 11571 19855 11577
rect 20162 11568 20168 11580
rect 20220 11568 20226 11620
rect 18598 11540 18604 11552
rect 15344 11512 16160 11540
rect 18559 11512 18604 11540
rect 15344 11500 15350 11512
rect 18598 11500 18604 11512
rect 18656 11500 18662 11552
rect 18782 11500 18788 11552
rect 18840 11540 18846 11552
rect 19429 11543 19487 11549
rect 19429 11540 19441 11543
rect 18840 11512 19441 11540
rect 18840 11500 18846 11512
rect 19429 11509 19441 11512
rect 19475 11509 19487 11543
rect 19429 11503 19487 11509
rect 19889 11543 19947 11549
rect 19889 11509 19901 11543
rect 19935 11540 19947 11543
rect 20257 11543 20315 11549
rect 20257 11540 20269 11543
rect 19935 11512 20269 11540
rect 19935 11509 19947 11512
rect 19889 11503 19947 11509
rect 20257 11509 20269 11512
rect 20303 11509 20315 11543
rect 20257 11503 20315 11509
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 2314 11296 2320 11348
rect 2372 11336 2378 11348
rect 2869 11339 2927 11345
rect 2869 11336 2881 11339
rect 2372 11308 2881 11336
rect 2372 11296 2378 11308
rect 2869 11305 2881 11308
rect 2915 11305 2927 11339
rect 2869 11299 2927 11305
rect 5166 11296 5172 11348
rect 5224 11336 5230 11348
rect 5721 11339 5779 11345
rect 5721 11336 5733 11339
rect 5224 11308 5733 11336
rect 5224 11296 5230 11308
rect 5721 11305 5733 11308
rect 5767 11305 5779 11339
rect 5721 11299 5779 11305
rect 5994 11296 6000 11348
rect 6052 11336 6058 11348
rect 6181 11339 6239 11345
rect 6181 11336 6193 11339
rect 6052 11308 6193 11336
rect 6052 11296 6058 11308
rect 6181 11305 6193 11308
rect 6227 11305 6239 11339
rect 6730 11336 6736 11348
rect 6691 11308 6736 11336
rect 6181 11299 6239 11305
rect 6730 11296 6736 11308
rect 6788 11296 6794 11348
rect 8573 11339 8631 11345
rect 7116 11308 8524 11336
rect 6362 11228 6368 11280
rect 6420 11268 6426 11280
rect 7116 11268 7144 11308
rect 6420 11240 7144 11268
rect 7193 11271 7251 11277
rect 6420 11228 6426 11240
rect 7193 11237 7205 11271
rect 7239 11268 7251 11271
rect 7239 11240 8432 11268
rect 7239 11237 7251 11240
rect 7193 11231 7251 11237
rect 1486 11200 1492 11212
rect 1447 11172 1492 11200
rect 1486 11160 1492 11172
rect 1544 11160 1550 11212
rect 1756 11203 1814 11209
rect 1756 11169 1768 11203
rect 1802 11200 1814 11203
rect 2590 11200 2596 11212
rect 1802 11172 2596 11200
rect 1802 11169 1814 11172
rect 1756 11163 1814 11169
rect 2590 11160 2596 11172
rect 2648 11160 2654 11212
rect 4062 11200 4068 11212
rect 4023 11172 4068 11200
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 4332 11203 4390 11209
rect 4332 11169 4344 11203
rect 4378 11200 4390 11203
rect 6086 11200 6092 11212
rect 4378 11172 5580 11200
rect 6047 11172 6092 11200
rect 4378 11169 4390 11172
rect 4332 11163 4390 11169
rect 5092 11144 5120 11172
rect 3142 11132 3148 11144
rect 3103 11104 3148 11132
rect 3142 11092 3148 11104
rect 3200 11092 3206 11144
rect 5074 11092 5080 11144
rect 5132 11092 5138 11144
rect 5552 11132 5580 11172
rect 6086 11160 6092 11172
rect 6144 11160 6150 11212
rect 7101 11203 7159 11209
rect 7101 11169 7113 11203
rect 7147 11200 7159 11203
rect 8294 11200 8300 11212
rect 7147 11172 8300 11200
rect 7147 11169 7159 11172
rect 7101 11163 7159 11169
rect 8294 11160 8300 11172
rect 8352 11160 8358 11212
rect 6365 11135 6423 11141
rect 6365 11132 6377 11135
rect 5552 11104 6377 11132
rect 6365 11101 6377 11104
rect 6411 11132 6423 11135
rect 6914 11132 6920 11144
rect 6411 11104 6920 11132
rect 6411 11101 6423 11104
rect 6365 11095 6423 11101
rect 6914 11092 6920 11104
rect 6972 11132 6978 11144
rect 7285 11135 7343 11141
rect 7285 11132 7297 11135
rect 6972 11104 7297 11132
rect 6972 11092 6978 11104
rect 7285 11101 7297 11104
rect 7331 11101 7343 11135
rect 7285 11095 7343 11101
rect 5442 11064 5448 11076
rect 5403 11036 5448 11064
rect 5442 11024 5448 11036
rect 5500 11024 5506 11076
rect 8404 11064 8432 11240
rect 8496 11200 8524 11308
rect 8573 11305 8585 11339
rect 8619 11305 8631 11339
rect 8573 11299 8631 11305
rect 8941 11339 8999 11345
rect 8941 11305 8953 11339
rect 8987 11336 8999 11339
rect 9398 11336 9404 11348
rect 8987 11308 9404 11336
rect 8987 11305 8999 11308
rect 8941 11299 8999 11305
rect 8588 11268 8616 11299
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 10413 11339 10471 11345
rect 10413 11305 10425 11339
rect 10459 11336 10471 11339
rect 12713 11339 12771 11345
rect 10459 11308 11928 11336
rect 10459 11305 10471 11308
rect 10413 11299 10471 11305
rect 9214 11268 9220 11280
rect 8588 11240 9220 11268
rect 9214 11228 9220 11240
rect 9272 11228 9278 11280
rect 9582 11228 9588 11280
rect 9640 11268 9646 11280
rect 11900 11268 11928 11308
rect 12713 11305 12725 11339
rect 12759 11336 12771 11339
rect 13357 11339 13415 11345
rect 13357 11336 13369 11339
rect 12759 11308 13369 11336
rect 12759 11305 12771 11308
rect 12713 11299 12771 11305
rect 13357 11305 13369 11308
rect 13403 11305 13415 11339
rect 13357 11299 13415 11305
rect 13725 11339 13783 11345
rect 13725 11305 13737 11339
rect 13771 11336 13783 11339
rect 16022 11336 16028 11348
rect 13771 11308 16028 11336
rect 13771 11305 13783 11308
rect 13725 11299 13783 11305
rect 16022 11296 16028 11308
rect 16080 11296 16086 11348
rect 17310 11296 17316 11348
rect 17368 11336 17374 11348
rect 17405 11339 17463 11345
rect 17405 11336 17417 11339
rect 17368 11308 17417 11336
rect 17368 11296 17374 11308
rect 17405 11305 17417 11308
rect 17451 11305 17463 11339
rect 17405 11299 17463 11305
rect 17954 11296 17960 11348
rect 18012 11336 18018 11348
rect 18417 11339 18475 11345
rect 18417 11336 18429 11339
rect 18012 11308 18429 11336
rect 18012 11296 18018 11308
rect 18417 11305 18429 11308
rect 18463 11305 18475 11339
rect 18782 11336 18788 11348
rect 18743 11308 18788 11336
rect 18417 11299 18475 11305
rect 18782 11296 18788 11308
rect 18840 11296 18846 11348
rect 18877 11339 18935 11345
rect 18877 11305 18889 11339
rect 18923 11336 18935 11339
rect 19245 11339 19303 11345
rect 19245 11336 19257 11339
rect 18923 11308 19257 11336
rect 18923 11305 18935 11308
rect 18877 11299 18935 11305
rect 19245 11305 19257 11308
rect 19291 11305 19303 11339
rect 19245 11299 19303 11305
rect 19889 11339 19947 11345
rect 19889 11305 19901 11339
rect 19935 11336 19947 11339
rect 20070 11336 20076 11348
rect 19935 11308 20076 11336
rect 19935 11305 19947 11308
rect 19889 11299 19947 11305
rect 20070 11296 20076 11308
rect 20128 11296 20134 11348
rect 12805 11271 12863 11277
rect 12805 11268 12817 11271
rect 9640 11240 11836 11268
rect 11900 11240 12817 11268
rect 9640 11228 9646 11240
rect 9033 11203 9091 11209
rect 9033 11200 9045 11203
rect 8496 11172 9045 11200
rect 9033 11169 9045 11172
rect 9079 11200 9091 11203
rect 9950 11200 9956 11212
rect 9079 11172 9956 11200
rect 9079 11169 9091 11172
rect 9033 11163 9091 11169
rect 9950 11160 9956 11172
rect 10008 11160 10014 11212
rect 10042 11160 10048 11212
rect 10100 11200 10106 11212
rect 10686 11200 10692 11212
rect 10100 11172 10692 11200
rect 10100 11160 10106 11172
rect 10686 11160 10692 11172
rect 10744 11200 10750 11212
rect 10781 11203 10839 11209
rect 10781 11200 10793 11203
rect 10744 11172 10793 11200
rect 10744 11160 10750 11172
rect 10781 11169 10793 11172
rect 10827 11169 10839 11203
rect 10781 11163 10839 11169
rect 9217 11135 9275 11141
rect 9217 11101 9229 11135
rect 9263 11132 9275 11135
rect 9766 11132 9772 11144
rect 9263 11104 9772 11132
rect 9263 11101 9275 11104
rect 9217 11095 9275 11101
rect 9766 11092 9772 11104
rect 9824 11092 9830 11144
rect 10134 11092 10140 11144
rect 10192 11132 10198 11144
rect 10502 11132 10508 11144
rect 10192 11104 10508 11132
rect 10192 11092 10198 11104
rect 10502 11092 10508 11104
rect 10560 11132 10566 11144
rect 10873 11135 10931 11141
rect 10873 11132 10885 11135
rect 10560 11104 10885 11132
rect 10560 11092 10566 11104
rect 10873 11101 10885 11104
rect 10919 11101 10931 11135
rect 10873 11095 10931 11101
rect 10962 11092 10968 11144
rect 11020 11132 11026 11144
rect 11698 11132 11704 11144
rect 11020 11104 11704 11132
rect 11020 11092 11026 11104
rect 11698 11092 11704 11104
rect 11756 11092 11762 11144
rect 11808 11132 11836 11240
rect 12805 11237 12817 11240
rect 12851 11237 12863 11271
rect 12805 11231 12863 11237
rect 12986 11228 12992 11280
rect 13044 11268 13050 11280
rect 14090 11268 14096 11280
rect 13044 11240 14096 11268
rect 13044 11228 13050 11240
rect 14090 11228 14096 11240
rect 14148 11268 14154 11280
rect 19058 11268 19064 11280
rect 14148 11240 14596 11268
rect 14148 11228 14154 11240
rect 14568 11209 14596 11240
rect 17604 11240 19064 11268
rect 12253 11203 12311 11209
rect 12253 11169 12265 11203
rect 12299 11200 12311 11203
rect 14553 11203 14611 11209
rect 12299 11172 14320 11200
rect 12299 11169 12311 11172
rect 12253 11163 12311 11169
rect 12710 11132 12716 11144
rect 11808 11104 12716 11132
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 12986 11132 12992 11144
rect 12947 11104 12992 11132
rect 12986 11092 12992 11104
rect 13044 11092 13050 11144
rect 13262 11092 13268 11144
rect 13320 11132 13326 11144
rect 13722 11132 13728 11144
rect 13320 11104 13728 11132
rect 13320 11092 13326 11104
rect 13722 11092 13728 11104
rect 13780 11132 13786 11144
rect 13817 11135 13875 11141
rect 13817 11132 13829 11135
rect 13780 11104 13829 11132
rect 13780 11092 13786 11104
rect 13817 11101 13829 11104
rect 13863 11101 13875 11135
rect 13817 11095 13875 11101
rect 13906 11092 13912 11144
rect 13964 11132 13970 11144
rect 14182 11132 14188 11144
rect 13964 11104 14188 11132
rect 13964 11092 13970 11104
rect 14182 11092 14188 11104
rect 14240 11092 14246 11144
rect 9674 11064 9680 11076
rect 8404 11036 9680 11064
rect 9674 11024 9680 11036
rect 9732 11024 9738 11076
rect 12345 11067 12403 11073
rect 12345 11033 12357 11067
rect 12391 11064 12403 11067
rect 12618 11064 12624 11076
rect 12391 11036 12624 11064
rect 12391 11033 12403 11036
rect 12345 11027 12403 11033
rect 12618 11024 12624 11036
rect 12676 11024 12682 11076
rect 14292 11064 14320 11172
rect 14553 11169 14565 11203
rect 14599 11169 14611 11203
rect 15286 11200 15292 11212
rect 15247 11172 15292 11200
rect 14553 11163 14611 11169
rect 15286 11160 15292 11172
rect 15344 11160 15350 11212
rect 15378 11160 15384 11212
rect 15436 11200 15442 11212
rect 15545 11203 15603 11209
rect 15545 11200 15557 11203
rect 15436 11172 15557 11200
rect 15436 11160 15442 11172
rect 15545 11169 15557 11172
rect 15591 11200 15603 11203
rect 17313 11203 17371 11209
rect 15591 11172 17080 11200
rect 15591 11169 15603 11172
rect 15545 11163 15603 11169
rect 17052 11132 17080 11172
rect 17313 11169 17325 11203
rect 17359 11200 17371 11203
rect 17604 11200 17632 11240
rect 19058 11228 19064 11240
rect 19116 11228 19122 11280
rect 19797 11271 19855 11277
rect 19797 11237 19809 11271
rect 19843 11268 19855 11271
rect 20898 11268 20904 11280
rect 19843 11240 20904 11268
rect 19843 11237 19855 11240
rect 19797 11231 19855 11237
rect 20898 11228 20904 11240
rect 20956 11228 20962 11280
rect 17359 11172 17632 11200
rect 17696 11172 19012 11200
rect 17359 11169 17371 11172
rect 17313 11163 17371 11169
rect 17494 11132 17500 11144
rect 17052 11104 17500 11132
rect 17494 11092 17500 11104
rect 17552 11092 17558 11144
rect 14369 11067 14427 11073
rect 14369 11064 14381 11067
rect 14292 11036 14381 11064
rect 14369 11033 14381 11036
rect 14415 11064 14427 11067
rect 15102 11064 15108 11076
rect 14415 11036 15108 11064
rect 14415 11033 14427 11036
rect 14369 11027 14427 11033
rect 15102 11024 15108 11036
rect 15160 11024 15166 11076
rect 16482 11024 16488 11076
rect 16540 11064 16546 11076
rect 16669 11067 16727 11073
rect 16669 11064 16681 11067
rect 16540 11036 16681 11064
rect 16540 11024 16546 11036
rect 16669 11033 16681 11036
rect 16715 11064 16727 11067
rect 17696 11064 17724 11172
rect 18984 11144 19012 11172
rect 17954 11132 17960 11144
rect 17915 11104 17960 11132
rect 17954 11092 17960 11104
rect 18012 11092 18018 11144
rect 18966 11132 18972 11144
rect 18927 11104 18972 11132
rect 18966 11092 18972 11104
rect 19024 11092 19030 11144
rect 19978 11132 19984 11144
rect 19939 11104 19984 11132
rect 19978 11092 19984 11104
rect 20036 11092 20042 11144
rect 16715 11036 17724 11064
rect 16715 11033 16727 11036
rect 16669 11027 16727 11033
rect 18690 11024 18696 11076
rect 18748 11064 18754 11076
rect 19429 11067 19487 11073
rect 19429 11064 19441 11067
rect 18748 11036 19441 11064
rect 18748 11024 18754 11036
rect 19429 11033 19441 11036
rect 19475 11033 19487 11067
rect 19429 11027 19487 11033
rect 3234 10956 3240 11008
rect 3292 10996 3298 11008
rect 10226 10996 10232 11008
rect 3292 10968 10232 10996
rect 3292 10956 3298 10968
rect 10226 10956 10232 10968
rect 10284 10956 10290 11008
rect 11882 10956 11888 11008
rect 11940 10996 11946 11008
rect 12069 10999 12127 11005
rect 12069 10996 12081 10999
rect 11940 10968 12081 10996
rect 11940 10956 11946 10968
rect 12069 10965 12081 10968
rect 12115 10965 12127 10999
rect 12069 10959 12127 10965
rect 12526 10956 12532 11008
rect 12584 10996 12590 11008
rect 16758 10996 16764 11008
rect 12584 10968 16764 10996
rect 12584 10956 12590 10968
rect 16758 10956 16764 10968
rect 16816 10956 16822 11008
rect 16942 10996 16948 11008
rect 16903 10968 16948 10996
rect 16942 10956 16948 10968
rect 17000 10956 17006 11008
rect 18874 10956 18880 11008
rect 18932 10996 18938 11008
rect 19245 10999 19303 11005
rect 19245 10996 19257 10999
rect 18932 10968 19257 10996
rect 18932 10956 18938 10968
rect 19245 10965 19257 10968
rect 19291 10965 19303 10999
rect 19245 10959 19303 10965
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 1765 10795 1823 10801
rect 1765 10761 1777 10795
rect 1811 10792 1823 10795
rect 2130 10792 2136 10804
rect 1811 10764 2136 10792
rect 1811 10761 1823 10764
rect 1765 10755 1823 10761
rect 2130 10752 2136 10764
rect 2188 10752 2194 10804
rect 3970 10792 3976 10804
rect 3931 10764 3976 10792
rect 3970 10752 3976 10764
rect 4028 10752 4034 10804
rect 4706 10752 4712 10804
rect 4764 10792 4770 10804
rect 4893 10795 4951 10801
rect 4893 10792 4905 10795
rect 4764 10764 4905 10792
rect 4764 10752 4770 10764
rect 4893 10761 4905 10764
rect 4939 10792 4951 10795
rect 4982 10792 4988 10804
rect 4939 10764 4988 10792
rect 4939 10761 4951 10764
rect 4893 10755 4951 10761
rect 4982 10752 4988 10764
rect 5040 10752 5046 10804
rect 7006 10752 7012 10804
rect 7064 10792 7070 10804
rect 8389 10795 8447 10801
rect 8389 10792 8401 10795
rect 7064 10764 8401 10792
rect 7064 10752 7070 10764
rect 8389 10761 8401 10764
rect 8435 10761 8447 10795
rect 12158 10792 12164 10804
rect 8389 10755 8447 10761
rect 8496 10764 12164 10792
rect 3418 10684 3424 10736
rect 3476 10684 3482 10736
rect 4062 10684 4068 10736
rect 4120 10724 4126 10736
rect 8496 10724 8524 10764
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 12437 10795 12495 10801
rect 12437 10761 12449 10795
rect 12483 10792 12495 10795
rect 12526 10792 12532 10804
rect 12483 10764 12532 10792
rect 12483 10761 12495 10764
rect 12437 10755 12495 10761
rect 12526 10752 12532 10764
rect 12584 10752 12590 10804
rect 14921 10795 14979 10801
rect 14921 10761 14933 10795
rect 14967 10792 14979 10795
rect 15010 10792 15016 10804
rect 14967 10764 15016 10792
rect 14967 10761 14979 10764
rect 14921 10755 14979 10761
rect 15010 10752 15016 10764
rect 15068 10752 15074 10804
rect 16117 10795 16175 10801
rect 16117 10761 16129 10795
rect 16163 10792 16175 10795
rect 18509 10795 18567 10801
rect 16163 10764 18000 10792
rect 16163 10761 16175 10764
rect 16117 10755 16175 10761
rect 4120 10696 8524 10724
rect 4120 10684 4126 10696
rect 11790 10684 11796 10736
rect 11848 10724 11854 10736
rect 11848 10696 15608 10724
rect 11848 10684 11854 10696
rect 2314 10656 2320 10668
rect 2275 10628 2320 10656
rect 2314 10616 2320 10628
rect 2372 10616 2378 10668
rect 2590 10616 2596 10668
rect 2648 10656 2654 10668
rect 3329 10659 3387 10665
rect 3329 10656 3341 10659
rect 2648 10628 3341 10656
rect 2648 10616 2654 10628
rect 3329 10625 3341 10628
rect 3375 10656 3387 10659
rect 3436 10656 3464 10684
rect 3375 10628 3464 10656
rect 3375 10625 3387 10628
rect 3329 10619 3387 10625
rect 3510 10616 3516 10668
rect 3568 10656 3574 10668
rect 3970 10656 3976 10668
rect 3568 10628 3976 10656
rect 3568 10616 3574 10628
rect 3970 10616 3976 10628
rect 4028 10616 4034 10668
rect 4617 10659 4675 10665
rect 4617 10625 4629 10659
rect 4663 10656 4675 10659
rect 5442 10656 5448 10668
rect 4663 10628 5448 10656
rect 4663 10625 4675 10628
rect 4617 10619 4675 10625
rect 5442 10616 5448 10628
rect 5500 10616 5506 10668
rect 5626 10656 5632 10668
rect 5587 10628 5632 10656
rect 5626 10616 5632 10628
rect 5684 10616 5690 10668
rect 7098 10616 7104 10668
rect 7156 10656 7162 10668
rect 7466 10656 7472 10668
rect 7156 10628 7472 10656
rect 7156 10616 7162 10628
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 7742 10616 7748 10668
rect 7800 10656 7806 10668
rect 7929 10659 7987 10665
rect 7929 10656 7941 10659
rect 7800 10628 7941 10656
rect 7800 10616 7806 10628
rect 7929 10625 7941 10628
rect 7975 10625 7987 10659
rect 7929 10619 7987 10625
rect 8113 10659 8171 10665
rect 8113 10625 8125 10659
rect 8159 10656 8171 10659
rect 8202 10656 8208 10668
rect 8159 10628 8208 10656
rect 8159 10625 8171 10628
rect 8113 10619 8171 10625
rect 8202 10616 8208 10628
rect 8260 10616 8266 10668
rect 9214 10656 9220 10668
rect 9175 10628 9220 10656
rect 9214 10616 9220 10628
rect 9272 10616 9278 10668
rect 9306 10616 9312 10668
rect 9364 10656 9370 10668
rect 9364 10628 9409 10656
rect 9364 10616 9370 10628
rect 12618 10616 12624 10668
rect 12676 10656 12682 10668
rect 12897 10659 12955 10665
rect 12897 10656 12909 10659
rect 12676 10628 12909 10656
rect 12676 10616 12682 10628
rect 12897 10625 12909 10628
rect 12943 10625 12955 10659
rect 12897 10619 12955 10625
rect 12989 10659 13047 10665
rect 12989 10625 13001 10659
rect 13035 10625 13047 10659
rect 12989 10619 13047 10625
rect 3142 10588 3148 10600
rect 3103 10560 3148 10588
rect 3142 10548 3148 10560
rect 3200 10548 3206 10600
rect 3418 10548 3424 10600
rect 3476 10588 3482 10600
rect 10962 10597 10968 10600
rect 8389 10591 8447 10597
rect 3476 10560 7972 10588
rect 3476 10548 3482 10560
rect 2133 10523 2191 10529
rect 2133 10489 2145 10523
rect 2179 10520 2191 10523
rect 4433 10523 4491 10529
rect 4433 10520 4445 10523
rect 2179 10492 2820 10520
rect 2179 10489 2191 10492
rect 2133 10483 2191 10489
rect 1946 10412 1952 10464
rect 2004 10452 2010 10464
rect 2792 10461 2820 10492
rect 3160 10492 4445 10520
rect 3160 10464 3188 10492
rect 4433 10489 4445 10492
rect 4479 10489 4491 10523
rect 4433 10483 4491 10489
rect 4893 10523 4951 10529
rect 4893 10489 4905 10523
rect 4939 10520 4951 10523
rect 5445 10523 5503 10529
rect 5445 10520 5457 10523
rect 4939 10492 5457 10520
rect 4939 10489 4951 10492
rect 4893 10483 4951 10489
rect 5445 10489 5457 10492
rect 5491 10489 5503 10523
rect 7944 10520 7972 10560
rect 8389 10557 8401 10591
rect 8435 10588 8447 10591
rect 8665 10591 8723 10597
rect 8665 10588 8677 10591
rect 8435 10560 8677 10588
rect 8435 10557 8447 10560
rect 8389 10551 8447 10557
rect 8665 10557 8677 10560
rect 8711 10557 8723 10591
rect 8665 10551 8723 10557
rect 10689 10591 10747 10597
rect 10689 10557 10701 10591
rect 10735 10557 10747 10591
rect 10956 10588 10968 10597
rect 10923 10560 10968 10588
rect 10689 10551 10747 10557
rect 10956 10551 10968 10560
rect 10704 10520 10732 10551
rect 10962 10548 10968 10551
rect 11020 10548 11026 10600
rect 12342 10548 12348 10600
rect 12400 10588 12406 10600
rect 13004 10588 13032 10619
rect 13078 10616 13084 10668
rect 13136 10656 13142 10668
rect 14001 10659 14059 10665
rect 14001 10656 14013 10659
rect 13136 10628 14013 10656
rect 13136 10616 13142 10628
rect 14001 10625 14013 10628
rect 14047 10625 14059 10659
rect 15470 10656 15476 10668
rect 15431 10628 15476 10656
rect 14001 10619 14059 10625
rect 15470 10616 15476 10628
rect 15528 10616 15534 10668
rect 15580 10656 15608 10696
rect 16482 10684 16488 10736
rect 16540 10724 16546 10736
rect 17972 10724 18000 10764
rect 18509 10761 18521 10795
rect 18555 10792 18567 10795
rect 18598 10792 18604 10804
rect 18555 10764 18604 10792
rect 18555 10761 18567 10764
rect 18509 10755 18567 10761
rect 18598 10752 18604 10764
rect 18656 10752 18662 10804
rect 19518 10792 19524 10804
rect 19479 10764 19524 10792
rect 19518 10752 19524 10764
rect 19576 10752 19582 10804
rect 19794 10724 19800 10736
rect 16540 10696 16712 10724
rect 17972 10696 19800 10724
rect 16540 10684 16546 10696
rect 16684 10665 16712 10696
rect 19794 10684 19800 10696
rect 19852 10684 19858 10736
rect 16577 10659 16635 10665
rect 16577 10656 16589 10659
rect 15580 10628 16589 10656
rect 16577 10625 16589 10628
rect 16623 10625 16635 10659
rect 16577 10619 16635 10625
rect 16669 10659 16727 10665
rect 16669 10625 16681 10659
rect 16715 10625 16727 10659
rect 16669 10619 16727 10625
rect 16850 10616 16856 10668
rect 16908 10656 16914 10668
rect 16908 10628 17071 10656
rect 16908 10616 16914 10628
rect 12400 10560 13032 10588
rect 16485 10591 16543 10597
rect 12400 10548 12406 10560
rect 16485 10557 16497 10591
rect 16531 10588 16543 10591
rect 16942 10588 16948 10600
rect 16531 10560 16948 10588
rect 16531 10557 16543 10560
rect 16485 10551 16543 10557
rect 16942 10548 16948 10560
rect 17000 10548 17006 10600
rect 17043 10588 17071 10628
rect 17494 10616 17500 10668
rect 17552 10656 17558 10668
rect 19061 10659 19119 10665
rect 19061 10656 19073 10659
rect 17552 10628 19073 10656
rect 17552 10616 17558 10628
rect 19061 10625 19073 10628
rect 19107 10656 19119 10659
rect 19978 10656 19984 10668
rect 19107 10628 19984 10656
rect 19107 10625 19119 10628
rect 19061 10619 19119 10625
rect 19978 10616 19984 10628
rect 20036 10656 20042 10668
rect 20073 10659 20131 10665
rect 20073 10656 20085 10659
rect 20036 10628 20085 10656
rect 20036 10616 20042 10628
rect 20073 10625 20085 10628
rect 20119 10625 20131 10659
rect 20073 10619 20131 10625
rect 19150 10588 19156 10600
rect 17043 10560 19156 10588
rect 19150 10548 19156 10560
rect 19208 10548 19214 10600
rect 19794 10548 19800 10600
rect 19852 10588 19858 10600
rect 20533 10591 20591 10597
rect 20533 10588 20545 10591
rect 19852 10560 20545 10588
rect 19852 10548 19858 10560
rect 20533 10557 20545 10560
rect 20579 10557 20591 10591
rect 20533 10551 20591 10557
rect 11146 10520 11152 10532
rect 7944 10492 8800 10520
rect 10704 10492 11152 10520
rect 5445 10483 5503 10489
rect 2225 10455 2283 10461
rect 2225 10452 2237 10455
rect 2004 10424 2237 10452
rect 2004 10412 2010 10424
rect 2225 10421 2237 10424
rect 2271 10421 2283 10455
rect 2225 10415 2283 10421
rect 2777 10455 2835 10461
rect 2777 10421 2789 10455
rect 2823 10421 2835 10455
rect 2777 10415 2835 10421
rect 3142 10412 3148 10464
rect 3200 10412 3206 10464
rect 3237 10455 3295 10461
rect 3237 10421 3249 10455
rect 3283 10452 3295 10455
rect 3694 10452 3700 10464
rect 3283 10424 3700 10452
rect 3283 10421 3295 10424
rect 3237 10415 3295 10421
rect 3694 10412 3700 10424
rect 3752 10412 3758 10464
rect 4154 10412 4160 10464
rect 4212 10452 4218 10464
rect 4341 10455 4399 10461
rect 4341 10452 4353 10455
rect 4212 10424 4353 10452
rect 4212 10412 4218 10424
rect 4341 10421 4353 10424
rect 4387 10421 4399 10455
rect 4341 10415 4399 10421
rect 4798 10412 4804 10464
rect 4856 10452 4862 10464
rect 4985 10455 5043 10461
rect 4985 10452 4997 10455
rect 4856 10424 4997 10452
rect 4856 10412 4862 10424
rect 4985 10421 4997 10424
rect 5031 10421 5043 10455
rect 5350 10452 5356 10464
rect 5311 10424 5356 10452
rect 4985 10415 5043 10421
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 5994 10452 6000 10464
rect 5955 10424 6000 10452
rect 5994 10412 6000 10424
rect 6052 10412 6058 10464
rect 7466 10452 7472 10464
rect 7427 10424 7472 10452
rect 7466 10412 7472 10424
rect 7524 10412 7530 10464
rect 7558 10412 7564 10464
rect 7616 10452 7622 10464
rect 7837 10455 7895 10461
rect 7837 10452 7849 10455
rect 7616 10424 7849 10452
rect 7616 10412 7622 10424
rect 7837 10421 7849 10424
rect 7883 10421 7895 10455
rect 8478 10452 8484 10464
rect 8439 10424 8484 10452
rect 7837 10415 7895 10421
rect 8478 10412 8484 10424
rect 8536 10412 8542 10464
rect 8772 10461 8800 10492
rect 11146 10480 11152 10492
rect 11204 10480 11210 10532
rect 12805 10523 12863 10529
rect 12805 10489 12817 10523
rect 12851 10520 12863 10523
rect 12851 10492 13492 10520
rect 12851 10489 12863 10492
rect 12805 10483 12863 10489
rect 8757 10455 8815 10461
rect 8757 10421 8769 10455
rect 8803 10421 8815 10455
rect 9122 10452 9128 10464
rect 9083 10424 9128 10452
rect 8757 10415 8815 10421
rect 9122 10412 9128 10424
rect 9180 10412 9186 10464
rect 11790 10412 11796 10464
rect 11848 10452 11854 10464
rect 12069 10455 12127 10461
rect 12069 10452 12081 10455
rect 11848 10424 12081 10452
rect 11848 10412 11854 10424
rect 12069 10421 12081 10424
rect 12115 10452 12127 10455
rect 12986 10452 12992 10464
rect 12115 10424 12992 10452
rect 12115 10421 12127 10424
rect 12069 10415 12127 10421
rect 12986 10412 12992 10424
rect 13044 10412 13050 10464
rect 13464 10461 13492 10492
rect 13630 10480 13636 10532
rect 13688 10520 13694 10532
rect 15289 10523 15347 10529
rect 15289 10520 15301 10523
rect 13688 10492 15301 10520
rect 13688 10480 13694 10492
rect 15289 10489 15301 10492
rect 15335 10520 15347 10523
rect 16206 10520 16212 10532
rect 15335 10492 16212 10520
rect 15335 10489 15347 10492
rect 15289 10483 15347 10489
rect 16206 10480 16212 10492
rect 16264 10480 16270 10532
rect 18598 10480 18604 10532
rect 18656 10520 18662 10532
rect 18969 10523 19027 10529
rect 18969 10520 18981 10523
rect 18656 10492 18981 10520
rect 18656 10480 18662 10492
rect 18969 10489 18981 10492
rect 19015 10489 19027 10523
rect 18969 10483 19027 10489
rect 19889 10523 19947 10529
rect 19889 10489 19901 10523
rect 19935 10520 19947 10523
rect 20070 10520 20076 10532
rect 19935 10492 20076 10520
rect 19935 10489 19947 10492
rect 19889 10483 19947 10489
rect 20070 10480 20076 10492
rect 20128 10520 20134 10532
rect 20438 10520 20444 10532
rect 20128 10492 20444 10520
rect 20128 10480 20134 10492
rect 20438 10480 20444 10492
rect 20496 10480 20502 10532
rect 20714 10480 20720 10532
rect 20772 10520 20778 10532
rect 20809 10523 20867 10529
rect 20809 10520 20821 10523
rect 20772 10492 20821 10520
rect 20772 10480 20778 10492
rect 20809 10489 20821 10492
rect 20855 10489 20867 10523
rect 20809 10483 20867 10489
rect 13449 10455 13507 10461
rect 13449 10421 13461 10455
rect 13495 10421 13507 10455
rect 13449 10415 13507 10421
rect 13538 10412 13544 10464
rect 13596 10452 13602 10464
rect 13817 10455 13875 10461
rect 13817 10452 13829 10455
rect 13596 10424 13829 10452
rect 13596 10412 13602 10424
rect 13817 10421 13829 10424
rect 13863 10421 13875 10455
rect 13817 10415 13875 10421
rect 13906 10412 13912 10464
rect 13964 10452 13970 10464
rect 15381 10455 15439 10461
rect 13964 10424 14009 10452
rect 13964 10412 13970 10424
rect 15381 10421 15393 10455
rect 15427 10452 15439 10455
rect 18414 10452 18420 10464
rect 15427 10424 18420 10452
rect 15427 10421 15439 10424
rect 15381 10415 15439 10421
rect 18414 10412 18420 10424
rect 18472 10412 18478 10464
rect 18506 10412 18512 10464
rect 18564 10452 18570 10464
rect 18782 10452 18788 10464
rect 18564 10424 18788 10452
rect 18564 10412 18570 10424
rect 18782 10412 18788 10424
rect 18840 10452 18846 10464
rect 18877 10455 18935 10461
rect 18877 10452 18889 10455
rect 18840 10424 18889 10452
rect 18840 10412 18846 10424
rect 18877 10421 18889 10424
rect 18923 10421 18935 10455
rect 18877 10415 18935 10421
rect 19518 10412 19524 10464
rect 19576 10452 19582 10464
rect 19981 10455 20039 10461
rect 19981 10452 19993 10455
rect 19576 10424 19993 10452
rect 19576 10412 19582 10424
rect 19981 10421 19993 10424
rect 20027 10421 20039 10455
rect 19981 10415 20039 10421
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 1946 10248 1952 10260
rect 1907 10220 1952 10248
rect 1946 10208 1952 10220
rect 2004 10208 2010 10260
rect 3418 10248 3424 10260
rect 3379 10220 3424 10248
rect 3418 10208 3424 10220
rect 3476 10208 3482 10260
rect 4154 10248 4160 10260
rect 4115 10220 4160 10248
rect 4154 10208 4160 10220
rect 4212 10208 4218 10260
rect 4525 10251 4583 10257
rect 4525 10217 4537 10251
rect 4571 10248 4583 10251
rect 5994 10248 6000 10260
rect 4571 10220 6000 10248
rect 4571 10217 4583 10220
rect 4525 10211 4583 10217
rect 5994 10208 6000 10220
rect 6052 10208 6058 10260
rect 6914 10248 6920 10260
rect 6875 10220 6920 10248
rect 6914 10208 6920 10220
rect 6972 10208 6978 10260
rect 7282 10208 7288 10260
rect 7340 10248 7346 10260
rect 7742 10248 7748 10260
rect 7340 10220 7748 10248
rect 7340 10208 7346 10220
rect 7742 10208 7748 10220
rect 7800 10208 7806 10260
rect 7837 10251 7895 10257
rect 7837 10217 7849 10251
rect 7883 10248 7895 10251
rect 8478 10248 8484 10260
rect 7883 10220 8484 10248
rect 7883 10217 7895 10220
rect 7837 10211 7895 10217
rect 8478 10208 8484 10220
rect 8536 10248 8542 10260
rect 8662 10248 8668 10260
rect 8536 10220 8668 10248
rect 8536 10208 8542 10220
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 9122 10208 9128 10260
rect 9180 10248 9186 10260
rect 9677 10251 9735 10257
rect 9677 10248 9689 10251
rect 9180 10220 9689 10248
rect 9180 10208 9186 10220
rect 9677 10217 9689 10220
rect 9723 10217 9735 10251
rect 9677 10211 9735 10217
rect 9858 10208 9864 10260
rect 9916 10248 9922 10260
rect 10045 10251 10103 10257
rect 10045 10248 10057 10251
rect 9916 10220 10057 10248
rect 9916 10208 9922 10220
rect 10045 10217 10057 10220
rect 10091 10248 10103 10251
rect 12986 10248 12992 10260
rect 10091 10220 12992 10248
rect 10091 10217 10103 10220
rect 10045 10211 10103 10217
rect 12986 10208 12992 10220
rect 13044 10208 13050 10260
rect 13081 10251 13139 10257
rect 13081 10217 13093 10251
rect 13127 10248 13139 10251
rect 13538 10248 13544 10260
rect 13127 10220 13544 10248
rect 13127 10217 13139 10220
rect 13081 10211 13139 10217
rect 13538 10208 13544 10220
rect 13596 10208 13602 10260
rect 13633 10251 13691 10257
rect 13633 10217 13645 10251
rect 13679 10248 13691 10251
rect 13906 10248 13912 10260
rect 13679 10220 13912 10248
rect 13679 10217 13691 10220
rect 13633 10211 13691 10217
rect 13906 10208 13912 10220
rect 13964 10208 13970 10260
rect 14001 10251 14059 10257
rect 14001 10217 14013 10251
rect 14047 10248 14059 10251
rect 14274 10248 14280 10260
rect 14047 10220 14280 10248
rect 14047 10217 14059 10220
rect 14001 10211 14059 10217
rect 14274 10208 14280 10220
rect 14332 10208 14338 10260
rect 17494 10208 17500 10260
rect 17552 10248 17558 10260
rect 17681 10251 17739 10257
rect 17681 10248 17693 10251
rect 17552 10220 17693 10248
rect 17552 10208 17558 10220
rect 17681 10217 17693 10220
rect 17727 10248 17739 10251
rect 18693 10251 18751 10257
rect 17727 10220 18184 10248
rect 17727 10217 17739 10220
rect 17681 10211 17739 10217
rect 4617 10183 4675 10189
rect 4617 10149 4629 10183
rect 4663 10180 4675 10183
rect 4706 10180 4712 10192
rect 4663 10152 4712 10180
rect 4663 10149 4675 10152
rect 4617 10143 4675 10149
rect 4706 10140 4712 10152
rect 4764 10140 4770 10192
rect 7466 10180 7472 10192
rect 5276 10152 7472 10180
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10072 1458 10124
rect 2314 10112 2320 10124
rect 2275 10084 2320 10112
rect 2314 10072 2320 10084
rect 2372 10072 2378 10124
rect 2409 10115 2467 10121
rect 2409 10081 2421 10115
rect 2455 10112 2467 10115
rect 3329 10115 3387 10121
rect 2455 10084 3280 10112
rect 2455 10081 2467 10084
rect 2409 10075 2467 10081
rect 2590 10044 2596 10056
rect 2551 10016 2596 10044
rect 2590 10004 2596 10016
rect 2648 10004 2654 10056
rect 3252 10044 3280 10084
rect 3329 10081 3341 10115
rect 3375 10112 3387 10115
rect 5276 10112 5304 10152
rect 7466 10140 7472 10152
rect 7524 10140 7530 10192
rect 11600 10183 11658 10189
rect 7576 10152 11560 10180
rect 3375 10084 5304 10112
rect 5353 10115 5411 10121
rect 3375 10081 3387 10084
rect 3329 10075 3387 10081
rect 5353 10081 5365 10115
rect 5399 10081 5411 10115
rect 5534 10112 5540 10124
rect 5495 10084 5540 10112
rect 5353 10075 5411 10081
rect 3510 10044 3516 10056
rect 3252 10016 3516 10044
rect 3510 10004 3516 10016
rect 3568 10004 3574 10056
rect 3605 10047 3663 10053
rect 3605 10013 3617 10047
rect 3651 10044 3663 10047
rect 4614 10044 4620 10056
rect 3651 10016 4620 10044
rect 3651 10013 3663 10016
rect 3605 10007 3663 10013
rect 4614 10004 4620 10016
rect 4672 10004 4678 10056
rect 4801 10047 4859 10053
rect 4801 10013 4813 10047
rect 4847 10044 4859 10047
rect 5074 10044 5080 10056
rect 4847 10016 5080 10044
rect 4847 10013 4859 10016
rect 4801 10007 4859 10013
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 1581 9979 1639 9985
rect 1581 9945 1593 9979
rect 1627 9976 1639 9979
rect 2866 9976 2872 9988
rect 1627 9948 2872 9976
rect 1627 9945 1639 9948
rect 1581 9939 1639 9945
rect 2866 9936 2872 9948
rect 2924 9936 2930 9988
rect 2961 9979 3019 9985
rect 2961 9945 2973 9979
rect 3007 9976 3019 9979
rect 4338 9976 4344 9988
rect 3007 9948 4344 9976
rect 3007 9945 3019 9948
rect 2961 9939 3019 9945
rect 4338 9936 4344 9948
rect 4396 9936 4402 9988
rect 5368 9976 5396 10075
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 5626 10072 5632 10124
rect 5684 10112 5690 10124
rect 5804 10115 5862 10121
rect 5804 10112 5816 10115
rect 5684 10084 5816 10112
rect 5684 10072 5690 10084
rect 5804 10081 5816 10084
rect 5850 10112 5862 10115
rect 6178 10112 6184 10124
rect 5850 10084 6184 10112
rect 5850 10081 5862 10084
rect 5804 10075 5862 10081
rect 6178 10072 6184 10084
rect 6236 10072 6242 10124
rect 6362 10072 6368 10124
rect 6420 10112 6426 10124
rect 7576 10112 7604 10152
rect 6420 10084 7604 10112
rect 6420 10072 6426 10084
rect 7742 10072 7748 10124
rect 7800 10112 7806 10124
rect 8185 10115 8243 10121
rect 8185 10112 8197 10115
rect 7800 10084 8197 10112
rect 7800 10072 7806 10084
rect 8185 10081 8197 10084
rect 8231 10112 8243 10115
rect 9766 10112 9772 10124
rect 8231 10084 9772 10112
rect 8231 10081 8243 10084
rect 8185 10075 8243 10081
rect 9766 10072 9772 10084
rect 9824 10072 9830 10124
rect 10137 10115 10195 10121
rect 10137 10081 10149 10115
rect 10183 10112 10195 10115
rect 10594 10112 10600 10124
rect 10183 10084 10600 10112
rect 10183 10081 10195 10084
rect 10137 10075 10195 10081
rect 10594 10072 10600 10084
rect 10652 10072 10658 10124
rect 11532 10112 11560 10152
rect 11600 10149 11612 10183
rect 11646 10180 11658 10183
rect 11790 10180 11796 10192
rect 11646 10152 11796 10180
rect 11646 10149 11658 10152
rect 11600 10143 11658 10149
rect 11790 10140 11796 10152
rect 11848 10140 11854 10192
rect 18046 10180 18052 10192
rect 11992 10152 18052 10180
rect 11992 10112 12020 10152
rect 18046 10140 18052 10152
rect 18104 10140 18110 10192
rect 11532 10084 12020 10112
rect 14090 10072 14096 10124
rect 14148 10112 14154 10124
rect 15102 10112 15108 10124
rect 14148 10084 14193 10112
rect 15063 10084 15108 10112
rect 14148 10072 14154 10084
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 15286 10072 15292 10124
rect 15344 10112 15350 10124
rect 15657 10115 15715 10121
rect 15657 10112 15669 10115
rect 15344 10084 15669 10112
rect 15344 10072 15350 10084
rect 15657 10081 15669 10084
rect 15703 10081 15715 10115
rect 16206 10112 16212 10124
rect 15657 10075 15715 10081
rect 15948 10084 16212 10112
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10044 7895 10047
rect 7926 10044 7932 10056
rect 7883 10016 7932 10044
rect 7883 10013 7895 10016
rect 7837 10007 7895 10013
rect 7926 10004 7932 10016
rect 7984 10004 7990 10056
rect 9784 9976 9812 10072
rect 10229 10047 10287 10053
rect 10229 10013 10241 10047
rect 10275 10013 10287 10047
rect 10229 10007 10287 10013
rect 10244 9976 10272 10007
rect 11330 10004 11336 10056
rect 11388 10044 11394 10056
rect 11388 10016 11433 10044
rect 11388 10004 11394 10016
rect 12434 10004 12440 10056
rect 12492 10044 12498 10056
rect 13630 10044 13636 10056
rect 12492 10016 13636 10044
rect 12492 10004 12498 10016
rect 13630 10004 13636 10016
rect 13688 10004 13694 10056
rect 14182 10044 14188 10056
rect 14143 10016 14188 10044
rect 14182 10004 14188 10016
rect 14240 10004 14246 10056
rect 15746 10044 15752 10056
rect 15707 10016 15752 10044
rect 15746 10004 15752 10016
rect 15804 10004 15810 10056
rect 15948 10053 15976 10084
rect 16206 10072 16212 10084
rect 16264 10112 16270 10124
rect 16557 10115 16615 10121
rect 16557 10112 16569 10115
rect 16264 10084 16569 10112
rect 16264 10072 16270 10084
rect 16557 10081 16569 10084
rect 16603 10081 16615 10115
rect 17957 10115 18015 10121
rect 17957 10112 17969 10115
rect 16557 10075 16615 10081
rect 17328 10084 17969 10112
rect 15933 10047 15991 10053
rect 15933 10013 15945 10047
rect 15979 10013 15991 10047
rect 15933 10007 15991 10013
rect 16114 10004 16120 10056
rect 16172 10044 16178 10056
rect 16298 10044 16304 10056
rect 16172 10016 16304 10044
rect 16172 10004 16178 10016
rect 16298 10004 16304 10016
rect 16356 10004 16362 10056
rect 5368 9948 5580 9976
rect 9784 9948 10272 9976
rect 14921 9979 14979 9985
rect 3602 9868 3608 9920
rect 3660 9908 3666 9920
rect 5169 9911 5227 9917
rect 5169 9908 5181 9911
rect 3660 9880 5181 9908
rect 3660 9868 3666 9880
rect 5169 9877 5181 9880
rect 5215 9908 5227 9911
rect 5442 9908 5448 9920
rect 5215 9880 5448 9908
rect 5215 9877 5227 9880
rect 5169 9871 5227 9877
rect 5442 9868 5448 9880
rect 5500 9868 5506 9920
rect 5552 9908 5580 9948
rect 14921 9945 14933 9979
rect 14967 9976 14979 9979
rect 15378 9976 15384 9988
rect 14967 9948 15384 9976
rect 14967 9945 14979 9948
rect 14921 9939 14979 9945
rect 15378 9936 15384 9948
rect 15436 9976 15442 9988
rect 16132 9976 16160 10004
rect 15436 9948 16160 9976
rect 15436 9936 15442 9948
rect 7006 9908 7012 9920
rect 5552 9880 7012 9908
rect 7006 9868 7012 9880
rect 7064 9868 7070 9920
rect 8202 9868 8208 9920
rect 8260 9908 8266 9920
rect 9306 9908 9312 9920
rect 8260 9880 9312 9908
rect 8260 9868 8266 9880
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 12342 9868 12348 9920
rect 12400 9908 12406 9920
rect 12713 9911 12771 9917
rect 12713 9908 12725 9911
rect 12400 9880 12725 9908
rect 12400 9868 12406 9880
rect 12713 9877 12725 9880
rect 12759 9877 12771 9911
rect 12713 9871 12771 9877
rect 15289 9911 15347 9917
rect 15289 9877 15301 9911
rect 15335 9908 15347 9911
rect 17328 9908 17356 10084
rect 17957 10081 17969 10084
rect 18003 10081 18015 10115
rect 17957 10075 18015 10081
rect 18156 10044 18184 10220
rect 18693 10217 18705 10251
rect 18739 10248 18751 10251
rect 18874 10248 18880 10260
rect 18739 10220 18880 10248
rect 18739 10217 18751 10220
rect 18693 10211 18751 10217
rect 18874 10208 18880 10220
rect 18932 10208 18938 10260
rect 19153 10251 19211 10257
rect 19153 10217 19165 10251
rect 19199 10248 19211 10251
rect 19242 10248 19248 10260
rect 19199 10220 19248 10248
rect 19199 10217 19211 10220
rect 19153 10211 19211 10217
rect 19242 10208 19248 10220
rect 19300 10208 19306 10260
rect 18233 10183 18291 10189
rect 18233 10149 18245 10183
rect 18279 10180 18291 10183
rect 19334 10180 19340 10192
rect 18279 10152 19340 10180
rect 18279 10149 18291 10152
rect 18233 10143 18291 10149
rect 19334 10140 19340 10152
rect 19392 10140 19398 10192
rect 18414 10072 18420 10124
rect 18472 10112 18478 10124
rect 18874 10112 18880 10124
rect 18472 10084 18880 10112
rect 18472 10072 18478 10084
rect 18874 10072 18880 10084
rect 18932 10112 18938 10124
rect 19061 10115 19119 10121
rect 19061 10112 19073 10115
rect 18932 10084 19073 10112
rect 18932 10072 18938 10084
rect 19061 10081 19073 10084
rect 19107 10112 19119 10115
rect 20073 10115 20131 10121
rect 20073 10112 20085 10115
rect 19107 10084 20085 10112
rect 19107 10081 19119 10084
rect 19061 10075 19119 10081
rect 20073 10081 20085 10084
rect 20119 10081 20131 10115
rect 20073 10075 20131 10081
rect 19245 10047 19303 10053
rect 19245 10044 19257 10047
rect 18156 10016 19257 10044
rect 19245 10013 19257 10016
rect 19291 10013 19303 10047
rect 19245 10007 19303 10013
rect 20165 10047 20223 10053
rect 20165 10013 20177 10047
rect 20211 10013 20223 10047
rect 20346 10044 20352 10056
rect 20307 10016 20352 10044
rect 20165 10007 20223 10013
rect 20070 9936 20076 9988
rect 20128 9976 20134 9988
rect 20180 9976 20208 10007
rect 20346 10004 20352 10016
rect 20404 10004 20410 10056
rect 20128 9948 20208 9976
rect 20128 9936 20134 9948
rect 19702 9908 19708 9920
rect 15335 9880 17356 9908
rect 19663 9880 19708 9908
rect 15335 9877 15347 9880
rect 15289 9871 15347 9877
rect 19702 9868 19708 9880
rect 19760 9868 19766 9920
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 3142 9664 3148 9716
rect 3200 9704 3206 9716
rect 4433 9707 4491 9713
rect 4433 9704 4445 9707
rect 3200 9676 4445 9704
rect 3200 9664 3206 9676
rect 4433 9673 4445 9676
rect 4479 9673 4491 9707
rect 7926 9704 7932 9716
rect 4433 9667 4491 9673
rect 7760 9676 7932 9704
rect 4157 9639 4215 9645
rect 4157 9605 4169 9639
rect 4203 9636 4215 9639
rect 4203 9608 6132 9636
rect 4203 9605 4215 9608
rect 4157 9599 4215 9605
rect 1854 9528 1860 9580
rect 1912 9568 1918 9580
rect 1949 9571 2007 9577
rect 1949 9568 1961 9571
rect 1912 9540 1961 9568
rect 1912 9528 1918 9540
rect 1949 9537 1961 9540
rect 1995 9537 2007 9571
rect 5074 9568 5080 9580
rect 1949 9531 2007 9537
rect 4632 9540 4936 9568
rect 5035 9540 5080 9568
rect 1765 9503 1823 9509
rect 1765 9469 1777 9503
rect 1811 9500 1823 9503
rect 2222 9500 2228 9512
rect 1811 9472 2228 9500
rect 1811 9469 1823 9472
rect 1765 9463 1823 9469
rect 2222 9460 2228 9472
rect 2280 9460 2286 9512
rect 2777 9503 2835 9509
rect 2777 9469 2789 9503
rect 2823 9500 2835 9503
rect 2823 9472 3372 9500
rect 2823 9469 2835 9472
rect 2777 9463 2835 9469
rect 2866 9392 2872 9444
rect 2924 9432 2930 9444
rect 3022 9435 3080 9441
rect 3022 9432 3034 9435
rect 2924 9404 3034 9432
rect 2924 9392 2930 9404
rect 3022 9401 3034 9404
rect 3068 9401 3080 9435
rect 3022 9395 3080 9401
rect 3142 9392 3148 9444
rect 3200 9432 3206 9444
rect 3344 9432 3372 9472
rect 3418 9460 3424 9512
rect 3476 9500 3482 9512
rect 4632 9500 4660 9540
rect 4798 9500 4804 9512
rect 3476 9472 4660 9500
rect 4759 9472 4804 9500
rect 3476 9460 3482 9472
rect 4798 9460 4804 9472
rect 4856 9460 4862 9512
rect 4908 9500 4936 9540
rect 5074 9528 5080 9540
rect 5132 9528 5138 9580
rect 6104 9577 6132 9608
rect 6089 9571 6147 9577
rect 6089 9537 6101 9571
rect 6135 9568 6147 9571
rect 6178 9568 6184 9580
rect 6135 9540 6184 9568
rect 6135 9537 6147 9540
rect 6089 9531 6147 9537
rect 6178 9528 6184 9540
rect 6236 9528 6242 9580
rect 7285 9571 7343 9577
rect 7285 9537 7297 9571
rect 7331 9568 7343 9571
rect 7558 9568 7564 9580
rect 7331 9540 7564 9568
rect 7331 9537 7343 9540
rect 7285 9531 7343 9537
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 7760 9577 7788 9676
rect 7926 9664 7932 9676
rect 7984 9664 7990 9716
rect 9784 9676 10824 9704
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9537 7803 9571
rect 7745 9531 7803 9537
rect 5905 9503 5963 9509
rect 5905 9500 5917 9503
rect 4908 9472 5917 9500
rect 5905 9469 5917 9472
rect 5951 9500 5963 9503
rect 7466 9500 7472 9512
rect 5951 9472 7472 9500
rect 5951 9469 5963 9472
rect 5905 9463 5963 9469
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 9784 9500 9812 9676
rect 10796 9636 10824 9676
rect 12986 9664 12992 9716
rect 13044 9704 13050 9716
rect 16206 9704 16212 9716
rect 13044 9676 16068 9704
rect 16167 9676 16212 9704
rect 13044 9664 13050 9676
rect 14274 9636 14280 9648
rect 10796 9608 14280 9636
rect 14274 9596 14280 9608
rect 14332 9596 14338 9648
rect 16040 9636 16068 9676
rect 16206 9664 16212 9676
rect 16264 9664 16270 9716
rect 18506 9704 18512 9716
rect 16316 9676 18512 9704
rect 16316 9636 16344 9676
rect 18506 9664 18512 9676
rect 18564 9664 18570 9716
rect 19242 9664 19248 9716
rect 19300 9664 19306 9716
rect 16040 9608 16344 9636
rect 16390 9596 16396 9648
rect 16448 9636 16454 9648
rect 16448 9608 17172 9636
rect 16448 9596 16454 9608
rect 10870 9528 10876 9580
rect 10928 9568 10934 9580
rect 12897 9571 12955 9577
rect 12897 9568 12909 9571
rect 10928 9540 12909 9568
rect 10928 9528 10934 9540
rect 12897 9537 12909 9540
rect 12943 9537 12955 9571
rect 13078 9568 13084 9580
rect 13039 9540 13084 9568
rect 12897 9531 12955 9537
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 16942 9528 16948 9580
rect 17000 9568 17006 9580
rect 17037 9571 17095 9577
rect 17037 9568 17049 9571
rect 17000 9540 17049 9568
rect 17000 9528 17006 9540
rect 17037 9537 17049 9540
rect 17083 9537 17095 9571
rect 17144 9568 17172 9608
rect 17402 9596 17408 9648
rect 17460 9636 17466 9648
rect 18233 9639 18291 9645
rect 18233 9636 18245 9639
rect 17460 9608 18245 9636
rect 17460 9596 17466 9608
rect 18233 9605 18245 9608
rect 18279 9605 18291 9639
rect 19260 9636 19288 9664
rect 18233 9599 18291 9605
rect 18331 9608 19288 9636
rect 18331 9568 18359 9608
rect 19334 9596 19340 9648
rect 19392 9596 19398 9648
rect 19426 9596 19432 9648
rect 19484 9596 19490 9648
rect 19521 9639 19579 9645
rect 19521 9605 19533 9639
rect 19567 9636 19579 9639
rect 20530 9636 20536 9648
rect 19567 9608 20536 9636
rect 19567 9605 19579 9608
rect 19521 9599 19579 9605
rect 20530 9596 20536 9608
rect 20588 9596 20594 9648
rect 18690 9568 18696 9580
rect 17144 9540 18359 9568
rect 18651 9540 18696 9568
rect 17037 9531 17095 9537
rect 18690 9528 18696 9540
rect 18748 9528 18754 9580
rect 18877 9571 18935 9577
rect 18877 9537 18889 9571
rect 18923 9568 18935 9571
rect 18966 9568 18972 9580
rect 18923 9540 18972 9568
rect 18923 9537 18935 9540
rect 18877 9531 18935 9537
rect 18966 9528 18972 9540
rect 19024 9528 19030 9580
rect 7852 9472 9812 9500
rect 9861 9503 9919 9509
rect 3602 9432 3608 9444
rect 3200 9404 3608 9432
rect 3200 9392 3206 9404
rect 3602 9392 3608 9404
rect 3660 9392 3666 9444
rect 4062 9392 4068 9444
rect 4120 9432 4126 9444
rect 7852 9432 7880 9472
rect 9861 9469 9873 9503
rect 9907 9469 9919 9503
rect 9861 9463 9919 9469
rect 10128 9503 10186 9509
rect 10128 9469 10140 9503
rect 10174 9500 10186 9503
rect 12342 9500 12348 9512
rect 10174 9472 12348 9500
rect 10174 9469 10186 9472
rect 10128 9463 10186 9469
rect 4120 9404 7880 9432
rect 8012 9435 8070 9441
rect 4120 9392 4126 9404
rect 8012 9401 8024 9435
rect 8058 9432 8070 9435
rect 8202 9432 8208 9444
rect 8058 9404 8208 9432
rect 8058 9401 8070 9404
rect 8012 9395 8070 9401
rect 8202 9392 8208 9404
rect 8260 9392 8266 9444
rect 8662 9392 8668 9444
rect 8720 9432 8726 9444
rect 9876 9432 9904 9463
rect 12342 9460 12348 9472
rect 12400 9460 12406 9512
rect 13262 9500 13268 9512
rect 12544 9472 13268 9500
rect 8720 9404 9904 9432
rect 8720 9392 8726 9404
rect 10226 9392 10232 9444
rect 10284 9432 10290 9444
rect 12544 9432 12572 9472
rect 13262 9460 13268 9472
rect 13320 9460 13326 9512
rect 14829 9503 14887 9509
rect 14829 9469 14841 9503
rect 14875 9500 14887 9503
rect 15378 9500 15384 9512
rect 14875 9472 15384 9500
rect 14875 9469 14887 9472
rect 14829 9463 14887 9469
rect 15378 9460 15384 9472
rect 15436 9460 15442 9512
rect 15930 9460 15936 9512
rect 15988 9500 15994 9512
rect 15988 9472 16988 9500
rect 15988 9460 15994 9472
rect 10284 9404 12572 9432
rect 10284 9392 10290 9404
rect 12618 9392 12624 9444
rect 12676 9432 12682 9444
rect 12805 9435 12863 9441
rect 12805 9432 12817 9435
rect 12676 9404 12817 9432
rect 12676 9392 12682 9404
rect 12805 9401 12817 9404
rect 12851 9401 12863 9435
rect 12805 9395 12863 9401
rect 15010 9392 15016 9444
rect 15068 9441 15074 9444
rect 15068 9435 15132 9441
rect 15068 9401 15086 9435
rect 15120 9401 15132 9435
rect 16853 9435 16911 9441
rect 16853 9432 16865 9435
rect 15068 9395 15132 9401
rect 15764 9404 16865 9432
rect 15068 9392 15074 9395
rect 4893 9367 4951 9373
rect 4893 9333 4905 9367
rect 4939 9364 4951 9367
rect 5445 9367 5503 9373
rect 5445 9364 5457 9367
rect 4939 9336 5457 9364
rect 4939 9333 4951 9336
rect 4893 9327 4951 9333
rect 5445 9333 5457 9336
rect 5491 9333 5503 9367
rect 5445 9327 5503 9333
rect 5626 9324 5632 9376
rect 5684 9364 5690 9376
rect 5813 9367 5871 9373
rect 5813 9364 5825 9367
rect 5684 9336 5825 9364
rect 5684 9324 5690 9336
rect 5813 9333 5825 9336
rect 5859 9333 5871 9367
rect 5813 9327 5871 9333
rect 5902 9324 5908 9376
rect 5960 9364 5966 9376
rect 6730 9364 6736 9376
rect 5960 9336 6736 9364
rect 5960 9324 5966 9336
rect 6730 9324 6736 9336
rect 6788 9364 6794 9376
rect 9125 9367 9183 9373
rect 9125 9364 9137 9367
rect 6788 9336 9137 9364
rect 6788 9324 6794 9336
rect 9125 9333 9137 9336
rect 9171 9333 9183 9367
rect 9125 9327 9183 9333
rect 10962 9324 10968 9376
rect 11020 9364 11026 9376
rect 11241 9367 11299 9373
rect 11241 9364 11253 9367
rect 11020 9336 11253 9364
rect 11020 9324 11026 9336
rect 11241 9333 11253 9336
rect 11287 9333 11299 9367
rect 11241 9327 11299 9333
rect 12437 9367 12495 9373
rect 12437 9333 12449 9367
rect 12483 9364 12495 9367
rect 12526 9364 12532 9376
rect 12483 9336 12532 9364
rect 12483 9333 12495 9336
rect 12437 9327 12495 9333
rect 12526 9324 12532 9336
rect 12584 9324 12590 9376
rect 14369 9367 14427 9373
rect 14369 9333 14381 9367
rect 14415 9364 14427 9367
rect 15764 9364 15792 9404
rect 16853 9401 16865 9404
rect 16899 9401 16911 9435
rect 16960 9432 16988 9472
rect 17954 9460 17960 9512
rect 18012 9500 18018 9512
rect 19352 9509 19380 9596
rect 18601 9503 18659 9509
rect 18601 9500 18613 9503
rect 18012 9472 18613 9500
rect 18012 9460 18018 9472
rect 18601 9469 18613 9472
rect 18647 9469 18659 9503
rect 18601 9463 18659 9469
rect 19337 9503 19395 9509
rect 19337 9469 19349 9503
rect 19383 9469 19395 9503
rect 19337 9463 19395 9469
rect 18046 9432 18052 9444
rect 16960 9404 18052 9432
rect 16853 9395 16911 9401
rect 18046 9392 18052 9404
rect 18104 9392 18110 9444
rect 19444 9432 19472 9596
rect 20346 9528 20352 9580
rect 20404 9568 20410 9580
rect 20441 9571 20499 9577
rect 20441 9568 20453 9571
rect 20404 9540 20453 9568
rect 20404 9528 20410 9540
rect 20441 9537 20453 9540
rect 20487 9537 20499 9571
rect 20441 9531 20499 9537
rect 20349 9435 20407 9441
rect 20349 9432 20361 9435
rect 19444 9404 20361 9432
rect 20349 9401 20361 9404
rect 20395 9401 20407 9435
rect 20349 9395 20407 9401
rect 16482 9364 16488 9376
rect 14415 9336 15792 9364
rect 16443 9336 16488 9364
rect 14415 9333 14427 9336
rect 14369 9327 14427 9333
rect 16482 9324 16488 9336
rect 16540 9324 16546 9376
rect 16666 9324 16672 9376
rect 16724 9364 16730 9376
rect 16945 9367 17003 9373
rect 16945 9364 16957 9367
rect 16724 9336 16957 9364
rect 16724 9324 16730 9336
rect 16945 9333 16957 9336
rect 16991 9333 17003 9367
rect 19886 9364 19892 9376
rect 19847 9336 19892 9364
rect 16945 9327 17003 9333
rect 19886 9324 19892 9336
rect 19944 9324 19950 9376
rect 20254 9364 20260 9376
rect 20215 9336 20260 9364
rect 20254 9324 20260 9336
rect 20312 9324 20318 9376
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 2222 9160 2228 9172
rect 2183 9132 2228 9160
rect 2222 9120 2228 9132
rect 2280 9120 2286 9172
rect 4525 9163 4583 9169
rect 4525 9129 4537 9163
rect 4571 9160 4583 9163
rect 4706 9160 4712 9172
rect 4571 9132 4712 9160
rect 4571 9129 4583 9132
rect 4525 9123 4583 9129
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 5166 9120 5172 9172
rect 5224 9160 5230 9172
rect 5445 9163 5503 9169
rect 5445 9160 5457 9163
rect 5224 9132 5457 9160
rect 5224 9120 5230 9132
rect 5445 9129 5457 9132
rect 5491 9129 5503 9163
rect 5445 9123 5503 9129
rect 5537 9163 5595 9169
rect 5537 9129 5549 9163
rect 5583 9160 5595 9163
rect 6086 9160 6092 9172
rect 5583 9132 6092 9160
rect 5583 9129 5595 9132
rect 5537 9123 5595 9129
rect 6086 9120 6092 9132
rect 6144 9120 6150 9172
rect 7282 9160 7288 9172
rect 7243 9132 7288 9160
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 7466 9120 7472 9172
rect 7524 9160 7530 9172
rect 7745 9163 7803 9169
rect 7745 9160 7757 9163
rect 7524 9132 7757 9160
rect 7524 9120 7530 9132
rect 7745 9129 7757 9132
rect 7791 9129 7803 9163
rect 8294 9160 8300 9172
rect 8255 9132 8300 9160
rect 7745 9123 7803 9129
rect 8294 9120 8300 9132
rect 8352 9120 8358 9172
rect 8570 9120 8576 9172
rect 8628 9160 8634 9172
rect 8665 9163 8723 9169
rect 8665 9160 8677 9163
rect 8628 9132 8677 9160
rect 8628 9120 8634 9132
rect 8665 9129 8677 9132
rect 8711 9129 8723 9163
rect 8665 9123 8723 9129
rect 8757 9163 8815 9169
rect 8757 9129 8769 9163
rect 8803 9160 8815 9163
rect 10226 9160 10232 9172
rect 8803 9132 10232 9160
rect 8803 9129 8815 9132
rect 8757 9123 8815 9129
rect 3970 9092 3976 9104
rect 1504 9064 3976 9092
rect 1504 9033 1532 9064
rect 3970 9052 3976 9064
rect 4028 9052 4034 9104
rect 7653 9095 7711 9101
rect 7653 9092 7665 9095
rect 5000 9064 7665 9092
rect 1489 9027 1547 9033
rect 1489 8993 1501 9027
rect 1535 8993 1547 9027
rect 2590 9024 2596 9036
rect 2551 8996 2596 9024
rect 1489 8987 1547 8993
rect 2590 8984 2596 8996
rect 2648 8984 2654 9036
rect 3694 8984 3700 9036
rect 3752 9024 3758 9036
rect 4893 9027 4951 9033
rect 4893 9024 4905 9027
rect 3752 8996 4905 9024
rect 3752 8984 3758 8996
rect 4893 8993 4905 8996
rect 4939 8993 4951 9027
rect 4893 8987 4951 8993
rect 1394 8916 1400 8968
rect 1452 8956 1458 8968
rect 1673 8959 1731 8965
rect 1673 8956 1685 8959
rect 1452 8928 1685 8956
rect 1452 8916 1458 8928
rect 1673 8925 1685 8928
rect 1719 8925 1731 8959
rect 1673 8919 1731 8925
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8925 2743 8959
rect 2866 8956 2872 8968
rect 2827 8928 2872 8956
rect 2685 8919 2743 8925
rect 2700 8888 2728 8919
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 4154 8916 4160 8968
rect 4212 8956 4218 8968
rect 5000 8965 5028 9064
rect 7653 9061 7665 9064
rect 7699 9061 7711 9095
rect 7653 9055 7711 9061
rect 5166 9024 5172 9036
rect 5092 8996 5172 9024
rect 5092 8965 5120 8996
rect 5166 8984 5172 8996
rect 5224 8984 5230 9036
rect 5902 9024 5908 9036
rect 5863 8996 5908 9024
rect 5902 8984 5908 8996
rect 5960 9024 5966 9036
rect 6638 9024 6644 9036
rect 5960 8996 6644 9024
rect 5960 8984 5966 8996
rect 6638 8984 6644 8996
rect 6696 8984 6702 9036
rect 8680 9024 8708 9123
rect 10226 9120 10232 9132
rect 10284 9120 10290 9172
rect 10870 9160 10876 9172
rect 10831 9132 10876 9160
rect 10870 9120 10876 9132
rect 10928 9120 10934 9172
rect 11698 9120 11704 9172
rect 11756 9160 11762 9172
rect 12158 9160 12164 9172
rect 11756 9132 12164 9160
rect 11756 9120 11762 9132
rect 12158 9120 12164 9132
rect 12216 9120 12222 9172
rect 14921 9163 14979 9169
rect 14921 9129 14933 9163
rect 14967 9160 14979 9163
rect 15010 9160 15016 9172
rect 14967 9132 15016 9160
rect 14967 9129 14979 9132
rect 14921 9123 14979 9129
rect 15010 9120 15016 9132
rect 15068 9120 15074 9172
rect 15286 9160 15292 9172
rect 15247 9132 15292 9160
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 15749 9163 15807 9169
rect 15749 9129 15761 9163
rect 15795 9160 15807 9163
rect 16301 9163 16359 9169
rect 16301 9160 16313 9163
rect 15795 9132 16313 9160
rect 15795 9129 15807 9132
rect 15749 9123 15807 9129
rect 16301 9129 16313 9132
rect 16347 9129 16359 9163
rect 16301 9123 16359 9129
rect 16574 9120 16580 9172
rect 16632 9160 16638 9172
rect 16669 9163 16727 9169
rect 16669 9160 16681 9163
rect 16632 9132 16681 9160
rect 16632 9120 16638 9132
rect 16669 9129 16681 9132
rect 16715 9129 16727 9163
rect 16669 9123 16727 9129
rect 16758 9120 16764 9172
rect 16816 9160 16822 9172
rect 19613 9163 19671 9169
rect 19613 9160 19625 9163
rect 16816 9132 19625 9160
rect 16816 9120 16822 9132
rect 19613 9129 19625 9132
rect 19659 9129 19671 9163
rect 19794 9160 19800 9172
rect 19755 9132 19800 9160
rect 19613 9123 19671 9129
rect 19794 9120 19800 9132
rect 19852 9120 19858 9172
rect 20254 9120 20260 9172
rect 20312 9160 20318 9172
rect 20901 9163 20959 9169
rect 20901 9160 20913 9163
rect 20312 9132 20913 9160
rect 20312 9120 20318 9132
rect 20901 9129 20913 9132
rect 20947 9129 20959 9163
rect 20901 9123 20959 9129
rect 10042 9092 10048 9104
rect 10003 9064 10048 9092
rect 10042 9052 10048 9064
rect 10100 9052 10106 9104
rect 10134 9052 10140 9104
rect 10192 9092 10198 9104
rect 11241 9095 11299 9101
rect 10192 9064 10237 9092
rect 10192 9052 10198 9064
rect 11241 9061 11253 9095
rect 11287 9092 11299 9095
rect 11974 9092 11980 9104
rect 11287 9064 11980 9092
rect 11287 9061 11299 9064
rect 11241 9055 11299 9061
rect 11974 9052 11980 9064
rect 12032 9052 12038 9104
rect 12802 9052 12808 9104
rect 12860 9092 12866 9104
rect 12986 9092 12992 9104
rect 12860 9064 12992 9092
rect 12860 9052 12866 9064
rect 12986 9052 12992 9064
rect 13044 9092 13050 9104
rect 15657 9095 15715 9101
rect 13044 9064 15056 9092
rect 13044 9052 13050 9064
rect 10870 9024 10876 9036
rect 6748 8996 8055 9024
rect 8680 8996 10876 9024
rect 4985 8959 5043 8965
rect 4985 8956 4997 8959
rect 4212 8928 4997 8956
rect 4212 8916 4218 8928
rect 4985 8925 4997 8928
rect 5031 8925 5043 8959
rect 4985 8919 5043 8925
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8925 5135 8959
rect 5442 8956 5448 8968
rect 5355 8928 5448 8956
rect 5077 8919 5135 8925
rect 5442 8916 5448 8928
rect 5500 8956 5506 8968
rect 5997 8959 6055 8965
rect 5997 8956 6009 8959
rect 5500 8928 6009 8956
rect 5500 8916 5506 8928
rect 5997 8925 6009 8928
rect 6043 8925 6055 8959
rect 6178 8956 6184 8968
rect 6091 8928 6184 8956
rect 5997 8919 6055 8925
rect 6178 8916 6184 8928
rect 6236 8956 6242 8968
rect 6748 8956 6776 8996
rect 6236 8928 6776 8956
rect 6236 8916 6242 8928
rect 7834 8916 7840 8968
rect 7892 8956 7898 8968
rect 8027 8956 8055 8996
rect 10870 8984 10876 8996
rect 10928 8984 10934 9036
rect 12141 9027 12199 9033
rect 12141 9024 12153 9027
rect 11532 8996 12153 9024
rect 11532 8965 11560 8996
rect 12141 8993 12153 8996
rect 12187 9024 12199 9027
rect 12894 9024 12900 9036
rect 12187 8996 12900 9024
rect 12187 8993 12199 8996
rect 12141 8987 12199 8993
rect 12894 8984 12900 8996
rect 12952 8984 12958 9036
rect 13078 8984 13084 9036
rect 13136 9024 13142 9036
rect 13808 9027 13866 9033
rect 13808 9024 13820 9027
rect 13136 8996 13820 9024
rect 13136 8984 13142 8996
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 7892 8928 7937 8956
rect 8027 8928 8953 8956
rect 7892 8916 7898 8928
rect 8941 8925 8953 8928
rect 8987 8956 8999 8959
rect 10229 8959 10287 8965
rect 10229 8956 10241 8959
rect 8987 8928 10241 8956
rect 8987 8925 8999 8928
rect 8941 8919 8999 8925
rect 10229 8925 10241 8928
rect 10275 8925 10287 8959
rect 11333 8959 11391 8965
rect 11333 8956 11345 8959
rect 10229 8919 10287 8925
rect 10336 8928 11345 8956
rect 3234 8888 3240 8900
rect 2700 8860 3240 8888
rect 3234 8848 3240 8860
rect 3292 8848 3298 8900
rect 4798 8848 4804 8900
rect 4856 8888 4862 8900
rect 5902 8888 5908 8900
rect 4856 8860 5908 8888
rect 4856 8848 4862 8860
rect 5902 8848 5908 8860
rect 5960 8848 5966 8900
rect 6822 8848 6828 8900
rect 6880 8888 6886 8900
rect 9674 8888 9680 8900
rect 6880 8860 7420 8888
rect 9635 8860 9680 8888
rect 6880 8848 6886 8860
rect 4706 8780 4712 8832
rect 4764 8820 4770 8832
rect 7190 8820 7196 8832
rect 4764 8792 7196 8820
rect 4764 8780 4770 8792
rect 7190 8780 7196 8792
rect 7248 8780 7254 8832
rect 7392 8820 7420 8860
rect 9674 8848 9680 8860
rect 9732 8848 9738 8900
rect 10336 8820 10364 8928
rect 11333 8925 11345 8928
rect 11379 8925 11391 8959
rect 11333 8919 11391 8925
rect 11517 8959 11575 8965
rect 11517 8925 11529 8959
rect 11563 8925 11575 8959
rect 11882 8956 11888 8968
rect 11795 8928 11888 8956
rect 11517 8919 11575 8925
rect 11348 8888 11376 8919
rect 11882 8916 11888 8928
rect 11940 8916 11946 8968
rect 11790 8888 11796 8900
rect 11348 8860 11796 8888
rect 11790 8848 11796 8860
rect 11848 8848 11854 8900
rect 7392 8792 10364 8820
rect 11146 8780 11152 8832
rect 11204 8820 11210 8832
rect 11900 8820 11928 8916
rect 13280 8897 13308 8996
rect 13808 8993 13820 8996
rect 13854 9024 13866 9027
rect 15028 9024 15056 9064
rect 15657 9061 15669 9095
rect 15703 9092 15715 9095
rect 16482 9092 16488 9104
rect 15703 9064 16488 9092
rect 15703 9061 15715 9064
rect 15657 9055 15715 9061
rect 16482 9052 16488 9064
rect 16540 9052 16546 9104
rect 18322 9092 18328 9104
rect 16592 9064 18328 9092
rect 16592 9024 16620 9064
rect 18322 9052 18328 9064
rect 18380 9092 18386 9104
rect 18690 9092 18696 9104
rect 18380 9064 18696 9092
rect 18380 9052 18386 9064
rect 18690 9052 18696 9064
rect 18748 9052 18754 9104
rect 18874 9052 18880 9104
rect 18932 9092 18938 9104
rect 19058 9092 19064 9104
rect 18932 9064 19064 9092
rect 18932 9052 18938 9064
rect 19058 9052 19064 9064
rect 19116 9052 19122 9104
rect 13854 8996 14964 9024
rect 15028 8996 16620 9024
rect 16761 9027 16819 9033
rect 13854 8993 13866 8996
rect 13808 8987 13866 8993
rect 13541 8959 13599 8965
rect 13541 8925 13553 8959
rect 13587 8925 13599 8959
rect 13541 8919 13599 8925
rect 13265 8891 13323 8897
rect 13265 8857 13277 8891
rect 13311 8857 13323 8891
rect 13265 8851 13323 8857
rect 12250 8820 12256 8832
rect 11204 8792 12256 8820
rect 11204 8780 11210 8792
rect 12250 8780 12256 8792
rect 12308 8820 12314 8832
rect 13556 8820 13584 8919
rect 14936 8888 14964 8996
rect 16761 8993 16773 9027
rect 16807 9024 16819 9027
rect 17770 9024 17776 9036
rect 16807 8996 17776 9024
rect 16807 8993 16819 8996
rect 16761 8987 16819 8993
rect 17770 8984 17776 8996
rect 17828 8984 17834 9036
rect 18408 9027 18466 9033
rect 18408 8993 18420 9027
rect 18454 9024 18466 9027
rect 19334 9024 19340 9036
rect 18454 8996 19340 9024
rect 18454 8993 18466 8996
rect 18408 8987 18466 8993
rect 19334 8984 19340 8996
rect 19392 8984 19398 9036
rect 19426 8984 19432 9036
rect 19484 9024 19490 9036
rect 20165 9027 20223 9033
rect 20165 9024 20177 9027
rect 19484 8996 20177 9024
rect 19484 8984 19490 8996
rect 20165 8993 20177 8996
rect 20211 8993 20223 9027
rect 20165 8987 20223 8993
rect 15013 8959 15071 8965
rect 15013 8925 15025 8959
rect 15059 8956 15071 8959
rect 15378 8956 15384 8968
rect 15059 8928 15384 8956
rect 15059 8925 15071 8928
rect 15013 8919 15071 8925
rect 15378 8916 15384 8928
rect 15436 8956 15442 8968
rect 15841 8959 15899 8965
rect 15841 8956 15853 8959
rect 15436 8928 15853 8956
rect 15436 8916 15442 8928
rect 15841 8925 15853 8928
rect 15887 8925 15899 8959
rect 15841 8919 15899 8925
rect 16298 8916 16304 8968
rect 16356 8956 16362 8968
rect 16574 8956 16580 8968
rect 16356 8928 16580 8956
rect 16356 8916 16362 8928
rect 16574 8916 16580 8928
rect 16632 8916 16638 8968
rect 16942 8956 16948 8968
rect 16903 8928 16948 8956
rect 16942 8916 16948 8928
rect 17000 8916 17006 8968
rect 17862 8916 17868 8968
rect 17920 8956 17926 8968
rect 18141 8959 18199 8965
rect 18141 8956 18153 8959
rect 17920 8928 18153 8956
rect 17920 8916 17926 8928
rect 18141 8925 18153 8928
rect 18187 8925 18199 8959
rect 18141 8919 18199 8925
rect 19518 8916 19524 8968
rect 19576 8956 19582 8968
rect 19613 8959 19671 8965
rect 19613 8956 19625 8959
rect 19576 8928 19625 8956
rect 19576 8916 19582 8928
rect 19613 8925 19625 8928
rect 19659 8925 19671 8959
rect 20254 8956 20260 8968
rect 20215 8928 20260 8956
rect 19613 8919 19671 8925
rect 20254 8916 20260 8928
rect 20312 8916 20318 8968
rect 20349 8959 20407 8965
rect 20349 8925 20361 8959
rect 20395 8925 20407 8959
rect 20349 8919 20407 8925
rect 16960 8888 16988 8916
rect 20364 8888 20392 8919
rect 14936 8860 16988 8888
rect 19536 8860 20392 8888
rect 12308 8792 13584 8820
rect 12308 8780 12314 8792
rect 15102 8780 15108 8832
rect 15160 8820 15166 8832
rect 19536 8829 19564 8860
rect 19521 8823 19579 8829
rect 19521 8820 19533 8823
rect 15160 8792 19533 8820
rect 15160 8780 15166 8792
rect 19521 8789 19533 8792
rect 19567 8789 19579 8823
rect 19521 8783 19579 8789
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 2866 8576 2872 8628
rect 2924 8616 2930 8628
rect 2961 8619 3019 8625
rect 2961 8616 2973 8619
rect 2924 8588 2973 8616
rect 2924 8576 2930 8588
rect 2961 8585 2973 8588
rect 3007 8585 3019 8619
rect 3234 8616 3240 8628
rect 3195 8588 3240 8616
rect 2961 8579 3019 8585
rect 3234 8576 3240 8588
rect 3292 8576 3298 8628
rect 4062 8576 4068 8628
rect 4120 8616 4126 8628
rect 12434 8616 12440 8628
rect 4120 8588 12440 8616
rect 4120 8576 4126 8588
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 14829 8619 14887 8625
rect 14829 8585 14841 8619
rect 14875 8616 14887 8619
rect 15746 8616 15752 8628
rect 14875 8588 15752 8616
rect 14875 8585 14887 8588
rect 14829 8579 14887 8585
rect 15746 8576 15752 8588
rect 15804 8576 15810 8628
rect 16945 8619 17003 8625
rect 16945 8585 16957 8619
rect 16991 8616 17003 8619
rect 16991 8588 19104 8616
rect 16991 8585 17003 8588
rect 16945 8579 17003 8585
rect 7653 8551 7711 8557
rect 7653 8548 7665 8551
rect 3712 8520 7665 8548
rect 3712 8489 3740 8520
rect 7653 8517 7665 8520
rect 7699 8517 7711 8551
rect 7653 8511 7711 8517
rect 10045 8551 10103 8557
rect 10045 8517 10057 8551
rect 10091 8548 10103 8551
rect 11333 8551 11391 8557
rect 11333 8548 11345 8551
rect 10091 8520 10180 8548
rect 10091 8517 10103 8520
rect 10045 8511 10103 8517
rect 3697 8483 3755 8489
rect 3697 8449 3709 8483
rect 3743 8449 3755 8483
rect 3697 8443 3755 8449
rect 3881 8483 3939 8489
rect 3881 8449 3893 8483
rect 3927 8449 3939 8483
rect 4706 8480 4712 8492
rect 4667 8452 4712 8480
rect 3881 8443 3939 8449
rect 1578 8412 1584 8424
rect 1539 8384 1584 8412
rect 1578 8372 1584 8384
rect 1636 8372 1642 8424
rect 1848 8347 1906 8353
rect 1848 8313 1860 8347
rect 1894 8344 1906 8347
rect 3786 8344 3792 8356
rect 1894 8316 3792 8344
rect 1894 8313 1906 8316
rect 1848 8307 1906 8313
rect 3786 8304 3792 8316
rect 3844 8344 3850 8356
rect 3896 8344 3924 8443
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 4893 8483 4951 8489
rect 4893 8449 4905 8483
rect 4939 8480 4951 8483
rect 5350 8480 5356 8492
rect 4939 8452 5356 8480
rect 4939 8449 4951 8452
rect 4893 8443 4951 8449
rect 5350 8440 5356 8452
rect 5408 8440 5414 8492
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8480 5963 8483
rect 7098 8480 7104 8492
rect 5951 8452 7104 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 7561 8483 7619 8489
rect 7561 8449 7573 8483
rect 7607 8480 7619 8483
rect 8202 8480 8208 8492
rect 7607 8452 8208 8480
rect 7607 8449 7619 8452
rect 7561 8443 7619 8449
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 8312 8452 8800 8480
rect 4157 8415 4215 8421
rect 4157 8381 4169 8415
rect 4203 8412 4215 8415
rect 6546 8412 6552 8424
rect 4203 8384 6552 8412
rect 4203 8381 4215 8384
rect 4157 8375 4215 8381
rect 6546 8372 6552 8384
rect 6604 8372 6610 8424
rect 8312 8412 8340 8452
rect 8662 8412 8668 8424
rect 6748 8384 8340 8412
rect 8623 8384 8668 8412
rect 3844 8316 3924 8344
rect 3844 8304 3850 8316
rect 3970 8304 3976 8356
rect 4028 8344 4034 8356
rect 4617 8347 4675 8353
rect 4028 8316 4568 8344
rect 4028 8304 4034 8316
rect 3602 8276 3608 8288
rect 3563 8248 3608 8276
rect 3602 8236 3608 8248
rect 3660 8236 3666 8288
rect 4157 8279 4215 8285
rect 4157 8245 4169 8279
rect 4203 8276 4215 8279
rect 4249 8279 4307 8285
rect 4249 8276 4261 8279
rect 4203 8248 4261 8276
rect 4203 8245 4215 8248
rect 4157 8239 4215 8245
rect 4249 8245 4261 8248
rect 4295 8245 4307 8279
rect 4540 8276 4568 8316
rect 4617 8313 4629 8347
rect 4663 8344 4675 8347
rect 4798 8344 4804 8356
rect 4663 8316 4804 8344
rect 4663 8313 4675 8316
rect 4617 8307 4675 8313
rect 4798 8304 4804 8316
rect 4856 8304 4862 8356
rect 5166 8304 5172 8356
rect 5224 8344 5230 8356
rect 5629 8347 5687 8353
rect 5629 8344 5641 8347
rect 5224 8316 5641 8344
rect 5224 8304 5230 8316
rect 5629 8313 5641 8316
rect 5675 8313 5687 8347
rect 5629 8307 5687 8313
rect 5721 8347 5779 8353
rect 5721 8313 5733 8347
rect 5767 8344 5779 8347
rect 6178 8344 6184 8356
rect 5767 8316 6184 8344
rect 5767 8313 5779 8316
rect 5721 8307 5779 8313
rect 6178 8304 6184 8316
rect 6236 8304 6242 8356
rect 6748 8344 6776 8384
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 8772 8412 8800 8452
rect 10152 8412 10180 8520
rect 10796 8520 11345 8548
rect 10796 8489 10824 8520
rect 11333 8517 11345 8520
rect 11379 8517 11391 8551
rect 11333 8511 11391 8517
rect 10781 8483 10839 8489
rect 10781 8449 10793 8483
rect 10827 8449 10839 8483
rect 10781 8443 10839 8449
rect 10873 8483 10931 8489
rect 10873 8449 10885 8483
rect 10919 8449 10931 8483
rect 10873 8443 10931 8449
rect 10888 8412 10916 8443
rect 10962 8440 10968 8492
rect 11020 8480 11026 8492
rect 11885 8483 11943 8489
rect 11885 8480 11897 8483
rect 11020 8452 11897 8480
rect 11020 8440 11026 8452
rect 11885 8449 11897 8452
rect 11931 8449 11943 8483
rect 11885 8443 11943 8449
rect 12250 8440 12256 8492
rect 12308 8480 12314 8492
rect 12437 8483 12495 8489
rect 12437 8480 12449 8483
rect 12308 8452 12449 8480
rect 12308 8440 12314 8452
rect 12437 8449 12449 8452
rect 12483 8449 12495 8483
rect 15378 8480 15384 8492
rect 15339 8452 15384 8480
rect 12437 8443 12495 8449
rect 15378 8440 15384 8452
rect 15436 8440 15442 8492
rect 16485 8483 16543 8489
rect 16485 8449 16497 8483
rect 16531 8480 16543 8483
rect 16942 8480 16948 8492
rect 16531 8452 16948 8480
rect 16531 8449 16543 8452
rect 16485 8443 16543 8449
rect 16942 8440 16948 8452
rect 17000 8440 17006 8492
rect 17589 8483 17647 8489
rect 17589 8449 17601 8483
rect 17635 8480 17647 8483
rect 19076 8480 19104 8588
rect 19334 8576 19340 8628
rect 19392 8616 19398 8628
rect 19429 8619 19487 8625
rect 19429 8616 19441 8619
rect 19392 8588 19441 8616
rect 19392 8576 19398 8588
rect 19429 8585 19441 8588
rect 19475 8585 19487 8619
rect 19429 8579 19487 8585
rect 19705 8619 19763 8625
rect 19705 8585 19717 8619
rect 19751 8616 19763 8619
rect 20254 8616 20260 8628
rect 19751 8588 20260 8616
rect 19751 8585 19763 8588
rect 19705 8579 19763 8585
rect 19444 8548 19472 8579
rect 20254 8576 20260 8588
rect 20312 8576 20318 8628
rect 20622 8576 20628 8628
rect 20680 8616 20686 8628
rect 20901 8619 20959 8625
rect 20901 8616 20913 8619
rect 20680 8588 20913 8616
rect 20680 8576 20686 8588
rect 20901 8585 20913 8588
rect 20947 8585 20959 8619
rect 20901 8579 20959 8585
rect 19978 8548 19984 8560
rect 19444 8520 19984 8548
rect 19978 8508 19984 8520
rect 20036 8548 20042 8560
rect 20036 8520 20300 8548
rect 20036 8508 20042 8520
rect 20272 8489 20300 8520
rect 20165 8483 20223 8489
rect 20165 8480 20177 8483
rect 17635 8452 18184 8480
rect 19076 8452 20177 8480
rect 17635 8449 17647 8452
rect 17589 8443 17647 8449
rect 8772 8384 10916 8412
rect 11701 8415 11759 8421
rect 11701 8381 11713 8415
rect 11747 8412 11759 8415
rect 11974 8412 11980 8424
rect 11747 8384 11980 8412
rect 11747 8381 11759 8384
rect 11701 8375 11759 8381
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 12526 8372 12532 8424
rect 12584 8412 12590 8424
rect 15289 8415 15347 8421
rect 15289 8412 15301 8415
rect 12584 8384 15301 8412
rect 12584 8372 12590 8384
rect 15289 8381 15301 8384
rect 15335 8381 15347 8415
rect 15289 8375 15347 8381
rect 16209 8415 16267 8421
rect 16209 8381 16221 8415
rect 16255 8412 16267 8415
rect 16390 8412 16396 8424
rect 16255 8384 16396 8412
rect 16255 8381 16267 8384
rect 16209 8375 16267 8381
rect 16390 8372 16396 8384
rect 16448 8372 16454 8424
rect 16574 8372 16580 8424
rect 16632 8412 16638 8424
rect 17862 8412 17868 8424
rect 16632 8384 17868 8412
rect 16632 8372 16638 8384
rect 17862 8372 17868 8384
rect 17920 8412 17926 8424
rect 18056 8415 18114 8421
rect 18056 8412 18068 8415
rect 17920 8384 18068 8412
rect 17920 8372 17926 8384
rect 18056 8381 18068 8384
rect 18102 8381 18114 8415
rect 18156 8412 18184 8452
rect 20165 8449 20177 8452
rect 20211 8449 20223 8483
rect 20165 8443 20223 8449
rect 20257 8483 20315 8489
rect 20257 8449 20269 8483
rect 20303 8449 20315 8483
rect 20257 8443 20315 8449
rect 18156 8384 18276 8412
rect 18056 8375 18114 8381
rect 6288 8316 6776 8344
rect 5261 8279 5319 8285
rect 5261 8276 5273 8279
rect 4540 8248 5273 8276
rect 4249 8239 4307 8245
rect 5261 8245 5273 8248
rect 5307 8245 5319 8279
rect 5261 8239 5319 8245
rect 5350 8236 5356 8288
rect 5408 8276 5414 8288
rect 6288 8276 6316 8316
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 7561 8347 7619 8353
rect 7561 8344 7573 8347
rect 6972 8316 7573 8344
rect 6972 8304 6978 8316
rect 7561 8313 7573 8316
rect 7607 8313 7619 8347
rect 7561 8307 7619 8313
rect 7650 8304 7656 8356
rect 7708 8344 7714 8356
rect 8018 8344 8024 8356
rect 7708 8316 8024 8344
rect 7708 8304 7714 8316
rect 8018 8304 8024 8316
rect 8076 8304 8082 8356
rect 8113 8347 8171 8353
rect 8113 8313 8125 8347
rect 8159 8344 8171 8347
rect 8570 8344 8576 8356
rect 8159 8316 8576 8344
rect 8159 8313 8171 8316
rect 8113 8307 8171 8313
rect 8570 8304 8576 8316
rect 8628 8304 8634 8356
rect 8846 8304 8852 8356
rect 8904 8353 8910 8356
rect 8904 8347 8968 8353
rect 8904 8313 8922 8347
rect 8956 8313 8968 8347
rect 11790 8344 11796 8356
rect 11751 8316 11796 8344
rect 8904 8307 8968 8313
rect 8904 8304 8910 8307
rect 11790 8304 11796 8316
rect 11848 8304 11854 8356
rect 12704 8347 12762 8353
rect 12704 8313 12716 8347
rect 12750 8344 12762 8347
rect 15102 8344 15108 8356
rect 12750 8316 15108 8344
rect 12750 8313 12762 8316
rect 12704 8307 12762 8313
rect 15102 8304 15108 8316
rect 15160 8304 15166 8356
rect 15197 8347 15255 8353
rect 15197 8313 15209 8347
rect 15243 8344 15255 8347
rect 15243 8316 15884 8344
rect 15243 8313 15255 8316
rect 15197 8307 15255 8313
rect 5408 8248 6316 8276
rect 5408 8236 5414 8248
rect 8202 8236 8208 8288
rect 8260 8276 8266 8288
rect 9214 8276 9220 8288
rect 8260 8248 9220 8276
rect 8260 8236 8266 8248
rect 9214 8236 9220 8248
rect 9272 8236 9278 8288
rect 10318 8276 10324 8288
rect 10279 8248 10324 8276
rect 10318 8236 10324 8248
rect 10376 8236 10382 8288
rect 10686 8276 10692 8288
rect 10647 8248 10692 8276
rect 10686 8236 10692 8248
rect 10744 8236 10750 8288
rect 12894 8236 12900 8288
rect 12952 8276 12958 8288
rect 15856 8285 15884 8316
rect 16022 8304 16028 8356
rect 16080 8344 16086 8356
rect 16301 8347 16359 8353
rect 16301 8344 16313 8347
rect 16080 8316 16313 8344
rect 16080 8304 16086 8316
rect 16301 8313 16313 8316
rect 16347 8344 16359 8347
rect 16758 8344 16764 8356
rect 16347 8316 16764 8344
rect 16347 8313 16359 8316
rect 16301 8307 16359 8313
rect 16758 8304 16764 8316
rect 16816 8304 16822 8356
rect 17313 8347 17371 8353
rect 17313 8313 17325 8347
rect 17359 8344 17371 8347
rect 18138 8344 18144 8356
rect 17359 8316 18144 8344
rect 17359 8313 17371 8316
rect 17313 8307 17371 8313
rect 18138 8304 18144 8316
rect 18196 8304 18202 8356
rect 18248 8344 18276 8384
rect 19702 8372 19708 8424
rect 19760 8412 19766 8424
rect 20073 8415 20131 8421
rect 20073 8412 20085 8415
rect 19760 8384 20085 8412
rect 19760 8372 19766 8384
rect 20073 8381 20085 8384
rect 20119 8381 20131 8415
rect 20714 8412 20720 8424
rect 20675 8384 20720 8412
rect 20073 8375 20131 8381
rect 20714 8372 20720 8384
rect 20772 8372 20778 8424
rect 18316 8347 18374 8353
rect 18316 8344 18328 8347
rect 18248 8316 18328 8344
rect 18248 8288 18276 8316
rect 18316 8313 18328 8316
rect 18362 8344 18374 8347
rect 20346 8344 20352 8356
rect 18362 8316 20352 8344
rect 18362 8313 18374 8316
rect 18316 8307 18374 8313
rect 20346 8304 20352 8316
rect 20404 8304 20410 8356
rect 13817 8279 13875 8285
rect 13817 8276 13829 8279
rect 12952 8248 13829 8276
rect 12952 8236 12958 8248
rect 13817 8245 13829 8248
rect 13863 8245 13875 8279
rect 13817 8239 13875 8245
rect 15841 8279 15899 8285
rect 15841 8245 15853 8279
rect 15887 8245 15899 8279
rect 17402 8276 17408 8288
rect 17363 8248 17408 8276
rect 15841 8239 15899 8245
rect 17402 8236 17408 8248
rect 17460 8236 17466 8288
rect 18230 8236 18236 8288
rect 18288 8236 18294 8288
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 3602 8032 3608 8084
rect 3660 8072 3666 8084
rect 4065 8075 4123 8081
rect 4065 8072 4077 8075
rect 3660 8044 4077 8072
rect 3660 8032 3666 8044
rect 4065 8041 4077 8044
rect 4111 8041 4123 8075
rect 4065 8035 4123 8041
rect 4246 8032 4252 8084
rect 4304 8072 4310 8084
rect 4525 8075 4583 8081
rect 4525 8072 4537 8075
rect 4304 8044 4537 8072
rect 4304 8032 4310 8044
rect 4525 8041 4537 8044
rect 4571 8041 4583 8075
rect 4525 8035 4583 8041
rect 5629 8075 5687 8081
rect 5629 8041 5641 8075
rect 5675 8072 5687 8075
rect 6914 8072 6920 8084
rect 5675 8044 6920 8072
rect 5675 8041 5687 8044
rect 5629 8035 5687 8041
rect 6914 8032 6920 8044
rect 6972 8032 6978 8084
rect 7098 8072 7104 8084
rect 7059 8044 7104 8072
rect 7098 8032 7104 8044
rect 7156 8032 7162 8084
rect 7745 8075 7803 8081
rect 7745 8041 7757 8075
rect 7791 8072 7803 8075
rect 8662 8072 8668 8084
rect 7791 8044 8668 8072
rect 7791 8041 7803 8044
rect 7745 8035 7803 8041
rect 8662 8032 8668 8044
rect 8720 8032 8726 8084
rect 9214 8072 9220 8084
rect 9175 8044 9220 8072
rect 9214 8032 9220 8044
rect 9272 8032 9278 8084
rect 10413 8075 10471 8081
rect 10413 8041 10425 8075
rect 10459 8072 10471 8075
rect 10686 8072 10692 8084
rect 10459 8044 10692 8072
rect 10459 8041 10471 8044
rect 10413 8035 10471 8041
rect 10686 8032 10692 8044
rect 10744 8032 10750 8084
rect 10873 8075 10931 8081
rect 10873 8041 10885 8075
rect 10919 8072 10931 8075
rect 12158 8072 12164 8084
rect 10919 8044 12164 8072
rect 10919 8041 10931 8044
rect 10873 8035 10931 8041
rect 12158 8032 12164 8044
rect 12216 8072 12222 8084
rect 12345 8075 12403 8081
rect 12216 8044 12296 8072
rect 12216 8032 12222 8044
rect 3142 8004 3148 8016
rect 2332 7976 3148 8004
rect 1578 7828 1584 7880
rect 1636 7868 1642 7880
rect 2332 7877 2360 7976
rect 3142 7964 3148 7976
rect 3200 7964 3206 8016
rect 3970 7964 3976 8016
rect 4028 8004 4034 8016
rect 12268 8004 12296 8044
rect 12345 8041 12357 8075
rect 12391 8072 12403 8075
rect 12618 8072 12624 8084
rect 12391 8044 12624 8072
rect 12391 8041 12403 8044
rect 12345 8035 12403 8041
rect 12618 8032 12624 8044
rect 12676 8032 12682 8084
rect 12713 8075 12771 8081
rect 12713 8041 12725 8075
rect 12759 8072 12771 8075
rect 12986 8072 12992 8084
rect 12759 8044 12992 8072
rect 12759 8041 12771 8044
rect 12713 8035 12771 8041
rect 12986 8032 12992 8044
rect 13044 8032 13050 8084
rect 18138 8032 18144 8084
rect 18196 8072 18202 8084
rect 18417 8075 18475 8081
rect 18417 8072 18429 8075
rect 18196 8044 18429 8072
rect 18196 8032 18202 8044
rect 18417 8041 18429 8044
rect 18463 8041 18475 8075
rect 19426 8072 19432 8084
rect 19387 8044 19432 8072
rect 18417 8035 18475 8041
rect 19426 8032 19432 8044
rect 19484 8032 19490 8084
rect 19797 8075 19855 8081
rect 19797 8041 19809 8075
rect 19843 8072 19855 8075
rect 19886 8072 19892 8084
rect 19843 8044 19892 8072
rect 19843 8041 19855 8044
rect 19797 8035 19855 8041
rect 19886 8032 19892 8044
rect 19944 8032 19950 8084
rect 12805 8007 12863 8013
rect 12805 8004 12817 8007
rect 4028 7976 10916 8004
rect 12268 7976 12817 8004
rect 4028 7964 4034 7976
rect 2584 7939 2642 7945
rect 2584 7905 2596 7939
rect 2630 7936 2642 7939
rect 3602 7936 3608 7948
rect 2630 7908 3608 7936
rect 2630 7905 2642 7908
rect 2584 7899 2642 7905
rect 3602 7896 3608 7908
rect 3660 7936 3666 7948
rect 4433 7939 4491 7945
rect 3660 7908 4384 7936
rect 3660 7896 3666 7908
rect 2317 7871 2375 7877
rect 2317 7868 2329 7871
rect 1636 7840 2329 7868
rect 1636 7828 1642 7840
rect 2317 7837 2329 7840
rect 2363 7837 2375 7871
rect 2317 7831 2375 7837
rect 3697 7803 3755 7809
rect 3697 7769 3709 7803
rect 3743 7800 3755 7803
rect 3786 7800 3792 7812
rect 3743 7772 3792 7800
rect 3743 7769 3755 7772
rect 3697 7763 3755 7769
rect 3786 7760 3792 7772
rect 3844 7760 3850 7812
rect 4356 7800 4384 7908
rect 4433 7905 4445 7939
rect 4479 7936 4491 7939
rect 4982 7936 4988 7948
rect 4479 7908 4988 7936
rect 4479 7905 4491 7908
rect 4433 7899 4491 7905
rect 4982 7896 4988 7908
rect 5040 7936 5046 7948
rect 5442 7936 5448 7948
rect 5040 7908 5448 7936
rect 5040 7896 5046 7908
rect 5442 7896 5448 7908
rect 5500 7896 5506 7948
rect 5988 7939 6046 7945
rect 5988 7905 6000 7939
rect 6034 7936 6046 7939
rect 6362 7936 6368 7948
rect 6034 7908 6368 7936
rect 6034 7905 6046 7908
rect 5988 7899 6046 7905
rect 6362 7896 6368 7908
rect 6420 7896 6426 7948
rect 8110 7945 8116 7948
rect 8104 7899 8116 7945
rect 8168 7936 8174 7948
rect 8168 7908 8204 7936
rect 8110 7896 8116 7899
rect 8168 7896 8174 7908
rect 10410 7896 10416 7948
rect 10468 7936 10474 7948
rect 10781 7939 10839 7945
rect 10781 7936 10793 7939
rect 10468 7908 10793 7936
rect 10468 7896 10474 7908
rect 10781 7905 10793 7908
rect 10827 7905 10839 7939
rect 10888 7936 10916 7976
rect 12805 7973 12817 7976
rect 12851 7973 12863 8007
rect 12805 7967 12863 7973
rect 15562 7936 15568 7948
rect 10888 7908 15568 7936
rect 10781 7899 10839 7905
rect 15562 7896 15568 7908
rect 15620 7896 15626 7948
rect 17028 7939 17086 7945
rect 17028 7905 17040 7939
rect 17074 7936 17086 7939
rect 17954 7936 17960 7948
rect 17074 7908 17960 7936
rect 17074 7905 17086 7908
rect 17028 7899 17086 7905
rect 17954 7896 17960 7908
rect 18012 7896 18018 7948
rect 18782 7936 18788 7948
rect 18743 7908 18788 7936
rect 18782 7896 18788 7908
rect 18840 7896 18846 7948
rect 18874 7896 18880 7948
rect 18932 7936 18938 7948
rect 18932 7908 18977 7936
rect 18932 7896 18938 7908
rect 4706 7868 4712 7880
rect 4619 7840 4712 7868
rect 4706 7828 4712 7840
rect 4764 7868 4770 7880
rect 5629 7871 5687 7877
rect 5629 7868 5641 7871
rect 4764 7840 5641 7868
rect 4764 7828 4770 7840
rect 5629 7837 5641 7840
rect 5675 7837 5687 7871
rect 5629 7831 5687 7837
rect 5721 7871 5779 7877
rect 5721 7837 5733 7871
rect 5767 7837 5779 7871
rect 5721 7831 5779 7837
rect 4724 7800 4752 7828
rect 4356 7772 4752 7800
rect 5258 7760 5264 7812
rect 5316 7800 5322 7812
rect 5736 7800 5764 7831
rect 6914 7828 6920 7880
rect 6972 7868 6978 7880
rect 7745 7871 7803 7877
rect 7745 7868 7757 7871
rect 6972 7840 7757 7868
rect 6972 7828 6978 7840
rect 7745 7837 7757 7840
rect 7791 7868 7803 7871
rect 7837 7871 7895 7877
rect 7837 7868 7849 7871
rect 7791 7840 7849 7868
rect 7791 7837 7803 7840
rect 7745 7831 7803 7837
rect 7837 7837 7849 7840
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 8846 7828 8852 7880
rect 8904 7868 8910 7880
rect 10962 7868 10968 7880
rect 8904 7840 10968 7868
rect 8904 7828 8910 7840
rect 10962 7828 10968 7840
rect 11020 7868 11026 7880
rect 12894 7868 12900 7880
rect 11020 7840 11113 7868
rect 12855 7840 12900 7868
rect 11020 7828 11026 7840
rect 12894 7828 12900 7840
rect 12952 7828 12958 7880
rect 16574 7828 16580 7880
rect 16632 7868 16638 7880
rect 16761 7871 16819 7877
rect 16761 7868 16773 7871
rect 16632 7840 16773 7868
rect 16632 7828 16638 7840
rect 16761 7837 16773 7840
rect 16807 7837 16819 7871
rect 18966 7868 18972 7880
rect 18927 7840 18972 7868
rect 16761 7831 16819 7837
rect 18966 7828 18972 7840
rect 19024 7828 19030 7880
rect 19886 7868 19892 7880
rect 19847 7840 19892 7868
rect 19886 7828 19892 7840
rect 19944 7828 19950 7880
rect 19978 7828 19984 7880
rect 20036 7868 20042 7880
rect 20036 7840 20081 7868
rect 20036 7828 20042 7840
rect 5316 7772 5764 7800
rect 18141 7803 18199 7809
rect 5316 7760 5322 7772
rect 18141 7769 18153 7803
rect 18187 7800 18199 7803
rect 18230 7800 18236 7812
rect 18187 7772 18236 7800
rect 18187 7769 18199 7772
rect 18141 7763 18199 7769
rect 18230 7760 18236 7772
rect 18288 7760 18294 7812
rect 4062 7692 4068 7744
rect 4120 7732 4126 7744
rect 15194 7732 15200 7744
rect 4120 7704 15200 7732
rect 4120 7692 4126 7704
rect 15194 7692 15200 7704
rect 15252 7692 15258 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 2501 7531 2559 7537
rect 2501 7497 2513 7531
rect 2547 7528 2559 7531
rect 2590 7528 2596 7540
rect 2547 7500 2596 7528
rect 2547 7497 2559 7500
rect 2501 7491 2559 7497
rect 2590 7488 2596 7500
rect 2648 7488 2654 7540
rect 3142 7488 3148 7540
rect 3200 7488 3206 7540
rect 5258 7528 5264 7540
rect 5000 7500 5264 7528
rect 3160 7460 3188 7488
rect 5000 7460 5028 7500
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 6362 7528 6368 7540
rect 6323 7500 6368 7528
rect 6362 7488 6368 7500
rect 6420 7488 6426 7540
rect 8110 7488 8116 7540
rect 8168 7528 8174 7540
rect 8297 7531 8355 7537
rect 8297 7528 8309 7531
rect 8168 7500 8309 7528
rect 8168 7488 8174 7500
rect 8297 7497 8309 7500
rect 8343 7497 8355 7531
rect 8570 7528 8576 7540
rect 8531 7500 8576 7528
rect 8297 7491 8355 7497
rect 3160 7432 5028 7460
rect 3145 7395 3203 7401
rect 3145 7361 3157 7395
rect 3191 7392 3203 7395
rect 3786 7392 3792 7404
rect 3191 7364 3792 7392
rect 3191 7361 3203 7364
rect 3145 7355 3203 7361
rect 3786 7352 3792 7364
rect 3844 7352 3850 7404
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7392 4215 7395
rect 4706 7392 4712 7404
rect 4203 7364 4712 7392
rect 4203 7361 4215 7364
rect 4157 7355 4215 7361
rect 4706 7352 4712 7364
rect 4764 7352 4770 7404
rect 5000 7401 5028 7432
rect 4985 7395 5043 7401
rect 4985 7361 4997 7395
rect 5031 7361 5043 7395
rect 6914 7392 6920 7404
rect 6875 7364 6920 7392
rect 4985 7355 5043 7361
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 8312 7392 8340 7491
rect 8570 7488 8576 7500
rect 8628 7488 8634 7540
rect 16301 7531 16359 7537
rect 16301 7497 16313 7531
rect 16347 7528 16359 7531
rect 17402 7528 17408 7540
rect 16347 7500 17408 7528
rect 16347 7497 16359 7500
rect 16301 7491 16359 7497
rect 17402 7488 17408 7500
rect 17460 7488 17466 7540
rect 19797 7531 19855 7537
rect 19797 7497 19809 7531
rect 19843 7528 19855 7531
rect 19886 7528 19892 7540
rect 19843 7500 19892 7528
rect 19843 7497 19855 7500
rect 19797 7491 19855 7497
rect 19886 7488 19892 7500
rect 19944 7488 19950 7540
rect 11698 7420 11704 7472
rect 11756 7460 11762 7472
rect 11756 7432 20208 7460
rect 11756 7420 11762 7432
rect 9125 7395 9183 7401
rect 9125 7392 9137 7395
rect 8312 7364 9137 7392
rect 9125 7361 9137 7364
rect 9171 7361 9183 7395
rect 9125 7355 9183 7361
rect 16945 7395 17003 7401
rect 16945 7361 16957 7395
rect 16991 7392 17003 7395
rect 17954 7392 17960 7404
rect 16991 7364 17960 7392
rect 16991 7361 17003 7364
rect 16945 7355 17003 7361
rect 17954 7352 17960 7364
rect 18012 7352 18018 7404
rect 5258 7333 5264 7336
rect 5252 7324 5264 7333
rect 5219 7296 5264 7324
rect 5252 7287 5264 7296
rect 5258 7284 5264 7287
rect 5316 7284 5322 7336
rect 9030 7284 9036 7336
rect 9088 7324 9094 7336
rect 16761 7327 16819 7333
rect 16761 7324 16773 7327
rect 9088 7296 16773 7324
rect 9088 7284 9094 7296
rect 16761 7293 16773 7296
rect 16807 7293 16819 7327
rect 16761 7287 16819 7293
rect 19061 7327 19119 7333
rect 19061 7293 19073 7327
rect 19107 7324 19119 7327
rect 19794 7324 19800 7336
rect 19107 7296 19800 7324
rect 19107 7293 19119 7296
rect 19061 7287 19119 7293
rect 19794 7284 19800 7296
rect 19852 7284 19858 7336
rect 20180 7333 20208 7432
rect 20346 7392 20352 7404
rect 20307 7364 20352 7392
rect 20346 7352 20352 7364
rect 20404 7352 20410 7404
rect 20165 7327 20223 7333
rect 20165 7293 20177 7327
rect 20211 7293 20223 7327
rect 20165 7287 20223 7293
rect 2869 7259 2927 7265
rect 2869 7225 2881 7259
rect 2915 7256 2927 7259
rect 2915 7228 3556 7256
rect 2915 7225 2927 7228
rect 2869 7219 2927 7225
rect 2958 7188 2964 7200
rect 2919 7160 2964 7188
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 3528 7197 3556 7228
rect 3786 7216 3792 7268
rect 3844 7256 3850 7268
rect 3973 7259 4031 7265
rect 3973 7256 3985 7259
rect 3844 7228 3985 7256
rect 3844 7216 3850 7228
rect 3973 7225 3985 7228
rect 4019 7256 4031 7259
rect 4154 7256 4160 7268
rect 4019 7228 4160 7256
rect 4019 7225 4031 7228
rect 3973 7219 4031 7225
rect 4154 7216 4160 7228
rect 4212 7216 4218 7268
rect 7098 7216 7104 7268
rect 7156 7265 7162 7268
rect 7156 7259 7220 7265
rect 7156 7225 7174 7259
rect 7208 7225 7220 7259
rect 7156 7219 7220 7225
rect 8941 7259 8999 7265
rect 8941 7225 8953 7259
rect 8987 7256 8999 7259
rect 8987 7228 11100 7256
rect 8987 7225 8999 7228
rect 8941 7219 8999 7225
rect 7156 7216 7162 7219
rect 11072 7200 11100 7228
rect 11606 7216 11612 7268
rect 11664 7256 11670 7268
rect 19337 7259 19395 7265
rect 19337 7256 19349 7259
rect 11664 7228 19349 7256
rect 11664 7216 11670 7228
rect 19337 7225 19349 7228
rect 19383 7225 19395 7259
rect 19337 7219 19395 7225
rect 3513 7191 3571 7197
rect 3513 7157 3525 7191
rect 3559 7157 3571 7191
rect 3878 7188 3884 7200
rect 3839 7160 3884 7188
rect 3513 7151 3571 7157
rect 3878 7148 3884 7160
rect 3936 7148 3942 7200
rect 4525 7191 4583 7197
rect 4525 7157 4537 7191
rect 4571 7188 4583 7191
rect 5350 7188 5356 7200
rect 4571 7160 5356 7188
rect 4571 7157 4583 7160
rect 4525 7151 4583 7157
rect 5350 7148 5356 7160
rect 5408 7148 5414 7200
rect 9030 7188 9036 7200
rect 8991 7160 9036 7188
rect 9030 7148 9036 7160
rect 9088 7148 9094 7200
rect 11054 7148 11060 7200
rect 11112 7188 11118 7200
rect 16669 7191 16727 7197
rect 16669 7188 16681 7191
rect 11112 7160 16681 7188
rect 11112 7148 11118 7160
rect 16669 7157 16681 7160
rect 16715 7157 16727 7191
rect 16669 7151 16727 7157
rect 20162 7148 20168 7200
rect 20220 7188 20226 7200
rect 20257 7191 20315 7197
rect 20257 7188 20269 7191
rect 20220 7160 20269 7188
rect 20220 7148 20226 7160
rect 20257 7157 20269 7160
rect 20303 7188 20315 7191
rect 20438 7188 20444 7200
rect 20303 7160 20444 7188
rect 20303 7157 20315 7160
rect 20257 7151 20315 7157
rect 20438 7148 20444 7160
rect 20496 7148 20502 7200
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 3329 6987 3387 6993
rect 3329 6953 3341 6987
rect 3375 6984 3387 6987
rect 3878 6984 3884 6996
rect 3375 6956 3884 6984
rect 3375 6953 3387 6956
rect 3329 6947 3387 6953
rect 3878 6944 3884 6956
rect 3936 6944 3942 6996
rect 5534 6984 5540 6996
rect 4540 6956 5540 6984
rect 1578 6848 1584 6860
rect 1539 6820 1584 6848
rect 1578 6808 1584 6820
rect 1636 6808 1642 6860
rect 1848 6851 1906 6857
rect 1848 6817 1860 6851
rect 1894 6848 1906 6851
rect 2222 6848 2228 6860
rect 1894 6820 2228 6848
rect 1894 6817 1906 6820
rect 1848 6811 1906 6817
rect 2222 6808 2228 6820
rect 2280 6808 2286 6860
rect 3142 6808 3148 6860
rect 3200 6848 3206 6860
rect 4540 6857 4568 6956
rect 5534 6944 5540 6956
rect 5592 6944 5598 6996
rect 6546 6984 6552 6996
rect 6507 6956 6552 6984
rect 6546 6944 6552 6956
rect 6604 6944 6610 6996
rect 17954 6984 17960 6996
rect 17867 6956 17960 6984
rect 17954 6944 17960 6956
rect 18012 6984 18018 6996
rect 18966 6984 18972 6996
rect 18012 6956 18972 6984
rect 18012 6944 18018 6956
rect 18966 6944 18972 6956
rect 19024 6944 19030 6996
rect 5810 6876 5816 6928
rect 5868 6916 5874 6928
rect 6822 6916 6828 6928
rect 5868 6888 6828 6916
rect 5868 6876 5874 6888
rect 6822 6876 6828 6888
rect 6880 6916 6886 6928
rect 7561 6919 7619 6925
rect 7561 6916 7573 6919
rect 6880 6888 7573 6916
rect 6880 6876 6886 6888
rect 7561 6885 7573 6888
rect 7607 6885 7619 6919
rect 7561 6879 7619 6885
rect 10410 6876 10416 6928
rect 10468 6916 10474 6928
rect 18506 6916 18512 6928
rect 10468 6888 18512 6916
rect 10468 6876 10474 6888
rect 18506 6876 18512 6888
rect 18564 6876 18570 6928
rect 4525 6851 4583 6857
rect 4525 6848 4537 6851
rect 3200 6820 4537 6848
rect 3200 6808 3206 6820
rect 4525 6817 4537 6820
rect 4571 6817 4583 6851
rect 5534 6848 5540 6860
rect 5495 6820 5540 6848
rect 4525 6811 4583 6817
rect 5534 6808 5540 6820
rect 5592 6808 5598 6860
rect 6641 6851 6699 6857
rect 6641 6817 6653 6851
rect 6687 6848 6699 6851
rect 7653 6851 7711 6857
rect 6687 6820 6868 6848
rect 6687 6817 6699 6820
rect 6641 6811 6699 6817
rect 4246 6740 4252 6792
rect 4304 6780 4310 6792
rect 4617 6783 4675 6789
rect 4617 6780 4629 6783
rect 4304 6752 4629 6780
rect 4304 6740 4310 6752
rect 4617 6749 4629 6752
rect 4663 6749 4675 6783
rect 4617 6743 4675 6749
rect 4801 6783 4859 6789
rect 4801 6749 4813 6783
rect 4847 6780 4859 6783
rect 5258 6780 5264 6792
rect 4847 6752 5264 6780
rect 4847 6749 4859 6752
rect 4801 6743 4859 6749
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 5629 6783 5687 6789
rect 5629 6749 5641 6783
rect 5675 6749 5687 6783
rect 5629 6743 5687 6749
rect 5813 6783 5871 6789
rect 5813 6749 5825 6783
rect 5859 6780 5871 6783
rect 6362 6780 6368 6792
rect 5859 6752 6368 6780
rect 5859 6749 5871 6752
rect 5813 6743 5871 6749
rect 2774 6672 2780 6724
rect 2832 6712 2838 6724
rect 2961 6715 3019 6721
rect 2961 6712 2973 6715
rect 2832 6684 2973 6712
rect 2832 6672 2838 6684
rect 2961 6681 2973 6684
rect 3007 6681 3019 6715
rect 2961 6675 3019 6681
rect 4157 6715 4215 6721
rect 4157 6681 4169 6715
rect 4203 6712 4215 6715
rect 5644 6712 5672 6743
rect 6362 6740 6368 6752
rect 6420 6740 6426 6792
rect 6733 6783 6791 6789
rect 6733 6749 6745 6783
rect 6779 6749 6791 6783
rect 6733 6743 6791 6749
rect 6178 6712 6184 6724
rect 4203 6684 5672 6712
rect 6139 6684 6184 6712
rect 4203 6681 4215 6684
rect 4157 6675 4215 6681
rect 6178 6672 6184 6684
rect 6236 6672 6242 6724
rect 6380 6712 6408 6740
rect 6748 6712 6776 6743
rect 6380 6684 6776 6712
rect 6840 6712 6868 6820
rect 7653 6817 7665 6851
rect 7699 6848 7711 6851
rect 12066 6848 12072 6860
rect 7699 6820 12072 6848
rect 7699 6817 7711 6820
rect 7653 6811 7711 6817
rect 12066 6808 12072 6820
rect 12124 6808 12130 6860
rect 16844 6851 16902 6857
rect 16844 6817 16856 6851
rect 16890 6848 16902 6851
rect 19150 6848 19156 6860
rect 16890 6820 19156 6848
rect 16890 6817 16902 6820
rect 16844 6811 16902 6817
rect 19150 6808 19156 6820
rect 19208 6808 19214 6860
rect 19328 6851 19386 6857
rect 19328 6817 19340 6851
rect 19374 6848 19386 6851
rect 19610 6848 19616 6860
rect 19374 6820 19616 6848
rect 19374 6817 19386 6820
rect 19328 6811 19386 6817
rect 19610 6808 19616 6820
rect 19668 6808 19674 6860
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6780 7895 6783
rect 8846 6780 8852 6792
rect 7883 6752 8852 6780
rect 7883 6749 7895 6752
rect 7837 6743 7895 6749
rect 8846 6740 8852 6752
rect 8904 6740 8910 6792
rect 16574 6780 16580 6792
rect 16535 6752 16580 6780
rect 16574 6740 16580 6752
rect 16632 6740 16638 6792
rect 19058 6780 19064 6792
rect 19019 6752 19064 6780
rect 19058 6740 19064 6752
rect 19116 6740 19122 6792
rect 20162 6740 20168 6792
rect 20220 6780 20226 6792
rect 20901 6783 20959 6789
rect 20901 6780 20913 6783
rect 20220 6752 20913 6780
rect 20220 6740 20226 6752
rect 20901 6749 20913 6752
rect 20947 6749 20959 6783
rect 20901 6743 20959 6749
rect 10318 6712 10324 6724
rect 6840 6684 10324 6712
rect 10318 6672 10324 6684
rect 10376 6672 10382 6724
rect 5166 6644 5172 6656
rect 5127 6616 5172 6644
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 7190 6644 7196 6656
rect 7151 6616 7196 6644
rect 7190 6604 7196 6616
rect 7248 6604 7254 6656
rect 7374 6604 7380 6656
rect 7432 6644 7438 6656
rect 17954 6644 17960 6656
rect 7432 6616 17960 6644
rect 7432 6604 7438 6616
rect 17954 6604 17960 6616
rect 18012 6604 18018 6656
rect 20441 6647 20499 6653
rect 20441 6613 20453 6647
rect 20487 6644 20499 6647
rect 20622 6644 20628 6656
rect 20487 6616 20628 6644
rect 20487 6613 20499 6616
rect 20441 6607 20499 6613
rect 20622 6604 20628 6616
rect 20680 6604 20686 6656
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 2958 6440 2964 6452
rect 2919 6412 2964 6440
rect 2958 6400 2964 6412
rect 3016 6400 3022 6452
rect 4985 6443 5043 6449
rect 4985 6409 4997 6443
rect 5031 6440 5043 6443
rect 5534 6440 5540 6452
rect 5031 6412 5540 6440
rect 5031 6409 5043 6412
rect 4985 6403 5043 6409
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 19150 6400 19156 6452
rect 19208 6440 19214 6452
rect 20346 6440 20352 6452
rect 19208 6412 20352 6440
rect 19208 6400 19214 6412
rect 20346 6400 20352 6412
rect 20404 6440 20410 6452
rect 20625 6443 20683 6449
rect 20625 6440 20637 6443
rect 20404 6412 20637 6440
rect 20404 6400 20410 6412
rect 20625 6409 20637 6412
rect 20671 6409 20683 6443
rect 20625 6403 20683 6409
rect 4062 6332 4068 6384
rect 4120 6372 4126 6384
rect 7006 6372 7012 6384
rect 4120 6344 7012 6372
rect 4120 6332 4126 6344
rect 7006 6332 7012 6344
rect 7064 6332 7070 6384
rect 3602 6304 3608 6316
rect 3563 6276 3608 6304
rect 3602 6264 3608 6276
rect 3660 6264 3666 6316
rect 5258 6264 5264 6316
rect 5316 6304 5322 6316
rect 5537 6307 5595 6313
rect 5537 6304 5549 6307
rect 5316 6276 5549 6304
rect 5316 6264 5322 6276
rect 5537 6273 5549 6276
rect 5583 6273 5595 6307
rect 5537 6267 5595 6273
rect 16574 6264 16580 6316
rect 16632 6304 16638 6316
rect 19058 6304 19064 6316
rect 16632 6276 19064 6304
rect 16632 6264 16638 6276
rect 19058 6264 19064 6276
rect 19116 6304 19122 6316
rect 19245 6307 19303 6313
rect 19245 6304 19257 6307
rect 19116 6276 19257 6304
rect 19116 6264 19122 6276
rect 19245 6273 19257 6276
rect 19291 6273 19303 6307
rect 19245 6267 19303 6273
rect 3970 6196 3976 6248
rect 4028 6236 4034 6248
rect 5350 6236 5356 6248
rect 4028 6208 4936 6236
rect 5311 6208 5356 6236
rect 4028 6196 4034 6208
rect 2866 6128 2872 6180
rect 2924 6168 2930 6180
rect 3418 6168 3424 6180
rect 2924 6140 3424 6168
rect 2924 6128 2930 6140
rect 3418 6128 3424 6140
rect 3476 6128 3482 6180
rect 4798 6168 4804 6180
rect 3620 6140 4804 6168
rect 3234 6060 3240 6112
rect 3292 6100 3298 6112
rect 3329 6103 3387 6109
rect 3329 6100 3341 6103
rect 3292 6072 3341 6100
rect 3292 6060 3298 6072
rect 3329 6069 3341 6072
rect 3375 6100 3387 6103
rect 3620 6100 3648 6140
rect 4798 6128 4804 6140
rect 4856 6128 4862 6180
rect 4908 6168 4936 6208
rect 5350 6196 5356 6208
rect 5408 6196 5414 6248
rect 19512 6239 19570 6245
rect 19512 6205 19524 6239
rect 19558 6236 19570 6239
rect 20622 6236 20628 6248
rect 19558 6208 20628 6236
rect 19558 6205 19570 6208
rect 19512 6199 19570 6205
rect 20622 6196 20628 6208
rect 20680 6196 20686 6248
rect 10226 6168 10232 6180
rect 4908 6140 10232 6168
rect 10226 6128 10232 6140
rect 10284 6128 10290 6180
rect 3375 6072 3648 6100
rect 3375 6069 3387 6072
rect 3329 6063 3387 6069
rect 3694 6060 3700 6112
rect 3752 6100 3758 6112
rect 3970 6100 3976 6112
rect 3752 6072 3976 6100
rect 3752 6060 3758 6072
rect 3970 6060 3976 6072
rect 4028 6100 4034 6112
rect 5445 6103 5503 6109
rect 5445 6100 5457 6103
rect 4028 6072 5457 6100
rect 4028 6060 4034 6072
rect 5445 6069 5457 6072
rect 5491 6069 5503 6103
rect 5445 6063 5503 6069
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 19794 5896 19800 5908
rect 19755 5868 19800 5896
rect 19794 5856 19800 5868
rect 19852 5856 19858 5908
rect 20162 5896 20168 5908
rect 20123 5868 20168 5896
rect 20162 5856 20168 5868
rect 20220 5856 20226 5908
rect 20254 5692 20260 5704
rect 20215 5664 20260 5692
rect 20254 5652 20260 5664
rect 20312 5652 20318 5704
rect 20346 5652 20352 5704
rect 20404 5692 20410 5704
rect 20404 5664 20449 5692
rect 20404 5652 20410 5664
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 6086 5312 6092 5364
rect 6144 5352 6150 5364
rect 17954 5352 17960 5364
rect 6144 5324 17960 5352
rect 6144 5312 6150 5324
rect 17954 5312 17960 5324
rect 18012 5312 18018 5364
rect 20073 5355 20131 5361
rect 20073 5321 20085 5355
rect 20119 5352 20131 5355
rect 20254 5352 20260 5364
rect 20119 5324 20260 5352
rect 20119 5321 20131 5324
rect 20073 5315 20131 5321
rect 20254 5312 20260 5324
rect 20312 5312 20318 5364
rect 4062 5244 4068 5296
rect 4120 5284 4126 5296
rect 11698 5284 11704 5296
rect 4120 5256 11704 5284
rect 4120 5244 4126 5256
rect 11698 5244 11704 5256
rect 11756 5244 11762 5296
rect 20622 5216 20628 5228
rect 20583 5188 20628 5216
rect 20622 5176 20628 5188
rect 20680 5176 20686 5228
rect 4062 4972 4068 5024
rect 4120 5012 4126 5024
rect 19889 5015 19947 5021
rect 19889 5012 19901 5015
rect 4120 4984 19901 5012
rect 4120 4972 4126 4984
rect 19889 4981 19901 4984
rect 19935 5012 19947 5015
rect 20441 5015 20499 5021
rect 20441 5012 20453 5015
rect 19935 4984 20453 5012
rect 19935 4981 19947 4984
rect 19889 4975 19947 4981
rect 20441 4981 20453 4984
rect 20487 4981 20499 5015
rect 20441 4975 20499 4981
rect 20530 4972 20536 5024
rect 20588 5012 20594 5024
rect 20588 4984 20633 5012
rect 20588 4972 20594 4984
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 14476 3080 15424 3108
rect 14476 3040 14504 3080
rect 4632 3012 14504 3040
rect 15013 3043 15071 3049
rect 4632 2981 4660 3012
rect 15013 3009 15025 3043
rect 15059 3040 15071 3043
rect 15289 3043 15347 3049
rect 15289 3040 15301 3043
rect 15059 3012 15301 3040
rect 15059 3009 15071 3012
rect 15013 3003 15071 3009
rect 15289 3009 15301 3012
rect 15335 3009 15347 3043
rect 15396 3040 15424 3080
rect 20438 3040 20444 3052
rect 15396 3012 20444 3040
rect 15289 3003 15347 3009
rect 20438 3000 20444 3012
rect 20496 3000 20502 3052
rect 4617 2975 4675 2981
rect 4617 2941 4629 2975
rect 4663 2941 4675 2975
rect 4890 2972 4896 2984
rect 4851 2944 4896 2972
rect 4617 2935 4675 2941
rect 4890 2932 4896 2944
rect 4948 2932 4954 2984
rect 5537 2975 5595 2981
rect 5537 2941 5549 2975
rect 5583 2972 5595 2975
rect 11146 2972 11152 2984
rect 5583 2944 11152 2972
rect 5583 2941 5595 2944
rect 5537 2935 5595 2941
rect 11146 2932 11152 2944
rect 11204 2932 11210 2984
rect 15105 2975 15163 2981
rect 15105 2941 15117 2975
rect 15151 2972 15163 2975
rect 15838 2972 15844 2984
rect 15151 2944 15844 2972
rect 15151 2941 15163 2944
rect 15105 2935 15163 2941
rect 15838 2932 15844 2944
rect 15896 2932 15902 2984
rect 5718 2864 5724 2916
rect 5776 2904 5782 2916
rect 5813 2907 5871 2913
rect 5813 2904 5825 2907
rect 5776 2876 5825 2904
rect 5776 2864 5782 2876
rect 5813 2873 5825 2876
rect 5859 2873 5871 2907
rect 5813 2867 5871 2873
rect 5074 2796 5080 2848
rect 5132 2836 5138 2848
rect 15013 2839 15071 2845
rect 15013 2836 15025 2839
rect 5132 2808 15025 2836
rect 5132 2796 5138 2808
rect 15013 2805 15025 2808
rect 15059 2805 15071 2839
rect 15013 2799 15071 2805
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 2958 1300 2964 1352
rect 3016 1340 3022 1352
rect 5902 1340 5908 1352
rect 3016 1312 5908 1340
rect 3016 1300 3022 1312
rect 5902 1300 5908 1312
rect 5960 1300 5966 1352
rect 2774 1028 2780 1080
rect 2832 1068 2838 1080
rect 4982 1068 4988 1080
rect 2832 1040 4988 1068
rect 2832 1028 2838 1040
rect 4982 1028 4988 1040
rect 5040 1028 5046 1080
rect 3326 212 3332 264
rect 3384 252 3390 264
rect 6822 252 6828 264
rect 3384 224 6828 252
rect 3384 212 3390 224
rect 6822 212 6828 224
rect 6880 212 6886 264
<< via1 >>
rect 3884 20952 3936 21004
rect 5540 20952 5592 21004
rect 2228 20612 2280 20664
rect 8668 20612 8720 20664
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 2780 20000 2832 20052
rect 8668 20043 8720 20052
rect 8668 20009 8677 20043
rect 8677 20009 8711 20043
rect 8711 20009 8720 20043
rect 8668 20000 8720 20009
rect 10232 20000 10284 20052
rect 11612 20000 11664 20052
rect 12256 20000 12308 20052
rect 16672 20000 16724 20052
rect 17500 20000 17552 20052
rect 19616 20043 19668 20052
rect 19616 20009 19625 20043
rect 19625 20009 19659 20043
rect 19659 20009 19668 20043
rect 19616 20000 19668 20009
rect 20168 20043 20220 20052
rect 20168 20009 20177 20043
rect 20177 20009 20211 20043
rect 20211 20009 20220 20043
rect 20168 20000 20220 20009
rect 20628 20000 20680 20052
rect 17868 19932 17920 19984
rect 2320 19907 2372 19916
rect 2320 19873 2329 19907
rect 2329 19873 2363 19907
rect 2363 19873 2372 19907
rect 2320 19864 2372 19873
rect 2872 19907 2924 19916
rect 2872 19873 2881 19907
rect 2881 19873 2915 19907
rect 2915 19873 2924 19907
rect 2872 19864 2924 19873
rect 7288 19864 7340 19916
rect 8484 19864 8536 19916
rect 8668 19864 8720 19916
rect 10140 19864 10192 19916
rect 11152 19864 11204 19916
rect 11612 19864 11664 19916
rect 12072 19864 12124 19916
rect 13268 19907 13320 19916
rect 13268 19873 13277 19907
rect 13277 19873 13311 19907
rect 13311 19873 13320 19907
rect 13268 19864 13320 19873
rect 14280 19907 14332 19916
rect 14280 19873 14289 19907
rect 14289 19873 14323 19907
rect 14323 19873 14332 19907
rect 14280 19864 14332 19873
rect 3056 19796 3108 19848
rect 8760 19839 8812 19848
rect 8760 19805 8769 19839
rect 8769 19805 8803 19839
rect 8803 19805 8812 19839
rect 10416 19839 10468 19848
rect 8760 19796 8812 19805
rect 10416 19805 10425 19839
rect 10425 19805 10459 19839
rect 10459 19805 10468 19839
rect 10416 19796 10468 19805
rect 11888 19796 11940 19848
rect 13360 19839 13412 19848
rect 13360 19805 13369 19839
rect 13369 19805 13403 19839
rect 13403 19805 13412 19839
rect 13360 19796 13412 19805
rect 13544 19839 13596 19848
rect 13544 19805 13553 19839
rect 13553 19805 13587 19839
rect 13587 19805 13596 19839
rect 13544 19796 13596 19805
rect 2412 19728 2464 19780
rect 11796 19728 11848 19780
rect 13176 19728 13228 19780
rect 15292 19864 15344 19916
rect 17224 19907 17276 19916
rect 17224 19873 17233 19907
rect 17233 19873 17267 19907
rect 17267 19873 17276 19907
rect 17224 19864 17276 19873
rect 18604 19864 18656 19916
rect 18696 19864 18748 19916
rect 19432 19907 19484 19916
rect 19432 19873 19441 19907
rect 19441 19873 19475 19907
rect 19475 19873 19484 19907
rect 19432 19864 19484 19873
rect 19616 19864 19668 19916
rect 3056 19703 3108 19712
rect 3056 19669 3065 19703
rect 3065 19669 3099 19703
rect 3099 19669 3108 19703
rect 3056 19660 3108 19669
rect 8944 19660 8996 19712
rect 9404 19660 9456 19712
rect 11060 19660 11112 19712
rect 12164 19703 12216 19712
rect 12164 19669 12173 19703
rect 12173 19669 12207 19703
rect 12207 19669 12216 19703
rect 12164 19660 12216 19669
rect 14096 19660 14148 19712
rect 14188 19660 14240 19712
rect 17408 19839 17460 19848
rect 17408 19805 17417 19839
rect 17417 19805 17451 19839
rect 17451 19805 17460 19839
rect 17408 19796 17460 19805
rect 19340 19796 19392 19848
rect 17040 19728 17092 19780
rect 19064 19771 19116 19780
rect 19064 19737 19073 19771
rect 19073 19737 19107 19771
rect 19107 19737 19116 19771
rect 19064 19728 19116 19737
rect 16856 19703 16908 19712
rect 16856 19669 16865 19703
rect 16865 19669 16899 19703
rect 16899 19669 16908 19703
rect 16856 19660 16908 19669
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 1952 19499 2004 19508
rect 1952 19465 1961 19499
rect 1961 19465 1995 19499
rect 1995 19465 2004 19499
rect 1952 19456 2004 19465
rect 3424 19499 3476 19508
rect 3424 19465 3433 19499
rect 3433 19465 3467 19499
rect 3467 19465 3476 19499
rect 3424 19456 3476 19465
rect 2320 19388 2372 19440
rect 5356 19388 5408 19440
rect 8760 19456 8812 19508
rect 8852 19456 8904 19508
rect 12716 19456 12768 19508
rect 8576 19388 8628 19440
rect 9588 19388 9640 19440
rect 17224 19388 17276 19440
rect 18052 19388 18104 19440
rect 8852 19320 8904 19372
rect 8944 19320 8996 19372
rect 1768 19295 1820 19304
rect 1768 19261 1777 19295
rect 1777 19261 1811 19295
rect 1811 19261 1820 19295
rect 1768 19252 1820 19261
rect 2504 19252 2556 19304
rect 3424 19252 3476 19304
rect 3792 19252 3844 19304
rect 3976 19295 4028 19304
rect 3976 19261 3985 19295
rect 3985 19261 4019 19295
rect 4019 19261 4028 19295
rect 3976 19252 4028 19261
rect 5908 19295 5960 19304
rect 5908 19261 5917 19295
rect 5917 19261 5951 19295
rect 5951 19261 5960 19295
rect 5908 19252 5960 19261
rect 7104 19295 7156 19304
rect 7104 19261 7113 19295
rect 7113 19261 7147 19295
rect 7147 19261 7156 19295
rect 7104 19252 7156 19261
rect 7748 19252 7800 19304
rect 9128 19252 9180 19304
rect 14280 19363 14332 19372
rect 14280 19329 14289 19363
rect 14289 19329 14323 19363
rect 14323 19329 14332 19363
rect 14280 19320 14332 19329
rect 15476 19363 15528 19372
rect 15476 19329 15485 19363
rect 15485 19329 15519 19363
rect 15519 19329 15528 19363
rect 15476 19320 15528 19329
rect 16856 19320 16908 19372
rect 18512 19320 18564 19372
rect 19064 19320 19116 19372
rect 9312 19252 9364 19304
rect 9588 19252 9640 19304
rect 11704 19252 11756 19304
rect 14096 19295 14148 19304
rect 14096 19261 14105 19295
rect 14105 19261 14139 19295
rect 14139 19261 14148 19295
rect 14096 19252 14148 19261
rect 204 19184 256 19236
rect 2872 19184 2924 19236
rect 6552 19184 6604 19236
rect 2964 19116 3016 19168
rect 5540 19116 5592 19168
rect 6460 19116 6512 19168
rect 8484 19116 8536 19168
rect 8852 19116 8904 19168
rect 9128 19159 9180 19168
rect 9128 19125 9137 19159
rect 9137 19125 9171 19159
rect 9171 19125 9180 19159
rect 9128 19116 9180 19125
rect 9220 19116 9272 19168
rect 10508 19116 10560 19168
rect 11888 19184 11940 19236
rect 12716 19227 12768 19236
rect 12716 19193 12750 19227
rect 12750 19193 12768 19227
rect 12716 19184 12768 19193
rect 12808 19184 12860 19236
rect 11796 19116 11848 19168
rect 14556 19184 14608 19236
rect 13544 19116 13596 19168
rect 16856 19184 16908 19236
rect 15200 19159 15252 19168
rect 15200 19125 15209 19159
rect 15209 19125 15243 19159
rect 15243 19125 15252 19159
rect 15200 19116 15252 19125
rect 15936 19116 15988 19168
rect 18880 19295 18932 19304
rect 18880 19261 18889 19295
rect 18889 19261 18923 19295
rect 18923 19261 18932 19295
rect 18880 19252 18932 19261
rect 17500 19184 17552 19236
rect 20352 19252 20404 19304
rect 20536 19295 20588 19304
rect 20536 19261 20545 19295
rect 20545 19261 20579 19295
rect 20579 19261 20588 19295
rect 20536 19252 20588 19261
rect 17040 19116 17092 19168
rect 17776 19116 17828 19168
rect 22100 19184 22152 19236
rect 19248 19116 19300 19168
rect 20720 19159 20772 19168
rect 20720 19125 20729 19159
rect 20729 19125 20763 19159
rect 20763 19125 20772 19159
rect 20720 19116 20772 19125
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 1584 18912 1636 18964
rect 3240 18912 3292 18964
rect 1032 18844 1084 18896
rect 5816 18844 5868 18896
rect 5908 18844 5960 18896
rect 7288 18887 7340 18896
rect 7288 18853 7297 18887
rect 7297 18853 7331 18887
rect 7331 18853 7340 18887
rect 7288 18844 7340 18853
rect 8760 18844 8812 18896
rect 2136 18776 2188 18828
rect 3700 18776 3752 18828
rect 4804 18776 4856 18828
rect 7012 18819 7064 18828
rect 7012 18785 7021 18819
rect 7021 18785 7055 18819
rect 7055 18785 7064 18819
rect 7012 18776 7064 18785
rect 7104 18776 7156 18828
rect 9312 18912 9364 18964
rect 13360 18912 13412 18964
rect 18512 18955 18564 18964
rect 12348 18844 12400 18896
rect 12624 18887 12676 18896
rect 12624 18853 12633 18887
rect 12633 18853 12667 18887
rect 12667 18853 12676 18887
rect 12624 18844 12676 18853
rect 13544 18844 13596 18896
rect 15476 18844 15528 18896
rect 18512 18921 18521 18955
rect 18521 18921 18555 18955
rect 18555 18921 18564 18955
rect 18512 18912 18564 18921
rect 17408 18887 17460 18896
rect 17408 18853 17442 18887
rect 17442 18853 17460 18887
rect 17408 18844 17460 18853
rect 3148 18683 3200 18692
rect 3148 18649 3157 18683
rect 3157 18649 3191 18683
rect 3191 18649 3200 18683
rect 3148 18640 3200 18649
rect 3240 18640 3292 18692
rect 4988 18640 5040 18692
rect 5908 18708 5960 18760
rect 10876 18776 10928 18828
rect 11060 18776 11112 18828
rect 12164 18776 12216 18828
rect 9312 18708 9364 18760
rect 9680 18751 9732 18760
rect 9680 18717 9689 18751
rect 9689 18717 9723 18751
rect 9723 18717 9732 18751
rect 12716 18751 12768 18760
rect 9680 18708 9732 18717
rect 12716 18717 12725 18751
rect 12725 18717 12759 18751
rect 12759 18717 12768 18751
rect 12716 18708 12768 18717
rect 6460 18640 6512 18692
rect 12808 18640 12860 18692
rect 1400 18572 1452 18624
rect 2044 18572 2096 18624
rect 2228 18572 2280 18624
rect 3332 18572 3384 18624
rect 3516 18572 3568 18624
rect 8392 18572 8444 18624
rect 9680 18572 9732 18624
rect 18604 18776 18656 18828
rect 14556 18615 14608 18624
rect 14556 18581 14565 18615
rect 14565 18581 14599 18615
rect 14599 18581 14608 18615
rect 14556 18572 14608 18581
rect 16120 18572 16172 18624
rect 18512 18708 18564 18760
rect 16672 18572 16724 18624
rect 18972 18572 19024 18624
rect 20168 18615 20220 18624
rect 20168 18581 20177 18615
rect 20177 18581 20211 18615
rect 20211 18581 20220 18615
rect 20168 18572 20220 18581
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 2044 18368 2096 18420
rect 2872 18368 2924 18420
rect 3516 18368 3568 18420
rect 9128 18368 9180 18420
rect 9220 18368 9272 18420
rect 9956 18368 10008 18420
rect 3792 18343 3844 18352
rect 3792 18309 3801 18343
rect 3801 18309 3835 18343
rect 3835 18309 3844 18343
rect 3792 18300 3844 18309
rect 6828 18300 6880 18352
rect 10784 18368 10836 18420
rect 11704 18368 11756 18420
rect 13268 18368 13320 18420
rect 15476 18368 15528 18420
rect 15936 18411 15988 18420
rect 15936 18377 15945 18411
rect 15945 18377 15979 18411
rect 15979 18377 15988 18411
rect 15936 18368 15988 18377
rect 16028 18368 16080 18420
rect 17040 18368 17092 18420
rect 17132 18368 17184 18420
rect 19616 18368 19668 18420
rect 20444 18368 20496 18420
rect 20720 18411 20772 18420
rect 20720 18377 20729 18411
rect 20729 18377 20763 18411
rect 20763 18377 20772 18411
rect 20720 18368 20772 18377
rect 12808 18300 12860 18352
rect 13084 18300 13136 18352
rect 2136 18232 2188 18284
rect 4804 18275 4856 18284
rect 1768 18207 1820 18216
rect 1768 18173 1777 18207
rect 1777 18173 1811 18207
rect 1811 18173 1820 18207
rect 1768 18164 1820 18173
rect 2044 18164 2096 18216
rect 3240 18164 3292 18216
rect 572 18028 624 18080
rect 2228 18028 2280 18080
rect 4804 18241 4813 18275
rect 4813 18241 4847 18275
rect 4847 18241 4856 18275
rect 4804 18232 4856 18241
rect 7288 18232 7340 18284
rect 8760 18275 8812 18284
rect 8760 18241 8769 18275
rect 8769 18241 8803 18275
rect 8803 18241 8812 18275
rect 8760 18232 8812 18241
rect 8944 18232 8996 18284
rect 3884 18164 3936 18216
rect 4160 18164 4212 18216
rect 5816 18164 5868 18216
rect 3792 18096 3844 18148
rect 6828 18096 6880 18148
rect 8668 18164 8720 18216
rect 8852 18164 8904 18216
rect 9312 18164 9364 18216
rect 12716 18232 12768 18284
rect 15752 18300 15804 18352
rect 17224 18300 17276 18352
rect 20260 18300 20312 18352
rect 15844 18232 15896 18284
rect 17408 18232 17460 18284
rect 19248 18232 19300 18284
rect 20168 18275 20220 18284
rect 20168 18241 20177 18275
rect 20177 18241 20211 18275
rect 20211 18241 20220 18275
rect 20168 18232 20220 18241
rect 5264 18028 5316 18080
rect 5724 18028 5776 18080
rect 6920 18071 6972 18080
rect 6920 18037 6929 18071
rect 6929 18037 6963 18071
rect 6963 18037 6972 18071
rect 6920 18028 6972 18037
rect 8668 18071 8720 18080
rect 8668 18037 8677 18071
rect 8677 18037 8711 18071
rect 8711 18037 8720 18071
rect 8668 18028 8720 18037
rect 9680 18096 9732 18148
rect 9772 18096 9824 18148
rect 10968 18028 11020 18080
rect 14188 18164 14240 18216
rect 14556 18207 14608 18216
rect 14556 18173 14590 18207
rect 14590 18173 14608 18207
rect 14556 18164 14608 18173
rect 19432 18164 19484 18216
rect 20076 18164 20128 18216
rect 13360 18139 13412 18148
rect 13360 18105 13369 18139
rect 13369 18105 13403 18139
rect 13403 18105 13412 18139
rect 13360 18096 13412 18105
rect 14372 18096 14424 18148
rect 16028 18028 16080 18080
rect 16304 18139 16356 18148
rect 16304 18105 16313 18139
rect 16313 18105 16347 18139
rect 16347 18105 16356 18139
rect 16304 18096 16356 18105
rect 19064 18096 19116 18148
rect 20904 18096 20956 18148
rect 17408 18071 17460 18080
rect 17408 18037 17417 18071
rect 17417 18037 17451 18071
rect 17451 18037 17460 18071
rect 17408 18028 17460 18037
rect 17592 18028 17644 18080
rect 18788 18028 18840 18080
rect 18972 18071 19024 18080
rect 18972 18037 18981 18071
rect 18981 18037 19015 18071
rect 19015 18037 19024 18071
rect 18972 18028 19024 18037
rect 19524 18071 19576 18080
rect 19524 18037 19533 18071
rect 19533 18037 19567 18071
rect 19567 18037 19576 18071
rect 19524 18028 19576 18037
rect 20536 18028 20588 18080
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 1952 17867 2004 17876
rect 1952 17833 1961 17867
rect 1961 17833 1995 17867
rect 1995 17833 2004 17867
rect 1952 17824 2004 17833
rect 2780 17824 2832 17876
rect 4068 17824 4120 17876
rect 6644 17824 6696 17876
rect 7104 17824 7156 17876
rect 3332 17688 3384 17740
rect 3516 17756 3568 17808
rect 4068 17620 4120 17672
rect 4252 17688 4304 17740
rect 4804 17688 4856 17740
rect 5816 17731 5868 17740
rect 5816 17697 5850 17731
rect 5850 17697 5868 17731
rect 5816 17688 5868 17697
rect 7288 17688 7340 17740
rect 8116 17756 8168 17808
rect 9404 17824 9456 17876
rect 9772 17824 9824 17876
rect 11152 17824 11204 17876
rect 12808 17824 12860 17876
rect 14004 17824 14056 17876
rect 15200 17824 15252 17876
rect 16580 17867 16632 17876
rect 16580 17833 16589 17867
rect 16589 17833 16623 17867
rect 16623 17833 16632 17867
rect 16580 17824 16632 17833
rect 17960 17824 18012 17876
rect 18788 17824 18840 17876
rect 20904 17867 20956 17876
rect 20904 17833 20913 17867
rect 20913 17833 20947 17867
rect 20947 17833 20956 17867
rect 20904 17824 20956 17833
rect 7564 17731 7616 17740
rect 7564 17697 7573 17731
rect 7573 17697 7607 17731
rect 7607 17697 7616 17731
rect 7564 17688 7616 17697
rect 9128 17688 9180 17740
rect 4712 17663 4764 17672
rect 3240 17552 3292 17604
rect 4712 17629 4721 17663
rect 4721 17629 4755 17663
rect 4755 17629 4764 17663
rect 4712 17620 4764 17629
rect 5540 17663 5592 17672
rect 5540 17629 5549 17663
rect 5549 17629 5583 17663
rect 5583 17629 5592 17663
rect 5540 17620 5592 17629
rect 6828 17620 6880 17672
rect 7748 17663 7800 17672
rect 7748 17629 7757 17663
rect 7757 17629 7791 17663
rect 7791 17629 7800 17663
rect 9772 17688 9824 17740
rect 10416 17756 10468 17808
rect 11796 17799 11848 17808
rect 10232 17688 10284 17740
rect 11152 17688 11204 17740
rect 11796 17765 11805 17799
rect 11805 17765 11839 17799
rect 11839 17765 11848 17799
rect 11796 17756 11848 17765
rect 14188 17756 14240 17808
rect 16856 17756 16908 17808
rect 19248 17799 19300 17808
rect 7748 17620 7800 17629
rect 9312 17620 9364 17672
rect 9496 17620 9548 17672
rect 11796 17620 11848 17672
rect 12624 17620 12676 17672
rect 13544 17620 13596 17672
rect 13728 17620 13780 17672
rect 15292 17688 15344 17740
rect 15752 17731 15804 17740
rect 15752 17697 15761 17731
rect 15761 17697 15795 17731
rect 15795 17697 15804 17731
rect 15752 17688 15804 17697
rect 16948 17731 17000 17740
rect 14556 17620 14608 17672
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 16948 17697 16957 17731
rect 16957 17697 16991 17731
rect 16991 17697 17000 17731
rect 16948 17688 17000 17697
rect 19248 17765 19282 17799
rect 19282 17765 19300 17799
rect 19248 17756 19300 17765
rect 18420 17731 18472 17740
rect 18420 17697 18429 17731
rect 18429 17697 18463 17731
rect 18463 17697 18472 17731
rect 18420 17688 18472 17697
rect 3056 17527 3108 17536
rect 3056 17493 3065 17527
rect 3065 17493 3099 17527
rect 3099 17493 3108 17527
rect 3056 17484 3108 17493
rect 3976 17484 4028 17536
rect 5448 17552 5500 17604
rect 9404 17552 9456 17604
rect 7380 17484 7432 17536
rect 19616 17688 19668 17740
rect 18604 17620 18656 17672
rect 18788 17620 18840 17672
rect 13268 17484 13320 17536
rect 16764 17484 16816 17536
rect 18972 17484 19024 17536
rect 19892 17484 19944 17536
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 2780 17280 2832 17332
rect 3056 17280 3108 17332
rect 6828 17323 6880 17332
rect 4068 17212 4120 17264
rect 5816 17212 5868 17264
rect 6828 17289 6837 17323
rect 6837 17289 6871 17323
rect 6871 17289 6880 17323
rect 6828 17280 6880 17289
rect 7104 17280 7156 17332
rect 10876 17280 10928 17332
rect 11612 17280 11664 17332
rect 15108 17280 15160 17332
rect 15384 17323 15436 17332
rect 15384 17289 15393 17323
rect 15393 17289 15427 17323
rect 15427 17289 15436 17323
rect 15384 17280 15436 17289
rect 16672 17280 16724 17332
rect 16948 17280 17000 17332
rect 18880 17280 18932 17332
rect 19340 17280 19392 17332
rect 21732 17280 21784 17332
rect 14188 17212 14240 17264
rect 17408 17212 17460 17264
rect 3976 17187 4028 17196
rect 3976 17153 3985 17187
rect 3985 17153 4019 17187
rect 4019 17153 4028 17187
rect 3976 17144 4028 17153
rect 1860 17076 1912 17128
rect 2964 17076 3016 17128
rect 4528 17119 4580 17128
rect 4528 17085 4537 17119
rect 4537 17085 4571 17119
rect 4571 17085 4580 17119
rect 4528 17076 4580 17085
rect 2136 17008 2188 17060
rect 6920 17144 6972 17196
rect 7380 17187 7432 17196
rect 7380 17153 7389 17187
rect 7389 17153 7423 17187
rect 7423 17153 7432 17187
rect 7380 17144 7432 17153
rect 8116 17144 8168 17196
rect 9036 17144 9088 17196
rect 9220 17144 9272 17196
rect 9404 17187 9456 17196
rect 9404 17153 9413 17187
rect 9413 17153 9447 17187
rect 9447 17153 9456 17187
rect 9404 17144 9456 17153
rect 9864 17144 9916 17196
rect 6644 17076 6696 17128
rect 6828 17076 6880 17128
rect 7472 17076 7524 17128
rect 10600 17076 10652 17128
rect 10876 17076 10928 17128
rect 5448 17008 5500 17060
rect 1952 16983 2004 16992
rect 1952 16949 1961 16983
rect 1961 16949 1995 16983
rect 1995 16949 2004 16983
rect 1952 16940 2004 16949
rect 3056 16983 3108 16992
rect 3056 16949 3065 16983
rect 3065 16949 3099 16983
rect 3099 16949 3108 16983
rect 3056 16940 3108 16949
rect 3884 16983 3936 16992
rect 3884 16949 3893 16983
rect 3893 16949 3927 16983
rect 3927 16949 3936 16983
rect 3884 16940 3936 16949
rect 8024 17008 8076 17060
rect 10048 17008 10100 17060
rect 10232 17008 10284 17060
rect 10968 17008 11020 17060
rect 11520 17051 11572 17060
rect 11520 17017 11529 17051
rect 11529 17017 11563 17051
rect 11563 17017 11572 17051
rect 11520 17008 11572 17017
rect 11704 17076 11756 17128
rect 13820 17144 13872 17196
rect 19156 17212 19208 17264
rect 13268 17119 13320 17128
rect 13268 17085 13277 17119
rect 13277 17085 13311 17119
rect 13311 17085 13320 17119
rect 13268 17076 13320 17085
rect 13360 17119 13412 17128
rect 13360 17085 13369 17119
rect 13369 17085 13403 17119
rect 13403 17085 13412 17119
rect 13360 17076 13412 17085
rect 14004 17076 14056 17128
rect 14096 17076 14148 17128
rect 8392 16940 8444 16992
rect 8944 16983 8996 16992
rect 8944 16949 8953 16983
rect 8953 16949 8987 16983
rect 8987 16949 8996 16983
rect 8944 16940 8996 16949
rect 9036 16940 9088 16992
rect 9404 16940 9456 16992
rect 10784 16940 10836 16992
rect 11704 16940 11756 16992
rect 11888 16940 11940 16992
rect 14556 17008 14608 17060
rect 16028 17076 16080 17128
rect 18052 17076 18104 17128
rect 19156 17076 19208 17128
rect 19524 17076 19576 17128
rect 19800 17187 19852 17196
rect 19800 17153 19809 17187
rect 19809 17153 19843 17187
rect 19843 17153 19852 17187
rect 19800 17144 19852 17153
rect 17776 17008 17828 17060
rect 17868 17008 17920 17060
rect 20076 17008 20128 17060
rect 16764 16940 16816 16992
rect 17684 16983 17736 16992
rect 17684 16949 17693 16983
rect 17693 16949 17727 16983
rect 17727 16949 17736 16983
rect 17684 16940 17736 16949
rect 18420 16983 18472 16992
rect 18420 16949 18429 16983
rect 18429 16949 18463 16983
rect 18463 16949 18472 16983
rect 18420 16940 18472 16949
rect 19616 16940 19668 16992
rect 20260 16940 20312 16992
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 4068 16736 4120 16788
rect 5448 16779 5500 16788
rect 4712 16668 4764 16720
rect 5448 16745 5457 16779
rect 5457 16745 5491 16779
rect 5491 16745 5500 16779
rect 5448 16736 5500 16745
rect 7104 16736 7156 16788
rect 7748 16736 7800 16788
rect 9496 16736 9548 16788
rect 11612 16736 11664 16788
rect 11888 16779 11940 16788
rect 11888 16745 11897 16779
rect 11897 16745 11931 16779
rect 11931 16745 11940 16779
rect 11888 16736 11940 16745
rect 12348 16736 12400 16788
rect 13360 16736 13412 16788
rect 14096 16779 14148 16788
rect 14096 16745 14105 16779
rect 14105 16745 14139 16779
rect 14139 16745 14148 16779
rect 14096 16736 14148 16745
rect 14556 16779 14608 16788
rect 14556 16745 14565 16779
rect 14565 16745 14599 16779
rect 14599 16745 14608 16779
rect 14556 16736 14608 16745
rect 7380 16668 7432 16720
rect 9128 16668 9180 16720
rect 1768 16643 1820 16652
rect 1768 16609 1777 16643
rect 1777 16609 1811 16643
rect 1811 16609 1820 16643
rect 1768 16600 1820 16609
rect 3148 16600 3200 16652
rect 4620 16600 4672 16652
rect 7656 16600 7708 16652
rect 10876 16643 10928 16652
rect 10876 16609 10885 16643
rect 10885 16609 10919 16643
rect 10919 16609 10928 16643
rect 10876 16600 10928 16609
rect 14740 16668 14792 16720
rect 2320 16575 2372 16584
rect 2320 16541 2329 16575
rect 2329 16541 2363 16575
rect 2363 16541 2372 16575
rect 2320 16532 2372 16541
rect 7472 16532 7524 16584
rect 1952 16507 2004 16516
rect 1952 16473 1961 16507
rect 1961 16473 1995 16507
rect 1995 16473 2004 16507
rect 1952 16464 2004 16473
rect 2228 16396 2280 16448
rect 3424 16396 3476 16448
rect 4068 16396 4120 16448
rect 9036 16532 9088 16584
rect 11152 16575 11204 16584
rect 11152 16541 11161 16575
rect 11161 16541 11195 16575
rect 11195 16541 11204 16575
rect 11152 16532 11204 16541
rect 9864 16464 9916 16516
rect 11704 16600 11756 16652
rect 13728 16600 13780 16652
rect 12348 16532 12400 16584
rect 14096 16600 14148 16652
rect 14924 16668 14976 16720
rect 18052 16736 18104 16788
rect 19156 16736 19208 16788
rect 16672 16668 16724 16720
rect 16948 16668 17000 16720
rect 18972 16668 19024 16720
rect 19340 16668 19392 16720
rect 15200 16600 15252 16652
rect 17040 16600 17092 16652
rect 17224 16600 17276 16652
rect 12808 16464 12860 16516
rect 15476 16532 15528 16584
rect 13544 16464 13596 16516
rect 15108 16464 15160 16516
rect 16764 16532 16816 16584
rect 17132 16575 17184 16584
rect 17132 16541 17141 16575
rect 17141 16541 17175 16575
rect 17175 16541 17184 16575
rect 17132 16532 17184 16541
rect 17960 16600 18012 16652
rect 19248 16600 19300 16652
rect 9772 16439 9824 16448
rect 9772 16405 9781 16439
rect 9781 16405 9815 16439
rect 9815 16405 9824 16439
rect 9772 16396 9824 16405
rect 12440 16396 12492 16448
rect 14004 16396 14056 16448
rect 15292 16439 15344 16448
rect 15292 16405 15301 16439
rect 15301 16405 15335 16439
rect 15335 16405 15344 16439
rect 15292 16396 15344 16405
rect 17408 16396 17460 16448
rect 18604 16396 18656 16448
rect 18880 16396 18932 16448
rect 19156 16396 19208 16448
rect 19984 16600 20036 16652
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 4252 16192 4304 16244
rect 7564 16192 7616 16244
rect 9036 16192 9088 16244
rect 11152 16192 11204 16244
rect 13820 16235 13872 16244
rect 13820 16201 13829 16235
rect 13829 16201 13863 16235
rect 13863 16201 13872 16235
rect 13820 16192 13872 16201
rect 15476 16235 15528 16244
rect 15476 16201 15485 16235
rect 15485 16201 15519 16235
rect 15519 16201 15528 16235
rect 15476 16192 15528 16201
rect 16396 16192 16448 16244
rect 17592 16235 17644 16244
rect 4804 16124 4856 16176
rect 6920 16124 6972 16176
rect 3148 16099 3200 16108
rect 3148 16065 3157 16099
rect 3157 16065 3191 16099
rect 3191 16065 3200 16099
rect 3148 16056 3200 16065
rect 4068 16056 4120 16108
rect 7380 16099 7432 16108
rect 7380 16065 7389 16099
rect 7389 16065 7423 16099
rect 7423 16065 7432 16099
rect 7380 16056 7432 16065
rect 7748 16056 7800 16108
rect 8208 16056 8260 16108
rect 2228 15988 2280 16040
rect 3240 15988 3292 16040
rect 7104 15988 7156 16040
rect 6092 15920 6144 15972
rect 1400 15852 1452 15904
rect 3056 15895 3108 15904
rect 3056 15861 3065 15895
rect 3065 15861 3099 15895
rect 3099 15861 3108 15895
rect 3056 15852 3108 15861
rect 4988 15852 5040 15904
rect 7380 15852 7432 15904
rect 8208 15895 8260 15904
rect 8208 15861 8217 15895
rect 8217 15861 8251 15895
rect 8251 15861 8260 15895
rect 8208 15852 8260 15861
rect 9496 16099 9548 16108
rect 9496 16065 9505 16099
rect 9505 16065 9539 16099
rect 9539 16065 9548 16099
rect 9496 16056 9548 16065
rect 9772 16056 9824 16108
rect 12440 16124 12492 16176
rect 17592 16201 17601 16235
rect 17601 16201 17635 16235
rect 17635 16201 17644 16235
rect 17592 16192 17644 16201
rect 19248 16192 19300 16244
rect 18972 16124 19024 16176
rect 8944 15988 8996 16040
rect 9404 16031 9456 16040
rect 9404 15997 9413 16031
rect 9413 15997 9447 16031
rect 9447 15997 9456 16031
rect 9404 15988 9456 15997
rect 10048 15988 10100 16040
rect 11612 16031 11664 16040
rect 11612 15997 11621 16031
rect 11621 15997 11655 16031
rect 11655 15997 11664 16031
rect 11612 15988 11664 15997
rect 12440 16031 12492 16040
rect 12440 15997 12449 16031
rect 12449 15997 12483 16031
rect 12483 15997 12492 16031
rect 12440 15988 12492 15997
rect 13084 15988 13136 16040
rect 13544 15988 13596 16040
rect 14372 16031 14424 16040
rect 14372 15997 14395 16031
rect 14395 15997 14424 16031
rect 11980 15920 12032 15972
rect 12808 15920 12860 15972
rect 14372 15988 14424 15997
rect 16856 16056 16908 16108
rect 17684 16056 17736 16108
rect 17960 16056 18012 16108
rect 17500 15988 17552 16040
rect 17960 15920 18012 15972
rect 18604 15988 18656 16040
rect 19616 15988 19668 16040
rect 19432 15920 19484 15972
rect 17132 15895 17184 15904
rect 17132 15861 17141 15895
rect 17141 15861 17175 15895
rect 17175 15861 17184 15895
rect 17132 15852 17184 15861
rect 17316 15852 17368 15904
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 1952 15691 2004 15700
rect 1952 15657 1961 15691
rect 1961 15657 1995 15691
rect 1995 15657 2004 15691
rect 1952 15648 2004 15657
rect 3056 15648 3108 15700
rect 3884 15648 3936 15700
rect 5540 15648 5592 15700
rect 7380 15691 7432 15700
rect 7380 15657 7389 15691
rect 7389 15657 7423 15691
rect 7423 15657 7432 15691
rect 7380 15648 7432 15657
rect 7564 15648 7616 15700
rect 2872 15623 2924 15632
rect 2872 15589 2881 15623
rect 2881 15589 2915 15623
rect 2915 15589 2924 15623
rect 2872 15580 2924 15589
rect 3424 15580 3476 15632
rect 8208 15580 8260 15632
rect 9588 15648 9640 15700
rect 10876 15648 10928 15700
rect 14096 15691 14148 15700
rect 14096 15657 14105 15691
rect 14105 15657 14139 15691
rect 14139 15657 14148 15691
rect 14096 15648 14148 15657
rect 15292 15648 15344 15700
rect 7656 15512 7708 15564
rect 7748 15512 7800 15564
rect 10692 15555 10744 15564
rect 3240 15444 3292 15496
rect 4160 15444 4212 15496
rect 4712 15487 4764 15496
rect 4712 15453 4721 15487
rect 4721 15453 4755 15487
rect 4755 15453 4764 15487
rect 4712 15444 4764 15453
rect 5356 15444 5408 15496
rect 4068 15376 4120 15428
rect 7288 15444 7340 15496
rect 10692 15521 10701 15555
rect 10701 15521 10735 15555
rect 10735 15521 10744 15555
rect 10692 15512 10744 15521
rect 11244 15512 11296 15564
rect 8484 15444 8536 15496
rect 9036 15487 9088 15496
rect 9036 15453 9045 15487
rect 9045 15453 9079 15487
rect 9079 15453 9088 15487
rect 9036 15444 9088 15453
rect 6184 15376 6236 15428
rect 10048 15444 10100 15496
rect 11152 15444 11204 15496
rect 12624 15580 12676 15632
rect 17132 15580 17184 15632
rect 17408 15648 17460 15700
rect 18696 15691 18748 15700
rect 18696 15657 18705 15691
rect 18705 15657 18739 15691
rect 18739 15657 18748 15691
rect 18696 15648 18748 15657
rect 19984 15648 20036 15700
rect 17868 15580 17920 15632
rect 12440 15512 12492 15564
rect 14372 15512 14424 15564
rect 13176 15444 13228 15496
rect 14556 15487 14608 15496
rect 14556 15453 14565 15487
rect 14565 15453 14599 15487
rect 14599 15453 14608 15487
rect 14556 15444 14608 15453
rect 15200 15512 15252 15564
rect 19524 15580 19576 15632
rect 7564 15308 7616 15360
rect 10416 15376 10468 15428
rect 12808 15376 12860 15428
rect 18880 15512 18932 15564
rect 20076 15555 20128 15564
rect 20076 15521 20085 15555
rect 20085 15521 20119 15555
rect 20119 15521 20128 15555
rect 20076 15512 20128 15521
rect 16028 15487 16080 15496
rect 16028 15453 16037 15487
rect 16037 15453 16071 15487
rect 16071 15453 16080 15487
rect 16028 15444 16080 15453
rect 11704 15308 11756 15360
rect 11980 15308 12032 15360
rect 17040 15376 17092 15428
rect 17868 15444 17920 15496
rect 18696 15444 18748 15496
rect 19248 15487 19300 15496
rect 19248 15453 19257 15487
rect 19257 15453 19291 15487
rect 19291 15453 19300 15487
rect 20168 15487 20220 15496
rect 19248 15444 19300 15453
rect 17776 15376 17828 15428
rect 18604 15376 18656 15428
rect 19708 15419 19760 15428
rect 19708 15385 19717 15419
rect 19717 15385 19751 15419
rect 19751 15385 19760 15419
rect 19708 15376 19760 15385
rect 20168 15453 20177 15487
rect 20177 15453 20211 15487
rect 20211 15453 20220 15487
rect 20168 15444 20220 15453
rect 17684 15351 17736 15360
rect 17684 15317 17693 15351
rect 17693 15317 17727 15351
rect 17727 15317 17736 15351
rect 17684 15308 17736 15317
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 7656 15104 7708 15156
rect 3424 15036 3476 15088
rect 9772 15104 9824 15156
rect 10048 15104 10100 15156
rect 10692 15104 10744 15156
rect 11704 15104 11756 15156
rect 12164 15104 12216 15156
rect 13084 15104 13136 15156
rect 13544 15104 13596 15156
rect 14464 15104 14516 15156
rect 14556 15104 14608 15156
rect 17960 15104 18012 15156
rect 9956 15036 10008 15088
rect 11520 15036 11572 15088
rect 11612 15036 11664 15088
rect 12072 15036 12124 15088
rect 12716 15036 12768 15088
rect 12992 15036 13044 15088
rect 19248 15104 19300 15156
rect 19432 15147 19484 15156
rect 19432 15113 19441 15147
rect 19441 15113 19475 15147
rect 19475 15113 19484 15147
rect 19432 15104 19484 15113
rect 20168 15104 20220 15156
rect 20628 15104 20680 15156
rect 1860 15011 1912 15020
rect 1860 14977 1869 15011
rect 1869 14977 1903 15011
rect 1903 14977 1912 15011
rect 1860 14968 1912 14977
rect 5816 14968 5868 15020
rect 7012 14968 7064 15020
rect 7472 15011 7524 15020
rect 7472 14977 7481 15011
rect 7481 14977 7515 15011
rect 7515 14977 7524 15011
rect 7472 14968 7524 14977
rect 2320 14943 2372 14952
rect 2320 14909 2329 14943
rect 2329 14909 2363 14943
rect 2363 14909 2372 14943
rect 2320 14900 2372 14909
rect 3884 14900 3936 14952
rect 7380 14900 7432 14952
rect 8208 14900 8260 14952
rect 9864 14900 9916 14952
rect 12164 14968 12216 15020
rect 13452 14968 13504 15020
rect 15108 14968 15160 15020
rect 10324 14900 10376 14952
rect 10600 14900 10652 14952
rect 10784 14900 10836 14952
rect 11704 14900 11756 14952
rect 11888 14900 11940 14952
rect 12900 14900 12952 14952
rect 13820 14943 13872 14952
rect 13820 14909 13829 14943
rect 13829 14909 13863 14943
rect 13863 14909 13872 14943
rect 13820 14900 13872 14909
rect 17316 14968 17368 15020
rect 15660 14943 15712 14952
rect 15660 14909 15669 14943
rect 15669 14909 15703 14943
rect 15703 14909 15712 14943
rect 15660 14900 15712 14909
rect 17684 14900 17736 14952
rect 17776 14900 17828 14952
rect 18328 14943 18380 14952
rect 18328 14909 18351 14943
rect 18351 14909 18380 14943
rect 18328 14900 18380 14909
rect 18604 14900 18656 14952
rect 3240 14832 3292 14884
rect 5448 14832 5500 14884
rect 9956 14832 10008 14884
rect 10876 14832 10928 14884
rect 11244 14832 11296 14884
rect 15936 14832 15988 14884
rect 3148 14764 3200 14816
rect 5356 14764 5408 14816
rect 6828 14807 6880 14816
rect 6828 14773 6837 14807
rect 6837 14773 6871 14807
rect 6871 14773 6880 14807
rect 6828 14764 6880 14773
rect 10324 14764 10376 14816
rect 10784 14764 10836 14816
rect 11980 14807 12032 14816
rect 11980 14773 11989 14807
rect 11989 14773 12023 14807
rect 12023 14773 12032 14807
rect 11980 14764 12032 14773
rect 12624 14807 12676 14816
rect 12624 14773 12633 14807
rect 12633 14773 12667 14807
rect 12667 14773 12676 14807
rect 12624 14764 12676 14773
rect 12992 14807 13044 14816
rect 12992 14773 13001 14807
rect 13001 14773 13035 14807
rect 13035 14773 13044 14807
rect 12992 14764 13044 14773
rect 15476 14764 15528 14816
rect 16856 14832 16908 14884
rect 17500 14832 17552 14884
rect 16948 14764 17000 14816
rect 18604 14764 18656 14816
rect 19340 14764 19392 14816
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 1952 14603 2004 14612
rect 1952 14569 1961 14603
rect 1961 14569 1995 14603
rect 1995 14569 2004 14603
rect 1952 14560 2004 14569
rect 4160 14560 4212 14612
rect 4988 14560 5040 14612
rect 5264 14560 5316 14612
rect 5816 14603 5868 14612
rect 5816 14569 5825 14603
rect 5825 14569 5859 14603
rect 5859 14569 5868 14603
rect 5816 14560 5868 14569
rect 6920 14560 6972 14612
rect 9588 14560 9640 14612
rect 10784 14603 10836 14612
rect 10784 14569 10793 14603
rect 10793 14569 10827 14603
rect 10827 14569 10836 14603
rect 10784 14560 10836 14569
rect 11244 14603 11296 14612
rect 11244 14569 11253 14603
rect 11253 14569 11287 14603
rect 11287 14569 11296 14603
rect 11244 14560 11296 14569
rect 11520 14560 11572 14612
rect 12440 14560 12492 14612
rect 12532 14560 12584 14612
rect 12624 14560 12676 14612
rect 3148 14492 3200 14544
rect 1676 14424 1728 14476
rect 3056 14467 3108 14476
rect 3056 14433 3065 14467
rect 3065 14433 3099 14467
rect 3099 14433 3108 14467
rect 3056 14424 3108 14433
rect 2228 14356 2280 14408
rect 3884 14424 3936 14476
rect 5540 14492 5592 14544
rect 7012 14492 7064 14544
rect 5080 14424 5132 14476
rect 5264 14424 5316 14476
rect 11888 14492 11940 14544
rect 12072 14492 12124 14544
rect 17408 14560 17460 14612
rect 18328 14603 18380 14612
rect 18328 14569 18337 14603
rect 18337 14569 18371 14603
rect 18371 14569 18380 14603
rect 18328 14560 18380 14569
rect 18604 14603 18656 14612
rect 18604 14569 18613 14603
rect 18613 14569 18647 14603
rect 18647 14569 18656 14603
rect 18604 14560 18656 14569
rect 5540 14356 5592 14408
rect 7472 14356 7524 14408
rect 9036 14424 9088 14476
rect 10048 14356 10100 14408
rect 10416 14356 10468 14408
rect 10784 14356 10836 14408
rect 13544 14424 13596 14476
rect 3424 14288 3476 14340
rect 7104 14288 7156 14340
rect 14832 14492 14884 14544
rect 17040 14492 17092 14544
rect 17868 14492 17920 14544
rect 17960 14492 18012 14544
rect 19156 14560 19208 14612
rect 14096 14467 14148 14476
rect 14096 14433 14105 14467
rect 14105 14433 14139 14467
rect 14139 14433 14148 14467
rect 14096 14424 14148 14433
rect 15016 14424 15068 14476
rect 16212 14424 16264 14476
rect 17776 14424 17828 14476
rect 14372 14356 14424 14408
rect 2044 14220 2096 14272
rect 7012 14220 7064 14272
rect 7472 14263 7524 14272
rect 7472 14229 7481 14263
rect 7481 14229 7515 14263
rect 7515 14229 7524 14263
rect 7472 14220 7524 14229
rect 7748 14263 7800 14272
rect 7748 14229 7757 14263
rect 7757 14229 7791 14263
rect 7791 14229 7800 14263
rect 7748 14220 7800 14229
rect 8300 14220 8352 14272
rect 9036 14220 9088 14272
rect 10968 14220 11020 14272
rect 13820 14288 13872 14340
rect 15384 14288 15436 14340
rect 13452 14220 13504 14272
rect 16304 14356 16356 14408
rect 16580 14356 16632 14408
rect 16856 14356 16908 14408
rect 18420 14356 18472 14408
rect 18972 14356 19024 14408
rect 19248 14424 19300 14476
rect 19800 14356 19852 14408
rect 20168 14399 20220 14408
rect 20168 14365 20177 14399
rect 20177 14365 20211 14399
rect 20211 14365 20220 14399
rect 20168 14356 20220 14365
rect 16764 14288 16816 14340
rect 17316 14220 17368 14272
rect 17592 14220 17644 14272
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 1676 13923 1728 13932
rect 1676 13889 1685 13923
rect 1685 13889 1719 13923
rect 1719 13889 1728 13923
rect 1676 13880 1728 13889
rect 3884 14016 3936 14068
rect 5080 14059 5132 14068
rect 5080 14025 5089 14059
rect 5089 14025 5123 14059
rect 5123 14025 5132 14059
rect 5080 14016 5132 14025
rect 5356 14059 5408 14068
rect 5356 14025 5365 14059
rect 5365 14025 5399 14059
rect 5399 14025 5408 14059
rect 5356 14016 5408 14025
rect 7012 14016 7064 14068
rect 8760 14059 8812 14068
rect 8760 14025 8769 14059
rect 8769 14025 8803 14059
rect 8803 14025 8812 14059
rect 8760 14016 8812 14025
rect 6000 13880 6052 13932
rect 9404 13923 9456 13932
rect 9404 13889 9413 13923
rect 9413 13889 9447 13923
rect 9447 13889 9456 13923
rect 9404 13880 9456 13889
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 3608 13812 3660 13864
rect 5264 13812 5316 13864
rect 6828 13812 6880 13864
rect 7380 13855 7432 13864
rect 7380 13821 7389 13855
rect 7389 13821 7423 13855
rect 7423 13821 7432 13855
rect 7380 13812 7432 13821
rect 1584 13744 1636 13796
rect 7472 13744 7524 13796
rect 8944 13744 8996 13796
rect 10416 13880 10468 13932
rect 10968 13923 11020 13932
rect 10968 13889 10977 13923
rect 10977 13889 11011 13923
rect 11011 13889 11020 13923
rect 10968 13880 11020 13889
rect 11152 14016 11204 14068
rect 11980 14016 12032 14068
rect 14832 14016 14884 14068
rect 15016 14059 15068 14068
rect 15016 14025 15025 14059
rect 15025 14025 15059 14059
rect 15059 14025 15068 14059
rect 15016 14016 15068 14025
rect 16580 14016 16632 14068
rect 17040 14016 17092 14068
rect 20168 14016 20220 14068
rect 11520 13948 11572 14000
rect 12440 13948 12492 14000
rect 11152 13880 11204 13932
rect 12164 13880 12216 13932
rect 15108 13948 15160 14000
rect 18512 13948 18564 14000
rect 12072 13812 12124 13864
rect 13452 13812 13504 13864
rect 16396 13880 16448 13932
rect 17500 13923 17552 13932
rect 17500 13889 17509 13923
rect 17509 13889 17543 13923
rect 17543 13889 17552 13923
rect 17500 13880 17552 13889
rect 16488 13855 16540 13864
rect 16488 13821 16497 13855
rect 16497 13821 16531 13855
rect 16531 13821 16540 13855
rect 16488 13812 16540 13821
rect 16672 13812 16724 13864
rect 20168 13880 20220 13932
rect 10048 13787 10100 13796
rect 10048 13753 10057 13787
rect 10057 13753 10091 13787
rect 10091 13753 10100 13787
rect 10048 13744 10100 13753
rect 14556 13744 14608 13796
rect 15016 13744 15068 13796
rect 7748 13676 7800 13728
rect 9220 13719 9272 13728
rect 9220 13685 9229 13719
rect 9229 13685 9263 13719
rect 9263 13685 9272 13719
rect 9220 13676 9272 13685
rect 13820 13676 13872 13728
rect 14372 13676 14424 13728
rect 15292 13676 15344 13728
rect 16212 13744 16264 13796
rect 18144 13812 18196 13864
rect 18696 13812 18748 13864
rect 19432 13812 19484 13864
rect 18972 13744 19024 13796
rect 19064 13744 19116 13796
rect 18788 13676 18840 13728
rect 19892 13676 19944 13728
rect 20260 13719 20312 13728
rect 20260 13685 20269 13719
rect 20269 13685 20303 13719
rect 20303 13685 20312 13719
rect 20260 13676 20312 13685
rect 20444 13676 20496 13728
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 1768 13515 1820 13524
rect 1768 13481 1777 13515
rect 1777 13481 1811 13515
rect 1811 13481 1820 13515
rect 1768 13472 1820 13481
rect 6460 13472 6512 13524
rect 6920 13515 6972 13524
rect 6920 13481 6929 13515
rect 6929 13481 6963 13515
rect 6963 13481 6972 13515
rect 6920 13472 6972 13481
rect 7380 13472 7432 13524
rect 8852 13515 8904 13524
rect 8852 13481 8861 13515
rect 8861 13481 8895 13515
rect 8895 13481 8904 13515
rect 8852 13472 8904 13481
rect 9404 13472 9456 13524
rect 9864 13472 9916 13524
rect 10232 13472 10284 13524
rect 10876 13472 10928 13524
rect 2136 13404 2188 13456
rect 3148 13404 3200 13456
rect 4068 13404 4120 13456
rect 1584 13379 1636 13388
rect 1584 13345 1593 13379
rect 1593 13345 1627 13379
rect 1627 13345 1636 13379
rect 1584 13336 1636 13345
rect 2412 13336 2464 13388
rect 4252 13336 4304 13388
rect 6644 13336 6696 13388
rect 7840 13404 7892 13456
rect 8760 13404 8812 13456
rect 11888 13472 11940 13524
rect 12624 13472 12676 13524
rect 12992 13515 13044 13524
rect 12992 13481 13001 13515
rect 13001 13481 13035 13515
rect 13035 13481 13044 13515
rect 12992 13472 13044 13481
rect 11520 13379 11572 13388
rect 3424 13268 3476 13320
rect 4712 13268 4764 13320
rect 5264 13268 5316 13320
rect 5908 13311 5960 13320
rect 5908 13277 5917 13311
rect 5917 13277 5951 13311
rect 5951 13277 5960 13311
rect 5908 13268 5960 13277
rect 6000 13311 6052 13320
rect 6000 13277 6009 13311
rect 6009 13277 6043 13311
rect 6043 13277 6052 13311
rect 6000 13268 6052 13277
rect 7380 13268 7432 13320
rect 5448 13243 5500 13252
rect 5448 13209 5457 13243
rect 5457 13209 5491 13243
rect 5491 13209 5500 13243
rect 5448 13200 5500 13209
rect 5632 13200 5684 13252
rect 6828 13200 6880 13252
rect 8484 13268 8536 13320
rect 3148 13132 3200 13184
rect 7748 13132 7800 13184
rect 11520 13345 11529 13379
rect 11529 13345 11563 13379
rect 11563 13345 11572 13379
rect 11520 13336 11572 13345
rect 12900 13404 12952 13456
rect 15108 13472 15160 13524
rect 15292 13515 15344 13524
rect 15292 13481 15301 13515
rect 15301 13481 15335 13515
rect 15335 13481 15344 13515
rect 15292 13472 15344 13481
rect 15568 13472 15620 13524
rect 13820 13404 13872 13456
rect 16396 13472 16448 13524
rect 19616 13515 19668 13524
rect 19616 13481 19625 13515
rect 19625 13481 19659 13515
rect 19659 13481 19668 13515
rect 19616 13472 19668 13481
rect 16304 13404 16356 13456
rect 19892 13404 19944 13456
rect 11888 13132 11940 13184
rect 12808 13336 12860 13388
rect 13544 13268 13596 13320
rect 14280 13311 14332 13320
rect 13176 13200 13228 13252
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 14464 13311 14516 13320
rect 14464 13277 14473 13311
rect 14473 13277 14507 13311
rect 14507 13277 14516 13311
rect 14464 13268 14516 13277
rect 17868 13336 17920 13388
rect 15292 13268 15344 13320
rect 16304 13311 16356 13320
rect 16304 13277 16313 13311
rect 16313 13277 16347 13311
rect 16347 13277 16356 13311
rect 16304 13268 16356 13277
rect 17776 13268 17828 13320
rect 18052 13336 18104 13388
rect 18236 13379 18288 13388
rect 18236 13345 18270 13379
rect 18270 13345 18288 13379
rect 18236 13336 18288 13345
rect 19156 13336 19208 13388
rect 19616 13336 19668 13388
rect 18972 13268 19024 13320
rect 13728 13132 13780 13184
rect 17500 13132 17552 13184
rect 19432 13132 19484 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 2780 12928 2832 12980
rect 5908 12928 5960 12980
rect 9220 12928 9272 12980
rect 11704 12928 11756 12980
rect 12072 12928 12124 12980
rect 6000 12860 6052 12912
rect 7104 12860 7156 12912
rect 7472 12860 7524 12912
rect 8300 12860 8352 12912
rect 4252 12835 4304 12844
rect 4252 12801 4261 12835
rect 4261 12801 4295 12835
rect 4295 12801 4304 12835
rect 4252 12792 4304 12801
rect 5264 12835 5316 12844
rect 5264 12801 5273 12835
rect 5273 12801 5307 12835
rect 5307 12801 5316 12835
rect 5264 12792 5316 12801
rect 6276 12835 6328 12844
rect 6276 12801 6285 12835
rect 6285 12801 6319 12835
rect 6319 12801 6328 12835
rect 6276 12792 6328 12801
rect 7748 12792 7800 12844
rect 7840 12835 7892 12844
rect 7840 12801 7849 12835
rect 7849 12801 7883 12835
rect 7883 12801 7892 12835
rect 7840 12792 7892 12801
rect 8944 12792 8996 12844
rect 1860 12724 1912 12776
rect 2596 12724 2648 12776
rect 4988 12724 5040 12776
rect 5356 12724 5408 12776
rect 8760 12724 8812 12776
rect 13544 12860 13596 12912
rect 13728 12835 13780 12844
rect 13728 12801 13737 12835
rect 13737 12801 13771 12835
rect 13771 12801 13780 12835
rect 13728 12792 13780 12801
rect 15752 12928 15804 12980
rect 16028 12928 16080 12980
rect 16304 12928 16356 12980
rect 16764 12928 16816 12980
rect 17776 12928 17828 12980
rect 18972 12971 19024 12980
rect 18972 12937 18981 12971
rect 18981 12937 19015 12971
rect 19015 12937 19024 12971
rect 18972 12928 19024 12937
rect 20168 12928 20220 12980
rect 15476 12860 15528 12912
rect 16856 12860 16908 12912
rect 13636 12724 13688 12776
rect 16120 12792 16172 12844
rect 16396 12792 16448 12844
rect 14372 12767 14424 12776
rect 14372 12733 14406 12767
rect 14406 12733 14424 12767
rect 14372 12724 14424 12733
rect 2964 12656 3016 12708
rect 6184 12699 6236 12708
rect 2504 12588 2556 12640
rect 6184 12665 6193 12699
rect 6193 12665 6227 12699
rect 6227 12665 6236 12699
rect 6184 12656 6236 12665
rect 16672 12724 16724 12776
rect 19156 12860 19208 12912
rect 19340 12860 19392 12912
rect 17500 12835 17552 12844
rect 17500 12801 17509 12835
rect 17509 12801 17543 12835
rect 17543 12801 17552 12835
rect 17500 12792 17552 12801
rect 17868 12792 17920 12844
rect 19432 12792 19484 12844
rect 20168 12792 20220 12844
rect 20260 12724 20312 12776
rect 5080 12631 5132 12640
rect 5080 12597 5089 12631
rect 5089 12597 5123 12631
rect 5123 12597 5132 12631
rect 5080 12588 5132 12597
rect 5816 12588 5868 12640
rect 6552 12588 6604 12640
rect 12992 12588 13044 12640
rect 15568 12656 15620 12708
rect 17316 12699 17368 12708
rect 17316 12665 17325 12699
rect 17325 12665 17359 12699
rect 17359 12665 17368 12699
rect 17316 12656 17368 12665
rect 17592 12656 17644 12708
rect 19524 12656 19576 12708
rect 14004 12588 14056 12640
rect 15476 12631 15528 12640
rect 15476 12597 15485 12631
rect 15485 12597 15519 12631
rect 15519 12597 15528 12631
rect 15476 12588 15528 12597
rect 15844 12588 15896 12640
rect 16120 12588 16172 12640
rect 16672 12588 16724 12640
rect 18972 12588 19024 12640
rect 19984 12631 20036 12640
rect 19984 12597 19993 12631
rect 19993 12597 20027 12631
rect 20027 12597 20036 12631
rect 19984 12588 20036 12597
rect 20904 12656 20956 12708
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 2964 12427 3016 12436
rect 2964 12393 2973 12427
rect 2973 12393 3007 12427
rect 3007 12393 3016 12427
rect 2964 12384 3016 12393
rect 4068 12384 4120 12436
rect 11888 12384 11940 12436
rect 1492 12248 1544 12300
rect 2596 12316 2648 12368
rect 5448 12316 5500 12368
rect 10600 12359 10652 12368
rect 2320 12248 2372 12300
rect 3976 12248 4028 12300
rect 2596 12180 2648 12232
rect 4068 12180 4120 12232
rect 4528 12223 4580 12232
rect 4528 12189 4537 12223
rect 4537 12189 4571 12223
rect 4571 12189 4580 12223
rect 4528 12180 4580 12189
rect 5264 12044 5316 12096
rect 6184 12223 6236 12232
rect 6184 12189 6193 12223
rect 6193 12189 6227 12223
rect 6227 12189 6236 12223
rect 6184 12180 6236 12189
rect 9312 12248 9364 12300
rect 10600 12325 10609 12359
rect 10609 12325 10643 12359
rect 10643 12325 10652 12359
rect 10600 12316 10652 12325
rect 10876 12316 10928 12368
rect 12348 12316 12400 12368
rect 13636 12384 13688 12436
rect 15292 12427 15344 12436
rect 15292 12393 15301 12427
rect 15301 12393 15335 12427
rect 15335 12393 15344 12427
rect 15292 12384 15344 12393
rect 10784 12248 10836 12300
rect 7840 12223 7892 12232
rect 7840 12189 7849 12223
rect 7849 12189 7883 12223
rect 7883 12189 7892 12223
rect 7840 12180 7892 12189
rect 6092 12044 6144 12096
rect 6460 12044 6512 12096
rect 7196 12044 7248 12096
rect 12440 12248 12492 12300
rect 14464 12316 14516 12368
rect 15568 12316 15620 12368
rect 17500 12384 17552 12436
rect 19616 12427 19668 12436
rect 19616 12393 19625 12427
rect 19625 12393 19659 12427
rect 19659 12393 19668 12427
rect 19616 12384 19668 12393
rect 19984 12427 20036 12436
rect 19984 12393 19993 12427
rect 19993 12393 20027 12427
rect 20027 12393 20036 12427
rect 19984 12384 20036 12393
rect 20904 12427 20956 12436
rect 20904 12393 20913 12427
rect 20913 12393 20947 12427
rect 20947 12393 20956 12427
rect 20904 12384 20956 12393
rect 18512 12316 18564 12368
rect 11152 12180 11204 12232
rect 12716 12180 12768 12232
rect 16120 12248 16172 12300
rect 17040 12248 17092 12300
rect 10968 12112 11020 12164
rect 9220 12087 9272 12096
rect 9220 12053 9229 12087
rect 9229 12053 9263 12087
rect 9263 12053 9272 12087
rect 9220 12044 9272 12053
rect 14280 12044 14332 12096
rect 15476 12044 15528 12096
rect 16396 12180 16448 12232
rect 16396 12044 16448 12096
rect 19616 12248 19668 12300
rect 19340 12180 19392 12232
rect 20168 12223 20220 12232
rect 20168 12189 20177 12223
rect 20177 12189 20211 12223
rect 20211 12189 20220 12223
rect 20168 12180 20220 12189
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 1400 11840 1452 11892
rect 3608 11840 3660 11892
rect 2320 11772 2372 11824
rect 2964 11704 3016 11756
rect 3424 11772 3476 11824
rect 9220 11840 9272 11892
rect 11796 11840 11848 11892
rect 11888 11840 11940 11892
rect 5264 11704 5316 11756
rect 5448 11747 5500 11756
rect 5448 11713 5457 11747
rect 5457 11713 5491 11747
rect 5491 11713 5500 11747
rect 5448 11704 5500 11713
rect 9312 11772 9364 11824
rect 15108 11840 15160 11892
rect 15568 11840 15620 11892
rect 15752 11883 15804 11892
rect 15752 11849 15761 11883
rect 15761 11849 15795 11883
rect 15795 11849 15804 11883
rect 15752 11840 15804 11849
rect 9956 11704 10008 11756
rect 10416 11704 10468 11756
rect 10784 11747 10836 11756
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 10784 11704 10836 11713
rect 10876 11704 10928 11756
rect 15660 11772 15712 11824
rect 3148 11679 3200 11688
rect 3148 11645 3157 11679
rect 3157 11645 3191 11679
rect 3191 11645 3200 11679
rect 3148 11636 3200 11645
rect 8208 11636 8260 11688
rect 8392 11636 8444 11688
rect 8852 11636 8904 11688
rect 9404 11636 9456 11688
rect 10968 11636 11020 11688
rect 14464 11704 14516 11756
rect 15568 11704 15620 11756
rect 16396 11840 16448 11892
rect 17040 11840 17092 11892
rect 19248 11840 19300 11892
rect 17776 11772 17828 11824
rect 18972 11704 19024 11756
rect 19984 11747 20036 11756
rect 19984 11713 19993 11747
rect 19993 11713 20027 11747
rect 20027 11713 20036 11747
rect 19984 11704 20036 11713
rect 20352 11704 20404 11756
rect 2136 11543 2188 11552
rect 2136 11509 2145 11543
rect 2145 11509 2179 11543
rect 2179 11509 2188 11543
rect 2136 11500 2188 11509
rect 3976 11500 4028 11552
rect 5172 11543 5224 11552
rect 5172 11509 5181 11543
rect 5181 11509 5215 11543
rect 5215 11509 5224 11543
rect 5172 11500 5224 11509
rect 6736 11500 6788 11552
rect 7012 11543 7064 11552
rect 7012 11509 7021 11543
rect 7021 11509 7055 11543
rect 7055 11509 7064 11543
rect 7012 11500 7064 11509
rect 9588 11500 9640 11552
rect 9772 11500 9824 11552
rect 9956 11500 10008 11552
rect 11888 11568 11940 11620
rect 12348 11568 12400 11620
rect 13636 11636 13688 11688
rect 13912 11636 13964 11688
rect 11704 11500 11756 11552
rect 13912 11500 13964 11552
rect 15016 11568 15068 11620
rect 15384 11636 15436 11688
rect 16120 11679 16172 11688
rect 16120 11645 16129 11679
rect 16129 11645 16163 11679
rect 16163 11645 16172 11679
rect 16120 11636 16172 11645
rect 16764 11636 16816 11688
rect 15844 11568 15896 11620
rect 15292 11500 15344 11552
rect 16488 11568 16540 11620
rect 19524 11568 19576 11620
rect 19616 11568 19668 11620
rect 20168 11568 20220 11620
rect 18604 11543 18656 11552
rect 18604 11509 18613 11543
rect 18613 11509 18647 11543
rect 18647 11509 18656 11543
rect 18604 11500 18656 11509
rect 18788 11500 18840 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 2320 11296 2372 11348
rect 5172 11296 5224 11348
rect 6000 11296 6052 11348
rect 6736 11339 6788 11348
rect 6736 11305 6745 11339
rect 6745 11305 6779 11339
rect 6779 11305 6788 11339
rect 6736 11296 6788 11305
rect 6368 11228 6420 11280
rect 1492 11203 1544 11212
rect 1492 11169 1501 11203
rect 1501 11169 1535 11203
rect 1535 11169 1544 11203
rect 1492 11160 1544 11169
rect 2596 11160 2648 11212
rect 4068 11203 4120 11212
rect 4068 11169 4077 11203
rect 4077 11169 4111 11203
rect 4111 11169 4120 11203
rect 4068 11160 4120 11169
rect 6092 11203 6144 11212
rect 3148 11135 3200 11144
rect 3148 11101 3157 11135
rect 3157 11101 3191 11135
rect 3191 11101 3200 11135
rect 3148 11092 3200 11101
rect 5080 11092 5132 11144
rect 6092 11169 6101 11203
rect 6101 11169 6135 11203
rect 6135 11169 6144 11203
rect 6092 11160 6144 11169
rect 8300 11160 8352 11212
rect 6920 11092 6972 11144
rect 5448 11067 5500 11076
rect 5448 11033 5457 11067
rect 5457 11033 5491 11067
rect 5491 11033 5500 11067
rect 5448 11024 5500 11033
rect 9404 11296 9456 11348
rect 9220 11228 9272 11280
rect 9588 11228 9640 11280
rect 16028 11296 16080 11348
rect 17316 11296 17368 11348
rect 17960 11296 18012 11348
rect 18788 11339 18840 11348
rect 18788 11305 18797 11339
rect 18797 11305 18831 11339
rect 18831 11305 18840 11339
rect 18788 11296 18840 11305
rect 20076 11296 20128 11348
rect 9956 11160 10008 11212
rect 10048 11160 10100 11212
rect 10692 11160 10744 11212
rect 9772 11092 9824 11144
rect 10140 11092 10192 11144
rect 10508 11092 10560 11144
rect 10968 11135 11020 11144
rect 10968 11101 10977 11135
rect 10977 11101 11011 11135
rect 11011 11101 11020 11135
rect 10968 11092 11020 11101
rect 11704 11092 11756 11144
rect 12992 11228 13044 11280
rect 14096 11228 14148 11280
rect 12716 11092 12768 11144
rect 12992 11135 13044 11144
rect 12992 11101 13001 11135
rect 13001 11101 13035 11135
rect 13035 11101 13044 11135
rect 12992 11092 13044 11101
rect 13268 11092 13320 11144
rect 13728 11092 13780 11144
rect 13912 11135 13964 11144
rect 13912 11101 13921 11135
rect 13921 11101 13955 11135
rect 13955 11101 13964 11135
rect 13912 11092 13964 11101
rect 14188 11092 14240 11144
rect 9680 11024 9732 11076
rect 12624 11024 12676 11076
rect 15292 11203 15344 11212
rect 15292 11169 15301 11203
rect 15301 11169 15335 11203
rect 15335 11169 15344 11203
rect 15292 11160 15344 11169
rect 15384 11160 15436 11212
rect 19064 11228 19116 11280
rect 20904 11228 20956 11280
rect 17500 11135 17552 11144
rect 17500 11101 17509 11135
rect 17509 11101 17543 11135
rect 17543 11101 17552 11135
rect 17500 11092 17552 11101
rect 15108 11024 15160 11076
rect 16488 11024 16540 11076
rect 17960 11135 18012 11144
rect 17960 11101 17969 11135
rect 17969 11101 18003 11135
rect 18003 11101 18012 11135
rect 17960 11092 18012 11101
rect 18972 11135 19024 11144
rect 18972 11101 18981 11135
rect 18981 11101 19015 11135
rect 19015 11101 19024 11135
rect 18972 11092 19024 11101
rect 19984 11135 20036 11144
rect 19984 11101 19993 11135
rect 19993 11101 20027 11135
rect 20027 11101 20036 11135
rect 19984 11092 20036 11101
rect 18696 11024 18748 11076
rect 3240 10956 3292 11008
rect 10232 10956 10284 11008
rect 11888 10956 11940 11008
rect 12532 10956 12584 11008
rect 16764 10956 16816 11008
rect 16948 10999 17000 11008
rect 16948 10965 16957 10999
rect 16957 10965 16991 10999
rect 16991 10965 17000 10999
rect 16948 10956 17000 10965
rect 18880 10956 18932 11008
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 2136 10752 2188 10804
rect 3976 10795 4028 10804
rect 3976 10761 3985 10795
rect 3985 10761 4019 10795
rect 4019 10761 4028 10795
rect 3976 10752 4028 10761
rect 4712 10752 4764 10804
rect 4988 10752 5040 10804
rect 7012 10752 7064 10804
rect 3424 10684 3476 10736
rect 4068 10684 4120 10736
rect 12164 10752 12216 10804
rect 12532 10752 12584 10804
rect 15016 10752 15068 10804
rect 11796 10684 11848 10736
rect 2320 10659 2372 10668
rect 2320 10625 2329 10659
rect 2329 10625 2363 10659
rect 2363 10625 2372 10659
rect 2320 10616 2372 10625
rect 2596 10616 2648 10668
rect 3516 10616 3568 10668
rect 3976 10616 4028 10668
rect 5448 10616 5500 10668
rect 5632 10659 5684 10668
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 7104 10616 7156 10668
rect 7472 10616 7524 10668
rect 7748 10616 7800 10668
rect 8208 10616 8260 10668
rect 9220 10659 9272 10668
rect 9220 10625 9229 10659
rect 9229 10625 9263 10659
rect 9263 10625 9272 10659
rect 9220 10616 9272 10625
rect 9312 10659 9364 10668
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 12624 10616 12676 10668
rect 3148 10591 3200 10600
rect 3148 10557 3157 10591
rect 3157 10557 3191 10591
rect 3191 10557 3200 10591
rect 3148 10548 3200 10557
rect 3424 10548 3476 10600
rect 1952 10412 2004 10464
rect 10968 10591 11020 10600
rect 10968 10557 11002 10591
rect 11002 10557 11020 10591
rect 10968 10548 11020 10557
rect 12348 10548 12400 10600
rect 13084 10616 13136 10668
rect 15476 10659 15528 10668
rect 15476 10625 15485 10659
rect 15485 10625 15519 10659
rect 15519 10625 15528 10659
rect 15476 10616 15528 10625
rect 16488 10684 16540 10736
rect 18604 10752 18656 10804
rect 19524 10795 19576 10804
rect 19524 10761 19533 10795
rect 19533 10761 19567 10795
rect 19567 10761 19576 10795
rect 19524 10752 19576 10761
rect 19800 10684 19852 10736
rect 16856 10616 16908 10668
rect 16948 10548 17000 10600
rect 17500 10616 17552 10668
rect 19984 10616 20036 10668
rect 19156 10548 19208 10600
rect 19800 10548 19852 10600
rect 3148 10412 3200 10464
rect 3700 10412 3752 10464
rect 4160 10412 4212 10464
rect 4804 10412 4856 10464
rect 5356 10455 5408 10464
rect 5356 10421 5365 10455
rect 5365 10421 5399 10455
rect 5399 10421 5408 10455
rect 5356 10412 5408 10421
rect 6000 10455 6052 10464
rect 6000 10421 6009 10455
rect 6009 10421 6043 10455
rect 6043 10421 6052 10455
rect 6000 10412 6052 10421
rect 7472 10455 7524 10464
rect 7472 10421 7481 10455
rect 7481 10421 7515 10455
rect 7515 10421 7524 10455
rect 7472 10412 7524 10421
rect 7564 10412 7616 10464
rect 8484 10455 8536 10464
rect 8484 10421 8493 10455
rect 8493 10421 8527 10455
rect 8527 10421 8536 10455
rect 8484 10412 8536 10421
rect 11152 10480 11204 10532
rect 9128 10455 9180 10464
rect 9128 10421 9137 10455
rect 9137 10421 9171 10455
rect 9171 10421 9180 10455
rect 9128 10412 9180 10421
rect 11796 10412 11848 10464
rect 12992 10412 13044 10464
rect 13636 10480 13688 10532
rect 16212 10480 16264 10532
rect 18604 10480 18656 10532
rect 20076 10480 20128 10532
rect 20444 10480 20496 10532
rect 20720 10480 20772 10532
rect 13544 10412 13596 10464
rect 13912 10455 13964 10464
rect 13912 10421 13921 10455
rect 13921 10421 13955 10455
rect 13955 10421 13964 10455
rect 13912 10412 13964 10421
rect 18420 10412 18472 10464
rect 18512 10412 18564 10464
rect 18788 10412 18840 10464
rect 19524 10412 19576 10464
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 1952 10251 2004 10260
rect 1952 10217 1961 10251
rect 1961 10217 1995 10251
rect 1995 10217 2004 10251
rect 1952 10208 2004 10217
rect 3424 10251 3476 10260
rect 3424 10217 3433 10251
rect 3433 10217 3467 10251
rect 3467 10217 3476 10251
rect 3424 10208 3476 10217
rect 4160 10251 4212 10260
rect 4160 10217 4169 10251
rect 4169 10217 4203 10251
rect 4203 10217 4212 10251
rect 4160 10208 4212 10217
rect 6000 10208 6052 10260
rect 6920 10251 6972 10260
rect 6920 10217 6929 10251
rect 6929 10217 6963 10251
rect 6963 10217 6972 10251
rect 6920 10208 6972 10217
rect 7288 10208 7340 10260
rect 7748 10208 7800 10260
rect 8484 10208 8536 10260
rect 8668 10208 8720 10260
rect 9128 10208 9180 10260
rect 9864 10208 9916 10260
rect 12992 10208 13044 10260
rect 13544 10208 13596 10260
rect 13912 10208 13964 10260
rect 14280 10208 14332 10260
rect 17500 10208 17552 10260
rect 4712 10140 4764 10192
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 2320 10115 2372 10124
rect 2320 10081 2329 10115
rect 2329 10081 2363 10115
rect 2363 10081 2372 10115
rect 2320 10072 2372 10081
rect 2596 10047 2648 10056
rect 2596 10013 2605 10047
rect 2605 10013 2639 10047
rect 2639 10013 2648 10047
rect 2596 10004 2648 10013
rect 7472 10140 7524 10192
rect 5540 10115 5592 10124
rect 3516 10004 3568 10056
rect 4620 10004 4672 10056
rect 5080 10004 5132 10056
rect 2872 9936 2924 9988
rect 4344 9936 4396 9988
rect 5540 10081 5549 10115
rect 5549 10081 5583 10115
rect 5583 10081 5592 10115
rect 5540 10072 5592 10081
rect 5632 10072 5684 10124
rect 6184 10072 6236 10124
rect 6368 10072 6420 10124
rect 7748 10072 7800 10124
rect 9772 10072 9824 10124
rect 10600 10072 10652 10124
rect 11796 10140 11848 10192
rect 18052 10140 18104 10192
rect 14096 10115 14148 10124
rect 14096 10081 14105 10115
rect 14105 10081 14139 10115
rect 14139 10081 14148 10115
rect 15108 10115 15160 10124
rect 14096 10072 14148 10081
rect 15108 10081 15117 10115
rect 15117 10081 15151 10115
rect 15151 10081 15160 10115
rect 15108 10072 15160 10081
rect 15292 10072 15344 10124
rect 7932 10047 7984 10056
rect 7932 10013 7941 10047
rect 7941 10013 7975 10047
rect 7975 10013 7984 10047
rect 7932 10004 7984 10013
rect 11336 10047 11388 10056
rect 11336 10013 11345 10047
rect 11345 10013 11379 10047
rect 11379 10013 11388 10047
rect 11336 10004 11388 10013
rect 12440 10004 12492 10056
rect 13636 10004 13688 10056
rect 14188 10047 14240 10056
rect 14188 10013 14197 10047
rect 14197 10013 14231 10047
rect 14231 10013 14240 10047
rect 14188 10004 14240 10013
rect 15752 10047 15804 10056
rect 15752 10013 15761 10047
rect 15761 10013 15795 10047
rect 15795 10013 15804 10047
rect 15752 10004 15804 10013
rect 16212 10072 16264 10124
rect 16120 10004 16172 10056
rect 16304 10047 16356 10056
rect 16304 10013 16313 10047
rect 16313 10013 16347 10047
rect 16347 10013 16356 10047
rect 16304 10004 16356 10013
rect 3608 9868 3660 9920
rect 5448 9868 5500 9920
rect 15384 9936 15436 9988
rect 7012 9868 7064 9920
rect 8208 9868 8260 9920
rect 9312 9911 9364 9920
rect 9312 9877 9321 9911
rect 9321 9877 9355 9911
rect 9355 9877 9364 9911
rect 9312 9868 9364 9877
rect 12348 9868 12400 9920
rect 18880 10208 18932 10260
rect 19248 10208 19300 10260
rect 19340 10140 19392 10192
rect 18420 10072 18472 10124
rect 18880 10072 18932 10124
rect 20352 10047 20404 10056
rect 20076 9936 20128 9988
rect 20352 10013 20361 10047
rect 20361 10013 20395 10047
rect 20395 10013 20404 10047
rect 20352 10004 20404 10013
rect 19708 9911 19760 9920
rect 19708 9877 19717 9911
rect 19717 9877 19751 9911
rect 19751 9877 19760 9911
rect 19708 9868 19760 9877
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 3148 9664 3200 9716
rect 1860 9528 1912 9580
rect 5080 9571 5132 9580
rect 2228 9460 2280 9512
rect 2872 9392 2924 9444
rect 3148 9392 3200 9444
rect 3424 9460 3476 9512
rect 4804 9503 4856 9512
rect 4804 9469 4813 9503
rect 4813 9469 4847 9503
rect 4847 9469 4856 9503
rect 4804 9460 4856 9469
rect 5080 9537 5089 9571
rect 5089 9537 5123 9571
rect 5123 9537 5132 9571
rect 5080 9528 5132 9537
rect 6184 9528 6236 9580
rect 7564 9528 7616 9580
rect 7932 9664 7984 9716
rect 7472 9460 7524 9512
rect 12992 9664 13044 9716
rect 16212 9707 16264 9716
rect 14280 9596 14332 9648
rect 16212 9673 16221 9707
rect 16221 9673 16255 9707
rect 16255 9673 16264 9707
rect 16212 9664 16264 9673
rect 18512 9664 18564 9716
rect 19248 9664 19300 9716
rect 16396 9596 16448 9648
rect 10876 9528 10928 9580
rect 13084 9571 13136 9580
rect 13084 9537 13093 9571
rect 13093 9537 13127 9571
rect 13127 9537 13136 9571
rect 13084 9528 13136 9537
rect 16948 9528 17000 9580
rect 17408 9596 17460 9648
rect 19340 9596 19392 9648
rect 19432 9596 19484 9648
rect 20536 9596 20588 9648
rect 18696 9571 18748 9580
rect 18696 9537 18705 9571
rect 18705 9537 18739 9571
rect 18739 9537 18748 9571
rect 18696 9528 18748 9537
rect 18972 9528 19024 9580
rect 3608 9392 3660 9444
rect 4068 9392 4120 9444
rect 8208 9392 8260 9444
rect 8668 9392 8720 9444
rect 12348 9460 12400 9512
rect 10232 9392 10284 9444
rect 13268 9460 13320 9512
rect 15384 9460 15436 9512
rect 15936 9460 15988 9512
rect 12624 9392 12676 9444
rect 15016 9392 15068 9444
rect 5632 9324 5684 9376
rect 5908 9324 5960 9376
rect 6736 9324 6788 9376
rect 10968 9324 11020 9376
rect 12532 9324 12584 9376
rect 17960 9460 18012 9512
rect 18052 9392 18104 9444
rect 20352 9528 20404 9580
rect 16488 9367 16540 9376
rect 16488 9333 16497 9367
rect 16497 9333 16531 9367
rect 16531 9333 16540 9367
rect 16488 9324 16540 9333
rect 16672 9324 16724 9376
rect 19892 9367 19944 9376
rect 19892 9333 19901 9367
rect 19901 9333 19935 9367
rect 19935 9333 19944 9367
rect 19892 9324 19944 9333
rect 20260 9367 20312 9376
rect 20260 9333 20269 9367
rect 20269 9333 20303 9367
rect 20303 9333 20312 9367
rect 20260 9324 20312 9333
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 2228 9163 2280 9172
rect 2228 9129 2237 9163
rect 2237 9129 2271 9163
rect 2271 9129 2280 9163
rect 2228 9120 2280 9129
rect 4712 9120 4764 9172
rect 5172 9120 5224 9172
rect 6092 9120 6144 9172
rect 7288 9163 7340 9172
rect 7288 9129 7297 9163
rect 7297 9129 7331 9163
rect 7331 9129 7340 9163
rect 7288 9120 7340 9129
rect 7472 9120 7524 9172
rect 8300 9163 8352 9172
rect 8300 9129 8309 9163
rect 8309 9129 8343 9163
rect 8343 9129 8352 9163
rect 8300 9120 8352 9129
rect 8576 9120 8628 9172
rect 3976 9052 4028 9104
rect 2596 9027 2648 9036
rect 2596 8993 2605 9027
rect 2605 8993 2639 9027
rect 2639 8993 2648 9027
rect 2596 8984 2648 8993
rect 3700 8984 3752 9036
rect 1400 8916 1452 8968
rect 2872 8959 2924 8968
rect 2872 8925 2881 8959
rect 2881 8925 2915 8959
rect 2915 8925 2924 8959
rect 2872 8916 2924 8925
rect 4160 8916 4212 8968
rect 5172 8984 5224 9036
rect 5908 9027 5960 9036
rect 5908 8993 5917 9027
rect 5917 8993 5951 9027
rect 5951 8993 5960 9027
rect 5908 8984 5960 8993
rect 6644 8984 6696 9036
rect 10232 9120 10284 9172
rect 10876 9163 10928 9172
rect 10876 9129 10885 9163
rect 10885 9129 10919 9163
rect 10919 9129 10928 9163
rect 10876 9120 10928 9129
rect 11704 9120 11756 9172
rect 12164 9120 12216 9172
rect 15016 9163 15068 9172
rect 15016 9129 15025 9163
rect 15025 9129 15059 9163
rect 15059 9129 15068 9163
rect 15016 9120 15068 9129
rect 15292 9163 15344 9172
rect 15292 9129 15301 9163
rect 15301 9129 15335 9163
rect 15335 9129 15344 9163
rect 15292 9120 15344 9129
rect 16580 9120 16632 9172
rect 16764 9120 16816 9172
rect 19800 9163 19852 9172
rect 19800 9129 19809 9163
rect 19809 9129 19843 9163
rect 19843 9129 19852 9163
rect 19800 9120 19852 9129
rect 20260 9120 20312 9172
rect 10048 9095 10100 9104
rect 10048 9061 10057 9095
rect 10057 9061 10091 9095
rect 10091 9061 10100 9095
rect 10048 9052 10100 9061
rect 10140 9095 10192 9104
rect 10140 9061 10149 9095
rect 10149 9061 10183 9095
rect 10183 9061 10192 9095
rect 10140 9052 10192 9061
rect 11980 9052 12032 9104
rect 12808 9052 12860 9104
rect 12992 9052 13044 9104
rect 5448 8959 5500 8968
rect 5448 8925 5457 8959
rect 5457 8925 5491 8959
rect 5491 8925 5500 8959
rect 5448 8916 5500 8925
rect 6184 8959 6236 8968
rect 6184 8925 6193 8959
rect 6193 8925 6227 8959
rect 6227 8925 6236 8959
rect 6184 8916 6236 8925
rect 7840 8959 7892 8968
rect 7840 8925 7849 8959
rect 7849 8925 7883 8959
rect 7883 8925 7892 8959
rect 10876 8984 10928 9036
rect 12900 8984 12952 9036
rect 13084 8984 13136 9036
rect 7840 8916 7892 8925
rect 3240 8848 3292 8900
rect 4804 8848 4856 8900
rect 5908 8848 5960 8900
rect 6828 8848 6880 8900
rect 9680 8891 9732 8900
rect 4712 8780 4764 8832
rect 7196 8780 7248 8832
rect 9680 8857 9689 8891
rect 9689 8857 9723 8891
rect 9723 8857 9732 8891
rect 9680 8848 9732 8857
rect 11888 8959 11940 8968
rect 11888 8925 11897 8959
rect 11897 8925 11931 8959
rect 11931 8925 11940 8959
rect 11888 8916 11940 8925
rect 11796 8848 11848 8900
rect 11152 8780 11204 8832
rect 16488 9052 16540 9104
rect 18328 9052 18380 9104
rect 18696 9052 18748 9104
rect 18880 9052 18932 9104
rect 19064 9052 19116 9104
rect 12256 8780 12308 8832
rect 17776 8984 17828 9036
rect 19340 8984 19392 9036
rect 19432 8984 19484 9036
rect 15384 8916 15436 8968
rect 16304 8916 16356 8968
rect 16580 8916 16632 8968
rect 16948 8959 17000 8968
rect 16948 8925 16957 8959
rect 16957 8925 16991 8959
rect 16991 8925 17000 8959
rect 16948 8916 17000 8925
rect 17868 8916 17920 8968
rect 19524 8916 19576 8968
rect 20260 8959 20312 8968
rect 20260 8925 20269 8959
rect 20269 8925 20303 8959
rect 20303 8925 20312 8959
rect 20260 8916 20312 8925
rect 15108 8780 15160 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 2872 8576 2924 8628
rect 3240 8619 3292 8628
rect 3240 8585 3249 8619
rect 3249 8585 3283 8619
rect 3283 8585 3292 8619
rect 3240 8576 3292 8585
rect 4068 8576 4120 8628
rect 12440 8576 12492 8628
rect 15752 8576 15804 8628
rect 4712 8483 4764 8492
rect 1584 8415 1636 8424
rect 1584 8381 1593 8415
rect 1593 8381 1627 8415
rect 1627 8381 1636 8415
rect 1584 8372 1636 8381
rect 3792 8304 3844 8356
rect 4712 8449 4721 8483
rect 4721 8449 4755 8483
rect 4755 8449 4764 8483
rect 4712 8440 4764 8449
rect 5356 8440 5408 8492
rect 7104 8440 7156 8492
rect 8208 8483 8260 8492
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 8208 8440 8260 8449
rect 6552 8372 6604 8424
rect 8668 8415 8720 8424
rect 3976 8304 4028 8356
rect 3608 8279 3660 8288
rect 3608 8245 3617 8279
rect 3617 8245 3651 8279
rect 3651 8245 3660 8279
rect 3608 8236 3660 8245
rect 4804 8304 4856 8356
rect 5172 8304 5224 8356
rect 6184 8304 6236 8356
rect 8668 8381 8677 8415
rect 8677 8381 8711 8415
rect 8711 8381 8720 8415
rect 8668 8372 8720 8381
rect 10968 8440 11020 8492
rect 12256 8440 12308 8492
rect 15384 8483 15436 8492
rect 15384 8449 15393 8483
rect 15393 8449 15427 8483
rect 15427 8449 15436 8483
rect 15384 8440 15436 8449
rect 16948 8440 17000 8492
rect 19340 8576 19392 8628
rect 20260 8576 20312 8628
rect 20628 8576 20680 8628
rect 19984 8508 20036 8560
rect 11980 8372 12032 8424
rect 12532 8372 12584 8424
rect 16396 8372 16448 8424
rect 16580 8372 16632 8424
rect 17868 8372 17920 8424
rect 5356 8236 5408 8288
rect 6920 8304 6972 8356
rect 7656 8304 7708 8356
rect 8024 8347 8076 8356
rect 8024 8313 8033 8347
rect 8033 8313 8067 8347
rect 8067 8313 8076 8347
rect 8024 8304 8076 8313
rect 8576 8304 8628 8356
rect 8852 8304 8904 8356
rect 11796 8347 11848 8356
rect 11796 8313 11805 8347
rect 11805 8313 11839 8347
rect 11839 8313 11848 8347
rect 11796 8304 11848 8313
rect 15108 8304 15160 8356
rect 8208 8236 8260 8288
rect 9220 8236 9272 8288
rect 10324 8279 10376 8288
rect 10324 8245 10333 8279
rect 10333 8245 10367 8279
rect 10367 8245 10376 8279
rect 10324 8236 10376 8245
rect 10692 8279 10744 8288
rect 10692 8245 10701 8279
rect 10701 8245 10735 8279
rect 10735 8245 10744 8279
rect 10692 8236 10744 8245
rect 12900 8236 12952 8288
rect 16028 8304 16080 8356
rect 16764 8304 16816 8356
rect 18144 8304 18196 8356
rect 19708 8372 19760 8424
rect 20720 8415 20772 8424
rect 20720 8381 20729 8415
rect 20729 8381 20763 8415
rect 20763 8381 20772 8415
rect 20720 8372 20772 8381
rect 20352 8304 20404 8356
rect 17408 8279 17460 8288
rect 17408 8245 17417 8279
rect 17417 8245 17451 8279
rect 17451 8245 17460 8279
rect 17408 8236 17460 8245
rect 18236 8236 18288 8288
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 3608 8032 3660 8084
rect 4252 8032 4304 8084
rect 6920 8032 6972 8084
rect 7104 8075 7156 8084
rect 7104 8041 7113 8075
rect 7113 8041 7147 8075
rect 7147 8041 7156 8075
rect 7104 8032 7156 8041
rect 8668 8032 8720 8084
rect 9220 8075 9272 8084
rect 9220 8041 9229 8075
rect 9229 8041 9263 8075
rect 9263 8041 9272 8075
rect 9220 8032 9272 8041
rect 10692 8032 10744 8084
rect 12164 8032 12216 8084
rect 1584 7828 1636 7880
rect 3148 7964 3200 8016
rect 3976 7964 4028 8016
rect 12624 8032 12676 8084
rect 12992 8032 13044 8084
rect 18144 8032 18196 8084
rect 19432 8075 19484 8084
rect 19432 8041 19441 8075
rect 19441 8041 19475 8075
rect 19475 8041 19484 8075
rect 19432 8032 19484 8041
rect 19892 8032 19944 8084
rect 3608 7896 3660 7948
rect 3792 7760 3844 7812
rect 4988 7896 5040 7948
rect 5448 7896 5500 7948
rect 6368 7896 6420 7948
rect 8116 7939 8168 7948
rect 8116 7905 8150 7939
rect 8150 7905 8168 7939
rect 8116 7896 8168 7905
rect 10416 7896 10468 7948
rect 15568 7896 15620 7948
rect 17960 7896 18012 7948
rect 18788 7939 18840 7948
rect 18788 7905 18797 7939
rect 18797 7905 18831 7939
rect 18831 7905 18840 7939
rect 18788 7896 18840 7905
rect 18880 7939 18932 7948
rect 18880 7905 18889 7939
rect 18889 7905 18923 7939
rect 18923 7905 18932 7939
rect 18880 7896 18932 7905
rect 4712 7871 4764 7880
rect 4712 7837 4721 7871
rect 4721 7837 4755 7871
rect 4755 7837 4764 7871
rect 4712 7828 4764 7837
rect 5264 7760 5316 7812
rect 6920 7828 6972 7880
rect 8852 7828 8904 7880
rect 10968 7871 11020 7880
rect 10968 7837 10977 7871
rect 10977 7837 11011 7871
rect 11011 7837 11020 7871
rect 12900 7871 12952 7880
rect 10968 7828 11020 7837
rect 12900 7837 12909 7871
rect 12909 7837 12943 7871
rect 12943 7837 12952 7871
rect 12900 7828 12952 7837
rect 16580 7828 16632 7880
rect 18972 7871 19024 7880
rect 18972 7837 18981 7871
rect 18981 7837 19015 7871
rect 19015 7837 19024 7871
rect 18972 7828 19024 7837
rect 19892 7871 19944 7880
rect 19892 7837 19901 7871
rect 19901 7837 19935 7871
rect 19935 7837 19944 7871
rect 19892 7828 19944 7837
rect 19984 7871 20036 7880
rect 19984 7837 19993 7871
rect 19993 7837 20027 7871
rect 20027 7837 20036 7871
rect 19984 7828 20036 7837
rect 18236 7760 18288 7812
rect 4068 7692 4120 7744
rect 15200 7692 15252 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 2596 7488 2648 7540
rect 3148 7488 3200 7540
rect 5264 7488 5316 7540
rect 6368 7531 6420 7540
rect 6368 7497 6377 7531
rect 6377 7497 6411 7531
rect 6411 7497 6420 7531
rect 6368 7488 6420 7497
rect 8116 7488 8168 7540
rect 8576 7531 8628 7540
rect 3792 7352 3844 7404
rect 4712 7352 4764 7404
rect 6920 7395 6972 7404
rect 6920 7361 6929 7395
rect 6929 7361 6963 7395
rect 6963 7361 6972 7395
rect 6920 7352 6972 7361
rect 8576 7497 8585 7531
rect 8585 7497 8619 7531
rect 8619 7497 8628 7531
rect 8576 7488 8628 7497
rect 17408 7488 17460 7540
rect 19892 7488 19944 7540
rect 11704 7420 11756 7472
rect 17960 7352 18012 7404
rect 5264 7327 5316 7336
rect 5264 7293 5298 7327
rect 5298 7293 5316 7327
rect 5264 7284 5316 7293
rect 9036 7284 9088 7336
rect 19800 7284 19852 7336
rect 20352 7395 20404 7404
rect 20352 7361 20361 7395
rect 20361 7361 20395 7395
rect 20395 7361 20404 7395
rect 20352 7352 20404 7361
rect 2964 7191 3016 7200
rect 2964 7157 2973 7191
rect 2973 7157 3007 7191
rect 3007 7157 3016 7191
rect 2964 7148 3016 7157
rect 3792 7216 3844 7268
rect 4160 7216 4212 7268
rect 7104 7216 7156 7268
rect 11612 7216 11664 7268
rect 3884 7191 3936 7200
rect 3884 7157 3893 7191
rect 3893 7157 3927 7191
rect 3927 7157 3936 7191
rect 3884 7148 3936 7157
rect 5356 7148 5408 7200
rect 9036 7191 9088 7200
rect 9036 7157 9045 7191
rect 9045 7157 9079 7191
rect 9079 7157 9088 7191
rect 9036 7148 9088 7157
rect 11060 7148 11112 7200
rect 20168 7148 20220 7200
rect 20444 7148 20496 7200
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 3884 6944 3936 6996
rect 1584 6851 1636 6860
rect 1584 6817 1593 6851
rect 1593 6817 1627 6851
rect 1627 6817 1636 6851
rect 1584 6808 1636 6817
rect 2228 6808 2280 6860
rect 3148 6808 3200 6860
rect 5540 6944 5592 6996
rect 6552 6987 6604 6996
rect 6552 6953 6561 6987
rect 6561 6953 6595 6987
rect 6595 6953 6604 6987
rect 6552 6944 6604 6953
rect 17960 6987 18012 6996
rect 17960 6953 17969 6987
rect 17969 6953 18003 6987
rect 18003 6953 18012 6987
rect 17960 6944 18012 6953
rect 18972 6944 19024 6996
rect 5816 6876 5868 6928
rect 6828 6876 6880 6928
rect 10416 6876 10468 6928
rect 18512 6876 18564 6928
rect 5540 6851 5592 6860
rect 5540 6817 5549 6851
rect 5549 6817 5583 6851
rect 5583 6817 5592 6851
rect 5540 6808 5592 6817
rect 4252 6740 4304 6792
rect 5264 6740 5316 6792
rect 2780 6672 2832 6724
rect 6368 6740 6420 6792
rect 6184 6715 6236 6724
rect 6184 6681 6193 6715
rect 6193 6681 6227 6715
rect 6227 6681 6236 6715
rect 6184 6672 6236 6681
rect 12072 6808 12124 6860
rect 19156 6808 19208 6860
rect 19616 6808 19668 6860
rect 8852 6740 8904 6792
rect 16580 6783 16632 6792
rect 16580 6749 16589 6783
rect 16589 6749 16623 6783
rect 16623 6749 16632 6783
rect 16580 6740 16632 6749
rect 19064 6783 19116 6792
rect 19064 6749 19073 6783
rect 19073 6749 19107 6783
rect 19107 6749 19116 6783
rect 19064 6740 19116 6749
rect 20168 6740 20220 6792
rect 10324 6672 10376 6724
rect 5172 6647 5224 6656
rect 5172 6613 5181 6647
rect 5181 6613 5215 6647
rect 5215 6613 5224 6647
rect 5172 6604 5224 6613
rect 7196 6647 7248 6656
rect 7196 6613 7205 6647
rect 7205 6613 7239 6647
rect 7239 6613 7248 6647
rect 7196 6604 7248 6613
rect 7380 6604 7432 6656
rect 17960 6604 18012 6656
rect 20628 6604 20680 6656
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 2964 6443 3016 6452
rect 2964 6409 2973 6443
rect 2973 6409 3007 6443
rect 3007 6409 3016 6443
rect 2964 6400 3016 6409
rect 5540 6400 5592 6452
rect 19156 6400 19208 6452
rect 20352 6400 20404 6452
rect 4068 6332 4120 6384
rect 7012 6332 7064 6384
rect 3608 6307 3660 6316
rect 3608 6273 3617 6307
rect 3617 6273 3651 6307
rect 3651 6273 3660 6307
rect 3608 6264 3660 6273
rect 5264 6264 5316 6316
rect 16580 6264 16632 6316
rect 19064 6264 19116 6316
rect 3976 6196 4028 6248
rect 5356 6239 5408 6248
rect 2872 6128 2924 6180
rect 3424 6171 3476 6180
rect 3424 6137 3433 6171
rect 3433 6137 3467 6171
rect 3467 6137 3476 6171
rect 3424 6128 3476 6137
rect 3240 6060 3292 6112
rect 4804 6128 4856 6180
rect 5356 6205 5365 6239
rect 5365 6205 5399 6239
rect 5399 6205 5408 6239
rect 5356 6196 5408 6205
rect 20628 6196 20680 6248
rect 10232 6128 10284 6180
rect 3700 6060 3752 6112
rect 3976 6060 4028 6112
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 19800 5899 19852 5908
rect 19800 5865 19809 5899
rect 19809 5865 19843 5899
rect 19843 5865 19852 5899
rect 19800 5856 19852 5865
rect 20168 5899 20220 5908
rect 20168 5865 20177 5899
rect 20177 5865 20211 5899
rect 20211 5865 20220 5899
rect 20168 5856 20220 5865
rect 20260 5695 20312 5704
rect 20260 5661 20269 5695
rect 20269 5661 20303 5695
rect 20303 5661 20312 5695
rect 20260 5652 20312 5661
rect 20352 5695 20404 5704
rect 20352 5661 20361 5695
rect 20361 5661 20395 5695
rect 20395 5661 20404 5695
rect 20352 5652 20404 5661
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 6092 5312 6144 5364
rect 17960 5312 18012 5364
rect 20260 5312 20312 5364
rect 4068 5244 4120 5296
rect 11704 5244 11756 5296
rect 20628 5219 20680 5228
rect 20628 5185 20637 5219
rect 20637 5185 20671 5219
rect 20671 5185 20680 5219
rect 20628 5176 20680 5185
rect 4068 4972 4120 5024
rect 20536 5015 20588 5024
rect 20536 4981 20545 5015
rect 20545 4981 20579 5015
rect 20579 4981 20588 5015
rect 20536 4972 20588 4981
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 20444 3000 20496 3052
rect 4896 2975 4948 2984
rect 4896 2941 4905 2975
rect 4905 2941 4939 2975
rect 4939 2941 4948 2975
rect 4896 2932 4948 2941
rect 11152 2932 11204 2984
rect 15844 2932 15896 2984
rect 5724 2864 5776 2916
rect 5080 2796 5132 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 2964 1300 3016 1352
rect 5908 1300 5960 1352
rect 2780 1028 2832 1080
rect 4988 1028 5040 1080
rect 3332 212 3384 264
rect 6828 212 6880 264
<< metal2 >>
rect 202 22320 258 22800
rect 570 22320 626 22800
rect 1030 22320 1086 22800
rect 1398 22320 1454 22800
rect 1858 22320 1914 22800
rect 2226 22320 2282 22800
rect 2686 22320 2742 22800
rect 3146 22320 3202 22800
rect 3238 22536 3294 22545
rect 3238 22471 3294 22480
rect 216 19242 244 22320
rect 204 19236 256 19242
rect 204 19178 256 19184
rect 584 18086 612 22320
rect 1044 18902 1072 22320
rect 1032 18896 1084 18902
rect 1032 18838 1084 18844
rect 1412 18630 1440 22320
rect 1768 19304 1820 19310
rect 1582 19272 1638 19281
rect 1768 19246 1820 19252
rect 1582 19207 1638 19216
rect 1596 18970 1624 19207
rect 1780 19145 1808 19246
rect 1766 19136 1822 19145
rect 1766 19071 1822 19080
rect 1872 19009 1900 22320
rect 2240 20670 2268 22320
rect 2228 20664 2280 20670
rect 2228 20606 2280 20612
rect 1950 19816 2006 19825
rect 1950 19751 2006 19760
rect 1964 19514 1992 19751
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 1858 19000 1914 19009
rect 1584 18964 1636 18970
rect 1858 18935 1914 18944
rect 1584 18906 1636 18912
rect 1950 18864 2006 18873
rect 1950 18799 2006 18808
rect 2136 18828 2188 18834
rect 1400 18624 1452 18630
rect 1400 18566 1452 18572
rect 1964 18426 1992 18799
rect 2136 18770 2188 18776
rect 2044 18624 2096 18630
rect 2044 18566 2096 18572
rect 2056 18426 2084 18566
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 2044 18420 2096 18426
rect 2044 18362 2096 18368
rect 2148 18290 2176 18770
rect 2240 18630 2268 20606
rect 2320 19916 2372 19922
rect 2320 19858 2372 19864
rect 2332 19446 2360 19858
rect 2412 19780 2464 19786
rect 2412 19722 2464 19728
rect 2320 19440 2372 19446
rect 2320 19382 2372 19388
rect 2228 18624 2280 18630
rect 2228 18566 2280 18572
rect 2136 18284 2188 18290
rect 2136 18226 2188 18232
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 2044 18216 2096 18222
rect 2044 18158 2096 18164
rect 572 18080 624 18086
rect 572 18022 624 18028
rect 1780 17785 1808 18158
rect 1950 17912 2006 17921
rect 1950 17847 1952 17856
rect 2004 17847 2006 17856
rect 1952 17818 2004 17824
rect 1766 17776 1822 17785
rect 1766 17711 1822 17720
rect 1860 17128 1912 17134
rect 1860 17070 1912 17076
rect 1768 16652 1820 16658
rect 1768 16594 1820 16600
rect 1400 15904 1452 15910
rect 1400 15846 1452 15852
rect 1412 15065 1440 15846
rect 1398 15056 1454 15065
rect 1398 14991 1454 15000
rect 1780 14770 1808 16594
rect 1872 15026 1900 17070
rect 1952 16992 2004 16998
rect 1950 16960 1952 16969
rect 2004 16960 2006 16969
rect 1950 16895 2006 16904
rect 1950 16552 2006 16561
rect 1950 16487 1952 16496
rect 2004 16487 2006 16496
rect 1952 16458 2004 16464
rect 1950 16008 2006 16017
rect 1950 15943 2006 15952
rect 1964 15706 1992 15943
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 1950 15600 2006 15609
rect 1950 15535 2006 15544
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 1780 14742 1900 14770
rect 1766 14648 1822 14657
rect 1766 14583 1822 14592
rect 1676 14476 1728 14482
rect 1676 14418 1728 14424
rect 1688 13938 1716 14418
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1412 11898 1440 13806
rect 1584 13796 1636 13802
rect 1584 13738 1636 13744
rect 1596 13394 1624 13738
rect 1780 13530 1808 14583
rect 1872 13977 1900 14742
rect 1964 14618 1992 15535
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 2056 14278 2084 18158
rect 2228 18080 2280 18086
rect 2228 18022 2280 18028
rect 2136 17060 2188 17066
rect 2136 17002 2188 17008
rect 2044 14272 2096 14278
rect 2044 14214 2096 14220
rect 1858 13968 1914 13977
rect 1858 13903 1914 13912
rect 1768 13524 1820 13530
rect 1768 13466 1820 13472
rect 2148 13462 2176 17002
rect 2240 16454 2268 18022
rect 2320 16584 2372 16590
rect 2424 16561 2452 19722
rect 2504 19304 2556 19310
rect 2504 19246 2556 19252
rect 2320 16526 2372 16532
rect 2410 16552 2466 16561
rect 2228 16448 2280 16454
rect 2228 16390 2280 16396
rect 2228 16040 2280 16046
rect 2228 15982 2280 15988
rect 2240 14414 2268 15982
rect 2332 14958 2360 16526
rect 2410 16487 2466 16496
rect 2320 14952 2372 14958
rect 2320 14894 2372 14900
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 2136 13456 2188 13462
rect 2136 13398 2188 13404
rect 2424 13394 2452 16487
rect 1584 13388 1636 13394
rect 1584 13330 1636 13336
rect 2412 13388 2464 13394
rect 2412 13330 2464 13336
rect 1860 12776 1912 12782
rect 1860 12718 1912 12724
rect 1492 12300 1544 12306
rect 1492 12242 1544 12248
rect 1400 11892 1452 11898
rect 1400 11834 1452 11840
rect 1504 11218 1532 12242
rect 1492 11212 1544 11218
rect 1492 11154 1544 11160
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1412 8974 1440 10066
rect 1872 9586 1900 12718
rect 2516 12646 2544 19246
rect 2700 17241 2728 22320
rect 3054 22128 3110 22137
rect 3054 22063 3110 22072
rect 2778 21584 2834 21593
rect 2778 21519 2834 21528
rect 2792 20058 2820 21519
rect 2962 20632 3018 20641
rect 2962 20567 3018 20576
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 2872 19916 2924 19922
rect 2872 19858 2924 19864
rect 2884 19242 2912 19858
rect 2872 19236 2924 19242
rect 2872 19178 2924 19184
rect 2976 19174 3004 20567
rect 3068 19854 3096 22063
rect 3056 19848 3108 19854
rect 3056 19790 3108 19796
rect 3056 19712 3108 19718
rect 3056 19654 3108 19660
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 3068 18873 3096 19654
rect 3054 18864 3110 18873
rect 3160 18850 3188 22320
rect 3252 18970 3280 22471
rect 3514 22320 3570 22800
rect 3974 22320 4030 22800
rect 4342 22320 4398 22800
rect 4802 22320 4858 22800
rect 5262 22320 5318 22800
rect 5630 22320 5686 22800
rect 6090 22320 6146 22800
rect 6458 22320 6514 22800
rect 6918 22320 6974 22800
rect 7378 22320 7434 22800
rect 7746 22320 7802 22800
rect 8206 22320 8262 22800
rect 8574 22320 8630 22800
rect 9034 22320 9090 22800
rect 9494 22320 9550 22800
rect 9862 22320 9918 22800
rect 10322 22320 10378 22800
rect 10690 22320 10746 22800
rect 11150 22320 11206 22800
rect 11610 22320 11666 22800
rect 11978 22320 12034 22800
rect 12438 22320 12494 22800
rect 12806 22320 12862 22800
rect 13266 22320 13322 22800
rect 13634 22320 13690 22800
rect 14094 22320 14150 22800
rect 14554 22320 14610 22800
rect 14922 22320 14978 22800
rect 15382 22320 15438 22800
rect 15750 22320 15806 22800
rect 16210 22320 16266 22800
rect 16670 22320 16726 22800
rect 17038 22320 17094 22800
rect 17498 22320 17554 22800
rect 17866 22320 17922 22800
rect 18326 22320 18382 22800
rect 18786 22320 18842 22800
rect 19154 22320 19210 22800
rect 19614 22320 19670 22800
rect 19982 22320 20038 22800
rect 20442 22320 20498 22800
rect 20718 22536 20774 22545
rect 20718 22471 20774 22480
rect 3422 20224 3478 20233
rect 3422 20159 3478 20168
rect 3436 19514 3464 20159
rect 3424 19508 3476 19514
rect 3424 19450 3476 19456
rect 3424 19304 3476 19310
rect 3424 19246 3476 19252
rect 3240 18964 3292 18970
rect 3240 18906 3292 18912
rect 3160 18822 3280 18850
rect 3054 18799 3110 18808
rect 3146 18728 3202 18737
rect 3252 18698 3280 18822
rect 3146 18663 3148 18672
rect 3200 18663 3202 18672
rect 3240 18692 3292 18698
rect 3148 18634 3200 18640
rect 3240 18634 3292 18640
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 2872 18420 2924 18426
rect 2872 18362 2924 18368
rect 2778 18320 2834 18329
rect 2778 18255 2834 18264
rect 2792 17882 2820 18255
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2778 17368 2834 17377
rect 2778 17303 2780 17312
rect 2832 17303 2834 17312
rect 2780 17274 2832 17280
rect 2686 17232 2742 17241
rect 2686 17167 2742 17176
rect 2884 15638 2912 18362
rect 3240 18216 3292 18222
rect 3238 18184 3240 18193
rect 3292 18184 3294 18193
rect 3238 18119 3294 18128
rect 3344 17898 3372 18566
rect 3252 17870 3372 17898
rect 3252 17610 3280 17870
rect 3332 17740 3384 17746
rect 3332 17682 3384 17688
rect 3240 17604 3292 17610
rect 3240 17546 3292 17552
rect 3056 17536 3108 17542
rect 3056 17478 3108 17484
rect 3068 17338 3096 17478
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 2964 17128 3016 17134
rect 2964 17070 3016 17076
rect 2872 15632 2924 15638
rect 2872 15574 2924 15580
rect 2778 14104 2834 14113
rect 2778 14039 2834 14048
rect 2792 12986 2820 14039
rect 2870 13696 2926 13705
rect 2870 13631 2926 13640
rect 2780 12980 2832 12986
rect 2780 12922 2832 12928
rect 2778 12880 2834 12889
rect 2778 12815 2834 12824
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 2608 12374 2636 12718
rect 2596 12368 2648 12374
rect 2596 12310 2648 12316
rect 2320 12300 2372 12306
rect 2320 12242 2372 12248
rect 2332 11830 2360 12242
rect 2608 12238 2636 12310
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2320 11824 2372 11830
rect 2320 11766 2372 11772
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2148 10810 2176 11494
rect 2332 11354 2360 11766
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2136 10804 2188 10810
rect 2136 10746 2188 10752
rect 2332 10674 2360 11290
rect 2596 11212 2648 11218
rect 2596 11154 2648 11160
rect 2608 10674 2636 11154
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 1964 10266 1992 10406
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 2320 10124 2372 10130
rect 2320 10066 2372 10072
rect 2332 9625 2360 10066
rect 2608 10062 2636 10610
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2318 9616 2374 9625
rect 1860 9580 1912 9586
rect 2318 9551 2374 9560
rect 1860 9522 1912 9528
rect 2228 9512 2280 9518
rect 2228 9454 2280 9460
rect 2240 9178 2268 9454
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 1400 8968 1452 8974
rect 1400 8910 1452 8916
rect 1584 8424 1636 8430
rect 1584 8366 1636 8372
rect 1596 7886 1624 8366
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1596 6866 1624 7822
rect 2608 7546 2636 8978
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 1584 6860 1636 6866
rect 1584 6802 1636 6808
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 2240 480 2268 6802
rect 2792 6730 2820 12815
rect 2884 9994 2912 13631
rect 2976 13297 3004 17070
rect 3056 16992 3108 16998
rect 3054 16960 3056 16969
rect 3108 16960 3110 16969
rect 3054 16895 3110 16904
rect 3148 16652 3200 16658
rect 3148 16594 3200 16600
rect 3160 16114 3188 16594
rect 3148 16108 3200 16114
rect 3148 16050 3200 16056
rect 3056 15904 3108 15910
rect 3056 15846 3108 15852
rect 3068 15706 3096 15846
rect 3056 15700 3108 15706
rect 3056 15642 3108 15648
rect 3160 14822 3188 16050
rect 3252 16046 3280 17546
rect 3240 16040 3292 16046
rect 3240 15982 3292 15988
rect 3240 15496 3292 15502
rect 3240 15438 3292 15444
rect 3252 14890 3280 15438
rect 3240 14884 3292 14890
rect 3240 14826 3292 14832
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 3160 14550 3188 14758
rect 3148 14544 3200 14550
rect 3148 14486 3200 14492
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 2962 13288 3018 13297
rect 2962 13223 3018 13232
rect 2964 12708 3016 12714
rect 2964 12650 3016 12656
rect 2976 12442 3004 12650
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 2976 11762 3004 12378
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2872 9988 2924 9994
rect 2872 9930 2924 9936
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2884 8974 2912 9386
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2884 8634 2912 8910
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2780 6724 2832 6730
rect 2780 6666 2832 6672
rect 2976 6458 3004 7142
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2872 6180 2924 6186
rect 2872 6122 2924 6128
rect 2884 1601 2912 6122
rect 3068 4321 3096 14418
rect 3148 13456 3200 13462
rect 3146 13424 3148 13433
rect 3200 13424 3202 13433
rect 3146 13359 3202 13368
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3160 11694 3188 13126
rect 3252 12889 3280 14826
rect 3238 12880 3294 12889
rect 3238 12815 3294 12824
rect 3148 11688 3200 11694
rect 3148 11630 3200 11636
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3160 10606 3188 11086
rect 3240 11008 3292 11014
rect 3240 10950 3292 10956
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3148 10464 3200 10470
rect 3148 10406 3200 10412
rect 3160 9722 3188 10406
rect 3252 10033 3280 10950
rect 3238 10024 3294 10033
rect 3238 9959 3294 9968
rect 3148 9716 3200 9722
rect 3148 9658 3200 9664
rect 3148 9444 3200 9450
rect 3148 9386 3200 9392
rect 3160 8022 3188 9386
rect 3240 8900 3292 8906
rect 3240 8842 3292 8848
rect 3252 8634 3280 8842
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3148 8016 3200 8022
rect 3148 7958 3200 7964
rect 3160 7546 3188 7958
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 3054 4312 3110 4321
rect 3054 4247 3110 4256
rect 3160 2961 3188 6802
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3146 2952 3202 2961
rect 3146 2887 3202 2896
rect 3252 2553 3280 6054
rect 3344 5817 3372 17682
rect 3436 16538 3464 19246
rect 3528 18630 3556 22320
rect 3882 21176 3938 21185
rect 3882 21111 3938 21120
rect 3896 21010 3924 21111
rect 3884 21004 3936 21010
rect 3884 20946 3936 20952
rect 3988 19310 4016 22320
rect 4356 19768 4384 22320
rect 4356 19740 4752 19768
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 3792 19304 3844 19310
rect 3790 19272 3792 19281
rect 3976 19304 4028 19310
rect 3844 19272 3846 19281
rect 3976 19246 4028 19252
rect 3790 19207 3846 19216
rect 3700 18828 3752 18834
rect 3700 18770 3752 18776
rect 3516 18624 3568 18630
rect 3516 18566 3568 18572
rect 3516 18420 3568 18426
rect 3516 18362 3568 18368
rect 3528 17814 3556 18362
rect 3516 17808 3568 17814
rect 3516 17750 3568 17756
rect 3436 16510 3556 16538
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 3436 15638 3464 16390
rect 3424 15632 3476 15638
rect 3424 15574 3476 15580
rect 3424 15088 3476 15094
rect 3424 15030 3476 15036
rect 3436 14346 3464 15030
rect 3424 14340 3476 14346
rect 3424 14282 3476 14288
rect 3424 13320 3476 13326
rect 3424 13262 3476 13268
rect 3436 11830 3464 13262
rect 3424 11824 3476 11830
rect 3424 11766 3476 11772
rect 3436 10742 3464 11766
rect 3424 10736 3476 10742
rect 3424 10678 3476 10684
rect 3528 10674 3556 16510
rect 3608 13864 3660 13870
rect 3608 13806 3660 13812
rect 3620 11898 3648 13806
rect 3608 11892 3660 11898
rect 3608 11834 3660 11840
rect 3712 11393 3740 18770
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 3792 18352 3844 18358
rect 3790 18320 3792 18329
rect 3844 18320 3846 18329
rect 3790 18255 3846 18264
rect 3884 18216 3936 18222
rect 3884 18158 3936 18164
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 3792 18148 3844 18154
rect 3792 18090 3844 18096
rect 3698 11384 3754 11393
rect 3698 11319 3754 11328
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3424 10600 3476 10606
rect 3424 10542 3476 10548
rect 3436 10266 3464 10542
rect 3700 10464 3752 10470
rect 3700 10406 3752 10412
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3514 10160 3570 10169
rect 3514 10095 3570 10104
rect 3528 10062 3556 10095
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3436 6186 3464 9454
rect 3620 9450 3648 9862
rect 3608 9444 3660 9450
rect 3608 9386 3660 9392
rect 3712 9042 3740 10406
rect 3804 9489 3832 18090
rect 3896 17082 3924 18158
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 4080 17678 4108 17818
rect 4068 17672 4120 17678
rect 4068 17614 4120 17620
rect 3976 17536 4028 17542
rect 3976 17478 4028 17484
rect 3988 17202 4016 17478
rect 4068 17264 4120 17270
rect 4172 17218 4200 18158
rect 4724 17898 4752 19740
rect 4816 18986 4844 22320
rect 4816 18958 5212 18986
rect 4804 18828 4856 18834
rect 4804 18770 4856 18776
rect 4816 18290 4844 18770
rect 4988 18692 5040 18698
rect 4988 18634 5040 18640
rect 4804 18284 4856 18290
rect 4804 18226 4856 18232
rect 4724 17870 4936 17898
rect 4252 17740 4304 17746
rect 4252 17682 4304 17688
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 4120 17212 4200 17218
rect 4068 17206 4200 17212
rect 3976 17196 4028 17202
rect 4080 17190 4200 17206
rect 3976 17138 4028 17144
rect 3896 17054 4016 17082
rect 3884 16992 3936 16998
rect 3884 16934 3936 16940
rect 3896 15706 3924 16934
rect 3884 15700 3936 15706
rect 3884 15642 3936 15648
rect 3884 14952 3936 14958
rect 3884 14894 3936 14900
rect 3896 14482 3924 14894
rect 3884 14476 3936 14482
rect 3884 14418 3936 14424
rect 3896 14074 3924 14418
rect 3884 14068 3936 14074
rect 3884 14010 3936 14016
rect 3988 13954 4016 17054
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 4080 16454 4108 16730
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 4264 16250 4292 17682
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 4528 17128 4580 17134
rect 4528 17070 4580 17076
rect 4540 16833 4568 17070
rect 4526 16824 4582 16833
rect 4526 16759 4582 16768
rect 4540 16640 4568 16759
rect 4724 16726 4752 17614
rect 4712 16720 4764 16726
rect 4712 16662 4764 16668
rect 4620 16652 4672 16658
rect 4540 16612 4620 16640
rect 4620 16594 4672 16600
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 4080 15434 4108 16050
rect 4724 15502 4752 16662
rect 4816 16182 4844 17682
rect 4804 16176 4856 16182
rect 4804 16118 4856 16124
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4068 15428 4120 15434
rect 4068 15370 4120 15376
rect 4172 14618 4200 15438
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 3896 13926 4016 13954
rect 3790 9480 3846 9489
rect 3790 9415 3846 9424
rect 3700 9036 3752 9042
rect 3700 8978 3752 8984
rect 3608 8288 3660 8294
rect 3608 8230 3660 8236
rect 3620 8090 3648 8230
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3608 7948 3660 7954
rect 3608 7890 3660 7896
rect 3620 6322 3648 7890
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 3712 6118 3740 8978
rect 3792 8356 3844 8362
rect 3792 8298 3844 8304
rect 3804 7818 3832 8298
rect 3792 7812 3844 7818
rect 3792 7754 3844 7760
rect 3804 7410 3832 7754
rect 3896 7585 3924 13926
rect 4068 13456 4120 13462
rect 4068 13398 4120 13404
rect 4080 12753 4108 13398
rect 4252 13388 4304 13394
rect 4252 13330 4304 13336
rect 4264 12850 4292 13330
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4066 12744 4122 12753
rect 4066 12679 4122 12688
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 4080 12345 4108 12378
rect 4066 12336 4122 12345
rect 3976 12300 4028 12306
rect 4066 12271 4122 12280
rect 3976 12242 4028 12248
rect 3988 11801 4016 12242
rect 4068 12232 4120 12238
rect 4528 12232 4580 12238
rect 4068 12174 4120 12180
rect 4526 12200 4528 12209
rect 4580 12200 4582 12209
rect 3974 11792 4030 11801
rect 3974 11727 4030 11736
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3988 10810 4016 11494
rect 4080 11218 4108 12174
rect 4526 12135 4582 12144
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4066 10840 4122 10849
rect 3976 10804 4028 10810
rect 4388 10832 4684 10852
rect 4724 10810 4752 13262
rect 4066 10775 4122 10784
rect 4712 10804 4764 10810
rect 3976 10746 4028 10752
rect 4080 10742 4108 10775
rect 4712 10746 4764 10752
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 3988 10305 4016 10610
rect 4160 10464 4212 10470
rect 4804 10464 4856 10470
rect 4160 10406 4212 10412
rect 4342 10432 4398 10441
rect 3974 10296 4030 10305
rect 4172 10266 4200 10406
rect 4804 10406 4856 10412
rect 4342 10367 4398 10376
rect 3974 10231 4030 10240
rect 4160 10260 4212 10266
rect 3988 9602 4016 10231
rect 4160 10202 4212 10208
rect 4356 9994 4384 10367
rect 4712 10192 4764 10198
rect 4712 10134 4764 10140
rect 4620 10056 4672 10062
rect 4618 10024 4620 10033
rect 4672 10024 4674 10033
rect 4344 9988 4396 9994
rect 4618 9959 4674 9968
rect 4344 9930 4396 9936
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 3988 9574 4292 9602
rect 4068 9444 4120 9450
rect 4068 9386 4120 9392
rect 3976 9104 4028 9110
rect 4080 9081 4108 9386
rect 3976 9046 4028 9052
rect 4066 9072 4122 9081
rect 3988 8362 4016 9046
rect 4066 9007 4122 9016
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4080 8537 4108 8570
rect 4066 8528 4122 8537
rect 4066 8463 4122 8472
rect 3976 8356 4028 8362
rect 3976 8298 4028 8304
rect 4066 8120 4122 8129
rect 4066 8055 4122 8064
rect 3976 8016 4028 8022
rect 3976 7958 4028 7964
rect 3882 7576 3938 7585
rect 3882 7511 3938 7520
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 3792 7268 3844 7274
rect 3792 7210 3844 7216
rect 3700 6112 3752 6118
rect 3700 6054 3752 6060
rect 3330 5808 3386 5817
rect 3330 5743 3386 5752
rect 3804 3505 3832 7210
rect 3884 7200 3936 7206
rect 3988 7177 4016 7958
rect 4080 7750 4108 8055
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 4172 7274 4200 8910
rect 4264 8090 4292 9574
rect 4724 9178 4752 10134
rect 4816 9518 4844 10406
rect 4804 9512 4856 9518
rect 4804 9454 4856 9460
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4804 8900 4856 8906
rect 4804 8842 4856 8848
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4342 8528 4398 8537
rect 4724 8498 4752 8774
rect 4342 8463 4398 8472
rect 4712 8492 4764 8498
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4356 7970 4384 8463
rect 4712 8434 4764 8440
rect 4816 8362 4844 8842
rect 4804 8356 4856 8362
rect 4804 8298 4856 8304
rect 4908 8265 4936 17870
rect 5000 17105 5028 18634
rect 4986 17096 5042 17105
rect 4986 17031 5042 17040
rect 5000 15910 5028 17031
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 5000 12782 5028 14554
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 5092 14074 5120 14418
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 4988 12776 5040 12782
rect 4988 12718 5040 12724
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 5092 11234 5120 12582
rect 5184 11642 5212 18958
rect 5276 18086 5304 22320
rect 5540 21004 5592 21010
rect 5540 20946 5592 20952
rect 5356 19440 5408 19446
rect 5356 19382 5408 19388
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 5368 15586 5396 19382
rect 5552 19174 5580 20946
rect 5540 19168 5592 19174
rect 5540 19110 5592 19116
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5448 17604 5500 17610
rect 5448 17546 5500 17552
rect 5460 17513 5488 17546
rect 5446 17504 5502 17513
rect 5446 17439 5502 17448
rect 5448 17060 5500 17066
rect 5448 17002 5500 17008
rect 5460 16794 5488 17002
rect 5552 16833 5580 17614
rect 5538 16824 5594 16833
rect 5448 16788 5500 16794
rect 5538 16759 5594 16768
rect 5448 16730 5500 16736
rect 5552 15706 5580 16759
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5276 15558 5396 15586
rect 5276 14618 5304 15558
rect 5356 15496 5408 15502
rect 5356 15438 5408 15444
rect 5368 15337 5396 15438
rect 5354 15328 5410 15337
rect 5354 15263 5410 15272
rect 5448 14884 5500 14890
rect 5448 14826 5500 14832
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 5276 13870 5304 14418
rect 5368 14074 5396 14758
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5264 13864 5316 13870
rect 5264 13806 5316 13812
rect 5276 13326 5304 13806
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5276 12850 5304 13262
rect 5460 13258 5488 14826
rect 5552 14550 5580 15642
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5552 14414 5580 14486
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5644 13258 5672 22320
rect 5908 19304 5960 19310
rect 5908 19246 5960 19252
rect 5722 19136 5778 19145
rect 5722 19071 5778 19080
rect 5736 18601 5764 19071
rect 5920 18902 5948 19246
rect 5816 18896 5868 18902
rect 5816 18838 5868 18844
rect 5908 18896 5960 18902
rect 5908 18838 5960 18844
rect 5722 18592 5778 18601
rect 5722 18527 5778 18536
rect 5828 18222 5856 18838
rect 5908 18760 5960 18766
rect 5908 18702 5960 18708
rect 5816 18216 5868 18222
rect 5816 18158 5868 18164
rect 5724 18080 5776 18086
rect 5724 18022 5776 18028
rect 5448 13252 5500 13258
rect 5448 13194 5500 13200
rect 5632 13252 5684 13258
rect 5632 13194 5684 13200
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 5276 11762 5304 12038
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5184 11614 5304 11642
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 5184 11354 5212 11494
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5092 11206 5212 11234
rect 5080 11144 5132 11150
rect 5080 11086 5132 11092
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 4894 8256 4950 8265
rect 4894 8191 4950 8200
rect 5000 8072 5028 10746
rect 5092 10062 5120 11086
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 5092 9586 5120 9998
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 5184 9178 5212 11206
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 5170 9072 5226 9081
rect 5170 9007 5172 9016
rect 5224 9007 5226 9016
rect 5172 8978 5224 8984
rect 5276 8480 5304 11614
rect 5368 10470 5396 12718
rect 5448 12368 5500 12374
rect 5448 12310 5500 12316
rect 5460 11762 5488 12310
rect 5538 12200 5594 12209
rect 5538 12135 5594 12144
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5460 11082 5488 11698
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5460 10674 5488 11018
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5368 9058 5396 10406
rect 5552 10130 5580 12135
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5644 10130 5672 10610
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5448 9920 5500 9926
rect 5552 9908 5580 10066
rect 5500 9880 5580 9908
rect 5448 9862 5500 9868
rect 5630 9616 5686 9625
rect 5630 9551 5686 9560
rect 5644 9382 5672 9551
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5368 9030 5580 9058
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 4264 7942 4384 7970
rect 4816 8044 5028 8072
rect 5092 8452 5304 8480
rect 5356 8492 5408 8498
rect 4160 7268 4212 7274
rect 4160 7210 4212 7216
rect 3884 7142 3936 7148
rect 3974 7168 4030 7177
rect 3896 7002 3924 7142
rect 3974 7103 4030 7112
rect 3884 6996 3936 7002
rect 3884 6938 3936 6944
rect 4264 6798 4292 7942
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4724 7410 4752 7822
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4252 6792 4304 6798
rect 3974 6760 4030 6769
rect 4252 6734 4304 6740
rect 3974 6695 4030 6704
rect 3988 6254 4016 6695
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 3976 6248 4028 6254
rect 4080 6225 4108 6326
rect 3976 6190 4028 6196
rect 4066 6216 4122 6225
rect 4066 6151 4122 6160
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3988 3913 4016 6054
rect 4068 5296 4120 5302
rect 4066 5264 4068 5273
rect 4120 5264 4122 5273
rect 4066 5199 4122 5208
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4080 4865 4108 4966
rect 4066 4856 4122 4865
rect 4066 4791 4122 4800
rect 3974 3904 4030 3913
rect 3974 3839 4030 3848
rect 3790 3496 3846 3505
rect 3790 3431 3846 3440
rect 3238 2544 3294 2553
rect 3238 2479 3294 2488
rect 4264 2009 4292 6734
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4816 6186 4844 8044
rect 4894 7984 4950 7993
rect 4894 7919 4950 7928
rect 4988 7948 5040 7954
rect 4804 6180 4856 6186
rect 4804 6122 4856 6128
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4908 2990 4936 7919
rect 4988 7890 5040 7896
rect 4896 2984 4948 2990
rect 4896 2926 4948 2932
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4250 2000 4306 2009
rect 4250 1935 4306 1944
rect 2870 1592 2926 1601
rect 2870 1527 2926 1536
rect 2964 1352 3016 1358
rect 2964 1294 3016 1300
rect 2780 1080 2832 1086
rect 2976 1057 3004 1294
rect 5000 1086 5028 7890
rect 5092 2854 5120 8452
rect 5356 8434 5408 8440
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 5184 6662 5212 8298
rect 5368 8294 5396 8434
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 5276 7546 5304 7754
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5368 7426 5396 8230
rect 5460 7954 5488 8910
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5276 7398 5396 7426
rect 5276 7342 5304 7398
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5276 6798 5304 7278
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5276 6322 5304 6734
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5368 6254 5396 7142
rect 5552 7002 5580 9030
rect 5644 8537 5672 9318
rect 5630 8528 5686 8537
rect 5630 8463 5686 8472
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5540 6860 5592 6866
rect 5540 6802 5592 6808
rect 5552 6458 5580 6802
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5736 2922 5764 18022
rect 5816 17740 5868 17746
rect 5816 17682 5868 17688
rect 5828 17270 5856 17682
rect 5816 17264 5868 17270
rect 5816 17206 5868 17212
rect 5816 15020 5868 15026
rect 5816 14962 5868 14968
rect 5828 14618 5856 14962
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5920 13410 5948 18702
rect 6104 17354 6132 22320
rect 6472 19174 6500 22320
rect 6932 19394 6960 22320
rect 7288 19916 7340 19922
rect 7288 19858 7340 19864
rect 6932 19366 7236 19394
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 6552 19236 6604 19242
rect 6552 19178 6604 19184
rect 6460 19168 6512 19174
rect 6460 19110 6512 19116
rect 6460 18692 6512 18698
rect 6460 18634 6512 18640
rect 6104 17326 6408 17354
rect 6092 15972 6144 15978
rect 6092 15914 6144 15920
rect 6000 13932 6052 13938
rect 6000 13874 6052 13880
rect 5828 13382 5948 13410
rect 5828 12866 5856 13382
rect 6012 13326 6040 13874
rect 5908 13320 5960 13326
rect 5908 13262 5960 13268
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 5920 12986 5948 13262
rect 5908 12980 5960 12986
rect 5908 12922 5960 12928
rect 6000 12912 6052 12918
rect 5828 12838 5948 12866
rect 6000 12854 6052 12860
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 5828 10169 5856 12582
rect 5920 10441 5948 12838
rect 6012 11354 6040 12854
rect 6104 12102 6132 15914
rect 6184 15428 6236 15434
rect 6184 15370 6236 15376
rect 6196 12714 6224 15370
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 6184 12708 6236 12714
rect 6184 12650 6236 12656
rect 6184 12232 6236 12238
rect 6182 12200 6184 12209
rect 6236 12200 6238 12209
rect 6182 12135 6238 12144
rect 6092 12096 6144 12102
rect 6092 12038 6144 12044
rect 6000 11348 6052 11354
rect 6000 11290 6052 11296
rect 6092 11212 6144 11218
rect 6092 11154 6144 11160
rect 6000 10464 6052 10470
rect 5906 10432 5962 10441
rect 6000 10406 6052 10412
rect 5906 10367 5962 10376
rect 6012 10266 6040 10406
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 5814 10160 5870 10169
rect 5814 10095 5870 10104
rect 5828 6934 5856 10095
rect 5906 10024 5962 10033
rect 5906 9959 5962 9968
rect 5920 9382 5948 9959
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 6104 9178 6132 11154
rect 6288 10146 6316 12786
rect 6380 11286 6408 17326
rect 6472 13530 6500 18634
rect 6460 13524 6512 13530
rect 6460 13466 6512 13472
rect 6564 12646 6592 19178
rect 6826 19000 6882 19009
rect 6826 18935 6882 18944
rect 6840 18358 6868 18935
rect 7116 18834 7144 19246
rect 7012 18828 7064 18834
rect 7012 18770 7064 18776
rect 7104 18828 7156 18834
rect 7104 18770 7156 18776
rect 6828 18352 6880 18358
rect 6828 18294 6880 18300
rect 6840 18154 6868 18294
rect 6828 18148 6880 18154
rect 6828 18090 6880 18096
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6644 17876 6696 17882
rect 6644 17818 6696 17824
rect 6656 17134 6684 17818
rect 6828 17672 6880 17678
rect 6828 17614 6880 17620
rect 6840 17338 6868 17614
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6932 17202 6960 18022
rect 7024 17898 7052 18770
rect 7024 17882 7144 17898
rect 7024 17876 7156 17882
rect 7024 17870 7104 17876
rect 7104 17818 7156 17824
rect 7208 17762 7236 19366
rect 7300 18902 7328 19858
rect 7288 18896 7340 18902
rect 7288 18838 7340 18844
rect 7288 18284 7340 18290
rect 7288 18226 7340 18232
rect 7024 17734 7236 17762
rect 7300 17746 7328 18226
rect 7288 17740 7340 17746
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 6644 17128 6696 17134
rect 6644 17070 6696 17076
rect 6828 17128 6880 17134
rect 6880 17076 6960 17082
rect 6828 17070 6960 17076
rect 6840 17054 6960 17070
rect 6932 16182 6960 17054
rect 6920 16176 6972 16182
rect 6920 16118 6972 16124
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6840 13870 6868 14758
rect 6932 14618 6960 16118
rect 7024 15026 7052 17734
rect 7288 17682 7340 17688
rect 7392 17626 7420 22320
rect 7760 19310 7788 22320
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 7748 19304 7800 19310
rect 8220 19292 8248 22320
rect 8484 19916 8536 19922
rect 8484 19858 8536 19864
rect 8220 19264 8340 19292
rect 8496 19281 8524 19858
rect 8588 19446 8616 22320
rect 8668 20664 8720 20670
rect 8668 20606 8720 20612
rect 8680 20058 8708 20606
rect 8668 20052 8720 20058
rect 8668 19994 8720 20000
rect 8668 19916 8720 19922
rect 8668 19858 8720 19864
rect 8576 19440 8628 19446
rect 8576 19382 8628 19388
rect 7748 19246 7800 19252
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 8116 17808 8168 17814
rect 8116 17750 8168 17756
rect 7564 17740 7616 17746
rect 7564 17682 7616 17688
rect 7208 17598 7420 17626
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 7116 16794 7144 17274
rect 7104 16788 7156 16794
rect 7104 16730 7156 16736
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 7012 15020 7064 15026
rect 7012 14962 7064 14968
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 7024 14550 7052 14962
rect 7012 14544 7064 14550
rect 7012 14486 7064 14492
rect 7116 14346 7144 15982
rect 7104 14340 7156 14346
rect 7104 14282 7156 14288
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 7024 14074 7052 14214
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6644 13388 6696 13394
rect 6644 13330 6696 13336
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 6368 11280 6420 11286
rect 6368 11222 6420 11228
rect 6366 10296 6422 10305
rect 6366 10231 6422 10240
rect 6196 10130 6316 10146
rect 6380 10130 6408 10231
rect 6184 10124 6316 10130
rect 6236 10118 6316 10124
rect 6368 10124 6420 10130
rect 6184 10066 6236 10072
rect 6368 10066 6420 10072
rect 6196 9586 6224 10066
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 6196 9081 6224 9522
rect 6182 9072 6238 9081
rect 5908 9036 5960 9042
rect 6182 9007 6238 9016
rect 5908 8978 5960 8984
rect 5920 8906 5948 8978
rect 6196 8974 6224 9007
rect 6184 8968 6236 8974
rect 6184 8910 6236 8916
rect 5908 8900 5960 8906
rect 5908 8842 5960 8848
rect 5816 6928 5868 6934
rect 5816 6870 5868 6876
rect 5724 2916 5776 2922
rect 5724 2858 5776 2864
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 5920 1358 5948 8842
rect 6472 8820 6500 12038
rect 6656 9042 6684 13330
rect 6828 13252 6880 13258
rect 6828 13194 6880 13200
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6748 11354 6776 11494
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6644 9036 6696 9042
rect 6644 8978 6696 8984
rect 6104 8792 6500 8820
rect 6104 5370 6132 8792
rect 6552 8424 6604 8430
rect 6552 8366 6604 8372
rect 6184 8356 6236 8362
rect 6184 8298 6236 8304
rect 6196 6730 6224 8298
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6380 7546 6408 7890
rect 6368 7540 6420 7546
rect 6368 7482 6420 7488
rect 6380 6798 6408 7482
rect 6564 7002 6592 8366
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6184 6724 6236 6730
rect 6184 6666 6236 6672
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 5908 1352 5960 1358
rect 5908 1294 5960 1300
rect 4988 1080 5040 1086
rect 2780 1022 2832 1028
rect 2962 1048 3018 1057
rect 2792 649 2820 1022
rect 4988 1022 5040 1028
rect 2962 983 3018 992
rect 2778 640 2834 649
rect 2778 575 2834 584
rect 6748 480 6776 9318
rect 6840 8906 6868 13194
rect 6932 12889 6960 13466
rect 7116 12918 7144 14282
rect 7104 12912 7156 12918
rect 6918 12880 6974 12889
rect 7104 12854 7156 12860
rect 6918 12815 6974 12824
rect 7208 12102 7236 17598
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 7392 17202 7420 17478
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7392 16726 7420 17138
rect 7472 17128 7524 17134
rect 7472 17070 7524 17076
rect 7484 16969 7512 17070
rect 7470 16960 7526 16969
rect 7470 16895 7526 16904
rect 7380 16720 7432 16726
rect 7380 16662 7432 16668
rect 7392 16114 7420 16662
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7380 16108 7432 16114
rect 7380 16050 7432 16056
rect 7380 15904 7432 15910
rect 7380 15846 7432 15852
rect 7392 15706 7420 15846
rect 7380 15700 7432 15706
rect 7380 15642 7432 15648
rect 7484 15586 7512 16526
rect 7576 16250 7604 17682
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 7760 16794 7788 17614
rect 8022 17232 8078 17241
rect 8128 17202 8156 17750
rect 8022 17167 8078 17176
rect 8116 17196 8168 17202
rect 8036 17066 8064 17167
rect 8116 17138 8168 17144
rect 8024 17060 8076 17066
rect 8128 17048 8156 17138
rect 8128 17020 8248 17048
rect 8024 17002 8076 17008
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 7656 16652 7708 16658
rect 7656 16594 7708 16600
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7392 15558 7512 15586
rect 7288 15496 7340 15502
rect 7288 15438 7340 15444
rect 7300 12594 7328 15438
rect 7392 14958 7420 15558
rect 7576 15366 7604 15642
rect 7668 15570 7696 16594
rect 8220 16114 8248 17020
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 7760 15570 7788 16050
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 8220 15638 8248 15846
rect 8208 15632 8260 15638
rect 8208 15574 8260 15580
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 7748 15564 7800 15570
rect 7748 15506 7800 15512
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7576 15042 7604 15302
rect 7668 15162 7696 15506
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 7472 15020 7524 15026
rect 7576 15014 7696 15042
rect 7472 14962 7524 14968
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 7392 13870 7420 14894
rect 7484 14414 7512 14962
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7380 13864 7432 13870
rect 7380 13806 7432 13812
rect 7392 13530 7420 13806
rect 7484 13802 7512 14214
rect 7472 13796 7524 13802
rect 7472 13738 7524 13744
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 7380 13320 7432 13326
rect 7484 13308 7512 13738
rect 7432 13280 7512 13308
rect 7380 13262 7432 13268
rect 7472 12912 7524 12918
rect 7472 12854 7524 12860
rect 7300 12566 7420 12594
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6932 10266 6960 11086
rect 7024 10810 7052 11494
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 7024 9926 7052 10746
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 7116 8616 7144 10610
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7300 9178 7328 10202
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7024 8588 7144 8616
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6932 8090 6960 8298
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6932 7410 6960 7822
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6828 6928 6880 6934
rect 6828 6870 6880 6876
rect 2226 0 2282 480
rect 3332 264 3384 270
rect 3330 232 3332 241
rect 3384 232 3386 241
rect 3330 167 3386 176
rect 6734 0 6790 480
rect 6840 270 6868 6870
rect 7024 6390 7052 8588
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7116 8090 7144 8434
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7116 7274 7144 8026
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 7208 6662 7236 8774
rect 7392 6662 7420 12566
rect 7484 10674 7512 12854
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7484 10198 7512 10406
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 7576 9586 7604 10406
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7484 9178 7512 9454
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7668 8362 7696 15014
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 7760 13734 7788 14214
rect 7748 13728 7800 13734
rect 7748 13670 7800 13676
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 7840 13456 7892 13462
rect 7840 13398 7892 13404
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7760 12850 7788 13126
rect 7852 12850 7880 13398
rect 8220 12900 8248 14894
rect 8312 14278 8340 19264
rect 8482 19272 8538 19281
rect 8482 19207 8538 19216
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 8392 18624 8444 18630
rect 8392 18566 8444 18572
rect 8404 17649 8432 18566
rect 8390 17640 8446 17649
rect 8390 17575 8446 17584
rect 8404 16998 8432 17575
rect 8392 16992 8444 16998
rect 8392 16934 8444 16940
rect 8496 15502 8524 19110
rect 8680 18222 8708 19858
rect 8760 19848 8812 19854
rect 8760 19790 8812 19796
rect 8772 19514 8800 19790
rect 8944 19712 8996 19718
rect 8944 19654 8996 19660
rect 8760 19508 8812 19514
rect 8760 19450 8812 19456
rect 8852 19508 8904 19514
rect 8852 19450 8904 19456
rect 8772 18902 8800 19450
rect 8864 19378 8892 19450
rect 8956 19378 8984 19654
rect 8852 19372 8904 19378
rect 8852 19314 8904 19320
rect 8944 19372 8996 19378
rect 8944 19314 8996 19320
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8760 18896 8812 18902
rect 8760 18838 8812 18844
rect 8772 18290 8800 18838
rect 8760 18284 8812 18290
rect 8760 18226 8812 18232
rect 8864 18222 8892 19110
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 8668 18216 8720 18222
rect 8668 18158 8720 18164
rect 8852 18216 8904 18222
rect 8852 18158 8904 18164
rect 8668 18080 8720 18086
rect 8956 18034 8984 18226
rect 8720 18028 8984 18034
rect 8668 18022 8984 18028
rect 8680 18006 8984 18022
rect 8680 16538 8708 18006
rect 9048 17202 9076 22320
rect 9404 19712 9456 19718
rect 9404 19654 9456 19660
rect 9128 19304 9180 19310
rect 9312 19304 9364 19310
rect 9180 19252 9260 19258
rect 9128 19246 9260 19252
rect 9312 19246 9364 19252
rect 9140 19230 9260 19246
rect 9232 19174 9260 19230
rect 9128 19168 9180 19174
rect 9128 19110 9180 19116
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9140 18426 9168 19110
rect 9324 18970 9352 19246
rect 9312 18964 9364 18970
rect 9312 18906 9364 18912
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9128 18420 9180 18426
rect 9128 18362 9180 18368
rect 9220 18420 9272 18426
rect 9220 18362 9272 18368
rect 9232 17785 9260 18362
rect 9324 18222 9352 18702
rect 9312 18216 9364 18222
rect 9312 18158 9364 18164
rect 9218 17776 9274 17785
rect 9128 17740 9180 17746
rect 9218 17711 9274 17720
rect 9128 17682 9180 17688
rect 9036 17196 9088 17202
rect 9036 17138 9088 17144
rect 9034 17096 9090 17105
rect 9034 17031 9090 17040
rect 9048 16998 9076 17031
rect 8944 16992 8996 16998
rect 8944 16934 8996 16940
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 8680 16510 8800 16538
rect 8772 15858 8800 16510
rect 8956 16046 8984 16934
rect 9140 16726 9168 17682
rect 9324 17678 9352 18158
rect 9416 17882 9444 19654
rect 9508 18714 9536 22320
rect 9588 19440 9640 19446
rect 9640 19388 9720 19394
rect 9588 19382 9720 19388
rect 9600 19366 9720 19382
rect 9588 19304 9640 19310
rect 9588 19246 9640 19252
rect 9600 18850 9628 19246
rect 9692 19009 9720 19366
rect 9678 19000 9734 19009
rect 9678 18935 9734 18944
rect 9600 18822 9720 18850
rect 9692 18766 9720 18822
rect 9680 18760 9732 18766
rect 9508 18686 9628 18714
rect 9680 18702 9732 18708
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 9312 17672 9364 17678
rect 9312 17614 9364 17620
rect 9496 17672 9548 17678
rect 9496 17614 9548 17620
rect 9404 17604 9456 17610
rect 9404 17546 9456 17552
rect 9416 17202 9444 17546
rect 9220 17196 9272 17202
rect 9404 17196 9456 17202
rect 9272 17156 9352 17184
rect 9220 17138 9272 17144
rect 9128 16720 9180 16726
rect 9128 16662 9180 16668
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 9048 16250 9076 16526
rect 9036 16244 9088 16250
rect 9036 16186 9088 16192
rect 8944 16040 8996 16046
rect 8944 15982 8996 15988
rect 8772 15830 9168 15858
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 9048 14482 9076 15438
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 8574 13968 8630 13977
rect 8574 13903 8630 13912
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 8300 12912 8352 12918
rect 8220 12872 8300 12900
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 7838 12336 7894 12345
rect 7838 12271 7894 12280
rect 7852 12238 7880 12271
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 8220 11694 8248 12872
rect 8300 12854 8352 12860
rect 8496 12345 8524 13262
rect 8482 12336 8538 12345
rect 8482 12271 8538 12280
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8392 11688 8444 11694
rect 8496 11676 8524 12271
rect 8444 11648 8524 11676
rect 8392 11630 8444 11636
rect 7820 11452 8116 11472
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 7760 10266 7788 10610
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7760 9058 7788 10066
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 7944 9722 7972 9998
rect 8220 9926 8248 10610
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 7932 9716 7984 9722
rect 7932 9658 7984 9664
rect 8220 9450 8248 9862
rect 8208 9444 8260 9450
rect 8208 9386 8260 9392
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 8312 9178 8340 11154
rect 8496 10470 8524 11648
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8496 10266 8524 10406
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8588 9178 8616 13903
rect 8772 13462 8800 14010
rect 8944 13796 8996 13802
rect 8944 13738 8996 13744
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8760 13456 8812 13462
rect 8760 13398 8812 13404
rect 8758 12880 8814 12889
rect 8758 12815 8814 12824
rect 8772 12782 8800 12815
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8864 11694 8892 13466
rect 8956 12850 8984 13738
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 8852 11688 8904 11694
rect 8852 11630 8904 11636
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8680 9450 8708 10202
rect 8668 9444 8720 9450
rect 8668 9386 8720 9392
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 7760 9030 7880 9058
rect 7852 8974 7880 9030
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 8022 8528 8078 8537
rect 8022 8463 8078 8472
rect 8208 8492 8260 8498
rect 8036 8362 8064 8463
rect 8208 8434 8260 8440
rect 7656 8356 7708 8362
rect 7656 8298 7708 8304
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 8220 8294 8248 8434
rect 8680 8430 8708 9386
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 8128 7546 8156 7890
rect 8588 7546 8616 8298
rect 8680 8090 8708 8366
rect 8852 8356 8904 8362
rect 8852 8298 8904 8304
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8864 7886 8892 8298
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 8864 6798 8892 7822
rect 9048 7342 9076 14214
rect 9140 10577 9168 15830
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 9232 12986 9260 13670
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9324 12424 9352 17156
rect 9404 17138 9456 17144
rect 9404 16992 9456 16998
rect 9404 16934 9456 16940
rect 9416 16046 9444 16934
rect 9508 16794 9536 17614
rect 9496 16788 9548 16794
rect 9496 16730 9548 16736
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 9404 16040 9456 16046
rect 9508 16017 9536 16050
rect 9404 15982 9456 15988
rect 9494 16008 9550 16017
rect 9494 15943 9550 15952
rect 9600 15706 9628 18686
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9692 18154 9720 18566
rect 9680 18148 9732 18154
rect 9680 18090 9732 18096
rect 9772 18148 9824 18154
rect 9772 18090 9824 18096
rect 9784 17882 9812 18090
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9784 17746 9812 17818
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 9678 17504 9734 17513
rect 9678 17439 9734 17448
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 9600 14618 9628 15642
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9692 14249 9720 17439
rect 9876 17320 9904 22320
rect 10232 20052 10284 20058
rect 10232 19994 10284 20000
rect 10140 19916 10192 19922
rect 10140 19858 10192 19864
rect 10152 18442 10180 19858
rect 9968 18426 10180 18442
rect 9956 18420 10180 18426
rect 10008 18414 10180 18420
rect 9956 18362 10008 18368
rect 9876 17292 9996 17320
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9876 16522 9904 17138
rect 9864 16516 9916 16522
rect 9864 16458 9916 16464
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9784 16114 9812 16390
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9784 14770 9812 15098
rect 9876 14958 9904 16458
rect 9968 15094 9996 17292
rect 10046 17232 10102 17241
rect 10046 17167 10102 17176
rect 10060 17066 10088 17167
rect 10048 17060 10100 17066
rect 10048 17002 10100 17008
rect 10152 16946 10180 18414
rect 10244 17746 10272 19994
rect 10232 17740 10284 17746
rect 10232 17682 10284 17688
rect 10244 17066 10272 17682
rect 10232 17060 10284 17066
rect 10232 17002 10284 17008
rect 10152 16918 10272 16946
rect 10138 16824 10194 16833
rect 10138 16759 10194 16768
rect 10048 16040 10100 16046
rect 10046 16008 10048 16017
rect 10100 16008 10102 16017
rect 10046 15943 10102 15952
rect 10060 15502 10088 15943
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 10060 15162 10088 15438
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 9956 15088 10008 15094
rect 9956 15030 10008 15036
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9968 14890 9996 15030
rect 9956 14884 10008 14890
rect 9956 14826 10008 14832
rect 9784 14742 9996 14770
rect 9678 14240 9734 14249
rect 9678 14175 9734 14184
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 9416 13530 9444 13874
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9324 12396 9444 12424
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9232 11898 9260 12038
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9324 11830 9352 12242
rect 9312 11824 9364 11830
rect 9312 11766 9364 11772
rect 9416 11694 9444 12396
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9416 11354 9444 11630
rect 9588 11552 9640 11558
rect 9588 11494 9640 11500
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9404 11348 9456 11354
rect 9404 11290 9456 11296
rect 9600 11286 9628 11494
rect 9220 11280 9272 11286
rect 9220 11222 9272 11228
rect 9588 11280 9640 11286
rect 9588 11222 9640 11228
rect 9232 10674 9260 11222
rect 9784 11150 9812 11494
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9220 10668 9272 10674
rect 9220 10610 9272 10616
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9126 10568 9182 10577
rect 9126 10503 9182 10512
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9140 10266 9168 10406
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9324 9926 9352 10610
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9692 8906 9720 11018
rect 9784 10130 9812 11086
rect 9876 10266 9904 13466
rect 9968 11762 9996 14742
rect 10048 14408 10100 14414
rect 10046 14376 10048 14385
rect 10100 14376 10102 14385
rect 10046 14311 10102 14320
rect 10046 14240 10102 14249
rect 10046 14175 10102 14184
rect 10060 13802 10088 14175
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 10060 12889 10088 13738
rect 10152 13410 10180 16759
rect 10244 13530 10272 16918
rect 10336 14958 10364 22320
rect 10416 19848 10468 19854
rect 10416 19790 10468 19796
rect 10428 17814 10456 19790
rect 10508 19168 10560 19174
rect 10508 19110 10560 19116
rect 10416 17808 10468 17814
rect 10416 17750 10468 17756
rect 10428 16697 10456 17750
rect 10414 16688 10470 16697
rect 10414 16623 10470 16632
rect 10416 15428 10468 15434
rect 10416 15370 10468 15376
rect 10324 14952 10376 14958
rect 10324 14894 10376 14900
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 10152 13382 10272 13410
rect 10046 12880 10102 12889
rect 10046 12815 10102 12824
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 9956 11552 10008 11558
rect 9956 11494 10008 11500
rect 9968 11218 9996 11494
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 10060 9110 10088 11154
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 10152 9110 10180 11086
rect 10244 11014 10272 13382
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 10244 10713 10272 10950
rect 10230 10704 10286 10713
rect 10230 10639 10286 10648
rect 10232 9444 10284 9450
rect 10232 9386 10284 9392
rect 10244 9178 10272 9386
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 10140 9104 10192 9110
rect 10140 9046 10192 9052
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 10336 8412 10364 14758
rect 10428 14657 10456 15370
rect 10414 14648 10470 14657
rect 10414 14583 10470 14592
rect 10416 14408 10468 14414
rect 10416 14350 10468 14356
rect 10428 13938 10456 14350
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10244 8384 10364 8412
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9232 8090 9260 8230
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 9048 7206 9076 7278
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 10244 6186 10272 8384
rect 10324 8288 10376 8294
rect 10324 8230 10376 8236
rect 10336 6730 10364 8230
rect 10428 7954 10456 11698
rect 10520 11150 10548 19110
rect 10598 17912 10654 17921
rect 10598 17847 10654 17856
rect 10612 17134 10640 17847
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10704 15722 10732 22320
rect 11164 20074 11192 22320
rect 11072 20046 11192 20074
rect 11624 20058 11652 22320
rect 11612 20052 11664 20058
rect 11072 19802 11100 20046
rect 11612 19994 11664 20000
rect 11152 19916 11204 19922
rect 11152 19858 11204 19864
rect 11612 19916 11664 19922
rect 11612 19858 11664 19864
rect 10980 19774 11100 19802
rect 10874 19000 10930 19009
rect 10874 18935 10930 18944
rect 10888 18834 10916 18935
rect 10876 18828 10928 18834
rect 10876 18770 10928 18776
rect 10980 18714 11008 19774
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 11072 18834 11100 19654
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 10980 18686 11100 18714
rect 10874 18592 10930 18601
rect 10874 18527 10930 18536
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10796 16998 10824 18362
rect 10888 17660 10916 18527
rect 10968 18080 11020 18086
rect 10968 18022 11020 18028
rect 10980 17785 11008 18022
rect 10966 17776 11022 17785
rect 10966 17711 11022 17720
rect 10888 17632 11008 17660
rect 10876 17332 10928 17338
rect 10876 17274 10928 17280
rect 10888 17134 10916 17274
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10980 17066 11008 17632
rect 10968 17060 11020 17066
rect 10968 17002 11020 17008
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10876 16652 10928 16658
rect 10876 16594 10928 16600
rect 10612 15694 10732 15722
rect 10888 15706 10916 16594
rect 10876 15700 10928 15706
rect 10612 15042 10640 15694
rect 10876 15642 10928 15648
rect 10692 15564 10744 15570
rect 10692 15506 10744 15512
rect 10704 15162 10732 15506
rect 10782 15328 10838 15337
rect 10782 15263 10838 15272
rect 10692 15156 10744 15162
rect 10692 15098 10744 15104
rect 10612 15014 10732 15042
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 10612 12374 10640 14894
rect 10600 12368 10652 12374
rect 10600 12310 10652 12316
rect 10598 11656 10654 11665
rect 10598 11591 10654 11600
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 10612 10130 10640 11591
rect 10704 11218 10732 15014
rect 10796 14958 10824 15263
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 10874 14920 10930 14929
rect 10874 14855 10876 14864
rect 10928 14855 10930 14864
rect 10876 14826 10928 14832
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10796 14618 10824 14758
rect 10874 14648 10930 14657
rect 10784 14612 10836 14618
rect 10874 14583 10930 14592
rect 10784 14554 10836 14560
rect 10784 14408 10836 14414
rect 10782 14376 10784 14385
rect 10836 14376 10838 14385
rect 10782 14311 10838 14320
rect 10888 13530 10916 14583
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10980 13938 11008 14214
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 10784 12300 10836 12306
rect 10784 12242 10836 12248
rect 10796 12209 10824 12242
rect 10782 12200 10838 12209
rect 10782 12135 10838 12144
rect 10888 11762 10916 12310
rect 10968 12164 11020 12170
rect 10968 12106 11020 12112
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10796 11257 10824 11698
rect 10980 11694 11008 12106
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 10782 11248 10838 11257
rect 10692 11212 10744 11218
rect 10782 11183 10838 11192
rect 10692 11154 10744 11160
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10980 10606 11008 11086
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 10888 9178 10916 9522
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10704 8090 10732 8230
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10416 7948 10468 7954
rect 10416 7890 10468 7896
rect 10428 6934 10456 7890
rect 10416 6928 10468 6934
rect 10416 6870 10468 6876
rect 10888 6769 10916 8978
rect 10980 8498 11008 9318
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10980 7886 11008 8434
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 11072 7206 11100 18686
rect 11164 17882 11192 19858
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 11152 17740 11204 17746
rect 11152 17682 11204 17688
rect 11164 16833 11192 17682
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 11624 17338 11652 19858
rect 11888 19848 11940 19854
rect 11888 19790 11940 19796
rect 11796 19780 11848 19786
rect 11796 19722 11848 19728
rect 11704 19304 11756 19310
rect 11704 19246 11756 19252
rect 11716 18426 11744 19246
rect 11808 19174 11836 19722
rect 11900 19242 11928 19790
rect 11888 19236 11940 19242
rect 11888 19178 11940 19184
rect 11796 19168 11848 19174
rect 11796 19110 11848 19116
rect 11886 19136 11942 19145
rect 11886 19071 11942 19080
rect 11900 18986 11928 19071
rect 11808 18958 11928 18986
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 11716 17660 11744 18362
rect 11808 17814 11836 18958
rect 11796 17808 11848 17814
rect 11796 17750 11848 17756
rect 11796 17672 11848 17678
rect 11716 17632 11796 17660
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11716 17134 11744 17632
rect 11796 17614 11848 17620
rect 11704 17128 11756 17134
rect 11704 17070 11756 17076
rect 11520 17060 11572 17066
rect 11520 17002 11572 17008
rect 11532 16969 11560 17002
rect 11704 16992 11756 16998
rect 11518 16960 11574 16969
rect 11704 16934 11756 16940
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11518 16895 11574 16904
rect 11150 16824 11206 16833
rect 11150 16759 11206 16768
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 11164 16250 11192 16526
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11164 15502 11192 16186
rect 11624 16046 11652 16730
rect 11716 16658 11744 16934
rect 11900 16794 11928 16934
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11992 16096 12020 22320
rect 12256 20052 12308 20058
rect 12256 19994 12308 20000
rect 12072 19916 12124 19922
rect 12072 19858 12124 19864
rect 11808 16068 12020 16096
rect 11612 16040 11664 16046
rect 11612 15982 11664 15988
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11256 15348 11284 15506
rect 11164 15320 11284 15348
rect 11704 15360 11756 15366
rect 11164 14074 11192 15320
rect 11704 15302 11756 15308
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 11716 15162 11744 15302
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11520 15088 11572 15094
rect 11520 15030 11572 15036
rect 11612 15088 11664 15094
rect 11612 15030 11664 15036
rect 11244 14884 11296 14890
rect 11244 14826 11296 14832
rect 11256 14618 11284 14826
rect 11532 14618 11560 15030
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 11520 14612 11572 14618
rect 11520 14554 11572 14560
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11520 14000 11572 14006
rect 11150 13968 11206 13977
rect 11520 13942 11572 13948
rect 11150 13903 11152 13912
rect 11204 13903 11206 13912
rect 11152 13874 11204 13880
rect 11532 13394 11560 13942
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 11152 12232 11204 12238
rect 11152 12174 11204 12180
rect 11164 10538 11192 12174
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11152 10532 11204 10538
rect 11152 10474 11204 10480
rect 11164 10010 11192 10474
rect 11336 10056 11388 10062
rect 11164 10004 11336 10010
rect 11164 9998 11388 10004
rect 11164 9982 11376 9998
rect 11164 8838 11192 9982
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11624 7274 11652 15030
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11716 12986 11744 14894
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11808 12050 11836 16068
rect 11980 15972 12032 15978
rect 11980 15914 12032 15920
rect 11992 15366 12020 15914
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 12084 15094 12112 19858
rect 12164 19712 12216 19718
rect 12164 19654 12216 19660
rect 12176 19417 12204 19654
rect 12162 19408 12218 19417
rect 12162 19343 12218 19352
rect 12164 18828 12216 18834
rect 12164 18770 12216 18776
rect 12176 15162 12204 18770
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 12072 15088 12124 15094
rect 12072 15030 12124 15036
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 11900 14550 11928 14894
rect 11980 14816 12032 14822
rect 11980 14758 12032 14764
rect 11888 14544 11940 14550
rect 11888 14486 11940 14492
rect 11992 14074 12020 14758
rect 12072 14544 12124 14550
rect 12072 14486 12124 14492
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 12084 13870 12112 14486
rect 12176 13938 12204 14962
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 12162 13832 12218 13841
rect 12162 13767 12218 13776
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11900 13190 11928 13466
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11716 12022 11836 12050
rect 11716 11665 11744 12022
rect 11900 11898 11928 12378
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11702 11656 11758 11665
rect 11702 11591 11758 11600
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11716 11150 11744 11494
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11808 10742 11836 11834
rect 11978 11792 12034 11801
rect 11978 11727 12034 11736
rect 11888 11620 11940 11626
rect 11888 11562 11940 11568
rect 11900 11014 11928 11562
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11796 10736 11848 10742
rect 11796 10678 11848 10684
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11808 10198 11836 10406
rect 11796 10192 11848 10198
rect 11796 10134 11848 10140
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11716 7478 11744 9114
rect 11900 8974 11928 10950
rect 11992 9110 12020 11727
rect 12084 10690 12112 12922
rect 12176 10810 12204 13767
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12084 10662 12204 10690
rect 12070 9888 12126 9897
rect 12070 9823 12126 9832
rect 11980 9104 12032 9110
rect 11980 9046 12032 9052
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 11796 8900 11848 8906
rect 11796 8842 11848 8848
rect 11808 8362 11836 8842
rect 11992 8430 12020 9046
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 11796 8356 11848 8362
rect 11796 8298 11848 8304
rect 11704 7472 11756 7478
rect 11704 7414 11756 7420
rect 11612 7268 11664 7274
rect 11612 7210 11664 7216
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 10874 6760 10930 6769
rect 10324 6724 10376 6730
rect 10874 6695 10930 6704
rect 10324 6666 10376 6672
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 10232 6180 10284 6186
rect 10232 6122 10284 6128
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11716 5302 11744 7414
rect 12084 6866 12112 9823
rect 12176 9178 12204 10662
rect 12164 9172 12216 9178
rect 12164 9114 12216 9120
rect 12268 8922 12296 19994
rect 12346 19136 12402 19145
rect 12346 19071 12402 19080
rect 12360 18902 12388 19071
rect 12348 18896 12400 18902
rect 12348 18838 12400 18844
rect 12452 17218 12480 22320
rect 12714 19544 12770 19553
rect 12714 19479 12716 19488
rect 12768 19479 12770 19488
rect 12716 19450 12768 19456
rect 12820 19394 12848 22320
rect 13280 20040 13308 22320
rect 13004 20012 13308 20040
rect 12820 19366 12940 19394
rect 12716 19236 12768 19242
rect 12716 19178 12768 19184
rect 12808 19236 12860 19242
rect 12808 19178 12860 19184
rect 12624 18896 12676 18902
rect 12624 18838 12676 18844
rect 12636 17678 12664 18838
rect 12728 18766 12756 19178
rect 12716 18760 12768 18766
rect 12716 18702 12768 18708
rect 12728 18290 12756 18702
rect 12820 18698 12848 19178
rect 12808 18692 12860 18698
rect 12808 18634 12860 18640
rect 12820 18358 12848 18634
rect 12808 18352 12860 18358
rect 12808 18294 12860 18300
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 12808 17876 12860 17882
rect 12808 17818 12860 17824
rect 12624 17672 12676 17678
rect 12820 17649 12848 17818
rect 12624 17614 12676 17620
rect 12806 17640 12862 17649
rect 12636 17377 12664 17614
rect 12806 17575 12862 17584
rect 12622 17368 12678 17377
rect 12622 17303 12678 17312
rect 12452 17190 12664 17218
rect 12346 17096 12402 17105
rect 12346 17031 12402 17040
rect 12360 16794 12388 17031
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12346 16688 12402 16697
rect 12346 16623 12402 16632
rect 12360 16590 12388 16623
rect 12348 16584 12400 16590
rect 12348 16526 12400 16532
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12452 16182 12480 16390
rect 12440 16176 12492 16182
rect 12440 16118 12492 16124
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 12452 15570 12480 15982
rect 12636 15638 12664 17190
rect 12808 16516 12860 16522
rect 12808 16458 12860 16464
rect 12820 15978 12848 16458
rect 12808 15972 12860 15978
rect 12808 15914 12860 15920
rect 12624 15632 12676 15638
rect 12624 15574 12676 15580
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12452 14618 12480 15506
rect 12636 14906 12664 15574
rect 12820 15434 12848 15914
rect 12808 15428 12860 15434
rect 12808 15370 12860 15376
rect 12716 15088 12768 15094
rect 12716 15030 12768 15036
rect 12544 14878 12664 14906
rect 12544 14618 12572 14878
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12636 14618 12664 14758
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12624 14612 12676 14618
rect 12624 14554 12676 14560
rect 12452 14006 12480 14554
rect 12440 14000 12492 14006
rect 12440 13942 12492 13948
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12636 13297 12664 13466
rect 12622 13288 12678 13297
rect 12622 13223 12678 13232
rect 12348 12368 12400 12374
rect 12348 12310 12400 12316
rect 12438 12336 12494 12345
rect 12360 11626 12388 12310
rect 12438 12271 12440 12280
rect 12492 12271 12494 12280
rect 12440 12242 12492 12248
rect 12728 12238 12756 15030
rect 12912 14958 12940 19366
rect 13004 15094 13032 20012
rect 13268 19916 13320 19922
rect 13268 19858 13320 19864
rect 13176 19780 13228 19786
rect 13176 19722 13228 19728
rect 13188 19145 13216 19722
rect 13174 19136 13230 19145
rect 13174 19071 13230 19080
rect 13280 18426 13308 19858
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 13372 18970 13400 19790
rect 13556 19174 13584 19790
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13360 18964 13412 18970
rect 13360 18906 13412 18912
rect 13556 18902 13584 19110
rect 13544 18896 13596 18902
rect 13544 18838 13596 18844
rect 13358 18456 13414 18465
rect 13268 18420 13320 18426
rect 13358 18391 13414 18400
rect 13268 18362 13320 18368
rect 13084 18352 13136 18358
rect 13084 18294 13136 18300
rect 13096 16046 13124 18294
rect 13372 18154 13400 18391
rect 13360 18148 13412 18154
rect 13360 18090 13412 18096
rect 13372 18057 13400 18090
rect 13358 18048 13414 18057
rect 13358 17983 13414 17992
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13280 17134 13308 17478
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13372 16794 13400 17070
rect 13360 16788 13412 16794
rect 13360 16730 13412 16736
rect 13556 16522 13584 17614
rect 13544 16516 13596 16522
rect 13544 16458 13596 16464
rect 13084 16040 13136 16046
rect 13084 15982 13136 15988
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 13176 15496 13228 15502
rect 13176 15438 13228 15444
rect 13084 15156 13136 15162
rect 13084 15098 13136 15104
rect 12992 15088 13044 15094
rect 12992 15030 13044 15036
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12912 13462 12940 14894
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 13004 13530 13032 14758
rect 12992 13524 13044 13530
rect 12992 13466 13044 13472
rect 12900 13456 12952 13462
rect 12900 13398 12952 13404
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 12348 11620 12400 11626
rect 12348 11562 12400 11568
rect 12728 11150 12756 12174
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12624 11076 12676 11082
rect 12624 11018 12676 11024
rect 12532 11008 12584 11014
rect 12532 10950 12584 10956
rect 12544 10810 12572 10950
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12636 10674 12664 11018
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 12360 9926 12388 10542
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12360 9518 12388 9862
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12176 8894 12296 8922
rect 12176 8090 12204 8894
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 12268 8498 12296 8774
rect 12452 8634 12480 9998
rect 12624 9444 12676 9450
rect 12624 9386 12676 9392
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12346 8528 12402 8537
rect 12256 8492 12308 8498
rect 12346 8463 12402 8472
rect 12256 8434 12308 8440
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 12360 6225 12388 8463
rect 12544 8430 12572 9318
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12636 8090 12664 9386
rect 12820 9110 12848 13330
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 13004 11286 13032 12582
rect 12992 11280 13044 11286
rect 12992 11222 13044 11228
rect 12992 11144 13044 11150
rect 13096 11121 13124 15098
rect 13188 13433 13216 15438
rect 13556 15162 13584 15982
rect 13544 15156 13596 15162
rect 13544 15098 13596 15104
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13464 14278 13492 14962
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13464 13870 13492 14214
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 13174 13424 13230 13433
rect 13174 13359 13230 13368
rect 13188 13258 13216 13359
rect 13556 13326 13584 14418
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13648 13274 13676 22320
rect 14108 19802 14136 22320
rect 14280 19916 14332 19922
rect 14280 19858 14332 19864
rect 14016 19774 14136 19802
rect 14016 19009 14044 19774
rect 14096 19712 14148 19718
rect 14096 19654 14148 19660
rect 14188 19712 14240 19718
rect 14188 19654 14240 19660
rect 14108 19310 14136 19654
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 14002 19000 14058 19009
rect 14002 18935 14058 18944
rect 14200 18306 14228 19654
rect 14292 19378 14320 19858
rect 14280 19372 14332 19378
rect 14280 19314 14332 19320
rect 14568 19242 14596 22320
rect 14936 20244 14964 22320
rect 14936 20216 15148 20244
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 14556 19236 14608 19242
rect 14556 19178 14608 19184
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 14556 18624 14608 18630
rect 14556 18566 14608 18572
rect 14016 18278 14228 18306
rect 14016 17882 14044 18278
rect 14568 18222 14596 18566
rect 14188 18216 14240 18222
rect 14188 18158 14240 18164
rect 14556 18216 14608 18222
rect 14556 18158 14608 18164
rect 14004 17876 14056 17882
rect 14004 17818 14056 17824
rect 14200 17814 14228 18158
rect 14372 18148 14424 18154
rect 14372 18090 14424 18096
rect 14188 17808 14240 17814
rect 13726 17776 13782 17785
rect 14188 17750 14240 17756
rect 13726 17711 13782 17720
rect 13740 17678 13768 17711
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13740 16658 13768 17614
rect 14188 17264 14240 17270
rect 14186 17232 14188 17241
rect 14240 17232 14242 17241
rect 13820 17196 13872 17202
rect 14186 17167 14242 17176
rect 13820 17138 13872 17144
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 13832 16250 13860 17138
rect 14004 17128 14056 17134
rect 14004 17070 14056 17076
rect 14096 17128 14148 17134
rect 14096 17070 14148 17076
rect 14186 17096 14242 17105
rect 14016 16454 14044 17070
rect 14108 16794 14136 17070
rect 14186 17031 14242 17040
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 14096 16652 14148 16658
rect 14096 16594 14148 16600
rect 14004 16448 14056 16454
rect 14004 16390 14056 16396
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 14108 15706 14136 16594
rect 14096 15700 14148 15706
rect 14096 15642 14148 15648
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13832 14346 13860 14894
rect 14096 14476 14148 14482
rect 14096 14418 14148 14424
rect 13820 14340 13872 14346
rect 13820 14282 13872 14288
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13832 13462 13860 13670
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13176 13252 13228 13258
rect 13648 13246 13860 13274
rect 13176 13194 13228 13200
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13544 12912 13596 12918
rect 13544 12854 13596 12860
rect 13556 12753 13584 12854
rect 13740 12850 13768 13126
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13636 12776 13688 12782
rect 13542 12744 13598 12753
rect 13832 12730 13860 13246
rect 13636 12718 13688 12724
rect 13542 12679 13598 12688
rect 13648 12442 13676 12718
rect 13740 12702 13860 12730
rect 13636 12436 13688 12442
rect 13636 12378 13688 12384
rect 13648 11694 13676 12378
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13740 11150 13768 12702
rect 14004 12640 14056 12646
rect 14004 12582 14056 12588
rect 14016 12322 14044 12582
rect 13924 12294 14044 12322
rect 13924 11694 13952 12294
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 13924 11150 13952 11494
rect 14108 11286 14136 14418
rect 14096 11280 14148 11286
rect 14096 11222 14148 11228
rect 14200 11234 14228 17031
rect 14384 16969 14412 18090
rect 14568 17678 14596 18158
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 15120 17338 15148 20216
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 15212 17882 15240 19110
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 15304 17746 15332 19858
rect 15292 17740 15344 17746
rect 15292 17682 15344 17688
rect 15396 17338 15424 22320
rect 15476 19372 15528 19378
rect 15476 19314 15528 19320
rect 15488 18902 15516 19314
rect 15476 18896 15528 18902
rect 15476 18838 15528 18844
rect 15488 18426 15516 18838
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15764 18358 15792 22320
rect 16224 19258 16252 22320
rect 16684 20058 16712 22320
rect 16672 20052 16724 20058
rect 16672 19994 16724 20000
rect 17052 19786 17080 22320
rect 17512 20058 17540 22320
rect 17500 20052 17552 20058
rect 17500 19994 17552 20000
rect 17880 19990 17908 22320
rect 17868 19984 17920 19990
rect 17868 19926 17920 19932
rect 17224 19916 17276 19922
rect 17224 19858 17276 19864
rect 17040 19780 17092 19786
rect 17040 19722 17092 19728
rect 16856 19712 16908 19718
rect 16856 19654 16908 19660
rect 16868 19378 16896 19654
rect 17236 19553 17264 19858
rect 17408 19848 17460 19854
rect 18340 19802 18368 22320
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 18696 19916 18748 19922
rect 18696 19858 18748 19864
rect 17408 19790 17460 19796
rect 17222 19544 17278 19553
rect 17222 19479 17278 19488
rect 17236 19446 17264 19479
rect 17224 19440 17276 19446
rect 17224 19382 17276 19388
rect 16856 19372 16908 19378
rect 16856 19314 16908 19320
rect 16224 19230 16620 19258
rect 15936 19168 15988 19174
rect 15936 19110 15988 19116
rect 15948 18426 15976 19110
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 16028 18420 16080 18426
rect 16028 18362 16080 18368
rect 15752 18352 15804 18358
rect 15752 18294 15804 18300
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15750 17776 15806 17785
rect 15750 17711 15752 17720
rect 15804 17711 15806 17720
rect 15752 17682 15804 17688
rect 15856 17678 15884 18226
rect 16040 18086 16068 18362
rect 16028 18080 16080 18086
rect 16028 18022 16080 18028
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15108 17332 15160 17338
rect 15108 17274 15160 17280
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 16028 17128 16080 17134
rect 16132 17116 16160 18566
rect 16304 18148 16356 18154
rect 16304 18090 16356 18096
rect 16080 17088 16160 17116
rect 16028 17070 16080 17076
rect 14556 17060 14608 17066
rect 14556 17002 14608 17008
rect 14370 16960 14426 16969
rect 14370 16895 14426 16904
rect 14568 16794 14596 17002
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14740 16720 14792 16726
rect 14924 16720 14976 16726
rect 14792 16668 14924 16674
rect 14740 16662 14976 16668
rect 14752 16646 14964 16662
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 15108 16516 15160 16522
rect 15108 16458 15160 16464
rect 14372 16040 14424 16046
rect 14372 15982 14424 15988
rect 14384 15570 14412 15982
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 14462 15600 14518 15609
rect 14372 15564 14424 15570
rect 14462 15535 14518 15544
rect 14372 15506 14424 15512
rect 14476 15162 14504 15535
rect 14556 15496 14608 15502
rect 14556 15438 14608 15444
rect 14568 15162 14596 15438
rect 14464 15156 14516 15162
rect 14464 15098 14516 15104
rect 14556 15156 14608 15162
rect 14556 15098 14608 15104
rect 15120 15026 15148 16458
rect 15212 15570 15240 16594
rect 15476 16584 15528 16590
rect 15476 16526 15528 16532
rect 15292 16448 15344 16454
rect 15292 16390 15344 16396
rect 15304 15706 15332 16390
rect 15488 16250 15516 16526
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 15200 15564 15252 15570
rect 15200 15506 15252 15512
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 14832 14544 14884 14550
rect 14832 14486 14884 14492
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14384 13734 14412 14350
rect 14844 14074 14872 14486
rect 15016 14476 15068 14482
rect 15016 14418 15068 14424
rect 15028 14074 15056 14418
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 15108 14000 15160 14006
rect 15108 13942 15160 13948
rect 14556 13796 14608 13802
rect 14556 13738 14608 13744
rect 15016 13796 15068 13802
rect 15016 13738 15068 13744
rect 14372 13728 14424 13734
rect 14372 13670 14424 13676
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14292 12102 14320 13262
rect 14384 12782 14412 13670
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14372 12776 14424 12782
rect 14372 12718 14424 12724
rect 14476 12374 14504 13262
rect 14464 12368 14516 12374
rect 14464 12310 14516 12316
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 14476 11762 14504 12310
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14200 11206 14320 11234
rect 13268 11144 13320 11150
rect 12992 11086 13044 11092
rect 13082 11112 13138 11121
rect 13004 10656 13032 11086
rect 13268 11086 13320 11092
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 13082 11047 13138 11056
rect 13084 10668 13136 10674
rect 13004 10628 13084 10656
rect 13004 10470 13032 10628
rect 13084 10610 13136 10616
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 12992 10260 13044 10266
rect 12992 10202 13044 10208
rect 13004 9722 13032 10202
rect 12992 9716 13044 9722
rect 12992 9658 13044 9664
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 12808 9104 12860 9110
rect 12808 9046 12860 9052
rect 12992 9104 13044 9110
rect 12992 9046 13044 9052
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12912 8294 12940 8978
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12912 7886 12940 8230
rect 13004 8090 13032 9046
rect 13096 9042 13124 9522
rect 13280 9518 13308 11086
rect 13636 10532 13688 10538
rect 13636 10474 13688 10480
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13556 10266 13584 10406
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13648 10062 13676 10474
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 13924 10266 13952 10406
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 13636 10056 13688 10062
rect 14108 10033 14136 10066
rect 14200 10062 14228 11086
rect 14292 10266 14320 11206
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 14188 10056 14240 10062
rect 13636 9998 13688 10004
rect 14094 10024 14150 10033
rect 14188 9998 14240 10004
rect 14094 9959 14150 9968
rect 14292 9654 14320 10202
rect 14568 10169 14596 13738
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 15028 11778 15056 13738
rect 15120 13530 15148 13942
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 15212 12594 15240 15506
rect 16040 15502 16068 17070
rect 16316 16561 16344 18090
rect 16592 17882 16620 19230
rect 16856 19236 16908 19242
rect 16856 19178 16908 19184
rect 16672 18624 16724 18630
rect 16672 18566 16724 18572
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 16684 17338 16712 18566
rect 16868 17814 16896 19178
rect 17040 19168 17092 19174
rect 17040 19110 17092 19116
rect 17052 18426 17080 19110
rect 17420 18902 17448 19790
rect 17972 19774 18368 19802
rect 17500 19236 17552 19242
rect 17500 19178 17552 19184
rect 17408 18896 17460 18902
rect 17408 18838 17460 18844
rect 17130 18456 17186 18465
rect 17040 18420 17092 18426
rect 17130 18391 17132 18400
rect 17040 18362 17092 18368
rect 17184 18391 17186 18400
rect 17132 18362 17184 18368
rect 17224 18352 17276 18358
rect 17224 18294 17276 18300
rect 16856 17808 16908 17814
rect 16856 17750 16908 17756
rect 16948 17740 17000 17746
rect 16948 17682 17000 17688
rect 16764 17536 16816 17542
rect 16764 17478 16816 17484
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16776 16998 16804 17478
rect 16960 17338 16988 17682
rect 16948 17332 17000 17338
rect 16948 17274 17000 17280
rect 16764 16992 16816 16998
rect 16764 16934 16816 16940
rect 16672 16720 16724 16726
rect 16672 16662 16724 16668
rect 16302 16552 16358 16561
rect 16302 16487 16358 16496
rect 16316 16266 16344 16487
rect 16316 16250 16436 16266
rect 16316 16244 16448 16250
rect 16316 16238 16396 16244
rect 16396 16186 16448 16192
rect 16028 15496 16080 15502
rect 16028 15438 16080 15444
rect 15660 14952 15712 14958
rect 15658 14920 15660 14929
rect 15712 14920 15714 14929
rect 15658 14855 15714 14864
rect 15936 14884 15988 14890
rect 15936 14826 15988 14832
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15384 14340 15436 14346
rect 15384 14282 15436 14288
rect 15292 13728 15344 13734
rect 15292 13670 15344 13676
rect 15304 13530 15332 13670
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15120 12566 15240 12594
rect 15120 11898 15148 12566
rect 15304 12442 15332 13262
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 15028 11750 15240 11778
rect 15016 11620 15068 11626
rect 15016 11562 15068 11568
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 15028 10810 15056 11562
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 14554 10160 14610 10169
rect 15120 10130 15148 11018
rect 14554 10095 14610 10104
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 15028 9178 15056 9386
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 13084 9036 13136 9042
rect 13084 8978 13136 8984
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15120 8362 15148 8774
rect 15108 8356 15160 8362
rect 15108 8298 15160 8304
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 15212 7750 15240 11750
rect 15396 11694 15424 14282
rect 15488 13161 15516 14758
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 15580 13410 15608 13466
rect 15580 13382 15700 13410
rect 15474 13152 15530 13161
rect 15474 13087 15530 13096
rect 15488 12918 15516 13087
rect 15476 12912 15528 12918
rect 15476 12854 15528 12860
rect 15568 12708 15620 12714
rect 15568 12650 15620 12656
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 15488 12345 15516 12582
rect 15580 12374 15608 12650
rect 15568 12368 15620 12374
rect 15474 12336 15530 12345
rect 15568 12310 15620 12316
rect 15474 12271 15530 12280
rect 15488 12102 15516 12271
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15304 11218 15332 11494
rect 15382 11248 15438 11257
rect 15292 11212 15344 11218
rect 15382 11183 15384 11192
rect 15292 11154 15344 11160
rect 15436 11183 15438 11192
rect 15384 11154 15436 11160
rect 15488 10674 15516 12038
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15580 11762 15608 11834
rect 15672 11830 15700 13382
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15764 11898 15792 12922
rect 15844 12640 15896 12646
rect 15844 12582 15896 12588
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15660 11824 15712 11830
rect 15660 11766 15712 11772
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 15304 9178 15332 10066
rect 15384 9988 15436 9994
rect 15384 9930 15436 9936
rect 15396 9518 15424 9930
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15384 8968 15436 8974
rect 15384 8910 15436 8916
rect 15396 8498 15424 8910
rect 15384 8492 15436 8498
rect 15384 8434 15436 8440
rect 15580 7954 15608 11698
rect 15856 11626 15884 12582
rect 15844 11620 15896 11626
rect 15844 11562 15896 11568
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15764 8634 15792 9998
rect 15948 9518 15976 14826
rect 16040 12986 16068 15438
rect 16684 14929 16712 16662
rect 16776 16590 16804 16934
rect 16948 16720 17000 16726
rect 16948 16662 17000 16668
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16762 16008 16818 16017
rect 16762 15943 16818 15952
rect 16670 14920 16726 14929
rect 16670 14855 16726 14864
rect 16302 14512 16358 14521
rect 16212 14476 16264 14482
rect 16302 14447 16358 14456
rect 16212 14418 16264 14424
rect 16224 14226 16252 14418
rect 16316 14414 16344 14447
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 16224 14198 16528 14226
rect 16500 13954 16528 14198
rect 16592 14074 16620 14350
rect 16776 14346 16804 15943
rect 16868 14890 16896 16050
rect 16856 14884 16908 14890
rect 16856 14826 16908 14832
rect 16960 14822 16988 16662
rect 17236 16658 17264 18294
rect 17420 18290 17448 18838
rect 17408 18284 17460 18290
rect 17408 18226 17460 18232
rect 17408 18080 17460 18086
rect 17408 18022 17460 18028
rect 17420 17270 17448 18022
rect 17408 17264 17460 17270
rect 17408 17206 17460 17212
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17052 15450 17080 16594
rect 17132 16584 17184 16590
rect 17420 16538 17448 17206
rect 17132 16526 17184 16532
rect 17144 15910 17172 16526
rect 17236 16510 17448 16538
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 17144 15638 17172 15846
rect 17132 15632 17184 15638
rect 17132 15574 17184 15580
rect 17052 15434 17172 15450
rect 17040 15428 17172 15434
rect 17092 15422 17172 15428
rect 17040 15370 17092 15376
rect 17052 15339 17080 15370
rect 17038 15056 17094 15065
rect 17038 14991 17094 15000
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 17052 14550 17080 14991
rect 17040 14544 17092 14550
rect 17040 14486 17092 14492
rect 16856 14408 16908 14414
rect 16856 14350 16908 14356
rect 16764 14340 16816 14346
rect 16764 14282 16816 14288
rect 16868 14226 16896 14350
rect 16776 14198 16896 14226
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16396 13932 16448 13938
rect 16500 13926 16620 13954
rect 16396 13874 16448 13880
rect 16212 13796 16264 13802
rect 16212 13738 16264 13744
rect 16118 13696 16174 13705
rect 16118 13631 16174 13640
rect 16132 13297 16160 13631
rect 16118 13288 16174 13297
rect 16118 13223 16174 13232
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 16132 12850 16160 13223
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 16132 12646 16160 12786
rect 16120 12640 16172 12646
rect 16120 12582 16172 12588
rect 16120 12300 16172 12306
rect 16120 12242 16172 12248
rect 16132 11694 16160 12242
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 16028 11348 16080 11354
rect 16028 11290 16080 11296
rect 15936 9512 15988 9518
rect 15936 9454 15988 9460
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 16040 8362 16068 11290
rect 16132 10062 16160 11630
rect 16224 10538 16252 13738
rect 16302 13560 16358 13569
rect 16408 13530 16436 13874
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16302 13495 16358 13504
rect 16396 13524 16448 13530
rect 16316 13462 16344 13495
rect 16396 13466 16448 13472
rect 16304 13456 16356 13462
rect 16304 13398 16356 13404
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16316 12986 16344 13262
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 16408 12238 16436 12786
rect 16396 12232 16448 12238
rect 16396 12174 16448 12180
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16408 11898 16436 12038
rect 16396 11892 16448 11898
rect 16396 11834 16448 11840
rect 16500 11778 16528 13806
rect 16408 11750 16528 11778
rect 16212 10532 16264 10538
rect 16212 10474 16264 10480
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 16224 9722 16252 10066
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16316 8974 16344 9998
rect 16408 9654 16436 11750
rect 16488 11620 16540 11626
rect 16488 11562 16540 11568
rect 16500 11082 16528 11562
rect 16488 11076 16540 11082
rect 16488 11018 16540 11024
rect 16500 10742 16528 11018
rect 16488 10736 16540 10742
rect 16488 10678 16540 10684
rect 16396 9648 16448 9654
rect 16396 9590 16448 9596
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16408 8430 16436 9590
rect 16488 9376 16540 9382
rect 16488 9318 16540 9324
rect 16500 9110 16528 9318
rect 16592 9178 16620 13926
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16684 12782 16712 13806
rect 16776 12986 16804 14198
rect 17040 14068 17092 14074
rect 17040 14010 17092 14016
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 16856 12912 16908 12918
rect 16856 12854 16908 12860
rect 16672 12776 16724 12782
rect 16672 12718 16724 12724
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16684 12209 16712 12582
rect 16670 12200 16726 12209
rect 16670 12135 16726 12144
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16776 11014 16804 11630
rect 16764 11008 16816 11014
rect 16764 10950 16816 10956
rect 16868 10674 16896 12854
rect 17052 12306 17080 14010
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 17052 11898 17080 12242
rect 17040 11892 17092 11898
rect 17040 11834 17092 11840
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16960 10606 16988 10950
rect 16948 10600 17000 10606
rect 16670 10568 16726 10577
rect 16948 10542 17000 10548
rect 16670 10503 16726 10512
rect 16684 9382 16712 10503
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 16764 9172 16816 9178
rect 16764 9114 16816 9120
rect 16488 9104 16540 9110
rect 16488 9046 16540 9052
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16592 8430 16620 8910
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16028 8356 16080 8362
rect 16028 8298 16080 8304
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 16592 7886 16620 8366
rect 16776 8362 16804 9114
rect 16960 8974 16988 9522
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 16960 8498 16988 8910
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 16764 8356 16816 8362
rect 16764 8298 16816 8304
rect 17144 8129 17172 15422
rect 17236 13569 17264 16510
rect 17408 16448 17460 16454
rect 17408 16390 17460 16396
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17328 15026 17356 15846
rect 17420 15706 17448 16390
rect 17512 16046 17540 19178
rect 17776 19168 17828 19174
rect 17776 19110 17828 19116
rect 17592 18080 17644 18086
rect 17592 18022 17644 18028
rect 17604 16250 17632 18022
rect 17788 17066 17816 19110
rect 17972 17882 18000 19774
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 18052 19440 18104 19446
rect 18052 19382 18104 19388
rect 18064 18873 18092 19382
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 18524 18970 18552 19314
rect 18512 18964 18564 18970
rect 18512 18906 18564 18912
rect 18050 18864 18106 18873
rect 18616 18834 18644 19858
rect 18708 19281 18736 19858
rect 18694 19272 18750 19281
rect 18694 19207 18750 19216
rect 18050 18799 18106 18808
rect 18604 18828 18656 18834
rect 18604 18770 18656 18776
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 18524 17796 18552 18702
rect 18694 18320 18750 18329
rect 18694 18255 18750 18264
rect 18524 17768 18644 17796
rect 18420 17740 18472 17746
rect 18472 17700 18552 17728
rect 18420 17682 18472 17688
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 18524 17320 18552 17700
rect 18616 17678 18644 17768
rect 18604 17672 18656 17678
rect 18604 17614 18656 17620
rect 18340 17292 18552 17320
rect 18052 17128 18104 17134
rect 17866 17096 17922 17105
rect 17776 17060 17828 17066
rect 18052 17070 18104 17076
rect 17866 17031 17868 17040
rect 17776 17002 17828 17008
rect 17920 17031 17922 17040
rect 17868 17002 17920 17008
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17958 16960 18014 16969
rect 17696 16697 17724 16934
rect 17958 16895 18014 16904
rect 17972 16810 18000 16895
rect 17880 16782 18000 16810
rect 18064 16794 18092 17070
rect 18052 16788 18104 16794
rect 17682 16688 17738 16697
rect 17682 16623 17738 16632
rect 17682 16552 17738 16561
rect 17682 16487 17738 16496
rect 17592 16244 17644 16250
rect 17592 16186 17644 16192
rect 17696 16114 17724 16487
rect 17684 16108 17736 16114
rect 17684 16050 17736 16056
rect 17500 16040 17552 16046
rect 17500 15982 17552 15988
rect 17408 15700 17460 15706
rect 17408 15642 17460 15648
rect 17880 15638 17908 16782
rect 18052 16730 18104 16736
rect 17960 16652 18012 16658
rect 17960 16594 18012 16600
rect 17972 16114 18000 16594
rect 18340 16572 18368 17292
rect 18708 17082 18736 18255
rect 18800 18086 18828 22320
rect 19168 22250 19196 22320
rect 18984 22222 19196 22250
rect 18880 19304 18932 19310
rect 18880 19246 18932 19252
rect 18788 18080 18840 18086
rect 18788 18022 18840 18028
rect 18786 17912 18842 17921
rect 18786 17847 18788 17856
rect 18840 17847 18842 17856
rect 18788 17818 18840 17824
rect 18788 17672 18840 17678
rect 18788 17614 18840 17620
rect 18800 17218 18828 17614
rect 18892 17338 18920 19246
rect 18984 18630 19012 22222
rect 19154 22128 19210 22137
rect 19154 22063 19210 22072
rect 19062 19816 19118 19825
rect 19062 19751 19064 19760
rect 19116 19751 19118 19760
rect 19064 19722 19116 19728
rect 19062 19408 19118 19417
rect 19062 19343 19064 19352
rect 19116 19343 19118 19352
rect 19064 19314 19116 19320
rect 18972 18624 19024 18630
rect 18972 18566 19024 18572
rect 19064 18148 19116 18154
rect 19064 18090 19116 18096
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 18984 17542 19012 18022
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18970 17368 19026 17377
rect 18880 17332 18932 17338
rect 18970 17303 19026 17312
rect 18880 17274 18932 17280
rect 18800 17190 18920 17218
rect 18708 17054 18828 17082
rect 18420 16992 18472 16998
rect 18420 16934 18472 16940
rect 18432 16640 18460 16934
rect 18432 16612 18736 16640
rect 18340 16544 18552 16572
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 17960 16108 18012 16114
rect 17960 16050 18012 16056
rect 17960 15972 18012 15978
rect 17960 15914 18012 15920
rect 17868 15632 17920 15638
rect 17868 15574 17920 15580
rect 17868 15496 17920 15502
rect 17868 15438 17920 15444
rect 17776 15428 17828 15434
rect 17776 15370 17828 15376
rect 17684 15360 17736 15366
rect 17684 15302 17736 15308
rect 17316 15020 17368 15026
rect 17316 14962 17368 14968
rect 17696 14958 17724 15302
rect 17788 14958 17816 15370
rect 17684 14952 17736 14958
rect 17684 14894 17736 14900
rect 17776 14952 17828 14958
rect 17776 14894 17828 14900
rect 17500 14884 17552 14890
rect 17500 14826 17552 14832
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 17316 14272 17368 14278
rect 17316 14214 17368 14220
rect 17222 13560 17278 13569
rect 17222 13495 17278 13504
rect 17328 12714 17356 14214
rect 17316 12708 17368 12714
rect 17316 12650 17368 12656
rect 17314 11656 17370 11665
rect 17314 11591 17370 11600
rect 17328 11354 17356 11591
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17420 9654 17448 14554
rect 17512 13938 17540 14826
rect 17788 14804 17816 14894
rect 17696 14776 17816 14804
rect 17592 14272 17644 14278
rect 17592 14214 17644 14220
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17500 13184 17552 13190
rect 17500 13126 17552 13132
rect 17512 12850 17540 13126
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17512 12442 17540 12786
rect 17604 12714 17632 14214
rect 17696 13308 17724 14776
rect 17880 14550 17908 15438
rect 17972 15162 18000 15914
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 17960 15156 18012 15162
rect 18524 15144 18552 16544
rect 18604 16448 18656 16454
rect 18604 16390 18656 16396
rect 18616 16046 18644 16390
rect 18604 16040 18656 16046
rect 18604 15982 18656 15988
rect 18616 15434 18644 15982
rect 18708 15706 18736 16612
rect 18696 15700 18748 15706
rect 18696 15642 18748 15648
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 18604 15428 18656 15434
rect 18604 15370 18656 15376
rect 17960 15098 18012 15104
rect 18432 15116 18552 15144
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 18340 14618 18368 14894
rect 18328 14612 18380 14618
rect 18328 14554 18380 14560
rect 17868 14544 17920 14550
rect 17960 14544 18012 14550
rect 17868 14486 17920 14492
rect 17958 14512 17960 14521
rect 18012 14512 18014 14521
rect 17776 14476 17828 14482
rect 17958 14447 18014 14456
rect 17776 14418 17828 14424
rect 17788 14362 17816 14418
rect 18432 14414 18460 15116
rect 18604 14952 18656 14958
rect 18602 14920 18604 14929
rect 18656 14920 18658 14929
rect 18602 14855 18658 14864
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 18510 14648 18566 14657
rect 18616 14618 18644 14758
rect 18510 14583 18566 14592
rect 18604 14612 18656 14618
rect 18420 14408 18472 14414
rect 17788 14334 18000 14362
rect 18420 14350 18472 14356
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17776 13320 17828 13326
rect 17696 13280 17776 13308
rect 17776 13262 17828 13268
rect 17788 12986 17816 13262
rect 17776 12980 17828 12986
rect 17776 12922 17828 12928
rect 17880 12850 17908 13330
rect 17868 12844 17920 12850
rect 17868 12786 17920 12792
rect 17592 12708 17644 12714
rect 17592 12650 17644 12656
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17776 11824 17828 11830
rect 17776 11766 17828 11772
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17512 10674 17540 11086
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17512 10266 17540 10610
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17788 10033 17816 11766
rect 17972 11354 18000 14334
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 18524 14006 18552 14583
rect 18604 14554 18656 14560
rect 18602 14512 18658 14521
rect 18602 14447 18658 14456
rect 18512 14000 18564 14006
rect 18512 13942 18564 13948
rect 18144 13864 18196 13870
rect 18064 13824 18144 13852
rect 18064 13394 18092 13824
rect 18144 13806 18196 13812
rect 18234 13424 18290 13433
rect 18052 13388 18104 13394
rect 18234 13359 18236 13368
rect 18052 13330 18104 13336
rect 18288 13359 18290 13368
rect 18236 13330 18288 13336
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 18512 12368 18564 12374
rect 18512 12310 18564 12316
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 17960 11144 18012 11150
rect 17960 11086 18012 11092
rect 17774 10024 17830 10033
rect 17774 9959 17830 9968
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 17788 9042 17816 9959
rect 17972 9518 18000 11086
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 18524 10470 18552 12310
rect 18616 11801 18644 14447
rect 18708 13870 18736 15438
rect 18696 13864 18748 13870
rect 18696 13806 18748 13812
rect 18800 13734 18828 17054
rect 18892 16454 18920 17190
rect 18984 16726 19012 17303
rect 18972 16720 19024 16726
rect 18972 16662 19024 16668
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18972 16176 19024 16182
rect 18972 16118 19024 16124
rect 18880 15564 18932 15570
rect 18880 15506 18932 15512
rect 18788 13728 18840 13734
rect 18788 13670 18840 13676
rect 18602 11792 18658 11801
rect 18602 11727 18658 11736
rect 18604 11552 18656 11558
rect 18604 11494 18656 11500
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18616 10810 18644 11494
rect 18800 11354 18828 11494
rect 18892 11393 18920 15506
rect 18984 14521 19012 16118
rect 19076 15745 19104 18090
rect 19168 17270 19196 22063
rect 19246 21176 19302 21185
rect 19246 21111 19302 21120
rect 19260 19174 19288 21111
rect 19628 20346 19656 22320
rect 19536 20318 19656 20346
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19260 17814 19288 18226
rect 19248 17808 19300 17814
rect 19352 17785 19380 19790
rect 19444 18222 19472 19858
rect 19432 18216 19484 18222
rect 19432 18158 19484 18164
rect 19536 18170 19564 20318
rect 19614 20224 19670 20233
rect 19614 20159 19670 20168
rect 19628 20058 19656 20159
rect 19616 20052 19668 20058
rect 19616 19994 19668 20000
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 19628 18426 19656 19858
rect 19616 18420 19668 18426
rect 19616 18362 19668 18368
rect 19536 18142 19656 18170
rect 19524 18080 19576 18086
rect 19524 18022 19576 18028
rect 19248 17750 19300 17756
rect 19338 17776 19394 17785
rect 19338 17711 19394 17720
rect 19340 17332 19392 17338
rect 19340 17274 19392 17280
rect 19156 17264 19208 17270
rect 19352 17241 19380 17274
rect 19156 17206 19208 17212
rect 19338 17232 19394 17241
rect 19338 17167 19394 17176
rect 19536 17134 19564 18022
rect 19628 17746 19656 18142
rect 19616 17740 19668 17746
rect 19616 17682 19668 17688
rect 19996 17649 20024 22320
rect 20166 20632 20222 20641
rect 20166 20567 20222 20576
rect 20180 20058 20208 20567
rect 20168 20052 20220 20058
rect 20168 19994 20220 20000
rect 20352 19304 20404 19310
rect 20352 19246 20404 19252
rect 20168 18624 20220 18630
rect 20168 18566 20220 18572
rect 20180 18290 20208 18566
rect 20260 18352 20312 18358
rect 20260 18294 20312 18300
rect 20168 18284 20220 18290
rect 20168 18226 20220 18232
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 19982 17640 20038 17649
rect 19982 17575 20038 17584
rect 19892 17536 19944 17542
rect 19812 17484 19892 17490
rect 19812 17478 19944 17484
rect 19812 17462 19932 17478
rect 19812 17202 19840 17462
rect 19800 17196 19852 17202
rect 19800 17138 19852 17144
rect 19156 17128 19208 17134
rect 19156 17070 19208 17076
rect 19524 17128 19576 17134
rect 19524 17070 19576 17076
rect 19168 16794 19196 17070
rect 19616 16992 19668 16998
rect 19616 16934 19668 16940
rect 19156 16788 19208 16794
rect 19156 16730 19208 16736
rect 19340 16720 19392 16726
rect 19340 16662 19392 16668
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19156 16448 19208 16454
rect 19156 16390 19208 16396
rect 19062 15736 19118 15745
rect 19062 15671 19118 15680
rect 19168 14618 19196 16390
rect 19260 16250 19288 16594
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19260 15502 19288 16186
rect 19248 15496 19300 15502
rect 19248 15438 19300 15444
rect 19352 15178 19380 16662
rect 19628 16130 19656 16934
rect 19628 16102 19748 16130
rect 19616 16040 19668 16046
rect 19616 15982 19668 15988
rect 19432 15972 19484 15978
rect 19432 15914 19484 15920
rect 19260 15162 19380 15178
rect 19444 15162 19472 15914
rect 19524 15632 19576 15638
rect 19524 15574 19576 15580
rect 19248 15156 19380 15162
rect 19300 15150 19380 15156
rect 19432 15156 19484 15162
rect 19248 15098 19300 15104
rect 19432 15098 19484 15104
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19156 14612 19208 14618
rect 19156 14554 19208 14560
rect 18970 14512 19026 14521
rect 18970 14447 19026 14456
rect 19248 14476 19300 14482
rect 19248 14418 19300 14424
rect 18972 14408 19024 14414
rect 18972 14350 19024 14356
rect 18984 13802 19012 14350
rect 18972 13796 19024 13802
rect 18972 13738 19024 13744
rect 19064 13796 19116 13802
rect 19064 13738 19116 13744
rect 18972 13320 19024 13326
rect 18972 13262 19024 13268
rect 18984 12986 19012 13262
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 18972 12640 19024 12646
rect 18970 12608 18972 12617
rect 19024 12608 19026 12617
rect 18970 12543 19026 12552
rect 18972 11756 19024 11762
rect 18972 11698 19024 11704
rect 18878 11384 18934 11393
rect 18788 11348 18840 11354
rect 18878 11319 18934 11328
rect 18788 11290 18840 11296
rect 18984 11150 19012 11698
rect 19076 11286 19104 13738
rect 19156 13388 19208 13394
rect 19156 13330 19208 13336
rect 19168 12918 19196 13330
rect 19156 12912 19208 12918
rect 19156 12854 19208 12860
rect 19260 11898 19288 14418
rect 19352 13025 19380 14758
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19444 13190 19472 13806
rect 19432 13184 19484 13190
rect 19432 13126 19484 13132
rect 19338 13016 19394 13025
rect 19338 12951 19394 12960
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 19352 12238 19380 12854
rect 19444 12850 19472 13126
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19536 12714 19564 15574
rect 19628 13530 19656 15982
rect 19720 15434 19748 16102
rect 19708 15428 19760 15434
rect 19708 15370 19760 15376
rect 19812 15314 19840 17138
rect 20088 17066 20116 18158
rect 20076 17060 20128 17066
rect 20076 17002 20128 17008
rect 20272 16998 20300 18294
rect 20260 16992 20312 16998
rect 20260 16934 20312 16940
rect 19984 16652 20036 16658
rect 19984 16594 20036 16600
rect 19996 15706 20024 16594
rect 19984 15700 20036 15706
rect 19984 15642 20036 15648
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 19720 15286 19840 15314
rect 19616 13524 19668 13530
rect 19616 13466 19668 13472
rect 19616 13388 19668 13394
rect 19616 13330 19668 13336
rect 19524 12708 19576 12714
rect 19524 12650 19576 12656
rect 19628 12442 19656 13330
rect 19616 12436 19668 12442
rect 19616 12378 19668 12384
rect 19616 12300 19668 12306
rect 19616 12242 19668 12248
rect 19340 12232 19392 12238
rect 19340 12174 19392 12180
rect 19248 11892 19300 11898
rect 19248 11834 19300 11840
rect 19628 11626 19656 12242
rect 19524 11620 19576 11626
rect 19524 11562 19576 11568
rect 19616 11620 19668 11626
rect 19616 11562 19668 11568
rect 19064 11280 19116 11286
rect 19064 11222 19116 11228
rect 18972 11144 19024 11150
rect 18972 11086 19024 11092
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18604 10804 18656 10810
rect 18604 10746 18656 10752
rect 18604 10532 18656 10538
rect 18604 10474 18656 10480
rect 18420 10464 18472 10470
rect 18050 10432 18106 10441
rect 18420 10406 18472 10412
rect 18512 10464 18564 10470
rect 18512 10406 18564 10412
rect 18050 10367 18106 10376
rect 18064 10198 18092 10367
rect 18052 10192 18104 10198
rect 18052 10134 18104 10140
rect 18432 10130 18460 10406
rect 18616 10248 18644 10474
rect 18524 10220 18644 10248
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 18524 9897 18552 10220
rect 18602 10160 18658 10169
rect 18602 10095 18658 10104
rect 18510 9888 18566 9897
rect 18116 9820 18412 9840
rect 18510 9823 18566 9832
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 18512 9716 18564 9722
rect 18512 9658 18564 9664
rect 18326 9616 18382 9625
rect 18326 9551 18382 9560
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 18050 9480 18106 9489
rect 18050 9415 18052 9424
rect 18104 9415 18106 9424
rect 18052 9386 18104 9392
rect 18340 9110 18368 9551
rect 18328 9104 18380 9110
rect 18524 9081 18552 9658
rect 18328 9046 18380 9052
rect 18510 9072 18566 9081
rect 17776 9036 17828 9042
rect 18510 9007 18566 9016
rect 17776 8978 17828 8984
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17130 8120 17186 8129
rect 17130 8055 17186 8064
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 16592 6798 16620 7822
rect 17420 7546 17448 8230
rect 17408 7540 17460 7546
rect 17408 7482 17460 7488
rect 16580 6792 16632 6798
rect 16580 6734 16632 6740
rect 16592 6322 16620 6734
rect 16580 6316 16632 6322
rect 16580 6258 16632 6264
rect 12346 6216 12402 6225
rect 12346 6151 12402 6160
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 11704 5296 11756 5302
rect 11704 5238 11756 5244
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 17788 3505 17816 8978
rect 17868 8968 17920 8974
rect 18616 8922 18644 10095
rect 18708 9586 18736 11018
rect 18880 11008 18932 11014
rect 18880 10950 18932 10956
rect 18788 10464 18840 10470
rect 18788 10406 18840 10412
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 18696 9104 18748 9110
rect 18696 9046 18748 9052
rect 17868 8910 17920 8916
rect 17880 8430 17908 8910
rect 18524 8894 18644 8922
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 18144 8356 18196 8362
rect 18144 8298 18196 8304
rect 18156 8090 18184 8298
rect 18236 8288 18288 8294
rect 18236 8230 18288 8236
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17972 7410 18000 7890
rect 18248 7818 18276 8230
rect 18236 7812 18288 7818
rect 18236 7754 18288 7760
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 18524 7585 18552 8894
rect 18510 7576 18566 7585
rect 18510 7511 18566 7520
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 17972 7002 18000 7346
rect 17960 6996 18012 7002
rect 17960 6938 18012 6944
rect 18512 6928 18564 6934
rect 18512 6870 18564 6876
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17972 5817 18000 6598
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 17958 5808 18014 5817
rect 17958 5743 18014 5752
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17972 4865 18000 5306
rect 18524 5273 18552 6870
rect 18510 5264 18566 5273
rect 18510 5199 18566 5208
rect 17958 4856 18014 4865
rect 17958 4791 18014 4800
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 17774 3496 17830 3505
rect 17774 3431 17830 3440
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 11152 2984 11204 2990
rect 11152 2926 11204 2932
rect 15844 2984 15896 2990
rect 15844 2926 15896 2932
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 11164 1442 11192 2926
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11164 1414 11376 1442
rect 11348 480 11376 1414
rect 15856 480 15884 2926
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 18708 649 18736 9046
rect 18800 7954 18828 10406
rect 18892 10266 18920 10950
rect 18880 10260 18932 10266
rect 18880 10202 18932 10208
rect 18880 10124 18932 10130
rect 18880 10066 18932 10072
rect 18892 9466 18920 10066
rect 18984 9586 19012 11086
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 18892 9438 19012 9466
rect 18880 9104 18932 9110
rect 18880 9046 18932 9052
rect 18892 7954 18920 9046
rect 18984 8480 19012 9438
rect 19076 9110 19104 11222
rect 19536 10810 19564 11562
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 19430 10704 19486 10713
rect 19430 10639 19486 10648
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 19064 9104 19116 9110
rect 19064 9046 19116 9052
rect 18984 8452 19104 8480
rect 18788 7948 18840 7954
rect 18788 7890 18840 7896
rect 18880 7948 18932 7954
rect 18880 7890 18932 7896
rect 18800 1057 18828 7890
rect 18786 1048 18842 1057
rect 18786 983 18842 992
rect 18694 640 18750 649
rect 18694 575 18750 584
rect 6828 264 6880 270
rect 6828 206 6880 212
rect 11334 0 11390 480
rect 15842 0 15898 480
rect 18892 241 18920 7890
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 18984 7002 19012 7822
rect 18972 6996 19024 7002
rect 18972 6938 19024 6944
rect 19076 6882 19104 8452
rect 19168 7177 19196 10542
rect 19248 10260 19300 10266
rect 19248 10202 19300 10208
rect 19260 9722 19288 10202
rect 19340 10192 19392 10198
rect 19340 10134 19392 10140
rect 19248 9716 19300 9722
rect 19248 9658 19300 9664
rect 19154 7168 19210 7177
rect 19154 7103 19210 7112
rect 18984 6854 19104 6882
rect 19156 6860 19208 6866
rect 18984 2961 19012 6854
rect 19156 6802 19208 6808
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 19076 6322 19104 6734
rect 19168 6458 19196 6802
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 19064 6316 19116 6322
rect 19064 6258 19116 6264
rect 18970 2952 19026 2961
rect 18970 2887 19026 2896
rect 19260 2553 19288 9658
rect 19352 9654 19380 10134
rect 19444 9654 19472 10639
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 19432 9648 19484 9654
rect 19432 9590 19484 9596
rect 19536 9194 19564 10406
rect 19720 10010 19748 15286
rect 19982 14784 20038 14793
rect 19982 14719 20038 14728
rect 19800 14408 19852 14414
rect 19800 14350 19852 14356
rect 19812 10742 19840 14350
rect 19892 13728 19944 13734
rect 19892 13670 19944 13676
rect 19904 13462 19932 13670
rect 19892 13456 19944 13462
rect 19892 13398 19944 13404
rect 19996 13138 20024 14719
rect 20088 13297 20116 15506
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 20180 15162 20208 15438
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 20180 14074 20208 14350
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 20168 13932 20220 13938
rect 20168 13874 20220 13880
rect 20074 13288 20130 13297
rect 20074 13223 20130 13232
rect 19996 13110 20116 13138
rect 19984 12640 20036 12646
rect 19984 12582 20036 12588
rect 19996 12442 20024 12582
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 19996 11150 20024 11698
rect 20088 11354 20116 13110
rect 20180 12986 20208 13874
rect 20260 13728 20312 13734
rect 20260 13670 20312 13676
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 20168 12844 20220 12850
rect 20168 12786 20220 12792
rect 20180 12238 20208 12786
rect 20272 12782 20300 13670
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 20364 11762 20392 19246
rect 20456 18737 20484 22320
rect 20626 21584 20682 21593
rect 20626 21519 20682 21528
rect 20640 20058 20668 21519
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 20536 19304 20588 19310
rect 20536 19246 20588 19252
rect 20626 19272 20682 19281
rect 20442 18728 20498 18737
rect 20442 18663 20498 18672
rect 20548 18465 20576 19246
rect 20626 19207 20682 19216
rect 20534 18456 20590 18465
rect 20444 18420 20496 18426
rect 20534 18391 20590 18400
rect 20444 18362 20496 18368
rect 20456 14362 20484 18362
rect 20548 18086 20576 18391
rect 20536 18080 20588 18086
rect 20536 18022 20588 18028
rect 20640 15162 20668 19207
rect 20732 19174 20760 22471
rect 20902 22320 20958 22800
rect 21270 22320 21326 22800
rect 21730 22320 21786 22800
rect 22098 22320 22154 22800
rect 22558 22320 22614 22800
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20718 18864 20774 18873
rect 20718 18799 20774 18808
rect 20732 18426 20760 18799
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 20916 18306 20944 22320
rect 20824 18278 20944 18306
rect 20824 18057 20852 18278
rect 21284 18193 21312 22320
rect 21270 18184 21326 18193
rect 20904 18148 20956 18154
rect 21270 18119 21326 18128
rect 20904 18090 20956 18096
rect 20810 18048 20866 18057
rect 20810 17983 20866 17992
rect 20916 17882 20944 18090
rect 20904 17876 20956 17882
rect 20904 17818 20956 17824
rect 21744 17338 21772 22320
rect 22112 19242 22140 22320
rect 22100 19236 22152 19242
rect 22100 19178 22152 19184
rect 22190 19000 22246 19009
rect 22572 18986 22600 22320
rect 22246 18958 22600 18986
rect 22190 18935 22246 18944
rect 21732 17332 21784 17338
rect 21732 17274 21784 17280
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20456 14334 20852 14362
rect 20534 14104 20590 14113
rect 20534 14039 20590 14048
rect 20444 13728 20496 13734
rect 20444 13670 20496 13676
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20168 11620 20220 11626
rect 20168 11562 20220 11568
rect 20076 11348 20128 11354
rect 20076 11290 20128 11296
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 19800 10736 19852 10742
rect 19800 10678 19852 10684
rect 19996 10674 20024 11086
rect 19984 10668 20036 10674
rect 19984 10610 20036 10616
rect 19800 10600 19852 10606
rect 19800 10542 19852 10548
rect 19527 9166 19564 9194
rect 19628 9982 19748 10010
rect 19527 9058 19555 9166
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19432 9036 19484 9042
rect 19527 9030 19564 9058
rect 19432 8978 19484 8984
rect 19352 8634 19380 8978
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19444 8090 19472 8978
rect 19536 8974 19564 9030
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19536 6780 19564 8910
rect 19628 6866 19656 9982
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 19720 8430 19748 9862
rect 19812 9178 19840 10542
rect 20076 10532 20128 10538
rect 20076 10474 20128 10480
rect 20088 9994 20116 10474
rect 20076 9988 20128 9994
rect 20076 9930 20128 9936
rect 19892 9376 19944 9382
rect 19892 9318 19944 9324
rect 19800 9172 19852 9178
rect 19800 9114 19852 9120
rect 19708 8424 19760 8430
rect 19708 8366 19760 8372
rect 19904 8090 19932 9318
rect 19984 8560 20036 8566
rect 19984 8502 20036 8508
rect 19892 8084 19944 8090
rect 19892 8026 19944 8032
rect 19996 7886 20024 8502
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 19904 7546 19932 7822
rect 19892 7540 19944 7546
rect 19892 7482 19944 7488
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 19616 6860 19668 6866
rect 19616 6802 19668 6808
rect 19444 6752 19564 6780
rect 19246 2544 19302 2553
rect 19246 2479 19302 2488
rect 19444 1601 19472 6752
rect 19812 5914 19840 7278
rect 19800 5908 19852 5914
rect 19800 5850 19852 5856
rect 20088 2009 20116 9930
rect 20180 7206 20208 11562
rect 20456 10538 20484 13670
rect 20444 10532 20496 10538
rect 20444 10474 20496 10480
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 20364 9586 20392 9998
rect 20548 9654 20576 14039
rect 20626 13696 20682 13705
rect 20626 13631 20682 13640
rect 20536 9648 20588 9654
rect 20536 9590 20588 9596
rect 20352 9580 20404 9586
rect 20352 9522 20404 9528
rect 20260 9376 20312 9382
rect 20260 9318 20312 9324
rect 20272 9178 20300 9318
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 20260 8968 20312 8974
rect 20260 8910 20312 8916
rect 20272 8634 20300 8910
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 20364 8362 20392 9522
rect 20640 8634 20668 13631
rect 20718 12880 20774 12889
rect 20718 12815 20774 12824
rect 20732 12050 20760 12815
rect 20824 12322 20852 14334
rect 20904 12708 20956 12714
rect 20904 12650 20956 12656
rect 20916 12442 20944 12650
rect 20904 12436 20956 12442
rect 20904 12378 20956 12384
rect 20824 12294 20944 12322
rect 20732 12022 20852 12050
rect 20720 10532 20772 10538
rect 20720 10474 20772 10480
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 20732 8430 20760 10474
rect 20824 8537 20852 12022
rect 20916 11286 20944 12294
rect 20904 11280 20956 11286
rect 20904 11222 20956 11228
rect 20810 8528 20866 8537
rect 20810 8463 20866 8472
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20352 8356 20404 8362
rect 20352 8298 20404 8304
rect 20364 7410 20392 8298
rect 20352 7404 20404 7410
rect 20352 7346 20404 7352
rect 20168 7200 20220 7206
rect 20168 7142 20220 7148
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 20180 5914 20208 6734
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 20168 5908 20220 5914
rect 20168 5850 20220 5856
rect 20364 5710 20392 6394
rect 20260 5704 20312 5710
rect 20260 5646 20312 5652
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 20272 5370 20300 5646
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 20456 3913 20484 7142
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20640 6254 20668 6598
rect 20628 6248 20680 6254
rect 20628 6190 20680 6196
rect 20640 5234 20668 6190
rect 20628 5228 20680 5234
rect 20628 5170 20680 5176
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 20548 4321 20576 4966
rect 20534 4312 20590 4321
rect 20534 4247 20590 4256
rect 20442 3904 20498 3913
rect 20442 3839 20498 3848
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 20074 2000 20130 2009
rect 20074 1935 20130 1944
rect 19430 1592 19486 1601
rect 19430 1527 19486 1536
rect 20456 480 20484 2994
rect 18878 232 18934 241
rect 18878 167 18934 176
rect 20442 0 20498 480
<< via2 >>
rect 3238 22480 3294 22536
rect 1582 19216 1638 19272
rect 1766 19080 1822 19136
rect 1950 19760 2006 19816
rect 1858 18944 1914 19000
rect 1950 18808 2006 18864
rect 1950 17876 2006 17912
rect 1950 17856 1952 17876
rect 1952 17856 2004 17876
rect 2004 17856 2006 17876
rect 1766 17720 1822 17776
rect 1398 15000 1454 15056
rect 1950 16940 1952 16960
rect 1952 16940 2004 16960
rect 2004 16940 2006 16960
rect 1950 16904 2006 16940
rect 1950 16516 2006 16552
rect 1950 16496 1952 16516
rect 1952 16496 2004 16516
rect 2004 16496 2006 16516
rect 1950 15952 2006 16008
rect 1950 15544 2006 15600
rect 1766 14592 1822 14648
rect 1858 13912 1914 13968
rect 2410 16496 2466 16552
rect 3054 22072 3110 22128
rect 2778 21528 2834 21584
rect 2962 20576 3018 20632
rect 3054 18808 3110 18864
rect 20718 22480 20774 22536
rect 3422 20168 3478 20224
rect 3146 18692 3202 18728
rect 3146 18672 3148 18692
rect 3148 18672 3200 18692
rect 3200 18672 3202 18692
rect 2778 18264 2834 18320
rect 2778 17332 2834 17368
rect 2778 17312 2780 17332
rect 2780 17312 2832 17332
rect 2832 17312 2834 17332
rect 2686 17176 2742 17232
rect 3238 18164 3240 18184
rect 3240 18164 3292 18184
rect 3292 18164 3294 18184
rect 3238 18128 3294 18164
rect 2778 14048 2834 14104
rect 2870 13640 2926 13696
rect 2778 12824 2834 12880
rect 2318 9560 2374 9616
rect 3054 16940 3056 16960
rect 3056 16940 3108 16960
rect 3108 16940 3110 16960
rect 3054 16904 3110 16940
rect 2962 13232 3018 13288
rect 3146 13404 3148 13424
rect 3148 13404 3200 13424
rect 3200 13404 3202 13424
rect 3146 13368 3202 13404
rect 3238 12824 3294 12880
rect 3238 9968 3294 10024
rect 3054 4256 3110 4312
rect 3146 2896 3202 2952
rect 3882 21120 3938 21176
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 3790 19252 3792 19272
rect 3792 19252 3844 19272
rect 3844 19252 3846 19272
rect 3790 19216 3846 19252
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 3790 18300 3792 18320
rect 3792 18300 3844 18320
rect 3844 18300 3846 18320
rect 3790 18264 3846 18300
rect 3698 11328 3754 11384
rect 3514 10104 3570 10160
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 4526 16768 4582 16824
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 3790 9424 3846 9480
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4066 12688 4122 12744
rect 4066 12280 4122 12336
rect 4526 12180 4528 12200
rect 4528 12180 4580 12200
rect 4580 12180 4582 12200
rect 3974 11736 4030 11792
rect 4526 12144 4582 12180
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4066 10784 4122 10840
rect 3974 10240 4030 10296
rect 4342 10376 4398 10432
rect 4618 10004 4620 10024
rect 4620 10004 4672 10024
rect 4672 10004 4674 10024
rect 4618 9968 4674 10004
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4066 9016 4122 9072
rect 4066 8472 4122 8528
rect 4066 8064 4122 8120
rect 3882 7520 3938 7576
rect 3330 5752 3386 5808
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 4342 8472 4398 8528
rect 4986 17040 5042 17096
rect 5446 17448 5502 17504
rect 5538 16768 5594 16824
rect 5354 15272 5410 15328
rect 5722 19080 5778 19136
rect 5722 18536 5778 18592
rect 4894 8200 4950 8256
rect 5170 9036 5226 9072
rect 5170 9016 5172 9036
rect 5172 9016 5224 9036
rect 5224 9016 5226 9036
rect 5538 12144 5594 12200
rect 5630 9560 5686 9616
rect 3974 7112 4030 7168
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 3974 6704 4030 6760
rect 4066 6160 4122 6216
rect 4066 5244 4068 5264
rect 4068 5244 4120 5264
rect 4120 5244 4122 5264
rect 4066 5208 4122 5244
rect 4066 4800 4122 4856
rect 3974 3848 4030 3904
rect 3790 3440 3846 3496
rect 3238 2488 3294 2544
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4894 7928 4950 7984
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 4250 1944 4306 2000
rect 2870 1536 2926 1592
rect 5630 8472 5686 8528
rect 6182 12180 6184 12200
rect 6184 12180 6236 12200
rect 6236 12180 6238 12200
rect 6182 12144 6238 12180
rect 5906 10376 5962 10432
rect 5814 10104 5870 10160
rect 5906 9968 5962 10024
rect 6826 18944 6882 19000
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 6366 10240 6422 10296
rect 6182 9016 6238 9072
rect 2962 992 3018 1048
rect 2778 584 2834 640
rect 6918 12824 6974 12880
rect 7470 16904 7526 16960
rect 8022 17176 8078 17232
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 3330 212 3332 232
rect 3332 212 3384 232
rect 3384 212 3386 232
rect 3330 176 3386 212
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 8482 19216 8538 19272
rect 8390 17584 8446 17640
rect 9218 17720 9274 17776
rect 9034 17040 9090 17096
rect 9678 18944 9734 19000
rect 8574 13912 8630 13968
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 7838 12280 7894 12336
rect 8482 12280 8538 12336
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 8758 12824 8814 12880
rect 8022 8472 8078 8528
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 9494 15952 9550 16008
rect 9678 17448 9734 17504
rect 10046 17176 10102 17232
rect 10138 16768 10194 16824
rect 10046 15988 10048 16008
rect 10048 15988 10100 16008
rect 10100 15988 10102 16008
rect 10046 15952 10102 15988
rect 9678 14184 9734 14240
rect 9126 10512 9182 10568
rect 10046 14356 10048 14376
rect 10048 14356 10100 14376
rect 10100 14356 10102 14376
rect 10046 14320 10102 14356
rect 10046 14184 10102 14240
rect 10414 16632 10470 16688
rect 10046 12824 10102 12880
rect 10230 10648 10286 10704
rect 10414 14592 10470 14648
rect 10598 17856 10654 17912
rect 10874 18944 10930 19000
rect 10874 18536 10930 18592
rect 10966 17720 11022 17776
rect 10782 15272 10838 15328
rect 10598 11600 10654 11656
rect 10874 14884 10930 14920
rect 10874 14864 10876 14884
rect 10876 14864 10928 14884
rect 10928 14864 10930 14884
rect 10874 14592 10930 14648
rect 10782 14356 10784 14376
rect 10784 14356 10836 14376
rect 10836 14356 10838 14376
rect 10782 14320 10838 14356
rect 10782 12144 10838 12200
rect 10782 11192 10838 11248
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 11886 19080 11942 19136
rect 11518 16904 11574 16960
rect 11150 16768 11206 16824
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 11150 13932 11206 13968
rect 11150 13912 11152 13932
rect 11152 13912 11204 13932
rect 11204 13912 11206 13932
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 12162 19352 12218 19408
rect 12162 13776 12218 13832
rect 11702 11600 11758 11656
rect 11978 11736 12034 11792
rect 12070 9832 12126 9888
rect 10874 6704 10930 6760
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 12346 19080 12402 19136
rect 12714 19508 12770 19544
rect 12714 19488 12716 19508
rect 12716 19488 12768 19508
rect 12768 19488 12770 19508
rect 12806 17584 12862 17640
rect 12622 17312 12678 17368
rect 12346 17040 12402 17096
rect 12346 16632 12402 16688
rect 12622 13232 12678 13288
rect 12438 12300 12494 12336
rect 12438 12280 12440 12300
rect 12440 12280 12492 12300
rect 12492 12280 12494 12300
rect 13174 19080 13230 19136
rect 13358 18400 13414 18456
rect 13358 17992 13414 18048
rect 12346 8472 12402 8528
rect 13174 13368 13230 13424
rect 14002 18944 14058 19000
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 13726 17720 13782 17776
rect 14186 17212 14188 17232
rect 14188 17212 14240 17232
rect 14240 17212 14242 17232
rect 14186 17176 14242 17212
rect 14186 17040 14242 17096
rect 13542 12688 13598 12744
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 17222 19488 17278 19544
rect 15750 17740 15806 17776
rect 15750 17720 15752 17740
rect 15752 17720 15804 17740
rect 15804 17720 15806 17740
rect 14370 16904 14426 16960
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 14462 15544 14518 15600
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 13082 11056 13138 11112
rect 14094 9968 14150 10024
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 17130 18420 17186 18456
rect 17130 18400 17132 18420
rect 17132 18400 17184 18420
rect 17184 18400 17186 18420
rect 16302 16496 16358 16552
rect 15658 14900 15660 14920
rect 15660 14900 15712 14920
rect 15712 14900 15714 14920
rect 15658 14864 15714 14900
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14554 10104 14610 10160
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 15474 13096 15530 13152
rect 15474 12280 15530 12336
rect 15382 11212 15438 11248
rect 15382 11192 15384 11212
rect 15384 11192 15436 11212
rect 15436 11192 15438 11212
rect 16762 15952 16818 16008
rect 16670 14864 16726 14920
rect 16302 14456 16358 14512
rect 17038 15000 17094 15056
rect 16118 13640 16174 13696
rect 16118 13232 16174 13288
rect 16302 13504 16358 13560
rect 16670 12144 16726 12200
rect 16670 10512 16726 10568
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 18050 18808 18106 18864
rect 18694 19216 18750 19272
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 18694 18264 18750 18320
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 17866 17060 17922 17096
rect 17866 17040 17868 17060
rect 17868 17040 17920 17060
rect 17920 17040 17922 17060
rect 17958 16904 18014 16960
rect 17682 16632 17738 16688
rect 17682 16496 17738 16552
rect 18786 17876 18842 17912
rect 18786 17856 18788 17876
rect 18788 17856 18840 17876
rect 18840 17856 18842 17876
rect 19154 22072 19210 22128
rect 19062 19780 19118 19816
rect 19062 19760 19064 19780
rect 19064 19760 19116 19780
rect 19116 19760 19118 19780
rect 19062 19372 19118 19408
rect 19062 19352 19064 19372
rect 19064 19352 19116 19372
rect 19116 19352 19118 19372
rect 18970 17312 19026 17368
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 17222 13504 17278 13560
rect 17314 11600 17370 11656
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 17958 14492 17960 14512
rect 17960 14492 18012 14512
rect 18012 14492 18014 14512
rect 17958 14456 18014 14492
rect 18602 14900 18604 14920
rect 18604 14900 18656 14920
rect 18656 14900 18658 14920
rect 18602 14864 18658 14900
rect 18510 14592 18566 14648
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18602 14456 18658 14512
rect 18234 13388 18290 13424
rect 18234 13368 18236 13388
rect 18236 13368 18288 13388
rect 18288 13368 18290 13388
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 17774 9968 17830 10024
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18602 11736 18658 11792
rect 19246 21120 19302 21176
rect 19614 20168 19670 20224
rect 19338 17720 19394 17776
rect 19338 17176 19394 17232
rect 20166 20576 20222 20632
rect 19982 17584 20038 17640
rect 19062 15680 19118 15736
rect 18970 14456 19026 14512
rect 18970 12588 18972 12608
rect 18972 12588 19024 12608
rect 19024 12588 19026 12608
rect 18970 12552 19026 12588
rect 18878 11328 18934 11384
rect 19338 12960 19394 13016
rect 18050 10376 18106 10432
rect 18602 10104 18658 10160
rect 18510 9832 18566 9888
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 18326 9560 18382 9616
rect 18050 9444 18106 9480
rect 18050 9424 18052 9444
rect 18052 9424 18104 9444
rect 18104 9424 18106 9444
rect 18510 9016 18566 9072
rect 17130 8064 17186 8120
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 12346 6160 12402 6216
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 18510 7520 18566 7576
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 17958 5752 18014 5808
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 18510 5208 18566 5264
rect 17958 4800 18014 4856
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 17774 3440 17830 3496
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 19430 10648 19486 10704
rect 18786 992 18842 1048
rect 18694 584 18750 640
rect 19154 7112 19210 7168
rect 18970 2896 19026 2952
rect 19982 14728 20038 14784
rect 20074 13232 20130 13288
rect 20626 21528 20682 21584
rect 20442 18672 20498 18728
rect 20626 19216 20682 19272
rect 20534 18400 20590 18456
rect 20718 18808 20774 18864
rect 21270 18128 21326 18184
rect 20810 17992 20866 18048
rect 22190 18944 22246 19000
rect 20534 14048 20590 14104
rect 19246 2488 19302 2544
rect 20626 13640 20682 13696
rect 20718 12824 20774 12880
rect 20810 8472 20866 8528
rect 20534 4256 20590 4312
rect 20442 3848 20498 3904
rect 20074 1944 20130 2000
rect 19430 1536 19486 1592
rect 18878 176 18934 232
<< metal3 >>
rect 0 22538 480 22568
rect 3233 22538 3299 22541
rect 0 22536 3299 22538
rect 0 22480 3238 22536
rect 3294 22480 3299 22536
rect 0 22478 3299 22480
rect 0 22448 480 22478
rect 3233 22475 3299 22478
rect 20713 22538 20779 22541
rect 22320 22538 22800 22568
rect 20713 22536 22800 22538
rect 20713 22480 20718 22536
rect 20774 22480 22800 22536
rect 20713 22478 22800 22480
rect 20713 22475 20779 22478
rect 22320 22448 22800 22478
rect 0 22130 480 22160
rect 3049 22130 3115 22133
rect 0 22128 3115 22130
rect 0 22072 3054 22128
rect 3110 22072 3115 22128
rect 0 22070 3115 22072
rect 0 22040 480 22070
rect 3049 22067 3115 22070
rect 19149 22130 19215 22133
rect 22320 22130 22800 22160
rect 19149 22128 22800 22130
rect 19149 22072 19154 22128
rect 19210 22072 22800 22128
rect 19149 22070 22800 22072
rect 19149 22067 19215 22070
rect 22320 22040 22800 22070
rect 0 21586 480 21616
rect 2773 21586 2839 21589
rect 0 21584 2839 21586
rect 0 21528 2778 21584
rect 2834 21528 2839 21584
rect 0 21526 2839 21528
rect 0 21496 480 21526
rect 2773 21523 2839 21526
rect 20621 21586 20687 21589
rect 22320 21586 22800 21616
rect 20621 21584 22800 21586
rect 20621 21528 20626 21584
rect 20682 21528 22800 21584
rect 20621 21526 22800 21528
rect 20621 21523 20687 21526
rect 22320 21496 22800 21526
rect 0 21178 480 21208
rect 3877 21178 3943 21181
rect 0 21176 3943 21178
rect 0 21120 3882 21176
rect 3938 21120 3943 21176
rect 0 21118 3943 21120
rect 0 21088 480 21118
rect 3877 21115 3943 21118
rect 19241 21178 19307 21181
rect 22320 21178 22800 21208
rect 19241 21176 22800 21178
rect 19241 21120 19246 21176
rect 19302 21120 22800 21176
rect 19241 21118 22800 21120
rect 19241 21115 19307 21118
rect 22320 21088 22800 21118
rect 0 20634 480 20664
rect 2957 20634 3023 20637
rect 0 20632 3023 20634
rect 0 20576 2962 20632
rect 3018 20576 3023 20632
rect 0 20574 3023 20576
rect 0 20544 480 20574
rect 2957 20571 3023 20574
rect 20161 20634 20227 20637
rect 22320 20634 22800 20664
rect 20161 20632 22800 20634
rect 20161 20576 20166 20632
rect 20222 20576 22800 20632
rect 20161 20574 22800 20576
rect 20161 20571 20227 20574
rect 22320 20544 22800 20574
rect 0 20226 480 20256
rect 3417 20226 3483 20229
rect 0 20224 3483 20226
rect 0 20168 3422 20224
rect 3478 20168 3483 20224
rect 0 20166 3483 20168
rect 0 20136 480 20166
rect 3417 20163 3483 20166
rect 19609 20226 19675 20229
rect 22320 20226 22800 20256
rect 19609 20224 22800 20226
rect 19609 20168 19614 20224
rect 19670 20168 22800 20224
rect 19609 20166 22800 20168
rect 19609 20163 19675 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 22320 20136 22800 20166
rect 14672 20095 14992 20096
rect 0 19818 480 19848
rect 1945 19818 2011 19821
rect 0 19816 2011 19818
rect 0 19760 1950 19816
rect 2006 19760 2011 19816
rect 0 19758 2011 19760
rect 0 19728 480 19758
rect 1945 19755 2011 19758
rect 19057 19818 19123 19821
rect 22320 19818 22800 19848
rect 19057 19816 22800 19818
rect 19057 19760 19062 19816
rect 19118 19760 22800 19816
rect 19057 19758 22800 19760
rect 19057 19755 19123 19758
rect 22320 19728 22800 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 12709 19546 12775 19549
rect 17217 19546 17283 19549
rect 12709 19544 17283 19546
rect 12709 19488 12714 19544
rect 12770 19488 17222 19544
rect 17278 19488 17283 19544
rect 12709 19486 17283 19488
rect 12709 19483 12775 19486
rect 17217 19483 17283 19486
rect 12157 19410 12223 19413
rect 19057 19410 19123 19413
rect 12157 19408 19123 19410
rect 12157 19352 12162 19408
rect 12218 19352 19062 19408
rect 19118 19352 19123 19408
rect 12157 19350 19123 19352
rect 12157 19347 12223 19350
rect 19057 19347 19123 19350
rect 0 19274 480 19304
rect 1577 19274 1643 19277
rect 0 19272 1643 19274
rect 0 19216 1582 19272
rect 1638 19216 1643 19272
rect 0 19214 1643 19216
rect 0 19184 480 19214
rect 1577 19211 1643 19214
rect 3785 19274 3851 19277
rect 8477 19274 8543 19277
rect 18689 19274 18755 19277
rect 3785 19272 8543 19274
rect 3785 19216 3790 19272
rect 3846 19216 8482 19272
rect 8538 19216 8543 19272
rect 3785 19214 8543 19216
rect 3785 19211 3851 19214
rect 8477 19211 8543 19214
rect 11884 19272 18755 19274
rect 11884 19216 18694 19272
rect 18750 19216 18755 19272
rect 11884 19214 18755 19216
rect 11884 19141 11944 19214
rect 18689 19211 18755 19214
rect 20621 19274 20687 19277
rect 22320 19274 22800 19304
rect 20621 19272 22800 19274
rect 20621 19216 20626 19272
rect 20682 19216 22800 19272
rect 20621 19214 22800 19216
rect 20621 19211 20687 19214
rect 22320 19184 22800 19214
rect 1761 19138 1827 19141
rect 5717 19138 5783 19141
rect 1761 19136 5783 19138
rect 1761 19080 1766 19136
rect 1822 19080 5722 19136
rect 5778 19080 5783 19136
rect 1761 19078 5783 19080
rect 1761 19075 1827 19078
rect 5717 19075 5783 19078
rect 11881 19136 11947 19141
rect 11881 19080 11886 19136
rect 11942 19080 11947 19136
rect 11881 19075 11947 19080
rect 12341 19138 12407 19141
rect 13169 19138 13235 19141
rect 12341 19136 13235 19138
rect 12341 19080 12346 19136
rect 12402 19080 13174 19136
rect 13230 19080 13235 19136
rect 12341 19078 13235 19080
rect 12341 19075 12407 19078
rect 13169 19075 13235 19078
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 1853 19002 1919 19005
rect 6821 19002 6887 19005
rect 1853 19000 6887 19002
rect 1853 18944 1858 19000
rect 1914 18944 6826 19000
rect 6882 18944 6887 19000
rect 1853 18942 6887 18944
rect 1853 18939 1919 18942
rect 6821 18939 6887 18942
rect 9673 19002 9739 19005
rect 9806 19002 9812 19004
rect 9673 19000 9812 19002
rect 9673 18944 9678 19000
rect 9734 18944 9812 19000
rect 9673 18942 9812 18944
rect 9673 18939 9739 18942
rect 9806 18940 9812 18942
rect 9876 18940 9882 19004
rect 10869 19002 10935 19005
rect 13997 19002 14063 19005
rect 22185 19002 22251 19005
rect 10869 19000 14063 19002
rect 10869 18944 10874 19000
rect 10930 18944 14002 19000
rect 14058 18944 14063 19000
rect 10869 18942 14063 18944
rect 10869 18939 10935 18942
rect 13997 18939 14063 18942
rect 17542 19000 22251 19002
rect 17542 18944 22190 19000
rect 22246 18944 22251 19000
rect 17542 18942 22251 18944
rect 0 18866 480 18896
rect 1945 18866 2011 18869
rect 0 18864 2011 18866
rect 0 18808 1950 18864
rect 2006 18808 2011 18864
rect 0 18806 2011 18808
rect 0 18776 480 18806
rect 1945 18803 2011 18806
rect 3049 18866 3115 18869
rect 17542 18866 17602 18942
rect 22185 18939 22251 18942
rect 3049 18864 17602 18866
rect 3049 18808 3054 18864
rect 3110 18808 17602 18864
rect 3049 18806 17602 18808
rect 18045 18866 18111 18869
rect 18638 18866 18644 18868
rect 18045 18864 18644 18866
rect 18045 18808 18050 18864
rect 18106 18808 18644 18864
rect 18045 18806 18644 18808
rect 3049 18803 3115 18806
rect 18045 18803 18111 18806
rect 18638 18804 18644 18806
rect 18708 18804 18714 18868
rect 20713 18866 20779 18869
rect 22320 18866 22800 18896
rect 20713 18864 22800 18866
rect 20713 18808 20718 18864
rect 20774 18808 22800 18864
rect 20713 18806 22800 18808
rect 20713 18803 20779 18806
rect 22320 18776 22800 18806
rect 3141 18730 3207 18733
rect 20437 18730 20503 18733
rect 3141 18728 20503 18730
rect 3141 18672 3146 18728
rect 3202 18672 20442 18728
rect 20498 18672 20503 18728
rect 3141 18670 20503 18672
rect 3141 18667 3207 18670
rect 20437 18667 20503 18670
rect 5717 18594 5783 18597
rect 10869 18594 10935 18597
rect 5717 18592 10935 18594
rect 5717 18536 5722 18592
rect 5778 18536 10874 18592
rect 10930 18536 10935 18592
rect 5717 18534 10935 18536
rect 5717 18531 5783 18534
rect 10869 18531 10935 18534
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 13353 18458 13419 18461
rect 17125 18458 17191 18461
rect 13353 18456 17191 18458
rect 13353 18400 13358 18456
rect 13414 18400 17130 18456
rect 17186 18400 17191 18456
rect 13353 18398 17191 18400
rect 13353 18395 13419 18398
rect 17125 18395 17191 18398
rect 19374 18396 19380 18460
rect 19444 18458 19450 18460
rect 20529 18458 20595 18461
rect 19444 18456 20595 18458
rect 19444 18400 20534 18456
rect 20590 18400 20595 18456
rect 19444 18398 20595 18400
rect 19444 18396 19450 18398
rect 20529 18395 20595 18398
rect 0 18322 480 18352
rect 2773 18322 2839 18325
rect 0 18320 2839 18322
rect 0 18264 2778 18320
rect 2834 18264 2839 18320
rect 0 18262 2839 18264
rect 0 18232 480 18262
rect 2773 18259 2839 18262
rect 3785 18322 3851 18325
rect 18689 18322 18755 18325
rect 22320 18322 22800 18352
rect 3785 18320 16866 18322
rect 3785 18264 3790 18320
rect 3846 18264 16866 18320
rect 3785 18262 16866 18264
rect 3785 18259 3851 18262
rect 3233 18186 3299 18189
rect 16806 18186 16866 18262
rect 18689 18320 22800 18322
rect 18689 18264 18694 18320
rect 18750 18264 22800 18320
rect 18689 18262 22800 18264
rect 18689 18259 18755 18262
rect 22320 18232 22800 18262
rect 21265 18186 21331 18189
rect 3233 18184 16682 18186
rect 3233 18128 3238 18184
rect 3294 18128 16682 18184
rect 3233 18126 16682 18128
rect 16806 18184 21331 18186
rect 16806 18128 21270 18184
rect 21326 18128 21331 18184
rect 16806 18126 21331 18128
rect 3233 18123 3299 18126
rect 13353 18052 13419 18053
rect 13302 17988 13308 18052
rect 13372 18050 13419 18052
rect 16622 18050 16682 18126
rect 21265 18123 21331 18126
rect 20805 18050 20871 18053
rect 13372 18048 13464 18050
rect 13414 17992 13464 18048
rect 13372 17990 13464 17992
rect 16622 18048 20871 18050
rect 16622 17992 20810 18048
rect 20866 17992 20871 18048
rect 16622 17990 20871 17992
rect 13372 17988 13419 17990
rect 13353 17987 13419 17988
rect 20805 17987 20871 17990
rect 7808 17984 8128 17985
rect 0 17914 480 17944
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 1945 17914 2011 17917
rect 0 17912 2011 17914
rect 0 17856 1950 17912
rect 2006 17856 2011 17912
rect 0 17854 2011 17856
rect 0 17824 480 17854
rect 1945 17851 2011 17854
rect 10593 17914 10659 17917
rect 18781 17914 18847 17917
rect 22320 17914 22800 17944
rect 10593 17912 13922 17914
rect 10593 17856 10598 17912
rect 10654 17856 13922 17912
rect 10593 17854 13922 17856
rect 10593 17851 10659 17854
rect 1761 17778 1827 17781
rect 9213 17778 9279 17781
rect 1761 17776 9279 17778
rect 1761 17720 1766 17776
rect 1822 17720 9218 17776
rect 9274 17720 9279 17776
rect 1761 17718 9279 17720
rect 1761 17715 1827 17718
rect 9213 17715 9279 17718
rect 10961 17778 11027 17781
rect 13721 17778 13787 17781
rect 10961 17776 13787 17778
rect 10961 17720 10966 17776
rect 11022 17720 13726 17776
rect 13782 17720 13787 17776
rect 10961 17718 13787 17720
rect 10961 17715 11027 17718
rect 13721 17715 13787 17718
rect 8385 17642 8451 17645
rect 12801 17642 12867 17645
rect 8385 17640 12867 17642
rect 8385 17584 8390 17640
rect 8446 17584 12806 17640
rect 12862 17584 12867 17640
rect 8385 17582 12867 17584
rect 13862 17642 13922 17854
rect 18781 17912 22800 17914
rect 18781 17856 18786 17912
rect 18842 17856 22800 17912
rect 18781 17854 22800 17856
rect 18781 17851 18847 17854
rect 22320 17824 22800 17854
rect 15745 17778 15811 17781
rect 19006 17778 19012 17780
rect 15745 17776 19012 17778
rect 15745 17720 15750 17776
rect 15806 17720 19012 17776
rect 15745 17718 19012 17720
rect 15745 17715 15811 17718
rect 19006 17716 19012 17718
rect 19076 17778 19082 17780
rect 19333 17778 19399 17781
rect 19076 17776 19399 17778
rect 19076 17720 19338 17776
rect 19394 17720 19399 17776
rect 19076 17718 19399 17720
rect 19076 17716 19082 17718
rect 19333 17715 19399 17718
rect 19977 17642 20043 17645
rect 13862 17640 20043 17642
rect 13862 17584 19982 17640
rect 20038 17584 20043 17640
rect 13862 17582 20043 17584
rect 8385 17579 8451 17582
rect 12801 17579 12867 17582
rect 19977 17579 20043 17582
rect 5441 17506 5507 17509
rect 9673 17506 9739 17509
rect 5441 17504 9739 17506
rect 5441 17448 5446 17504
rect 5502 17448 9678 17504
rect 9734 17448 9739 17504
rect 5441 17446 9739 17448
rect 5441 17443 5507 17446
rect 9673 17443 9739 17446
rect 4376 17440 4696 17441
rect 0 17370 480 17400
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 2773 17370 2839 17373
rect 0 17368 2839 17370
rect 0 17312 2778 17368
rect 2834 17312 2839 17368
rect 0 17310 2839 17312
rect 0 17280 480 17310
rect 2773 17307 2839 17310
rect 12617 17368 12683 17373
rect 12617 17312 12622 17368
rect 12678 17312 12683 17368
rect 12617 17307 12683 17312
rect 18965 17370 19031 17373
rect 22320 17370 22800 17400
rect 18965 17368 22800 17370
rect 18965 17312 18970 17368
rect 19026 17312 22800 17368
rect 18965 17310 22800 17312
rect 18965 17307 19031 17310
rect 2681 17234 2747 17237
rect 8017 17234 8083 17237
rect 2681 17232 8083 17234
rect 2681 17176 2686 17232
rect 2742 17176 8022 17232
rect 8078 17176 8083 17232
rect 2681 17174 8083 17176
rect 2681 17171 2747 17174
rect 8017 17171 8083 17174
rect 10041 17234 10107 17237
rect 12620 17234 12680 17307
rect 22320 17280 22800 17310
rect 10041 17232 12680 17234
rect 10041 17176 10046 17232
rect 10102 17176 12680 17232
rect 10041 17174 12680 17176
rect 14181 17234 14247 17237
rect 19333 17234 19399 17237
rect 14181 17232 19399 17234
rect 14181 17176 14186 17232
rect 14242 17176 19338 17232
rect 19394 17176 19399 17232
rect 14181 17174 19399 17176
rect 10041 17171 10107 17174
rect 14181 17171 14247 17174
rect 19333 17171 19399 17174
rect 4981 17098 5047 17101
rect 9029 17098 9095 17101
rect 12341 17098 12407 17101
rect 14181 17098 14247 17101
rect 17861 17098 17927 17101
rect 4981 17096 12266 17098
rect 4981 17040 4986 17096
rect 5042 17040 9034 17096
rect 9090 17040 12266 17096
rect 4981 17038 12266 17040
rect 4981 17035 5047 17038
rect 9029 17035 9095 17038
rect 0 16962 480 16992
rect 1945 16962 2011 16965
rect 0 16960 2011 16962
rect 0 16904 1950 16960
rect 2006 16904 2011 16960
rect 0 16902 2011 16904
rect 0 16872 480 16902
rect 1945 16899 2011 16902
rect 3049 16962 3115 16965
rect 7465 16962 7531 16965
rect 3049 16960 7531 16962
rect 3049 16904 3054 16960
rect 3110 16904 7470 16960
rect 7526 16904 7531 16960
rect 3049 16902 7531 16904
rect 3049 16899 3115 16902
rect 7465 16899 7531 16902
rect 11513 16962 11579 16965
rect 12014 16962 12020 16964
rect 11513 16960 12020 16962
rect 11513 16904 11518 16960
rect 11574 16904 12020 16960
rect 11513 16902 12020 16904
rect 11513 16899 11579 16902
rect 12014 16900 12020 16902
rect 12084 16900 12090 16964
rect 12206 16962 12266 17038
rect 12341 17096 17927 17098
rect 12341 17040 12346 17096
rect 12402 17040 14186 17096
rect 14242 17040 17866 17096
rect 17922 17040 17927 17096
rect 12341 17038 17927 17040
rect 12341 17035 12407 17038
rect 14181 17035 14247 17038
rect 17861 17035 17927 17038
rect 14365 16962 14431 16965
rect 12206 16960 14431 16962
rect 12206 16904 14370 16960
rect 14426 16904 14431 16960
rect 12206 16902 14431 16904
rect 14365 16899 14431 16902
rect 17953 16962 18019 16965
rect 22320 16962 22800 16992
rect 17953 16960 22800 16962
rect 17953 16904 17958 16960
rect 18014 16904 22800 16960
rect 17953 16902 22800 16904
rect 17953 16899 18019 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 22320 16872 22800 16902
rect 14672 16831 14992 16832
rect 4521 16826 4587 16829
rect 5533 16826 5599 16829
rect 4521 16824 5599 16826
rect 4521 16768 4526 16824
rect 4582 16768 5538 16824
rect 5594 16768 5599 16824
rect 4521 16766 5599 16768
rect 4521 16763 4587 16766
rect 5533 16763 5599 16766
rect 10133 16826 10199 16829
rect 11145 16826 11211 16829
rect 10133 16824 11211 16826
rect 10133 16768 10138 16824
rect 10194 16768 11150 16824
rect 11206 16768 11211 16824
rect 10133 16766 11211 16768
rect 10133 16763 10199 16766
rect 11145 16763 11211 16766
rect 10409 16690 10475 16693
rect 12341 16690 12407 16693
rect 17677 16690 17743 16693
rect 10409 16688 17743 16690
rect 10409 16632 10414 16688
rect 10470 16632 12346 16688
rect 12402 16632 17682 16688
rect 17738 16632 17743 16688
rect 10409 16630 17743 16632
rect 10409 16627 10475 16630
rect 12341 16627 12407 16630
rect 17677 16627 17743 16630
rect 0 16554 480 16584
rect 1945 16554 2011 16557
rect 0 16552 2011 16554
rect 0 16496 1950 16552
rect 2006 16496 2011 16552
rect 0 16494 2011 16496
rect 0 16464 480 16494
rect 1945 16491 2011 16494
rect 2405 16554 2471 16557
rect 16297 16554 16363 16557
rect 2405 16552 16363 16554
rect 2405 16496 2410 16552
rect 2466 16496 16302 16552
rect 16358 16496 16363 16552
rect 2405 16494 16363 16496
rect 2405 16491 2471 16494
rect 16297 16491 16363 16494
rect 17677 16554 17743 16557
rect 22320 16554 22800 16584
rect 17677 16552 22800 16554
rect 17677 16496 17682 16552
rect 17738 16496 22800 16552
rect 17677 16494 22800 16496
rect 17677 16491 17743 16494
rect 22320 16464 22800 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 0 16010 480 16040
rect 1945 16010 2011 16013
rect 0 16008 2011 16010
rect 0 15952 1950 16008
rect 2006 15952 2011 16008
rect 0 15950 2011 15952
rect 0 15920 480 15950
rect 1945 15947 2011 15950
rect 9489 16010 9555 16013
rect 10041 16010 10107 16013
rect 9489 16008 10107 16010
rect 9489 15952 9494 16008
rect 9550 15952 10046 16008
rect 10102 15952 10107 16008
rect 9489 15950 10107 15952
rect 9489 15947 9555 15950
rect 10041 15947 10107 15950
rect 16757 16010 16823 16013
rect 22320 16010 22800 16040
rect 16757 16008 22800 16010
rect 16757 15952 16762 16008
rect 16818 15952 22800 16008
rect 16757 15950 22800 15952
rect 16757 15947 16823 15950
rect 22320 15920 22800 15950
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 19057 15738 19123 15741
rect 19190 15738 19196 15740
rect 19057 15736 19196 15738
rect 19057 15680 19062 15736
rect 19118 15680 19196 15736
rect 19057 15678 19196 15680
rect 19057 15675 19123 15678
rect 19190 15676 19196 15678
rect 19260 15676 19266 15740
rect 0 15602 480 15632
rect 1945 15602 2011 15605
rect 0 15600 2011 15602
rect 0 15544 1950 15600
rect 2006 15544 2011 15600
rect 0 15542 2011 15544
rect 0 15512 480 15542
rect 1945 15539 2011 15542
rect 14457 15602 14523 15605
rect 22320 15602 22800 15632
rect 14457 15600 22800 15602
rect 14457 15544 14462 15600
rect 14518 15544 22800 15600
rect 14457 15542 22800 15544
rect 14457 15539 14523 15542
rect 22320 15512 22800 15542
rect 5349 15330 5415 15333
rect 10777 15330 10843 15333
rect 5349 15328 10843 15330
rect 5349 15272 5354 15328
rect 5410 15272 10782 15328
rect 10838 15272 10843 15328
rect 5349 15270 10843 15272
rect 5349 15267 5415 15270
rect 10777 15267 10843 15270
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 0 15058 480 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 480 14998
rect 1393 14995 1459 14998
rect 17033 15058 17099 15061
rect 22320 15058 22800 15088
rect 17033 15056 22800 15058
rect 17033 15000 17038 15056
rect 17094 15000 22800 15056
rect 17033 14998 22800 15000
rect 17033 14995 17099 14998
rect 22320 14968 22800 14998
rect 10869 14922 10935 14925
rect 15653 14922 15719 14925
rect 10869 14920 15719 14922
rect 10869 14864 10874 14920
rect 10930 14864 15658 14920
rect 15714 14864 15719 14920
rect 10869 14862 15719 14864
rect 10869 14859 10935 14862
rect 15653 14859 15719 14862
rect 16665 14922 16731 14925
rect 18597 14922 18663 14925
rect 16665 14920 18663 14922
rect 16665 14864 16670 14920
rect 16726 14864 18602 14920
rect 18658 14864 18663 14920
rect 16665 14862 18663 14864
rect 16665 14859 16731 14862
rect 18597 14859 18663 14862
rect 15656 14786 15716 14859
rect 19977 14786 20043 14789
rect 15656 14784 20043 14786
rect 15656 14728 19982 14784
rect 20038 14728 20043 14784
rect 15656 14726 20043 14728
rect 19977 14723 20043 14726
rect 7808 14720 8128 14721
rect 0 14650 480 14680
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 1761 14650 1827 14653
rect 0 14648 1827 14650
rect 0 14592 1766 14648
rect 1822 14592 1827 14648
rect 0 14590 1827 14592
rect 0 14560 480 14590
rect 1761 14587 1827 14590
rect 10409 14650 10475 14653
rect 10869 14650 10935 14653
rect 10409 14648 10935 14650
rect 10409 14592 10414 14648
rect 10470 14592 10874 14648
rect 10930 14592 10935 14648
rect 10409 14590 10935 14592
rect 10409 14587 10475 14590
rect 10869 14587 10935 14590
rect 18505 14650 18571 14653
rect 22320 14650 22800 14680
rect 18505 14648 22800 14650
rect 18505 14592 18510 14648
rect 18566 14592 22800 14648
rect 18505 14590 22800 14592
rect 18505 14587 18571 14590
rect 22320 14560 22800 14590
rect 16297 14514 16363 14517
rect 17953 14514 18019 14517
rect 16297 14512 18019 14514
rect 16297 14456 16302 14512
rect 16358 14456 17958 14512
rect 18014 14456 18019 14512
rect 16297 14454 18019 14456
rect 16297 14451 16363 14454
rect 17953 14451 18019 14454
rect 18597 14514 18663 14517
rect 18965 14514 19031 14517
rect 18597 14512 19031 14514
rect 18597 14456 18602 14512
rect 18658 14456 18970 14512
rect 19026 14456 19031 14512
rect 18597 14454 19031 14456
rect 18597 14451 18663 14454
rect 18965 14451 19031 14454
rect 10041 14378 10107 14381
rect 10777 14378 10843 14381
rect 10041 14376 10843 14378
rect 10041 14320 10046 14376
rect 10102 14320 10782 14376
rect 10838 14320 10843 14376
rect 10041 14318 10843 14320
rect 10041 14315 10107 14318
rect 10777 14315 10843 14318
rect 9673 14242 9739 14245
rect 10041 14242 10107 14245
rect 9673 14240 10107 14242
rect 9673 14184 9678 14240
rect 9734 14184 10046 14240
rect 10102 14184 10107 14240
rect 9673 14182 10107 14184
rect 9673 14179 9739 14182
rect 10041 14179 10107 14182
rect 4376 14176 4696 14177
rect 0 14106 480 14136
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 2773 14106 2839 14109
rect 0 14104 2839 14106
rect 0 14048 2778 14104
rect 2834 14048 2839 14104
rect 0 14046 2839 14048
rect 0 14016 480 14046
rect 2773 14043 2839 14046
rect 20529 14106 20595 14109
rect 22320 14106 22800 14136
rect 20529 14104 22800 14106
rect 20529 14048 20534 14104
rect 20590 14048 22800 14104
rect 20529 14046 22800 14048
rect 20529 14043 20595 14046
rect 22320 14016 22800 14046
rect 1853 13970 1919 13973
rect 8569 13970 8635 13973
rect 11145 13970 11211 13973
rect 1853 13968 11211 13970
rect 1853 13912 1858 13968
rect 1914 13912 8574 13968
rect 8630 13912 11150 13968
rect 11206 13912 11211 13968
rect 1853 13910 11211 13912
rect 1853 13907 1919 13910
rect 8569 13907 8635 13910
rect 11145 13907 11211 13910
rect 12157 13834 12223 13837
rect 13302 13834 13308 13836
rect 12157 13832 13308 13834
rect 12157 13776 12162 13832
rect 12218 13776 13308 13832
rect 12157 13774 13308 13776
rect 12157 13771 12223 13774
rect 13302 13772 13308 13774
rect 13372 13772 13378 13836
rect 0 13698 480 13728
rect 2865 13698 2931 13701
rect 0 13696 2931 13698
rect 0 13640 2870 13696
rect 2926 13640 2931 13696
rect 0 13638 2931 13640
rect 0 13608 480 13638
rect 2865 13635 2931 13638
rect 16113 13698 16179 13701
rect 19374 13698 19380 13700
rect 16113 13696 19380 13698
rect 16113 13640 16118 13696
rect 16174 13640 19380 13696
rect 16113 13638 19380 13640
rect 16113 13635 16179 13638
rect 19374 13636 19380 13638
rect 19444 13636 19450 13700
rect 20621 13698 20687 13701
rect 22320 13698 22800 13728
rect 20621 13696 22800 13698
rect 20621 13640 20626 13696
rect 20682 13640 22800 13696
rect 20621 13638 22800 13640
rect 20621 13635 20687 13638
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 22320 13608 22800 13638
rect 14672 13567 14992 13568
rect 16297 13562 16363 13565
rect 17217 13562 17283 13565
rect 16297 13560 17283 13562
rect 16297 13504 16302 13560
rect 16358 13504 17222 13560
rect 17278 13504 17283 13560
rect 16297 13502 17283 13504
rect 16297 13499 16363 13502
rect 17217 13499 17283 13502
rect 3141 13426 3207 13429
rect 13169 13426 13235 13429
rect 18229 13426 18295 13429
rect 3141 13424 12496 13426
rect 3141 13368 3146 13424
rect 3202 13368 12496 13424
rect 3141 13366 12496 13368
rect 3141 13363 3207 13366
rect 0 13290 480 13320
rect 2957 13290 3023 13293
rect 0 13288 3023 13290
rect 0 13232 2962 13288
rect 3018 13232 3023 13288
rect 0 13230 3023 13232
rect 0 13200 480 13230
rect 2957 13227 3023 13230
rect 12436 13154 12496 13366
rect 13169 13424 18295 13426
rect 13169 13368 13174 13424
rect 13230 13368 18234 13424
rect 18290 13368 18295 13424
rect 13169 13366 18295 13368
rect 13169 13363 13235 13366
rect 18229 13363 18295 13366
rect 12617 13290 12683 13293
rect 16113 13290 16179 13293
rect 12617 13288 16179 13290
rect 12617 13232 12622 13288
rect 12678 13232 16118 13288
rect 16174 13232 16179 13288
rect 12617 13230 16179 13232
rect 12617 13227 12683 13230
rect 16113 13227 16179 13230
rect 20069 13290 20135 13293
rect 22320 13290 22800 13320
rect 20069 13288 22800 13290
rect 20069 13232 20074 13288
rect 20130 13232 22800 13288
rect 20069 13230 22800 13232
rect 20069 13227 20135 13230
rect 22320 13200 22800 13230
rect 15469 13154 15535 13157
rect 12436 13152 15535 13154
rect 12436 13096 15474 13152
rect 15530 13096 15535 13152
rect 12436 13094 15535 13096
rect 15469 13091 15535 13094
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 19333 13018 19399 13021
rect 19333 13016 19442 13018
rect 19333 12960 19338 13016
rect 19394 12960 19442 13016
rect 19333 12955 19442 12960
rect 2773 12882 2839 12885
rect 3233 12882 3299 12885
rect 2773 12880 3299 12882
rect 2773 12824 2778 12880
rect 2834 12824 3238 12880
rect 3294 12824 3299 12880
rect 2773 12822 3299 12824
rect 2773 12819 2839 12822
rect 3233 12819 3299 12822
rect 6913 12882 6979 12885
rect 8753 12882 8819 12885
rect 6913 12880 8819 12882
rect 6913 12824 6918 12880
rect 6974 12824 8758 12880
rect 8814 12824 8819 12880
rect 6913 12822 8819 12824
rect 6913 12819 6979 12822
rect 8753 12819 8819 12822
rect 10041 12882 10107 12885
rect 19382 12882 19442 12955
rect 20713 12882 20779 12885
rect 10041 12880 20779 12882
rect 10041 12824 10046 12880
rect 10102 12824 20718 12880
rect 20774 12824 20779 12880
rect 10041 12822 20779 12824
rect 10041 12819 10107 12822
rect 20713 12819 20779 12822
rect 0 12746 480 12776
rect 4061 12746 4127 12749
rect 0 12744 4127 12746
rect 0 12688 4066 12744
rect 4122 12688 4127 12744
rect 0 12686 4127 12688
rect 0 12656 480 12686
rect 4061 12683 4127 12686
rect 13537 12746 13603 12749
rect 19190 12746 19196 12748
rect 13537 12744 19196 12746
rect 13537 12688 13542 12744
rect 13598 12688 19196 12744
rect 13537 12686 19196 12688
rect 13537 12683 13603 12686
rect 19190 12684 19196 12686
rect 19260 12746 19266 12748
rect 22320 12746 22800 12776
rect 19260 12686 22800 12746
rect 19260 12684 19266 12686
rect 22320 12656 22800 12686
rect 18965 12612 19031 12613
rect 18965 12608 19012 12612
rect 19076 12610 19082 12612
rect 18965 12552 18970 12608
rect 18965 12548 19012 12552
rect 19076 12550 19122 12610
rect 19076 12548 19082 12550
rect 18965 12547 19031 12548
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 0 12338 480 12368
rect 4061 12338 4127 12341
rect 0 12336 4127 12338
rect 0 12280 4066 12336
rect 4122 12280 4127 12336
rect 0 12278 4127 12280
rect 0 12248 480 12278
rect 4061 12275 4127 12278
rect 7833 12338 7899 12341
rect 8477 12338 8543 12341
rect 7833 12336 8543 12338
rect 7833 12280 7838 12336
rect 7894 12280 8482 12336
rect 8538 12280 8543 12336
rect 7833 12278 8543 12280
rect 7833 12275 7899 12278
rect 8477 12275 8543 12278
rect 12433 12338 12499 12341
rect 15469 12338 15535 12341
rect 12433 12336 15535 12338
rect 12433 12280 12438 12336
rect 12494 12280 15474 12336
rect 15530 12280 15535 12336
rect 12433 12278 15535 12280
rect 12433 12275 12499 12278
rect 15469 12275 15535 12278
rect 18638 12276 18644 12340
rect 18708 12338 18714 12340
rect 22320 12338 22800 12368
rect 18708 12278 22800 12338
rect 18708 12276 18714 12278
rect 22320 12248 22800 12278
rect 4521 12202 4587 12205
rect 5533 12202 5599 12205
rect 6177 12202 6243 12205
rect 4521 12200 6243 12202
rect 4521 12144 4526 12200
rect 4582 12144 5538 12200
rect 5594 12144 6182 12200
rect 6238 12144 6243 12200
rect 4521 12142 6243 12144
rect 4521 12139 4587 12142
rect 5533 12139 5599 12142
rect 6177 12139 6243 12142
rect 10777 12202 10843 12205
rect 16665 12202 16731 12205
rect 10777 12200 16731 12202
rect 10777 12144 10782 12200
rect 10838 12144 16670 12200
rect 16726 12144 16731 12200
rect 10777 12142 16731 12144
rect 10777 12139 10843 12142
rect 16665 12139 16731 12142
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 0 11794 480 11824
rect 3969 11794 4035 11797
rect 0 11792 4035 11794
rect 0 11736 3974 11792
rect 4030 11736 4035 11792
rect 0 11734 4035 11736
rect 0 11704 480 11734
rect 3969 11731 4035 11734
rect 9806 11732 9812 11796
rect 9876 11794 9882 11796
rect 11973 11794 12039 11797
rect 9876 11792 12039 11794
rect 9876 11736 11978 11792
rect 12034 11736 12039 11792
rect 9876 11734 12039 11736
rect 9876 11732 9882 11734
rect 11973 11731 12039 11734
rect 18597 11794 18663 11797
rect 22320 11794 22800 11824
rect 18597 11792 22800 11794
rect 18597 11736 18602 11792
rect 18658 11736 22800 11792
rect 18597 11734 22800 11736
rect 18597 11731 18663 11734
rect 22320 11704 22800 11734
rect 10593 11658 10659 11661
rect 11697 11658 11763 11661
rect 17309 11658 17375 11661
rect 10593 11656 17375 11658
rect 10593 11600 10598 11656
rect 10654 11600 11702 11656
rect 11758 11600 17314 11656
rect 17370 11600 17375 11656
rect 10593 11598 17375 11600
rect 10593 11595 10659 11598
rect 11697 11595 11763 11598
rect 17309 11595 17375 11598
rect 7808 11456 8128 11457
rect 0 11386 480 11416
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 3693 11386 3759 11389
rect 0 11384 3759 11386
rect 0 11328 3698 11384
rect 3754 11328 3759 11384
rect 0 11326 3759 11328
rect 0 11296 480 11326
rect 3693 11323 3759 11326
rect 18873 11386 18939 11389
rect 22320 11386 22800 11416
rect 18873 11384 22800 11386
rect 18873 11328 18878 11384
rect 18934 11328 22800 11384
rect 18873 11326 22800 11328
rect 18873 11323 18939 11326
rect 22320 11296 22800 11326
rect 10777 11250 10843 11253
rect 15377 11250 15443 11253
rect 10777 11248 15443 11250
rect 10777 11192 10782 11248
rect 10838 11192 15382 11248
rect 15438 11192 15443 11248
rect 10777 11190 15443 11192
rect 10777 11187 10843 11190
rect 15377 11187 15443 11190
rect 13077 11114 13143 11117
rect 13077 11112 18568 11114
rect 13077 11056 13082 11112
rect 13138 11056 18568 11112
rect 13077 11054 18568 11056
rect 13077 11051 13143 11054
rect 4376 10912 4696 10913
rect 0 10842 480 10872
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 4061 10842 4127 10845
rect 0 10840 4127 10842
rect 0 10784 4066 10840
rect 4122 10784 4127 10840
rect 0 10782 4127 10784
rect 18508 10842 18568 11054
rect 22320 10842 22800 10872
rect 18508 10782 22800 10842
rect 0 10752 480 10782
rect 4061 10779 4127 10782
rect 22320 10752 22800 10782
rect 10225 10706 10291 10709
rect 19425 10706 19491 10709
rect 10225 10704 19491 10706
rect 10225 10648 10230 10704
rect 10286 10648 19430 10704
rect 19486 10648 19491 10704
rect 10225 10646 19491 10648
rect 10225 10643 10291 10646
rect 19425 10643 19491 10646
rect 9121 10570 9187 10573
rect 16665 10570 16731 10573
rect 614 10568 16731 10570
rect 614 10512 9126 10568
rect 9182 10512 16670 10568
rect 16726 10512 16731 10568
rect 614 10510 16731 10512
rect 0 10434 480 10464
rect 614 10434 674 10510
rect 9121 10507 9187 10510
rect 16665 10507 16731 10510
rect 0 10374 674 10434
rect 4337 10434 4403 10437
rect 5901 10434 5967 10437
rect 4337 10432 5967 10434
rect 4337 10376 4342 10432
rect 4398 10376 5906 10432
rect 5962 10376 5967 10432
rect 4337 10374 5967 10376
rect 0 10344 480 10374
rect 4337 10371 4403 10374
rect 5901 10371 5967 10374
rect 18045 10434 18111 10437
rect 22320 10434 22800 10464
rect 18045 10432 22800 10434
rect 18045 10376 18050 10432
rect 18106 10376 22800 10432
rect 18045 10374 22800 10376
rect 18045 10371 18111 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 22320 10344 22800 10374
rect 14672 10303 14992 10304
rect 3969 10298 4035 10301
rect 6361 10298 6427 10301
rect 3969 10296 6427 10298
rect 3969 10240 3974 10296
rect 4030 10240 6366 10296
rect 6422 10240 6427 10296
rect 3969 10238 6427 10240
rect 3969 10235 4035 10238
rect 6361 10235 6427 10238
rect 3509 10162 3575 10165
rect 5809 10162 5875 10165
rect 3509 10160 5875 10162
rect 3509 10104 3514 10160
rect 3570 10104 5814 10160
rect 5870 10104 5875 10160
rect 3509 10102 5875 10104
rect 3509 10099 3575 10102
rect 5809 10099 5875 10102
rect 14549 10162 14615 10165
rect 18597 10162 18663 10165
rect 14549 10160 18663 10162
rect 14549 10104 14554 10160
rect 14610 10104 18602 10160
rect 18658 10104 18663 10160
rect 14549 10102 18663 10104
rect 14549 10099 14615 10102
rect 18597 10099 18663 10102
rect 0 10026 480 10056
rect 3233 10026 3299 10029
rect 0 10024 3299 10026
rect 0 9968 3238 10024
rect 3294 9968 3299 10024
rect 0 9966 3299 9968
rect 0 9936 480 9966
rect 3233 9963 3299 9966
rect 4613 10026 4679 10029
rect 5901 10026 5967 10029
rect 4613 10024 5967 10026
rect 4613 9968 4618 10024
rect 4674 9968 5906 10024
rect 5962 9968 5967 10024
rect 4613 9966 5967 9968
rect 4613 9963 4679 9966
rect 5901 9963 5967 9966
rect 14089 10026 14155 10029
rect 17769 10026 17835 10029
rect 22320 10026 22800 10056
rect 14089 10024 17835 10026
rect 14089 9968 14094 10024
rect 14150 9968 17774 10024
rect 17830 9968 17835 10024
rect 14089 9966 17835 9968
rect 14089 9963 14155 9966
rect 17769 9963 17835 9966
rect 17910 9966 22800 10026
rect 12065 9892 12131 9893
rect 12014 9890 12020 9892
rect 11938 9830 12020 9890
rect 12084 9890 12131 9892
rect 17910 9890 17970 9966
rect 22320 9936 22800 9966
rect 12084 9888 17970 9890
rect 12126 9832 17970 9888
rect 12014 9828 12020 9830
rect 12084 9830 17970 9832
rect 18505 9888 18571 9893
rect 18505 9832 18510 9888
rect 18566 9832 18571 9888
rect 12084 9828 12131 9830
rect 12065 9827 12131 9828
rect 18505 9827 18571 9832
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 2313 9618 2379 9621
rect 5625 9618 5691 9621
rect 2313 9616 5691 9618
rect 2313 9560 2318 9616
rect 2374 9560 5630 9616
rect 5686 9560 5691 9616
rect 2313 9558 5691 9560
rect 2313 9555 2379 9558
rect 5625 9555 5691 9558
rect 18321 9618 18387 9621
rect 18508 9618 18568 9827
rect 18321 9616 18568 9618
rect 18321 9560 18326 9616
rect 18382 9560 18568 9616
rect 18321 9558 18568 9560
rect 18321 9555 18387 9558
rect 0 9482 480 9512
rect 3785 9482 3851 9485
rect 0 9480 3851 9482
rect 0 9424 3790 9480
rect 3846 9424 3851 9480
rect 0 9422 3851 9424
rect 0 9392 480 9422
rect 3785 9419 3851 9422
rect 18045 9482 18111 9485
rect 22320 9482 22800 9512
rect 18045 9480 22800 9482
rect 18045 9424 18050 9480
rect 18106 9424 22800 9480
rect 18045 9422 22800 9424
rect 18045 9419 18111 9422
rect 22320 9392 22800 9422
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 0 9074 480 9104
rect 4061 9074 4127 9077
rect 0 9072 4127 9074
rect 0 9016 4066 9072
rect 4122 9016 4127 9072
rect 0 9014 4127 9016
rect 0 8984 480 9014
rect 4061 9011 4127 9014
rect 5165 9074 5231 9077
rect 6177 9074 6243 9077
rect 5165 9072 6243 9074
rect 5165 9016 5170 9072
rect 5226 9016 6182 9072
rect 6238 9016 6243 9072
rect 5165 9014 6243 9016
rect 5165 9011 5231 9014
rect 6177 9011 6243 9014
rect 18505 9074 18571 9077
rect 22320 9074 22800 9104
rect 18505 9072 22800 9074
rect 18505 9016 18510 9072
rect 18566 9016 22800 9072
rect 18505 9014 22800 9016
rect 18505 9011 18571 9014
rect 22320 8984 22800 9014
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 0 8530 480 8560
rect 4061 8530 4127 8533
rect 0 8528 4127 8530
rect 0 8472 4066 8528
rect 4122 8472 4127 8528
rect 0 8470 4127 8472
rect 0 8440 480 8470
rect 4061 8467 4127 8470
rect 4337 8530 4403 8533
rect 5625 8530 5691 8533
rect 4337 8528 5691 8530
rect 4337 8472 4342 8528
rect 4398 8472 5630 8528
rect 5686 8472 5691 8528
rect 4337 8470 5691 8472
rect 4337 8467 4403 8470
rect 5625 8467 5691 8470
rect 8017 8530 8083 8533
rect 12341 8530 12407 8533
rect 8017 8528 12407 8530
rect 8017 8472 8022 8528
rect 8078 8472 12346 8528
rect 12402 8472 12407 8528
rect 8017 8470 12407 8472
rect 8017 8467 8083 8470
rect 12341 8467 12407 8470
rect 20805 8530 20871 8533
rect 22320 8530 22800 8560
rect 20805 8528 22800 8530
rect 20805 8472 20810 8528
rect 20866 8472 22800 8528
rect 20805 8470 22800 8472
rect 20805 8467 20871 8470
rect 22320 8440 22800 8470
rect 4889 8258 4955 8261
rect 4846 8256 4955 8258
rect 4846 8200 4894 8256
rect 4950 8200 4955 8256
rect 4846 8195 4955 8200
rect 0 8122 480 8152
rect 4061 8122 4127 8125
rect 0 8120 4127 8122
rect 0 8064 4066 8120
rect 4122 8064 4127 8120
rect 0 8062 4127 8064
rect 0 8032 480 8062
rect 4061 8059 4127 8062
rect 4846 7989 4906 8195
rect 7808 8192 8128 8193
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 17125 8122 17191 8125
rect 22320 8122 22800 8152
rect 17125 8120 22800 8122
rect 17125 8064 17130 8120
rect 17186 8064 22800 8120
rect 17125 8062 22800 8064
rect 17125 8059 17191 8062
rect 22320 8032 22800 8062
rect 4846 7984 4955 7989
rect 4846 7928 4894 7984
rect 4950 7928 4955 7984
rect 4846 7926 4955 7928
rect 4889 7923 4955 7926
rect 4376 7648 4696 7649
rect 0 7578 480 7608
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 3877 7578 3943 7581
rect 0 7576 3943 7578
rect 0 7520 3882 7576
rect 3938 7520 3943 7576
rect 0 7518 3943 7520
rect 0 7488 480 7518
rect 3877 7515 3943 7518
rect 18505 7578 18571 7581
rect 22320 7578 22800 7608
rect 18505 7576 22800 7578
rect 18505 7520 18510 7576
rect 18566 7520 22800 7576
rect 18505 7518 22800 7520
rect 18505 7515 18571 7518
rect 22320 7488 22800 7518
rect 0 7170 480 7200
rect 3969 7170 4035 7173
rect 0 7168 4035 7170
rect 0 7112 3974 7168
rect 4030 7112 4035 7168
rect 0 7110 4035 7112
rect 0 7080 480 7110
rect 3969 7107 4035 7110
rect 19149 7170 19215 7173
rect 22320 7170 22800 7200
rect 19149 7168 22800 7170
rect 19149 7112 19154 7168
rect 19210 7112 22800 7168
rect 19149 7110 22800 7112
rect 19149 7107 19215 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 22320 7080 22800 7110
rect 14672 7039 14992 7040
rect 0 6762 480 6792
rect 3969 6762 4035 6765
rect 0 6760 4035 6762
rect 0 6704 3974 6760
rect 4030 6704 4035 6760
rect 0 6702 4035 6704
rect 0 6672 480 6702
rect 3969 6699 4035 6702
rect 10869 6762 10935 6765
rect 22320 6762 22800 6792
rect 10869 6760 22800 6762
rect 10869 6704 10874 6760
rect 10930 6704 22800 6760
rect 10869 6702 22800 6704
rect 10869 6699 10935 6702
rect 22320 6672 22800 6702
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 0 6218 480 6248
rect 4061 6218 4127 6221
rect 0 6216 4127 6218
rect 0 6160 4066 6216
rect 4122 6160 4127 6216
rect 0 6158 4127 6160
rect 0 6128 480 6158
rect 4061 6155 4127 6158
rect 12341 6218 12407 6221
rect 22320 6218 22800 6248
rect 12341 6216 22800 6218
rect 12341 6160 12346 6216
rect 12402 6160 22800 6216
rect 12341 6158 22800 6160
rect 12341 6155 12407 6158
rect 22320 6128 22800 6158
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 0 5810 480 5840
rect 3325 5810 3391 5813
rect 0 5808 3391 5810
rect 0 5752 3330 5808
rect 3386 5752 3391 5808
rect 0 5750 3391 5752
rect 0 5720 480 5750
rect 3325 5747 3391 5750
rect 17953 5810 18019 5813
rect 22320 5810 22800 5840
rect 17953 5808 22800 5810
rect 17953 5752 17958 5808
rect 18014 5752 22800 5808
rect 17953 5750 22800 5752
rect 17953 5747 18019 5750
rect 22320 5720 22800 5750
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 0 5266 480 5296
rect 4061 5266 4127 5269
rect 0 5264 4127 5266
rect 0 5208 4066 5264
rect 4122 5208 4127 5264
rect 0 5206 4127 5208
rect 0 5176 480 5206
rect 4061 5203 4127 5206
rect 18505 5266 18571 5269
rect 22320 5266 22800 5296
rect 18505 5264 22800 5266
rect 18505 5208 18510 5264
rect 18566 5208 22800 5264
rect 18505 5206 22800 5208
rect 18505 5203 18571 5206
rect 22320 5176 22800 5206
rect 7808 4928 8128 4929
rect 0 4858 480 4888
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 4061 4858 4127 4861
rect 0 4856 4127 4858
rect 0 4800 4066 4856
rect 4122 4800 4127 4856
rect 0 4798 4127 4800
rect 0 4768 480 4798
rect 4061 4795 4127 4798
rect 17953 4858 18019 4861
rect 22320 4858 22800 4888
rect 17953 4856 22800 4858
rect 17953 4800 17958 4856
rect 18014 4800 22800 4856
rect 17953 4798 22800 4800
rect 17953 4795 18019 4798
rect 22320 4768 22800 4798
rect 4376 4384 4696 4385
rect 0 4314 480 4344
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 3049 4314 3115 4317
rect 0 4312 3115 4314
rect 0 4256 3054 4312
rect 3110 4256 3115 4312
rect 0 4254 3115 4256
rect 0 4224 480 4254
rect 3049 4251 3115 4254
rect 20529 4314 20595 4317
rect 22320 4314 22800 4344
rect 20529 4312 22800 4314
rect 20529 4256 20534 4312
rect 20590 4256 22800 4312
rect 20529 4254 22800 4256
rect 20529 4251 20595 4254
rect 22320 4224 22800 4254
rect 0 3906 480 3936
rect 3969 3906 4035 3909
rect 0 3904 4035 3906
rect 0 3848 3974 3904
rect 4030 3848 4035 3904
rect 0 3846 4035 3848
rect 0 3816 480 3846
rect 3969 3843 4035 3846
rect 20437 3906 20503 3909
rect 22320 3906 22800 3936
rect 20437 3904 22800 3906
rect 20437 3848 20442 3904
rect 20498 3848 22800 3904
rect 20437 3846 22800 3848
rect 20437 3843 20503 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 22320 3816 22800 3846
rect 14672 3775 14992 3776
rect 0 3498 480 3528
rect 3785 3498 3851 3501
rect 0 3496 3851 3498
rect 0 3440 3790 3496
rect 3846 3440 3851 3496
rect 0 3438 3851 3440
rect 0 3408 480 3438
rect 3785 3435 3851 3438
rect 17769 3498 17835 3501
rect 22320 3498 22800 3528
rect 17769 3496 22800 3498
rect 17769 3440 17774 3496
rect 17830 3440 22800 3496
rect 17769 3438 22800 3440
rect 17769 3435 17835 3438
rect 22320 3408 22800 3438
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 0 2954 480 2984
rect 3141 2954 3207 2957
rect 0 2952 3207 2954
rect 0 2896 3146 2952
rect 3202 2896 3207 2952
rect 0 2894 3207 2896
rect 0 2864 480 2894
rect 3141 2891 3207 2894
rect 18965 2954 19031 2957
rect 22320 2954 22800 2984
rect 18965 2952 22800 2954
rect 18965 2896 18970 2952
rect 19026 2896 22800 2952
rect 18965 2894 22800 2896
rect 18965 2891 19031 2894
rect 22320 2864 22800 2894
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 0 2546 480 2576
rect 3233 2546 3299 2549
rect 0 2544 3299 2546
rect 0 2488 3238 2544
rect 3294 2488 3299 2544
rect 0 2486 3299 2488
rect 0 2456 480 2486
rect 3233 2483 3299 2486
rect 19241 2546 19307 2549
rect 22320 2546 22800 2576
rect 19241 2544 22800 2546
rect 19241 2488 19246 2544
rect 19302 2488 22800 2544
rect 19241 2486 22800 2488
rect 19241 2483 19307 2486
rect 22320 2456 22800 2486
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 0 2002 480 2032
rect 4245 2002 4311 2005
rect 0 2000 4311 2002
rect 0 1944 4250 2000
rect 4306 1944 4311 2000
rect 0 1942 4311 1944
rect 0 1912 480 1942
rect 4245 1939 4311 1942
rect 20069 2002 20135 2005
rect 22320 2002 22800 2032
rect 20069 2000 22800 2002
rect 20069 1944 20074 2000
rect 20130 1944 22800 2000
rect 20069 1942 22800 1944
rect 20069 1939 20135 1942
rect 22320 1912 22800 1942
rect 0 1594 480 1624
rect 2865 1594 2931 1597
rect 0 1592 2931 1594
rect 0 1536 2870 1592
rect 2926 1536 2931 1592
rect 0 1534 2931 1536
rect 0 1504 480 1534
rect 2865 1531 2931 1534
rect 19425 1594 19491 1597
rect 22320 1594 22800 1624
rect 19425 1592 22800 1594
rect 19425 1536 19430 1592
rect 19486 1536 22800 1592
rect 19425 1534 22800 1536
rect 19425 1531 19491 1534
rect 22320 1504 22800 1534
rect 0 1050 480 1080
rect 2957 1050 3023 1053
rect 0 1048 3023 1050
rect 0 992 2962 1048
rect 3018 992 3023 1048
rect 0 990 3023 992
rect 0 960 480 990
rect 2957 987 3023 990
rect 18781 1050 18847 1053
rect 22320 1050 22800 1080
rect 18781 1048 22800 1050
rect 18781 992 18786 1048
rect 18842 992 22800 1048
rect 18781 990 22800 992
rect 18781 987 18847 990
rect 22320 960 22800 990
rect 0 642 480 672
rect 2773 642 2839 645
rect 0 640 2839 642
rect 0 584 2778 640
rect 2834 584 2839 640
rect 0 582 2839 584
rect 0 552 480 582
rect 2773 579 2839 582
rect 18689 642 18755 645
rect 22320 642 22800 672
rect 18689 640 22800 642
rect 18689 584 18694 640
rect 18750 584 22800 640
rect 18689 582 22800 584
rect 18689 579 18755 582
rect 22320 552 22800 582
rect 0 234 480 264
rect 3325 234 3391 237
rect 0 232 3391 234
rect 0 176 3330 232
rect 3386 176 3391 232
rect 0 174 3391 176
rect 0 144 480 174
rect 3325 171 3391 174
rect 18873 234 18939 237
rect 22320 234 22800 264
rect 18873 232 22800 234
rect 18873 176 18878 232
rect 18934 176 22800 232
rect 18873 174 22800 176
rect 18873 171 18939 174
rect 22320 144 22800 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 9812 18940 9876 19004
rect 18644 18804 18708 18868
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 19380 18396 19444 18460
rect 13308 18048 13372 18052
rect 13308 17992 13358 18048
rect 13358 17992 13372 18048
rect 13308 17988 13372 17992
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 19012 17716 19076 17780
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 12020 16900 12084 16964
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 19196 15676 19260 15740
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 13308 13772 13372 13836
rect 19380 13636 19444 13700
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 19196 12684 19260 12748
rect 19012 12608 19076 12612
rect 19012 12552 19026 12608
rect 19026 12552 19076 12608
rect 19012 12548 19076 12552
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 18644 12276 18708 12340
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 9812 11732 9876 11796
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 12020 9888 12084 9892
rect 12020 9832 12070 9888
rect 12070 9832 12084 9888
rect 12020 9828 12084 9832
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 9811 19004 9877 19005
rect 9811 18940 9812 19004
rect 9876 18940 9877 19004
rect 9811 18939 9877 18940
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 9814 11797 9874 18939
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 13307 18052 13373 18053
rect 13307 17988 13308 18052
rect 13372 17988 13373 18052
rect 13307 17987 13373 17988
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 12019 16964 12085 16965
rect 12019 16900 12020 16964
rect 12084 16900 12085 16964
rect 12019 16899 12085 16900
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 9811 11796 9877 11797
rect 9811 11732 9812 11796
rect 9876 11732 9877 11796
rect 9811 11731 9877 11732
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 12022 9893 12082 16899
rect 13310 13837 13370 17987
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 13307 13836 13373 13837
rect 13307 13772 13308 13836
rect 13372 13772 13373 13836
rect 13307 13771 13373 13772
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 12019 9892 12085 9893
rect 12019 9828 12020 9892
rect 12084 9828 12085 9892
rect 12019 9827 12085 9828
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18643 18868 18709 18869
rect 18643 18804 18644 18868
rect 18708 18804 18709 18868
rect 18643 18803 18709 18804
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18646 12341 18706 18803
rect 19379 18460 19445 18461
rect 19379 18396 19380 18460
rect 19444 18396 19445 18460
rect 19379 18395 19445 18396
rect 19011 17780 19077 17781
rect 19011 17716 19012 17780
rect 19076 17716 19077 17780
rect 19011 17715 19077 17716
rect 19014 12613 19074 17715
rect 19195 15740 19261 15741
rect 19195 15676 19196 15740
rect 19260 15676 19261 15740
rect 19195 15675 19261 15676
rect 19198 12749 19258 15675
rect 19382 13701 19442 18395
rect 19379 13700 19445 13701
rect 19379 13636 19380 13700
rect 19444 13636 19445 13700
rect 19379 13635 19445 13636
rect 19195 12748 19261 12749
rect 19195 12684 19196 12748
rect 19260 12684 19261 12748
rect 19195 12683 19261 12684
rect 19011 12612 19077 12613
rect 19011 12548 19012 12612
rect 19076 12548 19077 12612
rect 19011 12547 19077 12548
rect 18643 12340 18709 12341
rect 18643 12276 18644 12340
rect 18708 12276 18709 12340
rect 18643 12275 18709 12276
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606821651
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1606821651
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1606821651
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1606821651
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  Test_en_N_FTB01 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 4600 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1606821651
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3588 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_35
timestamp 1606821651
transform 1 0 4324 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_N_FTB01
timestamp 1606821651
transform 1 0 5520 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606821651
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606821651
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1606821651
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_44
timestamp 1606821651
transform 1 0 5152 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_54
timestamp 1606821651
transform 1 0 6072 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 6624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1606821651
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1606821651
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1606821651
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1606821651
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606821651
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1606821651
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1606821651
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1606821651
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1606821651
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606821651
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606821651
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1606821651
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1606821651
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1606821651
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1606821651
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1606821651
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1606821651
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1606821651
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  clk_3_N_FTB01
timestamp 1606821651
transform 1 0 15088 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606821651
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1606821651
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1606821651
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_147
timestamp 1606821651
transform 1 0 14628 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_151
timestamp 1606821651
transform 1 0 14996 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_158
timestamp 1606821651
transform 1 0 15640 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606821651
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606821651
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1606821651
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1606821651
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1606821651
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_170
timestamp 1606821651
transform 1 0 16744 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_182
timestamp 1606821651
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1606821651
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1606821651
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1606821651
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1606821651
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606821651
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606821651
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606821651
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1606821651
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606821651
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1606821651
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1606821651
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606821651
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1606821651
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1606821651
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1606821651
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1606821651
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1606821651
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1606821651
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606821651
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1606821651
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1606821651
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1606821651
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1606821651
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1606821651
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606821651
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1606821651
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1606821651
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1606821651
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1606821651
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1606821651
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606821651
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606821651
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1606821651
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1606821651
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606821651
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1606821651
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1606821651
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1606821651
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1606821651
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606821651
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1606821651
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1606821651
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1606821651
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1606821651
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1606821651
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1606821651
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606821651
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1606821651
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1606821651
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1606821651
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1606821651
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1606821651
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606821651
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1606821651
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1606821651
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1606821651
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1606821651
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606821651
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606821651
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1606821651
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1606821651
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606821651
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1606821651
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1606821651
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1606821651
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1606821651
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1606821651
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1606821651
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606821651
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1606821651
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1606821651
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1606821651
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1606821651
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1606821651
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606821651
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1606821651
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1606821651
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1606821651
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1606821651
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1606821651
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606821651
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606821651
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1606821651
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1606821651
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606821651
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1606821651
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1606821651
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1606821651
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1606821651
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606821651
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1606821651
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1606821651
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1606821651
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1606821651
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1606821651
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1606821651
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606821651
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1606821651
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1606821651
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1606821651
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1606821651
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1606821651
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606821651
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1606821651
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1606821651
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 20056 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 19872 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_196
timestamp 1606821651
transform 1 0 19136 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606821651
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_215
timestamp 1606821651
transform 1 0 20884 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_219
timestamp 1606821651
transform 1 0 21252 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1606821651
transform 1 0 2944 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606821651
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606821651
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1606821651
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1606821651
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1606821651
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_15
timestamp 1606821651
transform 1 0 2484 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_19
timestamp 1606821651
transform 1 0 2852 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606821651
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606821651
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1606821651
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_29
timestamp 1606821651
transform 1 0 3772 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_41
timestamp 1606821651
transform 1 0 4876 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1606821651
transform 1 0 4968 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606821651
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1606821651
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1606821651
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1606821651
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1606821651
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1606821651
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1606821651
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1606821651
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1606821651
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606821651
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1606821651
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1606821651
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1606821651
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606821651
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1606821651
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1606821651
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1606821651
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1606821651
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1606821651
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1606821651
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1606821651
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606821651
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1606821651
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1606821651
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1606821651
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1606821651
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606821651
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1606821651
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1606821651
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1606821651
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 19228 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_38.mux_l2_in_0_
timestamp 1606821651
transform 1 0 19780 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1606821651
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_202
timestamp 1606821651
transform 1 0 19688 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_196
timestamp 1606821651
transform 1 0 19136 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606821651
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606821651
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606821651
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1606821651
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1606821651
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1606821651
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_213
timestamp 1606821651
transform 1 0 20700 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_219
timestamp 1606821651
transform 1 0 21252 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 1564 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606821651
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1606821651
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3312 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1606821651
transform 1 0 4140 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606821651
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_21
timestamp 1606821651
transform 1 0 3036 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606821651
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_32
timestamp 1606821651
transform 1 0 4048 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1606821651
transform 1 0 6164 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1606821651
transform 1 0 5152 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_42
timestamp 1606821651
transform 1 0 4968 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_53
timestamp 1606821651
transform 1 0 5980 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1606821651
transform 1 0 7176 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_64
timestamp 1606821651
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_75
timestamp 1606821651
transform 1 0 8004 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606821651
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_87
timestamp 1606821651
transform 1 0 9108 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1606821651
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1606821651
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1606821651
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1606821651
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1606821651
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1606821651
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606821651
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1606821651
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_166
timestamp 1606821651
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 16560 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_8_184
timestamp 1606821651
transform 1 0 18032 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 19044 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_8_192
timestamp 1606821651
transform 1 0 18768 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1606821651
transform 1 0 20884 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606821651
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606821651
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_211
timestamp 1606821651
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_218
timestamp 1606821651
transform 1 0 21160 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1606821651
transform 1 0 2484 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606821651
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1606821651
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1606821651
transform 1 0 4508 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1606821651
transform 1 0 3496 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_24
timestamp 1606821651
transform 1 0 3312 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_35
timestamp 1606821651
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_40
timestamp 1606821651
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 4968 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606821651
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_58
timestamp 1606821651
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_62
timestamp 1606821651
transform 1 0 6808 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6900 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8556 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_79
timestamp 1606821651
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_90
timestamp 1606821651
transform 1 0 9384 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_102
timestamp 1606821651
transform 1 0 10488 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606821651
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_114
timestamp 1606821651
transform 1 0 11592 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1606821651
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1606821651
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16284 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1606821651
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_159
timestamp 1606821651
transform 1 0 15732 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606821651
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_174
timestamp 1606821651
transform 1 0 17112 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1606821651
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_184
timestamp 1606821651
transform 1 0 18032 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1606821651
transform 1 0 19780 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19044 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_9_192
timestamp 1606821651
transform 1 0 18768 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_201
timestamp 1606821651
transform 1 0 19596 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606821651
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_212
timestamp 1606821651
transform 1 0 20608 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 2300 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606821651
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_3
timestamp 1606821651
transform 1 0 1380 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_11
timestamp 1606821651
transform 1 0 2116 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1606821651
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606821651
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1606821651
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_41
timestamp 1606821651
transform 1 0 4876 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 5704 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_49
timestamp 1606821651
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7820 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_10_66
timestamp 1606821651
transform 1 0 7176 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_72
timestamp 1606821651
transform 1 0 7728 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1606821651
transform 1 0 10396 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606821651
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_89
timestamp 1606821651
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_93
timestamp 1606821651
transform 1 0 9660 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1606821651
transform 1 0 12328 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_110
timestamp 1606821651
transform 1 0 11224 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_131
timestamp 1606821651
transform 1 0 13156 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_143
timestamp 1606821651
transform 1 0 14260 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606821651
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1606821651
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1606821651
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_166
timestamp 1606821651
transform 1 0 16376 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 16744 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_186
timestamp 1606821651
transform 1 0 18216 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1606821651
transform 1 0 18400 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1606821651
transform 1 0 19412 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1606821651
transform 1 0 19228 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_208
timestamp 1606821651
transform 1 0 20240 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606821651
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606821651
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1606821651
transform 1 0 20884 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1606821651
transform 1 0 21252 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 1564 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606821651
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1606821651
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1606821651
transform 1 0 4232 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1606821651
transform 1 0 3220 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_21
timestamp 1606821651
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_32
timestamp 1606821651
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1606821651
transform 1 0 5244 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606821651
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_43
timestamp 1606821651
transform 1 0 5060 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_54
timestamp 1606821651
transform 1 0 6072 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1606821651
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_62
timestamp 1606821651
transform 1 0 6808 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8648 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1606821651
transform 1 0 7636 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_11_70
timestamp 1606821651
transform 1 0 7544 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_80
timestamp 1606821651
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10304 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_98
timestamp 1606821651
transform 1 0 10120 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 12420 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11316 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606821651
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_109
timestamp 1606821651
transform 1 0 11132 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1606821651
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_139
timestamp 1606821651
transform 1 0 13892 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1606821651
transform 1 0 15824 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1606821651
transform 1 0 14812 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_147
timestamp 1606821651
transform 1 0 14628 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_158
timestamp 1606821651
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 18032 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16928 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606821651
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp 1606821651
transform 1 0 16652 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1606821651
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1606821651
transform 1 0 19688 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_200
timestamp 1606821651
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _096_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 20700 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606821651
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_211
timestamp 1606821651
transform 1 0 20516 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_217
timestamp 1606821651
transform 1 0 21068 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1472 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1606821651
transform 1 0 2208 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606821651
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1606821651
transform 1 0 1380 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_10
timestamp 1606821651
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1606821651
transform 1 0 4508 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606821651
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_21
timestamp 1606821651
transform 1 0 3036 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1606821651
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_32
timestamp 1606821651
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_36
timestamp 1606821651
transform 1 0 4416 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1606821651
transform 1 0 5520 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_46
timestamp 1606821651
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_57
timestamp 1606821651
transform 1 0 6348 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1606821651
transform 1 0 7268 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1606821651
transform 1 0 8280 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_65
timestamp 1606821651
transform 1 0 7084 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_76
timestamp 1606821651
transform 1 0 8096 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606821651
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_87
timestamp 1606821651
transform 1 0 9108 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1606821651
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_102
timestamp 1606821651
transform 1 0 10488 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 11868 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10856 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_115
timestamp 1606821651
transform 1 0 11684 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 13524 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_133
timestamp 1606821651
transform 1 0 13340 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1606821651
transform 1 0 16284 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1606821651
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606821651
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1606821651
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_163
timestamp 1606821651
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 18124 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_12_174
timestamp 1606821651
transform 1 0 17112 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_182
timestamp 1606821651
transform 1 0 17848 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1606821651
transform 1 0 19780 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_201
timestamp 1606821651
transform 1 0 19596 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1606821651
transform 1 0 20884 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606821651
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606821651
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1606821651
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_218
timestamp 1606821651
transform 1 0 21160 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_7
timestamp 1606821651
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1606821651
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606821651
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606821651
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1606821651
transform 1 0 1932 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1748 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1606821651
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_18
timestamp 1606821651
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_17
timestamp 1606821651
transform 1 0 2668 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_13
timestamp 1606821651
transform 1 0 2300 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1606821651
transform 1 0 2944 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2760 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1606821651
transform 1 0 4416 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1606821651
transform 1 0 4140 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606821651
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_34
timestamp 1606821651
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1606821651
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_32
timestamp 1606821651
transform 1 0 4048 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_47
timestamp 1606821651
transform 1 0 5428 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_42
timestamp 1606821651
transform 1 0 4968 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_45
timestamp 1606821651
transform 1 0 5244 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_left_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 5152 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1606821651
transform 1 0 5428 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_13_62
timestamp 1606821651
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_60
timestamp 1606821651
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_56
timestamp 1606821651
transform 1 0 6256 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606821651
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 5520 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1606821651
transform 1 0 7268 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7912 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7728 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_13_66
timestamp 1606821651
transform 1 0 7176 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_70
timestamp 1606821651
transform 1 0 7544 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_64
timestamp 1606821651
transform 1 0 6992 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_72
timestamp 1606821651
transform 1 0 7728 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9844 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1606821651
transform 1 0 9660 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606821651
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_88
timestamp 1606821651
transform 1 0 9200 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_94
timestamp 1606821651
transform 1 0 9752 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1606821651
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_102
timestamp 1606821651
transform 1 0 10488 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 11316 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606821651
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_111
timestamp 1606821651
transform 1 0 11316 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_119
timestamp 1606821651
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_110
timestamp 1606821651
transform 1 0 11224 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1606821651
transform 1 0 14352 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1606821651
transform 1 0 13064 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1606821651
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_13_132
timestamp 1606821651
transform 1 0 13248 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_127
timestamp 1606821651
transform 1 0 12788 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_133
timestamp 1606821651
transform 1 0 13340 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_145
timestamp 1606821651
transform 1 0 14444 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 14812 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 16284 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1606821651
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606821651
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_147
timestamp 1606821651
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_165
timestamp 1606821651
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_149
timestamp 1606821651
transform 1 0 14812 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_163
timestamp 1606821651
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1606821651
transform 1 0 16468 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 17940 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1606821651
transform 1 0 18216 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606821651
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_176
timestamp 1606821651
transform 1 0 17296 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1606821651
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_184
timestamp 1606821651
transform 1 0 18032 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_181
timestamp 1606821651
transform 1 0 17756 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1606821651
transform 1 0 19320 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1606821651
transform 1 0 19688 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1606821651
transform 1 0 19872 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1606821651
transform 1 0 18676 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_13_195
timestamp 1606821651
transform 1 0 19044 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_202
timestamp 1606821651
transform 1 0 19688 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_189
timestamp 1606821651
transform 1 0 18492 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_200
timestamp 1606821651
transform 1 0 19504 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606821651
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606821651
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606821651
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_213
timestamp 1606821651
transform 1 0 20700 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_219
timestamp 1606821651
transform 1 0 21252 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_211
timestamp 1606821651
transform 1 0 20516 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1606821651
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1606821651
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1606821651
transform 1 0 2760 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1606821651
transform 1 0 1748 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606821651
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1606821651
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_16
timestamp 1606821651
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1606821651
transform 1 0 3956 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1606821651
transform 1 0 3588 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_40
timestamp 1606821651
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1606821651
transform 1 0 5980 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1606821651
transform 1 0 4968 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606821651
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_51
timestamp 1606821651
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_56
timestamp 1606821651
transform 1 0 6256 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1606821651
transform 1 0 6624 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_62
timestamp 1606821651
transform 1 0 6808 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8740 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1606821651
transform 1 0 7452 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 8464 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_68
timestamp 1606821651
transform 1 0 7360 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_78
timestamp 1606821651
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10672 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_15_92
timestamp 1606821651
transform 1 0 9568 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606821651
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1606821651
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1606821651
transform 1 0 13432 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1606821651
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_143
timestamp 1606821651
transform 1 0 14260 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1606821651
transform 1 0 14904 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16100 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_149
timestamp 1606821651
transform 1 0 14812 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_159
timestamp 1606821651
transform 1 0 15732 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606821651
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_172
timestamp 1606821651
transform 1 0 16928 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_180
timestamp 1606821651
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_184
timestamp 1606821651
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1606821651
transform 1 0 18492 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1606821651
transform 1 0 19504 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_188
timestamp 1606821651
transform 1 0 18400 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_198
timestamp 1606821651
transform 1 0 19320 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 20516 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606821651
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_209
timestamp 1606821651
transform 1 0 20332 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_217
timestamp 1606821651
transform 1 0 21068 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 1472 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606821651
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1606821651
transform 1 0 1380 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_20
timestamp 1606821651
transform 1 0 2944 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1606821651
transform 1 0 3128 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 4048 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606821651
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_25
timestamp 1606821651
transform 1 0 3404 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6716 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1606821651
transform 1 0 5704 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_48
timestamp 1606821651
transform 1 0 5520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_59
timestamp 1606821651
transform 1 0 6532 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8556 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_70
timestamp 1606821651
transform 1 0 7544 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_78
timestamp 1606821651
transform 1 0 8280 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10396 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606821651
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1606821651
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_93
timestamp 1606821651
transform 1 0 9660 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12328 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 12052 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_110
timestamp 1606821651
transform 1 0 11224 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_118
timestamp 1606821651
transform 1 0 11960 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1606821651
transform 1 0 13340 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 14352 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_131
timestamp 1606821651
transform 1 0 13156 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_142
timestamp 1606821651
transform 1 0 14168 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15272 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606821651
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_147
timestamp 1606821651
transform 1 0 14628 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1606821651
transform 1 0 17940 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1606821651
transform 1 0 16928 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1606821651
transform 1 0 16744 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_181
timestamp 1606821651
transform 1 0 17756 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_186
timestamp 1606821651
transform 1 0 18216 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1606821651
transform 1 0 19412 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1606821651
transform 1 0 18400 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1606821651
transform 1 0 19228 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_208
timestamp 1606821651
transform 1 0 20240 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606821651
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606821651
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1606821651
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1606821651
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1606821651
transform 1 0 2760 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1606821651
transform 1 0 1748 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606821651
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1606821651
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_16
timestamp 1606821651
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4784 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1606821651
transform 1 0 3772 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_27
timestamp 1606821651
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_38
timestamp 1606821651
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606821651
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_49
timestamp 1606821651
transform 1 0 5612 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1606821651
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 8280 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1606821651
transform 1 0 7268 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 6992 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_76
timestamp 1606821651
transform 1 0 8096 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10120 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_94
timestamp 1606821651
transform 1 0 9752 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11132 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606821651
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_107
timestamp 1606821651
transform 1 0 10948 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1606821651
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_123
timestamp 1606821651
transform 1 0 12420 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13064 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_17_129
timestamp 1606821651
transform 1 0 12972 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 16100 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1606821651
transform 1 0 14720 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 15732 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_146
timestamp 1606821651
transform 1 0 14536 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_157
timestamp 1606821651
transform 1 0 15548 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_162
timestamp 1606821651
transform 1 0 16008 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1606821651
transform 1 0 18124 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606821651
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_179
timestamp 1606821651
transform 1 0 17572 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_184
timestamp 1606821651
transform 1 0 18032 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1606821651
transform 1 0 19412 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_194
timestamp 1606821651
transform 1 0 18952 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_198
timestamp 1606821651
transform 1 0 19320 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_208
timestamp 1606821651
transform 1 0 20240 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 20424 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606821651
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_216
timestamp 1606821651
transform 1 0 20976 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 1564 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606821651
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1606821651
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 4508 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606821651
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_21
timestamp 1606821651
transform 1 0 3036 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1606821651
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_32
timestamp 1606821651
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_36
timestamp 1606821651
transform 1 0 4416 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6164 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_53
timestamp 1606821651
transform 1 0 5980 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7820 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_71
timestamp 1606821651
transform 1 0 7636 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10212 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606821651
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_89
timestamp 1606821651
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_93
timestamp 1606821651
transform 1 0 9660 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 11224 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_108
timestamp 1606821651
transform 1 0 11040 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 12880 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_126
timestamp 1606821651
transform 1 0 12696 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_144
timestamp 1606821651
transform 1 0 14352 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1606821651
transform 1 0 14720 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1606821651
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606821651
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1606821651
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_163
timestamp 1606821651
transform 1 0 16100 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 16468 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_18_183
timestamp 1606821651
transform 1 0 17940 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1606821651
transform 1 0 18584 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1606821651
transform 1 0 19596 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_189
timestamp 1606821651
transform 1 0 18492 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_199
timestamp 1606821651
transform 1 0 19412 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1606821651
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606821651
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606821651
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_210
timestamp 1606821651
transform 1 0 20424 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_218
timestamp 1606821651
transform 1 0 21160 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_9
timestamp 1606821651
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1606821651
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1606821651
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606821651
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606821651
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1606821651
transform 1 0 1748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1606821651
transform 1 0 1564 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_11
timestamp 1606821651
transform 1 0 2116 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1606821651
transform 1 0 2116 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1606821651
transform 1 0 2300 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2484 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1606821651
transform 1 0 4232 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1606821651
transform 1 0 4692 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1606821651
transform 1 0 4416 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606821651
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_31
timestamp 1606821651
transform 1 0 3956 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_37
timestamp 1606821651
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_22
timestamp 1606821651
transform 1 0 3128 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1606821651
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_32
timestamp 1606821651
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1606821651
transform 1 0 5428 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1606821651
transform 1 0 6440 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1606821651
transform 1 0 5704 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606821651
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_48
timestamp 1606821651
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1606821651
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_62
timestamp 1606821651
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_45
timestamp 1606821651
transform 1 0 5244 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_56
timestamp 1606821651
transform 1 0 6256 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7452 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1606821651
transform 1 0 8188 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1606821651
transform 1 0 7176 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_75
timestamp 1606821651
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_67
timestamp 1606821651
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_93
timestamp 1606821651
transform 1 0 9660 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1606821651
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1606821651
transform 1 0 8924 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_91
timestamp 1606821651
transform 1 0 9476 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_86
timestamp 1606821651
transform 1 0 9016 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 9660 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606821651
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1606821651
transform 1 0 9200 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_100
timestamp 1606821651
transform 1 0 10304 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_96
timestamp 1606821651
transform 1 0 9936 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_left_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 10396 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10028 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 11500 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606821651
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1606821651
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_123
timestamp 1606821651
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 14076 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1606821651
transform 1 0 12972 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13800 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1606821651
transform 1 0 13248 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 12788 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_130
timestamp 1606821651
transform 1 0 13064 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1606821651
transform 1 0 14628 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 16284 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1606821651
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1606821651
transform 1 0 15916 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606821651
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1606821651
transform 1 0 15732 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_157
timestamp 1606821651
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1606821651
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_163
timestamp 1606821651
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 17940 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1606821651
transform 1 0 16928 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 18216 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606821651
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_170
timestamp 1606821651
transform 1 0 16744 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1606821651
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_184
timestamp 1606821651
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_181
timestamp 1606821651
transform 1 0 17756 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1606821651
transform 1 0 19964 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1606821651
transform 1 0 18952 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1606821651
transform 1 0 19596 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_192
timestamp 1606821651
transform 1 0 18768 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_203
timestamp 1606821651
transform 1 0 19780 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_199
timestamp 1606821651
transform 1 0 19412 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606821651
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606821651
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606821651
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_214
timestamp 1606821651
transform 1 0 20792 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_210
timestamp 1606821651
transform 1 0 20424 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1606821651
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1606821651
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2116 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1380 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606821651
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_9
timestamp 1606821651
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_17
timestamp 1606821651
transform 1 0 2668 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 3680 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_21_25
timestamp 1606821651
transform 1 0 3404 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5336 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606821651
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_44
timestamp 1606821651
transform 1 0 5152 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_55
timestamp 1606821651
transform 1 0 6164 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_21_62
timestamp 1606821651
transform 1 0 6808 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7360 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1606821651
transform 1 0 9660 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10488 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1606821651
transform 1 0 8832 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1606821651
transform 1 0 11316 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606821651
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1606821651
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_123
timestamp 1606821651
transform 1 0 12420 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1606821651
transform 1 0 12880 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 13340 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_21_127
timestamp 1606821651
transform 1 0 12788 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_131
timestamp 1606821651
transform 1 0 13156 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1606821651
transform 1 0 16008 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1606821651
transform 1 0 14996 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_149
timestamp 1606821651
transform 1 0 14812 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_160
timestamp 1606821651
transform 1 0 15824 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1606821651
transform 1 0 18032 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 17204 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606821651
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_171
timestamp 1606821651
transform 1 0 16836 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1606821651
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 18584 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1606821651
transform 1 0 20240 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_188
timestamp 1606821651
transform 1 0 18400 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_206
timestamp 1606821651
transform 1 0 20056 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606821651
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_217
timestamp 1606821651
transform 1 0 21068 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1606821651
transform 1 0 1748 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1606821651
transform 1 0 2668 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606821651
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1606821651
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_11
timestamp 1606821651
transform 1 0 2116 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 4416 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606821651
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_26
timestamp 1606821651
transform 1 0 3496 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_30
timestamp 1606821651
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_32
timestamp 1606821651
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6072 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_52
timestamp 1606821651
transform 1 0 5888 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1606821651
transform 1 0 7728 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_70
timestamp 1606821651
transform 1 0 7544 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_81
timestamp 1606821651
transform 1 0 8556 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606821651
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_89
timestamp 1606821651
transform 1 0 9292 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_102
timestamp 1606821651
transform 1 0 10488 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1606821651
transform 1 0 10764 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 12236 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11224 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_108
timestamp 1606821651
transform 1 0 11040 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_119
timestamp 1606821651
transform 1 0 12052 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1606821651
transform 1 0 14168 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 13892 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_137
timestamp 1606821651
transform 1 0 13708 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1606821651
transform 1 0 15364 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1606821651
transform 1 0 15916 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606821651
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1606821651
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_154
timestamp 1606821651
transform 1 0 15272 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_159
timestamp 1606821651
transform 1 0 15732 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 16928 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_170
timestamp 1606821651
transform 1 0 16744 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1606821651
transform 1 0 19596 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1606821651
transform 1 0 18584 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_188
timestamp 1606821651
transform 1 0 18400 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_199
timestamp 1606821651
transform 1 0 19412 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1606821651
transform 1 0 20884 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606821651
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606821651
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_210
timestamp 1606821651
transform 1 0 20424 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_218
timestamp 1606821651
transform 1 0 21160 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 2300 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1564 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606821651
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1606821651
transform 1 0 1380 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_11
timestamp 1606821651
transform 1 0 2116 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4508 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_29
timestamp 1606821651
transform 1 0 3772 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606821651
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_46
timestamp 1606821651
transform 1 0 5336 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_58
timestamp 1606821651
transform 1 0 6440 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8740 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 7820 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_71
timestamp 1606821651
transform 1 0 7636 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_76
timestamp 1606821651
transform 1 0 8096 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_82
timestamp 1606821651
transform 1 0 8648 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1606821651
transform 1 0 10580 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_99
timestamp 1606821651
transform 1 0 10212 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1606821651
transform 1 0 11776 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12604 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606821651
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_112
timestamp 1606821651
transform 1 0 11408 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_120
timestamp 1606821651
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_123
timestamp 1606821651
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1606821651
transform 1 0 14076 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 13616 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_134
timestamp 1606821651
transform 1 0 13432 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_139
timestamp 1606821651
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_145
timestamp 1606821651
transform 1 0 14444 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1606821651
transform 1 0 16192 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1606821651
transform 1 0 15640 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_2_
timestamp 1606821651
transform 1 0 14628 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_156
timestamp 1606821651
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_162
timestamp 1606821651
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 18032 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1606821651
transform 1 0 16744 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606821651
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_168
timestamp 1606821651
transform 1 0 16560 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_179
timestamp 1606821651
transform 1 0 17572 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1606821651
transform 1 0 19688 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_200
timestamp 1606821651
transform 1 0 19504 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1606821651
transform 1 0 20700 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606821651
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_211
timestamp 1606821651
transform 1 0 20516 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_217
timestamp 1606821651
transform 1 0 21068 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1606821651
transform 1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 2484 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606821651
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1606821651
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_11
timestamp 1606821651
transform 1 0 2116 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1606821651
transform 1 0 3496 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1606821651
transform 1 0 4048 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606821651
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_24
timestamp 1606821651
transform 1 0 3312 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1606821651
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_41
timestamp 1606821651
transform 1 0 4876 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1606821651
transform 1 0 5060 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 6072 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_52
timestamp 1606821651
transform 1 0 5888 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_57
timestamp 1606821651
transform 1 0 6348 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1606821651
transform 1 0 6900 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8556 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1606821651
transform 1 0 7360 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_66
timestamp 1606821651
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_77
timestamp 1606821651
transform 1 0 8188 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1606821651
transform 1 0 10304 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606821651
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_90
timestamp 1606821651
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_93
timestamp 1606821651
transform 1 0 9660 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_99
timestamp 1606821651
transform 1 0 10212 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 11316 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_109
timestamp 1606821651
transform 1 0 11132 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12972 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1606821651
transform 1 0 14076 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_127
timestamp 1606821651
transform 1 0 12788 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_138
timestamp 1606821651
transform 1 0 13800 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1606821651
transform 1 0 15456 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 16008 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606821651
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_150
timestamp 1606821651
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1606821651
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_160
timestamp 1606821651
transform 1 0 15824 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1606821651
transform 1 0 17664 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_178
timestamp 1606821651
transform 1 0 17480 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1606821651
transform 1 0 19688 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_1_
timestamp 1606821651
transform 1 0 18676 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_189
timestamp 1606821651
transform 1 0 18492 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_200
timestamp 1606821651
transform 1 0 19504 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606821651
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606821651
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_211
timestamp 1606821651
transform 1 0 20516 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1606821651
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1606821651
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1606821651
transform 1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 2576 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606821651
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1606821651
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_11
timestamp 1606821651
transform 1 0 2116 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_15
timestamp 1606821651
transform 1 0 2484 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1606821651
transform 1 0 4324 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_25_25
timestamp 1606821651
transform 1 0 3404 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_33
timestamp 1606821651
transform 1 0 4140 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1606821651
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606821651
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_44
timestamp 1606821651
transform 1 0 5152 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_56
timestamp 1606821651
transform 1 0 6256 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_60
timestamp 1606821651
transform 1 0 6624 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1606821651
transform 1 0 7820 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_71
timestamp 1606821651
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_82
timestamp 1606821651
transform 1 0 8648 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 9936 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8924 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_94
timestamp 1606821651
transform 1 0 9752 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 12420 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 11592 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606821651
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_112
timestamp 1606821651
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_120
timestamp 1606821651
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 14076 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_139
timestamp 1606821651
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15732 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_157
timestamp 1606821651
transform 1 0 15548 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1606821651
transform 1 0 17388 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 18032 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606821651
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1606821651
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_181
timestamp 1606821651
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 18952 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_190
timestamp 1606821651
transform 1 0 18584 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 20608 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606821651
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_210
timestamp 1606821651
transform 1 0 20424 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_218
timestamp 1606821651
transform 1 0 21160 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1606821651
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1606821651
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606821651
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606821651
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1606821651
transform 1 0 1748 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1606821651
transform 1 0 1748 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_17
timestamp 1606821651
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_11
timestamp 1606821651
transform 1 0 2116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_11
timestamp 1606821651
transform 1 0 2116 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1606821651
transform 1 0 2852 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1606821651
transform 1 0 2300 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 2300 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 4048 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4508 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1606821651
transform 1 0 3496 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606821651
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1606821651
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_23
timestamp 1606821651
transform 1 0 3220 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_35
timestamp 1606821651
transform 1 0 4324 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 6072 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606821651
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_48
timestamp 1606821651
transform 1 0 5520 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_53
timestamp 1606821651
transform 1 0 5980 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7728 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1606821651
transform 1 0 7820 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_70
timestamp 1606821651
transform 1 0 7544 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_71
timestamp 1606821651
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_82
timestamp 1606821651
transform 1 0 8648 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9936 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1606821651
transform 1 0 8924 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1606821651
transform 1 0 10488 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606821651
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_left_track_1.prog_clk
timestamp 1606821651
transform 1 0 9844 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_88
timestamp 1606821651
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1606821651
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_98
timestamp 1606821651
transform 1 0 10120 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_94
timestamp 1606821651
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1606821651
transform 1 0 12420 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_1_
timestamp 1606821651
transform 1 0 11500 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11132 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12512 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606821651
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_111
timestamp 1606821651
transform 1 0 11316 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_122
timestamp 1606821651
transform 1 0 12328 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_105
timestamp 1606821651
transform 1 0 10764 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_118
timestamp 1606821651
transform 1 0 11960 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_126
timestamp 1606821651
transform 1 0 12696 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_133
timestamp 1606821651
transform 1 0 13340 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12880 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_143
timestamp 1606821651
transform 1 0 14260 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_137
timestamp 1606821651
transform 1 0 13708 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_139
timestamp 1606821651
transform 1 0 13892 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1606821651
transform 1 0 14076 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1606821651
transform 1 0 13892 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1606821651
transform 1 0 13616 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 14444 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_27_151
timestamp 1606821651
transform 1 0 14996 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_150
timestamp 1606821651
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606821651
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_3_
timestamp 1606821651
transform 1 0 15272 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1606821651
transform 1 0 15180 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_163
timestamp 1606821651
transform 1 0 16100 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_157
timestamp 1606821651
transform 1 0 15548 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_163
timestamp 1606821651
transform 1 0 16100 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1606821651
transform 1 0 15732 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 16284 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1606821651
transform 1 0 17480 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 18216 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l3_in_0_
timestamp 1606821651
transform 1 0 18032 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16468 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606821651
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_176
timestamp 1606821651
transform 1 0 17296 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_182
timestamp 1606821651
transform 1 0 17848 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1606821651
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19872 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1606821651
transform 1 0 19228 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_202
timestamp 1606821651
transform 1 0 19688 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_193
timestamp 1606821651
transform 1 0 18860 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_206
timestamp 1606821651
transform 1 0 20056 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_210
timestamp 1606821651
transform 1 0 20424 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1606821651
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1606821651
transform 1 0 20516 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_215
timestamp 1606821651
transform 1 0 20884 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_218
timestamp 1606821651
transform 1 0 21160 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606821651
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1606821651
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_219
timestamp 1606821651
transform 1 0 21252 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606821651
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606821651
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1606821651
transform 1 0 2300 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1606821651
transform 1 0 1748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1606821651
transform 1 0 2852 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606821651
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1606821651
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_11
timestamp 1606821651
transform 1 0 2116 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_17
timestamp 1606821651
transform 1 0 2668 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4048 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606821651
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_23
timestamp 1606821651
transform 1 0 3220 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_41
timestamp 1606821651
transform 1 0 4876 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 5520 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_28_47
timestamp 1606821651
transform 1 0 5428 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8556 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1606821651
transform 1 0 7176 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_64
timestamp 1606821651
transform 1 0 6992 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_75
timestamp 1606821651
transform 1 0 8004 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9660 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606821651
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1606821651
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1606821651
transform 1 0 12328 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_1_
timestamp 1606821651
transform 1 0 11316 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_109
timestamp 1606821651
transform 1 0 11132 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_120
timestamp 1606821651
transform 1 0 12144 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_125
timestamp 1606821651
transform 1 0 12604 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1606821651
transform 1 0 13892 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 14444 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1606821651
transform 1 0 12788 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_28_136
timestamp 1606821651
transform 1 0 13616 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_143
timestamp 1606821651
transform 1 0 14260 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1606821651
transform 1 0 16376 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_1_
timestamp 1606821651
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606821651
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_151
timestamp 1606821651
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_163
timestamp 1606821651
transform 1 0 16100 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1606821651
transform 1 0 17664 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 16928 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_170
timestamp 1606821651
transform 1 0 16744 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_178
timestamp 1606821651
transform 1 0 17480 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_184
timestamp 1606821651
transform 1 0 18032 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1606821651
transform 1 0 18400 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 18952 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_192
timestamp 1606821651
transform 1 0 18768 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1606821651
transform 1 0 20884 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606821651
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606821651
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_210
timestamp 1606821651
transform 1 0 20424 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_218
timestamp 1606821651
transform 1 0 21160 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1606821651
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2300 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606821651
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1606821651
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_11
timestamp 1606821651
transform 1 0 2116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_19
timestamp 1606821651
transform 1 0 2852 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1606821651
transform 1 0 3588 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1606821651
transform 1 0 3036 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 4508 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_25
timestamp 1606821651
transform 1 0 3404 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_31
timestamp 1606821651
transform 1 0 3956 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606821651
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_43
timestamp 1606821651
transform 1 0 5060 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_55
timestamp 1606821651
transform 1 0 6164 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_62
timestamp 1606821651
transform 1 0 6808 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1606821651
transform 1 0 8188 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1606821651
transform 1 0 6900 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_72
timestamp 1606821651
transform 1 0 7728 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_76
timestamp 1606821651
transform 1 0 8096 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10028 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 9200 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_86
timestamp 1606821651
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_94
timestamp 1606821651
transform 1 0 9752 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1606821651
transform 1 0 11868 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1606821651
transform 1 0 12420 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606821651
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1606821651
transform 1 0 11500 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1606821651
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 14260 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_1_
timestamp 1606821651
transform 1 0 12880 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_126
timestamp 1606821651
transform 1 0 12696 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_137
timestamp 1606821651
transform 1 0 13708 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1606821651
transform 1 0 15916 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_159
timestamp 1606821651
transform 1 0 15732 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1606821651
transform 1 0 18032 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_1_
timestamp 1606821651
transform 1 0 16928 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606821651
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_170
timestamp 1606821651
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1606821651
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_187
timestamp 1606821651
transform 1 0 18308 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1606821651
transform 1 0 18492 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1606821651
transform 1 0 19504 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_198
timestamp 1606821651
transform 1 0 19320 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1606821651
transform 1 0 20516 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606821651
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_209
timestamp 1606821651
transform 1 0 20332 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_215
timestamp 1606821651
transform 1 0 20884 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_219
timestamp 1606821651
transform 1 0 21252 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1606821651
transform 1 0 2392 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1606821651
transform 1 0 1840 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1606821651
transform 1 0 2944 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606821651
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1606821651
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_7
timestamp 1606821651
transform 1 0 1748 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_12
timestamp 1606821651
transform 1 0 2208 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_18
timestamp 1606821651
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606821651
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_24
timestamp 1606821651
transform 1 0 3312 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_30
timestamp 1606821651
transform 1 0 3864 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1606821651
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1606821651
transform 1 0 5336 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 6256 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_44
timestamp 1606821651
transform 1 0 5152 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_50
timestamp 1606821651
transform 1 0 5704 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_62
timestamp 1606821651
transform 1 0 6808 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 7728 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 6992 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_70
timestamp 1606821651
transform 1 0 7544 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9660 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606821651
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_88
timestamp 1606821651
transform 1 0 9200 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 11408 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12144 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_30_109
timestamp 1606821651
transform 1 0 11132 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_118
timestamp 1606821651
transform 1 0 11960 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13156 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_129
timestamp 1606821651
transform 1 0 12972 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15456 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606821651
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_147
timestamp 1606821651
transform 1 0 14628 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_154
timestamp 1606821651
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 17112 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_172
timestamp 1606821651
transform 1 0 16928 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 18768 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_190
timestamp 1606821651
transform 1 0 18584 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_208
timestamp 1606821651
transform 1 0 20240 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606821651
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606821651
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1606821651
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1606821651
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1606821651
transform 1 0 2300 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1606821651
transform 1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606821651
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1606821651
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1606821651
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_17
timestamp 1606821651
transform 1 0 2668 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1606821651
transform 1 0 3220 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3772 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_27
timestamp 1606821651
transform 1 0 3588 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_41
timestamp 1606821651
transform 1 0 4876 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1606821651
transform 1 0 5888 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606821651
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_49
timestamp 1606821651
transform 1 0 5612 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_56
timestamp 1606821651
transform 1 0 6256 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_60
timestamp 1606821651
transform 1 0 6624 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_62
timestamp 1606821651
transform 1 0 6808 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7084 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8740 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_81
timestamp 1606821651
transform 1 0 8556 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10304 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_31_92
timestamp 1606821651
transform 1 0 9568 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 12420 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606821651
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_116
timestamp 1606821651
transform 1 0 11776 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 14076 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1606821651
transform 1 0 13892 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1606821651
transform 1 0 14812 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 15824 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_147
timestamp 1606821651
transform 1 0 14628 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_158
timestamp 1606821651
transform 1 0 15640 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_166
timestamp 1606821651
transform 1 0 16376 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16928 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 18032 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606821651
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1606821651
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1606821651
transform 1 0 19964 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 18860 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_31_190
timestamp 1606821651
transform 1 0 18584 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_199
timestamp 1606821651
transform 1 0 19412 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1606821651
transform 1 0 20516 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606821651
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_209
timestamp 1606821651
transform 1 0 20332 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1606821651
transform 1 0 20884 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_219
timestamp 1606821651
transform 1 0 21252 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1606821651
transform 1 0 2852 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1606821651
transform 1 0 2300 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1606821651
transform 1 0 1748 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606821651
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1606821651
transform 1 0 1380 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_11
timestamp 1606821651
transform 1 0 2116 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_17
timestamp 1606821651
transform 1 0 2668 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606821651
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_23
timestamp 1606821651
transform 1 0 3220 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1606821651
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606821651
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1606821651
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1606821651
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1606821651
transform 1 0 7636 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8188 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_32_63
timestamp 1606821651
transform 1 0 6900 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_75
timestamp 1606821651
transform 1 0 8004 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1606821651
transform 1 0 9200 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9844 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606821651
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_86
timestamp 1606821651
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_91
timestamp 1606821651
transform 1 0 9476 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_94
timestamp 1606821651
transform 1 0 9752 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_104
timestamp 1606821651
transform 1 0 10672 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1606821651
transform 1 0 11960 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10948 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606821651
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_116
timestamp 1606821651
transform 1 0 11776 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_122
timestamp 1606821651
transform 1 0 12328 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_125
timestamp 1606821651
transform 1 0 12604 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1606821651
transform 1 0 14260 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12880 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_32_137
timestamp 1606821651
transform 1 0 13708 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1606821651
transform 1 0 14812 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1606821651
transform 1 0 15824 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606821651
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_147
timestamp 1606821651
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_153
timestamp 1606821651
transform 1 0 15180 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_156
timestamp 1606821651
transform 1 0 15456 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_164
timestamp 1606821651
transform 1 0 16192 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1606821651
transform 1 0 18308 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16836 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606821651
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_170
timestamp 1606821651
transform 1 0 16744 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_180
timestamp 1606821651
transform 1 0 17664 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1606821651
transform 1 0 19964 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1606821651
transform 1 0 19412 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1606821651
transform 1 0 18860 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_191
timestamp 1606821651
transform 1 0 18676 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1606821651
transform 1 0 19228 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_203
timestamp 1606821651
transform 1 0 19780 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1606821651
transform 1 0 20516 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606821651
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606821651
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1606821651
transform 1 0 20332 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1606821651
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1606821651
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 202 22320 258 22800 6 SC_IN_TOP
port 0 nsew default input
rlabel metal2 s 22558 22320 22614 22800 6 SC_OUT_TOP
port 1 nsew default tristate
rlabel metal2 s 4342 22320 4398 22800 6 Test_en_N_out
port 2 nsew default tristate
rlabel metal2 s 20442 0 20498 480 6 Test_en_S_in
port 3 nsew default input
rlabel metal2 s 2226 0 2282 480 6 ccff_head
port 4 nsew default input
rlabel metal2 s 6734 0 6790 480 6 ccff_tail
port 5 nsew default tristate
rlabel metal3 s 0 4224 480 4344 6 chanx_left_in[0]
port 6 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[10]
port 7 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[11]
port 8 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[12]
port 9 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[13]
port 10 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[14]
port 11 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[15]
port 12 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[16]
port 13 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[17]
port 14 nsew default input
rlabel metal3 s 0 12656 480 12776 6 chanx_left_in[18]
port 15 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chanx_left_in[19]
port 16 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[1]
port 17 nsew default input
rlabel metal3 s 0 5176 480 5296 6 chanx_left_in[2]
port 18 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[3]
port 19 nsew default input
rlabel metal3 s 0 6128 480 6248 6 chanx_left_in[4]
port 20 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[5]
port 21 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[6]
port 22 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[7]
port 23 nsew default input
rlabel metal3 s 0 8032 480 8152 6 chanx_left_in[8]
port 24 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[9]
port 25 nsew default input
rlabel metal3 s 0 13608 480 13728 6 chanx_left_out[0]
port 26 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chanx_left_out[10]
port 27 nsew default tristate
rlabel metal3 s 0 18776 480 18896 6 chanx_left_out[11]
port 28 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chanx_left_out[12]
port 29 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_left_out[13]
port 30 nsew default tristate
rlabel metal3 s 0 20136 480 20256 6 chanx_left_out[14]
port 31 nsew default tristate
rlabel metal3 s 0 20544 480 20664 6 chanx_left_out[15]
port 32 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[16]
port 33 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[17]
port 34 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[18]
port 35 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[19]
port 36 nsew default tristate
rlabel metal3 s 0 14016 480 14136 6 chanx_left_out[1]
port 37 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[2]
port 38 nsew default tristate
rlabel metal3 s 0 14968 480 15088 6 chanx_left_out[3]
port 39 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[4]
port 40 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[5]
port 41 nsew default tristate
rlabel metal3 s 0 16464 480 16584 6 chanx_left_out[6]
port 42 nsew default tristate
rlabel metal3 s 0 16872 480 16992 6 chanx_left_out[7]
port 43 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[8]
port 44 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[9]
port 45 nsew default tristate
rlabel metal3 s 22320 4224 22800 4344 6 chanx_right_in[0]
port 46 nsew default input
rlabel metal3 s 22320 8984 22800 9104 6 chanx_right_in[10]
port 47 nsew default input
rlabel metal3 s 22320 9392 22800 9512 6 chanx_right_in[11]
port 48 nsew default input
rlabel metal3 s 22320 9936 22800 10056 6 chanx_right_in[12]
port 49 nsew default input
rlabel metal3 s 22320 10344 22800 10464 6 chanx_right_in[13]
port 50 nsew default input
rlabel metal3 s 22320 10752 22800 10872 6 chanx_right_in[14]
port 51 nsew default input
rlabel metal3 s 22320 11296 22800 11416 6 chanx_right_in[15]
port 52 nsew default input
rlabel metal3 s 22320 11704 22800 11824 6 chanx_right_in[16]
port 53 nsew default input
rlabel metal3 s 22320 12248 22800 12368 6 chanx_right_in[17]
port 54 nsew default input
rlabel metal3 s 22320 12656 22800 12776 6 chanx_right_in[18]
port 55 nsew default input
rlabel metal3 s 22320 13200 22800 13320 6 chanx_right_in[19]
port 56 nsew default input
rlabel metal3 s 22320 4768 22800 4888 6 chanx_right_in[1]
port 57 nsew default input
rlabel metal3 s 22320 5176 22800 5296 6 chanx_right_in[2]
port 58 nsew default input
rlabel metal3 s 22320 5720 22800 5840 6 chanx_right_in[3]
port 59 nsew default input
rlabel metal3 s 22320 6128 22800 6248 6 chanx_right_in[4]
port 60 nsew default input
rlabel metal3 s 22320 6672 22800 6792 6 chanx_right_in[5]
port 61 nsew default input
rlabel metal3 s 22320 7080 22800 7200 6 chanx_right_in[6]
port 62 nsew default input
rlabel metal3 s 22320 7488 22800 7608 6 chanx_right_in[7]
port 63 nsew default input
rlabel metal3 s 22320 8032 22800 8152 6 chanx_right_in[8]
port 64 nsew default input
rlabel metal3 s 22320 8440 22800 8560 6 chanx_right_in[9]
port 65 nsew default input
rlabel metal3 s 22320 13608 22800 13728 6 chanx_right_out[0]
port 66 nsew default tristate
rlabel metal3 s 22320 18232 22800 18352 6 chanx_right_out[10]
port 67 nsew default tristate
rlabel metal3 s 22320 18776 22800 18896 6 chanx_right_out[11]
port 68 nsew default tristate
rlabel metal3 s 22320 19184 22800 19304 6 chanx_right_out[12]
port 69 nsew default tristate
rlabel metal3 s 22320 19728 22800 19848 6 chanx_right_out[13]
port 70 nsew default tristate
rlabel metal3 s 22320 20136 22800 20256 6 chanx_right_out[14]
port 71 nsew default tristate
rlabel metal3 s 22320 20544 22800 20664 6 chanx_right_out[15]
port 72 nsew default tristate
rlabel metal3 s 22320 21088 22800 21208 6 chanx_right_out[16]
port 73 nsew default tristate
rlabel metal3 s 22320 21496 22800 21616 6 chanx_right_out[17]
port 74 nsew default tristate
rlabel metal3 s 22320 22040 22800 22160 6 chanx_right_out[18]
port 75 nsew default tristate
rlabel metal3 s 22320 22448 22800 22568 6 chanx_right_out[19]
port 76 nsew default tristate
rlabel metal3 s 22320 14016 22800 14136 6 chanx_right_out[1]
port 77 nsew default tristate
rlabel metal3 s 22320 14560 22800 14680 6 chanx_right_out[2]
port 78 nsew default tristate
rlabel metal3 s 22320 14968 22800 15088 6 chanx_right_out[3]
port 79 nsew default tristate
rlabel metal3 s 22320 15512 22800 15632 6 chanx_right_out[4]
port 80 nsew default tristate
rlabel metal3 s 22320 15920 22800 16040 6 chanx_right_out[5]
port 81 nsew default tristate
rlabel metal3 s 22320 16464 22800 16584 6 chanx_right_out[6]
port 82 nsew default tristate
rlabel metal3 s 22320 16872 22800 16992 6 chanx_right_out[7]
port 83 nsew default tristate
rlabel metal3 s 22320 17280 22800 17400 6 chanx_right_out[8]
port 84 nsew default tristate
rlabel metal3 s 22320 17824 22800 17944 6 chanx_right_out[9]
port 85 nsew default tristate
rlabel metal2 s 5630 22320 5686 22800 6 chany_top_in[0]
port 86 nsew default input
rlabel metal2 s 9862 22320 9918 22800 6 chany_top_in[10]
port 87 nsew default input
rlabel metal2 s 10322 22320 10378 22800 6 chany_top_in[11]
port 88 nsew default input
rlabel metal2 s 10690 22320 10746 22800 6 chany_top_in[12]
port 89 nsew default input
rlabel metal2 s 11150 22320 11206 22800 6 chany_top_in[13]
port 90 nsew default input
rlabel metal2 s 11610 22320 11666 22800 6 chany_top_in[14]
port 91 nsew default input
rlabel metal2 s 11978 22320 12034 22800 6 chany_top_in[15]
port 92 nsew default input
rlabel metal2 s 12438 22320 12494 22800 6 chany_top_in[16]
port 93 nsew default input
rlabel metal2 s 12806 22320 12862 22800 6 chany_top_in[17]
port 94 nsew default input
rlabel metal2 s 13266 22320 13322 22800 6 chany_top_in[18]
port 95 nsew default input
rlabel metal2 s 13634 22320 13690 22800 6 chany_top_in[19]
port 96 nsew default input
rlabel metal2 s 6090 22320 6146 22800 6 chany_top_in[1]
port 97 nsew default input
rlabel metal2 s 6458 22320 6514 22800 6 chany_top_in[2]
port 98 nsew default input
rlabel metal2 s 6918 22320 6974 22800 6 chany_top_in[3]
port 99 nsew default input
rlabel metal2 s 7378 22320 7434 22800 6 chany_top_in[4]
port 100 nsew default input
rlabel metal2 s 7746 22320 7802 22800 6 chany_top_in[5]
port 101 nsew default input
rlabel metal2 s 8206 22320 8262 22800 6 chany_top_in[6]
port 102 nsew default input
rlabel metal2 s 8574 22320 8630 22800 6 chany_top_in[7]
port 103 nsew default input
rlabel metal2 s 9034 22320 9090 22800 6 chany_top_in[8]
port 104 nsew default input
rlabel metal2 s 9494 22320 9550 22800 6 chany_top_in[9]
port 105 nsew default input
rlabel metal2 s 14094 22320 14150 22800 6 chany_top_out[0]
port 106 nsew default tristate
rlabel metal2 s 18326 22320 18382 22800 6 chany_top_out[10]
port 107 nsew default tristate
rlabel metal2 s 18786 22320 18842 22800 6 chany_top_out[11]
port 108 nsew default tristate
rlabel metal2 s 19154 22320 19210 22800 6 chany_top_out[12]
port 109 nsew default tristate
rlabel metal2 s 19614 22320 19670 22800 6 chany_top_out[13]
port 110 nsew default tristate
rlabel metal2 s 19982 22320 20038 22800 6 chany_top_out[14]
port 111 nsew default tristate
rlabel metal2 s 20442 22320 20498 22800 6 chany_top_out[15]
port 112 nsew default tristate
rlabel metal2 s 20902 22320 20958 22800 6 chany_top_out[16]
port 113 nsew default tristate
rlabel metal2 s 21270 22320 21326 22800 6 chany_top_out[17]
port 114 nsew default tristate
rlabel metal2 s 21730 22320 21786 22800 6 chany_top_out[18]
port 115 nsew default tristate
rlabel metal2 s 22098 22320 22154 22800 6 chany_top_out[19]
port 116 nsew default tristate
rlabel metal2 s 14554 22320 14610 22800 6 chany_top_out[1]
port 117 nsew default tristate
rlabel metal2 s 14922 22320 14978 22800 6 chany_top_out[2]
port 118 nsew default tristate
rlabel metal2 s 15382 22320 15438 22800 6 chany_top_out[3]
port 119 nsew default tristate
rlabel metal2 s 15750 22320 15806 22800 6 chany_top_out[4]
port 120 nsew default tristate
rlabel metal2 s 16210 22320 16266 22800 6 chany_top_out[5]
port 121 nsew default tristate
rlabel metal2 s 16670 22320 16726 22800 6 chany_top_out[6]
port 122 nsew default tristate
rlabel metal2 s 17038 22320 17094 22800 6 chany_top_out[7]
port 123 nsew default tristate
rlabel metal2 s 17498 22320 17554 22800 6 chany_top_out[8]
port 124 nsew default tristate
rlabel metal2 s 17866 22320 17922 22800 6 chany_top_out[9]
port 125 nsew default tristate
rlabel metal2 s 4802 22320 4858 22800 6 clk_3_N_out
port 126 nsew default tristate
rlabel metal2 s 15842 0 15898 480 6 clk_3_S_in
port 127 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_11_
port 128 nsew default input
rlabel metal3 s 0 2864 480 2984 6 left_bottom_grid_pin_13_
port 129 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_bottom_grid_pin_15_
port 130 nsew default input
rlabel metal3 s 0 3816 480 3936 6 left_bottom_grid_pin_17_
port 131 nsew default input
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_1_
port 132 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_3_
port 133 nsew default input
rlabel metal3 s 0 960 480 1080 6 left_bottom_grid_pin_5_
port 134 nsew default input
rlabel metal3 s 0 1504 480 1624 6 left_bottom_grid_pin_7_
port 135 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_9_
port 136 nsew default input
rlabel metal2 s 3974 22320 4030 22800 6 prog_clk_0_N_in
port 137 nsew default input
rlabel metal2 s 5262 22320 5318 22800 6 prog_clk_3_N_out
port 138 nsew default tristate
rlabel metal2 s 11334 0 11390 480 6 prog_clk_3_S_in
port 139 nsew default input
rlabel metal3 s 22320 2456 22800 2576 6 right_bottom_grid_pin_11_
port 140 nsew default input
rlabel metal3 s 22320 2864 22800 2984 6 right_bottom_grid_pin_13_
port 141 nsew default input
rlabel metal3 s 22320 3408 22800 3528 6 right_bottom_grid_pin_15_
port 142 nsew default input
rlabel metal3 s 22320 3816 22800 3936 6 right_bottom_grid_pin_17_
port 143 nsew default input
rlabel metal3 s 22320 144 22800 264 6 right_bottom_grid_pin_1_
port 144 nsew default input
rlabel metal3 s 22320 552 22800 672 6 right_bottom_grid_pin_3_
port 145 nsew default input
rlabel metal3 s 22320 960 22800 1080 6 right_bottom_grid_pin_5_
port 146 nsew default input
rlabel metal3 s 22320 1504 22800 1624 6 right_bottom_grid_pin_7_
port 147 nsew default input
rlabel metal3 s 22320 1912 22800 2032 6 right_bottom_grid_pin_9_
port 148 nsew default input
rlabel metal2 s 570 22320 626 22800 6 top_left_grid_pin_42_
port 149 nsew default input
rlabel metal2 s 1030 22320 1086 22800 6 top_left_grid_pin_43_
port 150 nsew default input
rlabel metal2 s 1398 22320 1454 22800 6 top_left_grid_pin_44_
port 151 nsew default input
rlabel metal2 s 1858 22320 1914 22800 6 top_left_grid_pin_45_
port 152 nsew default input
rlabel metal2 s 2226 22320 2282 22800 6 top_left_grid_pin_46_
port 153 nsew default input
rlabel metal2 s 2686 22320 2742 22800 6 top_left_grid_pin_47_
port 154 nsew default input
rlabel metal2 s 3146 22320 3202 22800 6 top_left_grid_pin_48_
port 155 nsew default input
rlabel metal2 s 3514 22320 3570 22800 6 top_left_grid_pin_49_
port 156 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 157 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 158 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22800
<< end >>
