* NGSPICE file created from sb_1__0_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand3_4 abstract view
.subckt scs8hd_nand3_4 A B C Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

.subckt sb_1__0_ address[0] address[1] address[2] address[3] address[4] address[5]
+ address[6] chanx_left_in[0] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4]
+ chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_out[0]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_right_in[0] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_out[0] chanx_right_out[1] chanx_right_out[2]
+ chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6] chanx_right_out[7]
+ chanx_right_out[8] chany_top_in[0] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_out[0] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] data_in enable
+ left_bottom_grid_pin_11_ left_bottom_grid_pin_13_ left_bottom_grid_pin_15_ left_bottom_grid_pin_1_
+ left_bottom_grid_pin_3_ left_bottom_grid_pin_5_ left_bottom_grid_pin_7_ left_bottom_grid_pin_9_
+ left_top_grid_pin_10_ right_bottom_grid_pin_11_ right_bottom_grid_pin_13_ right_bottom_grid_pin_15_
+ right_bottom_grid_pin_1_ right_bottom_grid_pin_3_ right_bottom_grid_pin_5_ right_bottom_grid_pin_7_
+ right_bottom_grid_pin_9_ right_top_grid_pin_10_ top_left_grid_pin_13_ top_right_grid_pin_11_
+ vpwr vgnd
XANTENNA_mem_top_track_2.LATCH_1_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_104 vgnd vpwr scs8hd_fill_1
XFILLER_9_159 vpwr vgnd scs8hd_fill_2
XFILLER_13_144 vpwr vgnd scs8hd_fill_2
XANTENNA__113__B _075_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 chanx_right_in[6] mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_107 vpwr vgnd scs8hd_fill_2
XFILLER_10_158 vgnd vpwr scs8hd_decap_4
XFILLER_12_32 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_76 vgnd vpwr scs8hd_decap_4
XFILLER_37_62 vgnd vpwr scs8hd_decap_12
XFILLER_18_247 vpwr vgnd scs8hd_fill_2
XFILLER_18_258 vgnd vpwr scs8hd_decap_12
XANTENNA__108__B _111_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_162 vpwr vgnd scs8hd_fill_2
XANTENNA__124__A _096_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_3_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_31 vgnd vpwr scs8hd_decap_12
X_062_ _060_/A address[2] address[0] _079_/A vgnd vpwr scs8hd_or3_4
X_131_ _131_/HI _131_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_110 vpwr vgnd scs8hd_fill_2
XFILLER_9_11 vgnd vpwr scs8hd_decap_12
XFILLER_9_77 vpwr vgnd scs8hd_fill_2
XANTENNA__119__A _091_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_97 vgnd vpwr scs8hd_decap_3
XFILLER_11_242 vpwr vgnd scs8hd_fill_2
XFILLER_11_253 vpwr vgnd scs8hd_fill_2
XFILLER_11_275 vpwr vgnd scs8hd_fill_2
X_114_ _075_/A address[3] _104_/X _060_/C _114_/Y vgnd vpwr scs8hd_nor4_4
X_045_ _045_/A _045_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__105__C address[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB _109_/Y vgnd vpwr scs8hd_diode_2
XFILLER_38_117 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_4_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_9.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__121__B _120_/B vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_track_0.LATCH_4_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
XANTENNA__116__B _075_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_14.LATCH_1_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_67 vpwr vgnd scs8hd_fill_2
XFILLER_13_3 vpwr vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_1_.latch data_in mem_right_track_8.LATCH_1_.latch/Q _073_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_219 vpwr vgnd scs8hd_fill_2
XANTENNA__042__A _042_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _131_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_175 vpwr vgnd scs8hd_fill_2
XFILLER_40_178 vgnd vpwr scs8hd_fill_1
XFILLER_31_86 vgnd vpwr scs8hd_decap_12
XFILLER_0_263 vpwr vgnd scs8hd_fill_2
XFILLER_0_252 vpwr vgnd scs8hd_fill_2
XFILLER_31_123 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB _092_/Y vgnd vpwr scs8hd_diode_2
XFILLER_16_120 vgnd vpwr scs8hd_decap_3
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_245 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_145 vgnd vpwr scs8hd_decap_8
XFILLER_22_101 vgnd vpwr scs8hd_fill_1
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_3_57 vpwr vgnd scs8hd_fill_2
XANTENNA__113__C _104_/X vgnd vpwr scs8hd_diode_2
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_5_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_top_track_0.INVTX1_3_.scs8hd_inv_1 chanx_left_in[0] mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_193 vpwr vgnd scs8hd_fill_2
XFILLER_27_226 vpwr vgnd scs8hd_fill_2
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A right_bottom_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_27_248 vpwr vgnd scs8hd_fill_2
XFILLER_27_237 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_115 vgnd vpwr scs8hd_fill_1
XFILLER_10_137 vgnd vpwr scs8hd_decap_4
XFILLER_12_88 vpwr vgnd scs8hd_fill_2
XFILLER_37_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_141 vpwr vgnd scs8hd_fill_2
XANTENNA__124__B _120_/B vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _140_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_251 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_4_.scs8hd_inv_1 right_bottom_grid_pin_7_ mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__050__A enable vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_43 vgnd vpwr scs8hd_decap_12
X_130_ _130_/HI _130_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_122 vpwr vgnd scs8hd_fill_2
X_061_ _067_/A _078_/A _061_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mem_right_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_47 vgnd vpwr scs8hd_decap_4
XFILLER_0_58 vpwr vgnd scs8hd_fill_2
XANTENNA__119__B _120_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_23 vgnd vpwr scs8hd_decap_12
XFILLER_20_232 vgnd vpwr scs8hd_fill_1
XANTENNA__045__A _045_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_254 vgnd vpwr scs8hd_fill_1
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
X_113_ address[4] _075_/B _104_/X address[0] _113_/Y vgnd vpwr scs8hd_nor4_4
X_044_ _044_/A _044_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB _089_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__105__D _082_/X vgnd vpwr scs8hd_diode_2
XFILLER_38_129 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.INVTX1_6_.scs8hd_inv_1 left_bottom_grid_pin_5_ mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_184 vgnd vpwr scs8hd_decap_12
XFILLER_4_228 vpwr vgnd scs8hd_fill_2
XFILLER_20_44 vgnd vpwr scs8hd_decap_12
XFILLER_29_97 vpwr vgnd scs8hd_fill_2
XANTENNA__116__C _104_/X vgnd vpwr scs8hd_diode_2
XFILLER_6_46 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB _081_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_162 vpwr vgnd scs8hd_fill_2
XFILLER_19_195 vpwr vgnd scs8hd_fill_2
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_165 vpwr vgnd scs8hd_fill_2
XFILLER_15_77 vpwr vgnd scs8hd_fill_2
XFILLER_31_98 vgnd vpwr scs8hd_decap_8
XFILLER_0_275 vpwr vgnd scs8hd_fill_2
XFILLER_31_135 vgnd vpwr scs8hd_fill_1
Xmux_right_track_16.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_113 vgnd vpwr scs8hd_decap_4
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_165 vpwr vgnd scs8hd_fill_2
XFILLER_16_187 vgnd vpwr scs8hd_decap_8
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_22_113 vpwr vgnd scs8hd_fill_2
XANTENNA__053__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_26_32 vgnd vpwr scs8hd_decap_12
Xmux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ _042_/Y mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_9_139 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_113 vpwr vgnd scs8hd_fill_2
XFILLER_13_179 vpwr vgnd scs8hd_fill_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
XANTENNA__113__D address[0] vgnd vpwr scs8hd_diode_2
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__138__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_8_161 vgnd vpwr scs8hd_decap_3
XFILLER_27_205 vpwr vgnd scs8hd_fill_2
XANTENNA__048__A address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_86 vgnd vpwr scs8hd_decap_12
XFILLER_37_31 vgnd vpwr scs8hd_decap_12
XFILLER_33_208 vgnd vpwr scs8hd_decap_12
XFILLER_5_175 vpwr vgnd scs8hd_fill_2
XFILLER_32_263 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.INVTX1_7_.scs8hd_inv_1 chanx_left_in[4] mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_55 vgnd vpwr scs8hd_decap_6
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_145 vpwr vgnd scs8hd_fill_2
X_060_ _060_/A address[2] _060_/C _078_/A vgnd vpwr scs8hd_or3_4
XFILLER_2_178 vgnd vpwr scs8hd_fill_1
XFILLER_0_15 vgnd vpwr scs8hd_decap_12
XFILLER_9_35 vgnd vpwr scs8hd_decap_6
XFILLER_14_241 vgnd vpwr scs8hd_decap_4
XFILLER_9_57 vpwr vgnd scs8hd_fill_2
XFILLER_36_3 vgnd vpwr scs8hd_decap_12
XANTENNA__151__A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _042_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_244 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XANTENNA__061__A _067_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_44 vgnd vpwr scs8hd_decap_12
XFILLER_34_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A _133_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_18_88 vpwr vgnd scs8hd_fill_2
X_043_ _043_/A _043_/Y vgnd vpwr scs8hd_inv_8
X_112_ address[4] _075_/B _104_/X _060_/C _112_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_7_248 vpwr vgnd scs8hd_fill_2
XFILLER_7_259 vpwr vgnd scs8hd_fill_2
XANTENNA__146__A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_6_270 vgnd vpwr scs8hd_decap_4
XFILLER_37_196 vgnd vpwr scs8hd_decap_12
XANTENNA__056__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_20_56 vgnd vpwr scs8hd_decap_12
XFILLER_28_163 vpwr vgnd scs8hd_fill_2
XFILLER_28_141 vpwr vgnd scs8hd_fill_2
XANTENNA__116__D _060_/C vgnd vpwr scs8hd_diode_2
XFILLER_3_273 vgnd vpwr scs8hd_decap_4
XFILLER_3_262 vpwr vgnd scs8hd_fill_2
XFILLER_3_251 vgnd vpwr scs8hd_decap_4
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_141 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_199 vpwr vgnd scs8hd_fill_2
XFILLER_0_243 vgnd vpwr scs8hd_decap_4
Xmux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _128_/HI mem_right_track_0.LATCH_2_.latch/Q
+ mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_31_158 vpwr vgnd scs8hd_fill_2
XFILLER_31_147 vgnd vpwr scs8hd_decap_8
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_9.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB _069_/Y vgnd vpwr scs8hd_diode_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_177 vgnd vpwr scs8hd_fill_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_258 vpwr vgnd scs8hd_fill_2
XFILLER_39_236 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_125 vgnd vpwr scs8hd_decap_3
XFILLER_26_44 vgnd vpwr scs8hd_decap_12
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_26_88 vgnd vpwr scs8hd_decap_4
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_169 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_3_15 vgnd vpwr scs8hd_decap_12
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
XANTENNA__154__A _154_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__064__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_12_46 vpwr vgnd scs8hd_fill_2
XFILLER_18_206 vpwr vgnd scs8hd_fill_2
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_98 vgnd vpwr scs8hd_decap_12
XFILLER_37_43 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _135_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_7 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_0_.latch data_in mem_top_track_0.LATCH_0_.latch/Q _111_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A left_bottom_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__149__A _149_/A vgnd vpwr scs8hd_diode_2
XANTENNA__059__A _067_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_168 vpwr vgnd scs8hd_fill_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
Xmem_left_track_17.LATCH_3_.latch data_in mem_left_track_17.LATCH_3_.latch/Q _100_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_3 vgnd vpwr scs8hd_decap_12
XANTENNA__061__B _078_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_56 vgnd vpwr scs8hd_decap_12
XFILLER_34_44 vgnd vpwr scs8hd_decap_12
X_111_ _096_/A _111_/B _111_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_238 vgnd vpwr scs8hd_decap_6
XFILLER_11_245 vgnd vpwr scs8hd_decap_8
X_042_ _042_/A _042_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB _065_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB _042_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__162__A _162_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_81 vpwr vgnd scs8hd_fill_2
XANTENNA__072__A _079_/A vgnd vpwr scs8hd_diode_2
XANTENNA__056__B _075_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_68 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_241 vgnd vpwr scs8hd_decap_3
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XANTENNA__157__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XFILLER_19_175 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_25_123 vgnd vpwr scs8hd_decap_4
XFILLER_25_112 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_145 vgnd vpwr scs8hd_decap_4
XANTENNA__067__A _067_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_145 vgnd vpwr scs8hd_decap_6
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_1_.latch data_in mem_left_track_1.LATCH_1_.latch/Q _088_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_67 vgnd vpwr scs8hd_decap_6
XFILLER_26_56 vpwr vgnd scs8hd_fill_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_13_148 vpwr vgnd scs8hd_fill_2
XFILLER_3_27 vgnd vpwr scs8hd_decap_12
Xmem_right_track_16.LATCH_2_.latch data_in mem_right_track_16.LATCH_2_.latch/Q _079_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__064__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_10_118 vpwr vgnd scs8hd_fill_2
XFILLER_12_36 vgnd vpwr scs8hd_fill_1
XANTENNA__080__A _080_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_55 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_16.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_26_273 vpwr vgnd scs8hd_fill_2
XFILLER_5_100 vpwr vgnd scs8hd_fill_2
XFILLER_17_240 vpwr vgnd scs8hd_fill_2
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XFILLER_23_243 vgnd vpwr scs8hd_fill_1
XFILLER_23_210 vgnd vpwr scs8hd_decap_4
XANTENNA__059__B _059_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__075__A _075_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_114 vpwr vgnd scs8hd_fill_2
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_224 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_68 vgnd vpwr scs8hd_decap_12
XFILLER_34_56 vgnd vpwr scs8hd_decap_12
XFILLER_11_213 vpwr vgnd scs8hd_fill_2
X_110_ _080_/A _111_/B _110_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_217 vpwr vgnd scs8hd_fill_2
XFILLER_7_228 vgnd vpwr scs8hd_decap_4
X_041_ _041_/A _041_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_110 vgnd vpwr scs8hd_decap_12
XANTENNA__056__C _075_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__072__B _070_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XFILLER_13_7 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB _095_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_105 vgnd vpwr scs8hd_decap_12
XFILLER_25_179 vpwr vgnd scs8hd_fill_2
XANTENNA__067__B _096_/A vgnd vpwr scs8hd_diode_2
XANTENNA__083__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_267 vgnd vpwr scs8hd_decap_8
XFILLER_0_256 vgnd vpwr scs8hd_decap_4
XFILLER_31_127 vpwr vgnd scs8hd_fill_2
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA__078__A _078_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_138 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_193 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_39 vgnd vpwr scs8hd_decap_12
XFILLER_12_182 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__064__C _060_/C vgnd vpwr scs8hd_diode_2
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
XFILLER_12_59 vpwr vgnd scs8hd_fill_2
XANTENNA__080__B _079_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_241 vgnd vpwr scs8hd_decap_12
Xmem_right_track_0.LATCH_1_.latch data_in mem_right_track_0.LATCH_1_.latch/Q _065_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_top_track_8.LATCH_1_.latch data_in _043_/A _114_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_123 vgnd vpwr scs8hd_decap_4
XFILLER_5_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_233 vpwr vgnd scs8hd_fill_2
XANTENNA__075__B _075_/B vgnd vpwr scs8hd_diode_2
XANTENNA__091__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_126 vpwr vgnd scs8hd_fill_2
XFILLER_14_211 vgnd vpwr scs8hd_fill_1
XFILLER_13_80 vgnd vpwr scs8hd_decap_4
XFILLER_1_181 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_258 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[0] mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_68 vgnd vpwr scs8hd_decap_12
XANTENNA__086__A _078_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_79 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_199 vpwr vgnd scs8hd_fill_2
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XFILLER_40_117 vgnd vpwr scs8hd_decap_12
XFILLER_25_169 vgnd vpwr scs8hd_decap_4
XFILLER_15_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__083__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_15_59 vpwr vgnd scs8hd_fill_2
XFILLER_0_213 vpwr vgnd scs8hd_fill_2
XFILLER_0_202 vgnd vpwr scs8hd_decap_4
XFILLER_16_103 vpwr vgnd scs8hd_fill_2
XFILLER_31_117 vgnd vpwr scs8hd_fill_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_125 vpwr vgnd scs8hd_fill_2
XFILLER_16_169 vgnd vpwr scs8hd_decap_8
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_80 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_3_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_228 vgnd vpwr scs8hd_decap_3
XPHY_0 vgnd vpwr scs8hd_decap_3
XFILLER_22_117 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_180 vgnd vpwr scs8hd_decap_3
Xmem_left_track_9.LATCH_2_.latch data_in mem_left_track_9.LATCH_2_.latch/Q _094_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_7_71 vpwr vgnd scs8hd_fill_2
XANTENNA__078__B _079_/B vgnd vpwr scs8hd_diode_2
XANTENNA__094__A _079_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_117 vpwr vgnd scs8hd_fill_2
Xmem_top_track_14.LATCH_0_.latch data_in _046_/A _117_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_154 vgnd vpwr scs8hd_decap_3
XFILLER_12_150 vgnd vpwr scs8hd_decap_3
XFILLER_27_209 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _041_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
Xmux_right_track_0.INVTX1_4_.scs8hd_inv_1 right_bottom_grid_pin_5_ mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_253 vgnd vpwr scs8hd_decap_12
Xmem_top_track_16.LATCH_3_.latch data_in mem_top_track_16.LATCH_3_.latch/Q _121_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__089__A _096_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_113 vgnd vpwr scs8hd_decap_4
XFILLER_5_179 vpwr vgnd scs8hd_fill_2
Xmux_top_track_14.tap_buf4_0_.scs8hd_inv_1 mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ _155_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_245 vgnd vpwr scs8hd_decap_12
XANTENNA__075__C _075_/C vgnd vpwr scs8hd_diode_2
XANTENNA__091__B _094_/B vgnd vpwr scs8hd_diode_2
XFILLER_2_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A left_bottom_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_204 vpwr vgnd scs8hd_fill_2
XFILLER_20_248 vgnd vpwr scs8hd_decap_6
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
XANTENNA__086__B _087_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_226 vpwr vgnd scs8hd_fill_2
XFILLER_11_259 vpwr vgnd scs8hd_fill_2
XFILLER_24_91 vgnd vpwr scs8hd_fill_1
XFILLER_24_80 vpwr vgnd scs8hd_fill_2
XFILLER_6_241 vgnd vpwr scs8hd_decap_8
XFILLER_6_274 vgnd vpwr scs8hd_fill_1
XFILLER_27_3 vgnd vpwr scs8hd_decap_12
X_099_ _059_/B _103_/B _099_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_123 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_1_62 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_5_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XFILLER_28_145 vpwr vgnd scs8hd_fill_2
XFILLER_28_189 vgnd vpwr scs8hd_decap_6
XFILLER_28_167 vgnd vpwr scs8hd_decap_12
XANTENNA__097__A _075_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_233 vpwr vgnd scs8hd_fill_2
XFILLER_3_222 vpwr vgnd scs8hd_fill_2
XFILLER_10_71 vgnd vpwr scs8hd_decap_4
XFILLER_10_93 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_101 vpwr vgnd scs8hd_fill_2
XFILLER_19_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB _072_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_129 vgnd vpwr scs8hd_decap_12
XFILLER_25_115 vpwr vgnd scs8hd_fill_2
XFILLER_25_104 vpwr vgnd scs8hd_fill_2
XFILLER_15_27 vgnd vpwr scs8hd_decap_12
XFILLER_31_59 vpwr vgnd scs8hd_fill_2
XFILLER_31_15 vgnd vpwr scs8hd_decap_12
XANTENNA__083__C _090_/C vgnd vpwr scs8hd_diode_2
XFILLER_0_247 vgnd vpwr scs8hd_fill_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_38_251 vgnd vpwr scs8hd_decap_12
XFILLER_26_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__094__B _094_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_162 vpwr vgnd scs8hd_fill_2
XFILLER_21_140 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB _084_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_80 vgnd vpwr scs8hd_decap_12
XFILLER_8_122 vgnd vpwr scs8hd_fill_1
XFILLER_8_166 vgnd vpwr scs8hd_decap_3
XFILLER_16_81 vpwr vgnd scs8hd_fill_2
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XANTENNA__089__B _087_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_4_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_26_265 vgnd vpwr scs8hd_decap_8
Xmem_right_track_8.LATCH_2_.latch data_in mem_right_track_8.LATCH_2_.latch/Q _072_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XFILLER_5_158 vpwr vgnd scs8hd_fill_2
XFILLER_17_221 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB _076_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_202 vgnd vpwr scs8hd_decap_12
XFILLER_17_254 vpwr vgnd scs8hd_fill_2
XFILLER_17_265 vgnd vpwr scs8hd_decap_12
XFILLER_4_84 vgnd vpwr scs8hd_decap_3
XFILLER_23_257 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.INVTX1_5_.scs8hd_inv_1 right_bottom_grid_pin_15_ mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_6_.scs8hd_inv_1 left_bottom_grid_pin_9_ mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_224 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_5_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _131_/HI mem_top_track_0.LATCH_5_.latch/Q
+ mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_14.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
XFILLER_10_271 vgnd vpwr scs8hd_decap_4
X_098_ _091_/A _103_/B _098_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_135 vgnd vpwr scs8hd_decap_12
XFILLER_1_85 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_59 vpwr vgnd scs8hd_fill_2
XFILLER_28_179 vgnd vpwr scs8hd_fill_1
XFILLER_28_124 vpwr vgnd scs8hd_fill_2
XANTENNA__097__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_36_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB _100_/Y vgnd vpwr scs8hd_diode_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _115_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_50 vpwr vgnd scs8hd_fill_2
XFILLER_34_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_19_81 vgnd vpwr scs8hd_decap_4
XFILLER_19_179 vpwr vgnd scs8hd_fill_2
XFILLER_33_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_25_149 vgnd vpwr scs8hd_fill_1
XFILLER_25_127 vgnd vpwr scs8hd_fill_1
XFILLER_15_39 vgnd vpwr scs8hd_decap_12
XFILLER_31_27 vgnd vpwr scs8hd_decap_12
XANTENNA__083__D _082_/X vgnd vpwr scs8hd_diode_2
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_182 vgnd vpwr scs8hd_fill_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_208 vgnd vpwr scs8hd_decap_12
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_15_171 vgnd vpwr scs8hd_decap_3
XFILLER_15_193 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_38_263 vgnd vpwr scs8hd_decap_12
XFILLER_26_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A right_bottom_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_230 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _126_/HI mem_left_track_17.LATCH_2_.latch/Q
+ mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_16_93 vgnd vpwr scs8hd_fill_1
XFILLER_8_145 vgnd vpwr scs8hd_decap_8
XFILLER_8_178 vgnd vpwr scs8hd_decap_6
XFILLER_8_189 vpwr vgnd scs8hd_fill_2
XFILLER_12_185 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_211 vgnd vpwr scs8hd_fill_1
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
XFILLER_17_211 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _144_/A vgnd vpwr scs8hd_inv_1
XFILLER_4_181 vgnd vpwr scs8hd_decap_8
XFILLER_23_225 vpwr vgnd scs8hd_fill_2
XFILLER_23_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.tap_buf4_0_.scs8hd_inv_1 mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ _161_/A vgnd vpwr scs8hd_inv_1
XFILLER_14_203 vpwr vgnd scs8hd_fill_2
XFILLER_14_247 vgnd vpwr scs8hd_decap_12
XFILLER_1_184 vgnd vpwr scs8hd_decap_3
XFILLER_1_162 vpwr vgnd scs8hd_fill_2
XFILLER_38_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _127_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
X_097_ _075_/A address[3] _090_/C _082_/X _103_/B vgnd vpwr scs8hd_or4_4
XFILLER_37_147 vgnd vpwr scs8hd_decap_12
XFILLER_1_42 vgnd vpwr scs8hd_decap_8
XFILLER_1_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_27 vgnd vpwr scs8hd_decap_12
XANTENNA__097__C _090_/C vgnd vpwr scs8hd_diode_2
XFILLER_10_84 vpwr vgnd scs8hd_fill_2
XFILLER_19_114 vpwr vgnd scs8hd_fill_2
XFILLER_34_117 vgnd vpwr scs8hd_decap_12
XFILLER_27_191 vgnd vpwr scs8hd_decap_3
XFILLER_19_158 vpwr vgnd scs8hd_fill_2
X_149_ _149_/A chanx_right_out[4] vgnd vpwr scs8hd_buf_2
XFILLER_32_3 vgnd vpwr scs8hd_decap_12
XFILLER_18_191 vgnd vpwr scs8hd_decap_8
XFILLER_31_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_227 vgnd vpwr scs8hd_decap_8
XFILLER_31_109 vpwr vgnd scs8hd_fill_2
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_194 vpwr vgnd scs8hd_fill_2
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_164 vgnd vpwr scs8hd_decap_12
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_15_150 vgnd vpwr scs8hd_decap_4
XFILLER_7_96 vpwr vgnd scs8hd_fill_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_21_175 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_242 vpwr vgnd scs8hd_fill_2
XFILLER_12_120 vpwr vgnd scs8hd_fill_2
XFILLER_12_142 vgnd vpwr scs8hd_decap_8
XFILLER_32_93 vgnd vpwr scs8hd_decap_12
XFILLER_8_135 vgnd vpwr scs8hd_decap_8
XFILLER_35_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_127 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_93 vgnd vpwr scs8hd_decap_4
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XFILLER_23_237 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_right_track_8.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A right_bottom_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_40 vpwr vgnd scs8hd_fill_2
XFILLER_14_259 vgnd vpwr scs8hd_decap_12
XFILLER_13_62 vgnd vpwr scs8hd_decap_3
XFILLER_13_95 vpwr vgnd scs8hd_fill_2
XANTENNA__100__A _078_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB _122_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_93 vgnd vpwr scs8hd_decap_12
X_096_ _096_/A _094_/B _096_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_37_159 vgnd vpwr scs8hd_decap_12
Xmem_top_track_0.LATCH_1_.latch data_in mem_top_track_0.LATCH_1_.latch/Q _110_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_39 vgnd vpwr scs8hd_decap_12
XANTENNA__097__D _082_/X vgnd vpwr scs8hd_diode_2
XFILLER_3_269 vpwr vgnd scs8hd_fill_2
XFILLER_3_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A chany_top_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_34_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_14.INVTX1_1_.scs8hd_inv_1 chanx_left_in[8] mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_148_ chanx_left_in[4] chanx_right_out[5] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_079_ _079_/A _079_/B _079_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_3 vgnd vpwr scs8hd_decap_12
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
Xmem_left_track_17.LATCH_4_.latch data_in mem_left_track_17.LATCH_4_.latch/Q _099_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_239 vpwr vgnd scs8hd_fill_2
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_107 vpwr vgnd scs8hd_fill_2
XFILLER_16_129 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_62 vgnd vpwr scs8hd_decap_3
XFILLER_21_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_5_.scs8hd_inv_1 left_bottom_grid_pin_1_ mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_30_176 vgnd vpwr scs8hd_decap_12
XFILLER_30_154 vgnd vpwr scs8hd_fill_1
XFILLER_30_121 vgnd vpwr scs8hd_fill_1
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_7_53 vpwr vgnd scs8hd_fill_2
XFILLER_7_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_110 vpwr vgnd scs8hd_fill_2
XFILLER_21_187 vgnd vpwr scs8hd_decap_4
XFILLER_21_154 vpwr vgnd scs8hd_fill_2
XFILLER_21_132 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB _042_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_103 vpwr vgnd scs8hd_fill_2
XFILLER_8_125 vgnd vpwr scs8hd_fill_1
XFILLER_12_110 vgnd vpwr scs8hd_fill_1
XFILLER_12_165 vgnd vpwr scs8hd_decap_8
XFILLER_12_176 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A left_bottom_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__103__A _096_/A vgnd vpwr scs8hd_diode_2
Xmux_right_track_0.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
XFILLER_26_224 vgnd vpwr scs8hd_decap_8
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XFILLER_23_19 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_120 vpwr vgnd scs8hd_fill_2
XFILLER_38_93 vgnd vpwr scs8hd_decap_12
XANTENNA__100__B _103_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_175 vgnd vpwr scs8hd_decap_4
Xmem_left_track_1.LATCH_2_.latch data_in mem_left_track_1.LATCH_2_.latch/Q _087_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_208 vgnd vpwr scs8hd_decap_4
XFILLER_9_231 vgnd vpwr scs8hd_fill_1
XFILLER_9_242 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.LATCH_3_.latch data_in mem_right_track_16.LATCH_3_.latch/Q _078_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_84 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_095_ _080_/A _094_/B _095_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__111__A _096_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_66 vgnd vpwr scs8hd_decap_4
Xmux_right_track_8.INVTX1_6_.scs8hd_inv_1 chanx_left_in[1] mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_28_149 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_237 vpwr vgnd scs8hd_fill_2
XFILLER_3_226 vpwr vgnd scs8hd_fill_2
XFILLER_10_97 vpwr vgnd scs8hd_fill_2
XFILLER_19_62 vgnd vpwr scs8hd_decap_12
XFILLER_27_182 vgnd vpwr scs8hd_fill_1
X_078_ _078_/A _079_/B _078_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__106__A _091_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_147_ chanx_left_in[5] chanx_right_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_119 vgnd vpwr scs8hd_decap_3
XFILLER_25_108 vgnd vpwr scs8hd_decap_4
XFILLER_18_171 vgnd vpwr scs8hd_decap_4
XFILLER_33_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_24_174 vgnd vpwr scs8hd_decap_8
XFILLER_24_163 vpwr vgnd scs8hd_fill_2
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_3_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB _087_/Y vgnd vpwr scs8hd_diode_2
XFILLER_30_188 vgnd vpwr scs8hd_decap_12
XFILLER_30_133 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_3_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_199 vpwr vgnd scs8hd_fill_2
XFILLER_16_85 vpwr vgnd scs8hd_fill_2
XANTENNA__103__B _103_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB _079_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_73 vpwr vgnd scs8hd_fill_2
XFILLER_27_62 vgnd vpwr scs8hd_decap_6
XFILLER_27_51 vgnd vpwr scs8hd_decap_8
XFILLER_17_236 vpwr vgnd scs8hd_fill_2
XFILLER_17_258 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_16.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.INVTX1_2_.scs8hd_inv_1 chany_top_in[7] mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_left_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_4_162 vgnd vpwr scs8hd_decap_4
XANTENNA__114__A _075_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_206 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_228 vgnd vpwr scs8hd_decap_4
XFILLER_22_272 vgnd vpwr scs8hd_decap_3
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_110 vpwr vgnd scs8hd_fill_2
XFILLER_1_154 vpwr vgnd scs8hd_fill_2
XFILLER_1_198 vpwr vgnd scs8hd_fill_2
XFILLER_9_210 vgnd vpwr scs8hd_decap_4
XANTENNA__109__A _079_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_209 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_094_ _079_/A _094_/B _094_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_224 vpwr vgnd scs8hd_fill_2
XANTENNA__111__B _111_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB _103_/Y vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_2_.latch data_in mem_right_track_0.LATCH_2_.latch/Q _063_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_128 vpwr vgnd scs8hd_fill_2
XFILLER_3_205 vpwr vgnd scs8hd_fill_2
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_10_54 vpwr vgnd scs8hd_fill_2
XFILLER_35_51 vgnd vpwr scs8hd_decap_8
XFILLER_19_74 vgnd vpwr scs8hd_fill_1
XFILLER_19_85 vgnd vpwr scs8hd_fill_1
XFILLER_19_128 vpwr vgnd scs8hd_fill_2
XFILLER_35_62 vgnd vpwr scs8hd_decap_12
X_146_ chanx_left_in[6] chanx_right_out[7] vgnd vpwr scs8hd_buf_2
X_077_ _059_/B _079_/B _077_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__122__A _079_/A vgnd vpwr scs8hd_diode_2
XANTENNA__106__B _111_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_0_208 vgnd vpwr scs8hd_decap_3
XFILLER_24_120 vgnd vpwr scs8hd_decap_8
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_15_131 vpwr vgnd scs8hd_fill_2
XFILLER_30_145 vgnd vpwr scs8hd_decap_8
XANTENNA__117__A _075_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_197 vpwr vgnd scs8hd_fill_2
XFILLER_30_3 vgnd vpwr scs8hd_decap_12
X_129_ _129_/HI _129_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_12
XFILLER_29_234 vgnd vpwr scs8hd_decap_8
XFILLER_29_223 vgnd vpwr scs8hd_decap_4
Xmux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_2_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_64 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_2_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _130_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_7_160 vpwr vgnd scs8hd_fill_2
XFILLER_7_171 vpwr vgnd scs8hd_fill_2
XFILLER_7_193 vpwr vgnd scs8hd_fill_2
XFILLER_37_19 vgnd vpwr scs8hd_decap_12
XFILLER_34_270 vgnd vpwr scs8hd_decap_4
XFILLER_5_119 vgnd vpwr scs8hd_decap_3
Xmux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__114__B address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_152 vgnd vpwr scs8hd_fill_1
XFILLER_4_89 vgnd vpwr scs8hd_decap_3
XFILLER_4_67 vgnd vpwr scs8hd_decap_6
XFILLER_4_56 vgnd vpwr scs8hd_decap_8
XFILLER_23_229 vpwr vgnd scs8hd_fill_2
XFILLER_14_207 vgnd vpwr scs8hd_decap_4
XFILLER_13_76 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_3_.latch data_in mem_left_track_9.LATCH_3_.latch/Q _093_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
Xmem_top_track_14.LATCH_1_.latch data_in _045_/A _116_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__109__B _111_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_192 vpwr vgnd scs8hd_fill_2
XFILLER_39_181 vpwr vgnd scs8hd_fill_2
X_162_ _162_/A chany_top_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_6_258 vgnd vpwr scs8hd_decap_12
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
X_093_ _078_/A _094_/B _093_/Y vgnd vpwr scs8hd_nor2_4
Xmem_top_track_16.LATCH_4_.latch data_in mem_top_track_16.LATCH_4_.latch/Q _120_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_1_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_107 vgnd vpwr scs8hd_decap_8
XFILLER_10_88 vgnd vpwr scs8hd_decap_4
XFILLER_19_118 vpwr vgnd scs8hd_fill_2
XFILLER_35_74 vgnd vpwr scs8hd_decap_12
XFILLER_27_173 vgnd vpwr scs8hd_decap_3
XFILLER_19_97 vpwr vgnd scs8hd_fill_2
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
X_145_ _145_/A chanx_right_out[8] vgnd vpwr scs8hd_buf_2
Xmux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_4_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__122__B _120_/B vgnd vpwr scs8hd_diode_2
X_076_ _091_/A _079_/B _076_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_18_151 vpwr vgnd scs8hd_fill_2
XFILLER_33_110 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.INVTX1_0_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_132 vpwr vgnd scs8hd_fill_2
XFILLER_24_110 vgnd vpwr scs8hd_fill_1
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_198 vgnd vpwr scs8hd_decap_4
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_113 vgnd vpwr scs8hd_decap_8
XFILLER_30_102 vgnd vpwr scs8hd_decap_3
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_15_176 vpwr vgnd scs8hd_fill_2
XFILLER_15_187 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB _061_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__117__B _075_/B vgnd vpwr scs8hd_diode_2
X_128_ _128_/HI _128_/LO vgnd vpwr scs8hd_conb_1
XFILLER_38_202 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_3 vpwr vgnd scs8hd_fill_2
X_059_ _067_/A _059_/B _059_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_21_179 vpwr vgnd scs8hd_fill_2
XANTENNA__043__A _043_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_257 vgnd vpwr scs8hd_decap_12
XFILLER_29_202 vpwr vgnd scs8hd_fill_2
XFILLER_12_102 vpwr vgnd scs8hd_fill_2
XFILLER_12_124 vpwr vgnd scs8hd_fill_2
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A left_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_2.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_190 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.INVTX1_2_.scs8hd_inv_1 chanx_right_in[8] mux_top_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XFILLER_26_205 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A left_bottom_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__114__C _104_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_2.LATCH_0_.latch_SLEEPB _113_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_252 vgnd vpwr scs8hd_decap_12
XFILLER_22_241 vgnd vpwr scs8hd_decap_8
XFILLER_13_99 vgnd vpwr scs8hd_decap_3
XFILLER_1_134 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_234 vgnd vpwr scs8hd_decap_8
XFILLER_9_245 vgnd vpwr scs8hd_decap_12
XANTENNA__141__A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__051__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_24_76 vpwr vgnd scs8hd_fill_2
XFILLER_24_32 vgnd vpwr scs8hd_decap_12
X_161_ _161_/A chany_top_out[1] vgnd vpwr scs8hd_buf_2
X_092_ _059_/B _094_/B _092_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_8.LATCH_3_.latch data_in mem_right_track_8.LATCH_3_.latch/Q _071_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__136__A _136_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_141 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__046__A _046_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_67 vpwr vgnd scs8hd_fill_2
XFILLER_35_86 vgnd vpwr scs8hd_decap_12
XFILLER_27_152 vpwr vgnd scs8hd_fill_2
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_144_ _144_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
X_075_ _075_/A _075_/B _075_/C _079_/B vgnd vpwr scs8hd_or3_4
XFILLER_18_130 vpwr vgnd scs8hd_fill_2
XFILLER_18_163 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB _110_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_2_.scs8hd_inv_1 chany_top_in[8] mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_11 vgnd vpwr scs8hd_decap_12
XFILLER_21_99 vgnd vpwr scs8hd_decap_3
XFILLER_30_125 vpwr vgnd scs8hd_fill_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XANTENNA__117__C _104_/X vgnd vpwr scs8hd_diode_2
XFILLER_15_111 vpwr vgnd scs8hd_fill_2
X_127_ _127_/HI _127_/LO vgnd vpwr scs8hd_conb_1
X_058_ address[1] _054_/B address[0] _059_/B vgnd vpwr scs8hd_or3_4
XFILLER_7_57 vpwr vgnd scs8hd_fill_2
XFILLER_16_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_158 vpwr vgnd scs8hd_fill_2
XFILLER_21_136 vgnd vpwr scs8hd_decap_4
XFILLER_21_114 vgnd vpwr scs8hd_decap_6
Xmux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_5_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_29_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_14.LATCH_0_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_107 vpwr vgnd scs8hd_fill_2
XFILLER_8_118 vgnd vpwr scs8hd_decap_4
XFILLER_16_44 vgnd vpwr scs8hd_decap_12
XFILLER_32_32 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__144__A _144_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_180 vgnd vpwr scs8hd_decap_3
Xmux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _045_/A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB _093_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__054__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_17_217 vpwr vgnd scs8hd_fill_2
XFILLER_4_198 vpwr vgnd scs8hd_fill_2
XFILLER_4_154 vpwr vgnd scs8hd_fill_2
XFILLER_4_132 vgnd vpwr scs8hd_decap_3
XFILLER_4_110 vpwr vgnd scs8hd_fill_2
XANTENNA__114__D _060_/C vgnd vpwr scs8hd_diode_2
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XANTENNA__139__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_16_261 vgnd vpwr scs8hd_decap_12
XANTENNA__049__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_22_264 vgnd vpwr scs8hd_decap_8
Xmux_top_track_0.INVTX1_2_.scs8hd_inv_1 chanx_right_in[7] mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_13_242 vpwr vgnd scs8hd_fill_2
XFILLER_9_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_160_ chanx_right_in[4] chany_top_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
XFILLER_24_88 vgnd vpwr scs8hd_fill_1
XFILLER_24_44 vgnd vpwr scs8hd_decap_12
X_091_ _091_/A _094_/B _091_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_8.INVTX1_3_.scs8hd_inv_1 right_bottom_grid_pin_1_ mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_205 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_2.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_15 vgnd vpwr scs8hd_decap_12
XANTENNA__152__A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__062__A _060_/A vgnd vpwr scs8hd_diode_2
XFILLER_10_46 vgnd vpwr scs8hd_fill_1
XFILLER_19_11 vgnd vpwr scs8hd_decap_12
XFILLER_19_77 vpwr vgnd scs8hd_fill_2
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
XFILLER_35_98 vgnd vpwr scs8hd_decap_12
X_074_ _096_/A _070_/B _074_/Y vgnd vpwr scs8hd_nor2_4
X_143_ chanx_right_in[0] chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XFILLER_33_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_175 vgnd vpwr scs8hd_fill_1
XANTENNA__147__A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_2_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_24_167 vgnd vpwr scs8hd_decap_4
XFILLER_24_145 vgnd vpwr scs8hd_decap_8
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_1.INVTX1_5_.scs8hd_inv_1 left_top_grid_pin_10_ mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__057__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_67 vpwr vgnd scs8hd_fill_2
XFILLER_21_23 vgnd vpwr scs8hd_decap_12
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_123 vgnd vpwr scs8hd_decap_3
XANTENNA__117__D address[0] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_156 vpwr vgnd scs8hd_fill_2
XFILLER_15_167 vpwr vgnd scs8hd_fill_2
X_126_ _126_/HI _126_/LO vgnd vpwr scs8hd_conb_1
X_057_ _091_/A _067_/A _057_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_21_104 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_32_44 vgnd vpwr scs8hd_decap_12
XFILLER_16_56 vgnd vpwr scs8hd_decap_8
XFILLER_16_89 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__160__A chanx_right_in[4] vgnd vpwr scs8hd_diode_2
X_109_ _079_/A _111_/B _109_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_19_270 vgnd vpwr scs8hd_decap_6
XFILLER_34_251 vgnd vpwr scs8hd_decap_4
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__054__B _054_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__070__A _059_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_99 vpwr vgnd scs8hd_fill_2
XFILLER_27_77 vgnd vpwr scs8hd_decap_3
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
XFILLER_4_144 vpwr vgnd scs8hd_fill_2
XFILLER_4_15 vgnd vpwr scs8hd_decap_12
XFILLER_31_232 vgnd vpwr scs8hd_decap_12
XANTENNA__155__A _155_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_251 vgnd vpwr scs8hd_fill_1
XFILLER_16_273 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XANTENNA__065__A _067_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_114 vgnd vpwr scs8hd_decap_4
XFILLER_1_158 vpwr vgnd scs8hd_fill_2
XFILLER_38_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_214 vgnd vpwr scs8hd_fill_1
XFILLER_13_210 vpwr vgnd scs8hd_fill_2
XFILLER_9_269 vgnd vpwr scs8hd_decap_8
XFILLER_39_184 vgnd vpwr scs8hd_decap_4
XFILLER_24_56 vgnd vpwr scs8hd_decap_12
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XFILLER_6_228 vgnd vpwr scs8hd_decap_4
XFILLER_10_224 vpwr vgnd scs8hd_fill_2
XFILLER_10_235 vgnd vpwr scs8hd_decap_12
X_090_ address[4] _075_/B _090_/C _082_/X _094_/B vgnd vpwr scs8hd_or4_4
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_0.INVTX1_6_.scs8hd_inv_1 chanx_left_in[0] mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_27 vgnd vpwr scs8hd_decap_12
XFILLER_36_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_209 vpwr vgnd scs8hd_fill_2
XANTENNA__062__B address[2] vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_132 vpwr vgnd scs8hd_fill_2
XFILLER_19_23 vgnd vpwr scs8hd_decap_12
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
XFILLER_27_187 vpwr vgnd scs8hd_fill_2
X_142_ chanx_right_in[1] chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_073_ _080_/A _070_/B _073_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_33_135 vgnd vpwr scs8hd_decap_12
XFILLER_24_102 vpwr vgnd scs8hd_fill_2
XFILLER_2_81 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_2.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_32_190 vgnd vpwr scs8hd_decap_12
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__057__B _067_/A vgnd vpwr scs8hd_diode_2
XANTENNA__073__A _080_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_35 vgnd vpwr scs8hd_decap_12
XFILLER_15_135 vpwr vgnd scs8hd_fill_2
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
X_125_ _125_/HI _125_/LO vgnd vpwr scs8hd_conb_1
X_056_ address[4] _075_/B _075_/C _067_/A vgnd vpwr scs8hd_or3_4
XFILLER_38_227 vgnd vpwr scs8hd_decap_12
XANTENNA__158__A _158_/A vgnd vpwr scs8hd_diode_2
XANTENNA__068__A _075_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_68 vpwr vgnd scs8hd_fill_2
XFILLER_32_56 vgnd vpwr scs8hd_decap_12
XFILLER_12_138 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_2_.latch data_in mem_top_track_0.LATCH_2_.latch/Q _109_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
XFILLER_28_271 vgnd vpwr scs8hd_decap_4
XFILLER_7_164 vpwr vgnd scs8hd_fill_2
XFILLER_7_175 vpwr vgnd scs8hd_fill_2
XFILLER_7_197 vpwr vgnd scs8hd_fill_2
X_108_ _078_/A _111_/B _108_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A right_bottom_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_34_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB _070_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__070__B _070_/B vgnd vpwr scs8hd_diode_2
XANTENNA__054__C _060_/C vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _158_/A vgnd vpwr scs8hd_inv_1
XFILLER_8_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_244 vgnd vpwr scs8hd_decap_12
Xmem_left_track_17.LATCH_5_.latch data_in mem_left_track_17.LATCH_5_.latch/Q _098_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_27 vgnd vpwr scs8hd_decap_4
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_13_36 vpwr vgnd scs8hd_fill_2
XANTENNA__065__B _080_/A vgnd vpwr scs8hd_diode_2
XANTENNA__081__A _096_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_44 vgnd vpwr scs8hd_decap_12
XFILLER_0_181 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_1.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_196 vgnd vpwr scs8hd_decap_12
XFILLER_24_68 vgnd vpwr scs8hd_decap_8
XANTENNA__076__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XFILLER_10_247 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_36_166 vgnd vpwr scs8hd_decap_12
XANTENNA__062__C address[0] vgnd vpwr scs8hd_diode_2
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_19_35 vgnd vpwr scs8hd_decap_12
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A right_bottom_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
X_141_ chanx_right_in[2] chanx_left_out[3] vgnd vpwr scs8hd_buf_2
X_072_ _079_/A _070_/B _072_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_16.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _043_/A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_33_147 vgnd vpwr scs8hd_decap_12
XFILLER_18_199 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_left_track_1.LATCH_3_.latch data_in mem_left_track_1.LATCH_3_.latch/Q _086_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB _067_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__073__B _070_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_47 vgnd vpwr scs8hd_decap_12
XFILLER_23_191 vpwr vgnd scs8hd_fill_2
XFILLER_7_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A left_bottom_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
X_124_ _096_/A _120_/B _124_/Y vgnd vpwr scs8hd_nor2_4
X_055_ enable address[5] _090_/C _075_/C vgnd vpwr scs8hd_nand3_4
XFILLER_23_7 vgnd vpwr scs8hd_decap_12
XFILLER_38_239 vgnd vpwr scs8hd_decap_12
Xmem_right_track_16.LATCH_4_.latch data_in mem_right_track_16.LATCH_4_.latch/Q _077_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_206 vpwr vgnd scs8hd_fill_2
XANTENNA__068__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_12_106 vpwr vgnd scs8hd_fill_2
XFILLER_32_68 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_128 vgnd vpwr scs8hd_fill_1
XANTENNA__084__A _091_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB _098_/Y vgnd vpwr scs8hd_diode_2
XFILLER_22_90 vpwr vgnd scs8hd_fill_2
XFILLER_7_143 vgnd vpwr scs8hd_decap_6
XFILLER_11_161 vpwr vgnd scs8hd_fill_2
XFILLER_11_172 vpwr vgnd scs8hd_fill_2
XFILLER_11_194 vpwr vgnd scs8hd_fill_2
X_107_ _059_/B _111_/B _107_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_8_81 vpwr vgnd scs8hd_fill_2
XANTENNA__079__A _079_/A vgnd vpwr scs8hd_diode_2
XFILLER_40_256 vgnd vpwr scs8hd_decap_12
XFILLER_25_242 vpwr vgnd scs8hd_fill_2
XFILLER_4_168 vpwr vgnd scs8hd_fill_2
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _044_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_3_190 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__081__B _079_/B vgnd vpwr scs8hd_diode_2
XFILLER_1_138 vgnd vpwr scs8hd_decap_3
XFILLER_38_56 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_227 vgnd vpwr scs8hd_decap_4
XFILLER_13_223 vpwr vgnd scs8hd_fill_2
XFILLER_13_234 vpwr vgnd scs8hd_fill_2
XFILLER_13_245 vgnd vpwr scs8hd_decap_12
XFILLER_8_271 vgnd vpwr scs8hd_decap_4
XFILLER_5_60 vgnd vpwr scs8hd_fill_1
XFILLER_39_131 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_259 vgnd vpwr scs8hd_decap_12
XANTENNA__076__B _079_/B vgnd vpwr scs8hd_diode_2
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XANTENNA__092__A _059_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_252 vpwr vgnd scs8hd_fill_2
XFILLER_5_263 vgnd vpwr scs8hd_decap_12
XFILLER_36_178 vgnd vpwr scs8hd_decap_12
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XFILLER_19_47 vgnd vpwr scs8hd_decap_12
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_27_178 vpwr vgnd scs8hd_fill_2
XFILLER_27_156 vpwr vgnd scs8hd_fill_2
XANTENNA__087__A _079_/A vgnd vpwr scs8hd_diode_2
X_071_ _078_/A _070_/B _071_/Y vgnd vpwr scs8hd_nor2_4
X_140_ _140_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_4_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_18_134 vpwr vgnd scs8hd_fill_2
XFILLER_18_145 vgnd vpwr scs8hd_decap_4
XFILLER_18_167 vpwr vgnd scs8hd_fill_2
XFILLER_33_159 vgnd vpwr scs8hd_decap_12
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_18_178 vpwr vgnd scs8hd_fill_2
XFILLER_21_59 vpwr vgnd scs8hd_fill_2
XFILLER_30_129 vgnd vpwr scs8hd_decap_4
XFILLER_30_107 vgnd vpwr scs8hd_decap_3
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_4_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_16.INVTX1_3_.scs8hd_inv_1 chanx_left_in[7] mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_15_115 vpwr vgnd scs8hd_fill_2
XFILLER_7_39 vgnd vpwr scs8hd_decap_3
X_054_ address[1] _054_/B _060_/C _091_/A vgnd vpwr scs8hd_or3_4
X_123_ _080_/A _120_/B _123_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_14_192 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_262 vgnd vpwr scs8hd_decap_12
XANTENNA__068__C _075_/C vgnd vpwr scs8hd_diode_2
XFILLER_16_15 vgnd vpwr scs8hd_decap_12
Xmem_right_track_0.LATCH_3_.latch data_in mem_right_track_0.LATCH_3_.latch/Q _061_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__084__B _087_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_140 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB _096_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_100 vgnd vpwr scs8hd_decap_3
XFILLER_11_184 vgnd vpwr scs8hd_decap_3
X_106_ _091_/A _111_/B _106_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_19_240 vpwr vgnd scs8hd_fill_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XFILLER_8_71 vgnd vpwr scs8hd_decap_8
XFILLER_8_93 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_top_track_14.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__079__B _079_/B vgnd vpwr scs8hd_diode_2
XFILLER_25_210 vpwr vgnd scs8hd_fill_2
XFILLER_40_268 vgnd vpwr scs8hd_decap_6
XFILLER_40_213 vgnd vpwr scs8hd_fill_1
XANTENNA__095__A _080_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_14.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_210 vgnd vpwr scs8hd_decap_4
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_257 vgnd vpwr scs8hd_decap_12
XFILLER_3_180 vgnd vpwr scs8hd_fill_1
XFILLER_22_224 vgnd vpwr scs8hd_decap_8
XFILLER_1_106 vpwr vgnd scs8hd_fill_2
XFILLER_38_68 vgnd vpwr scs8hd_decap_12
XFILLER_9_217 vgnd vpwr scs8hd_fill_1
XFILLER_13_257 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_83 vpwr vgnd scs8hd_fill_2
XFILLER_39_165 vpwr vgnd scs8hd_fill_2
XANTENNA__092__B _094_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_209 vgnd vpwr scs8hd_decap_3
XFILLER_39_6 vpwr vgnd scs8hd_fill_2
XFILLER_30_80 vgnd vpwr scs8hd_fill_1
XFILLER_5_275 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A chany_top_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__087__B _087_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_070_ _059_/B _070_/B _070_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.INVTX1_2_.scs8hd_inv_1 chany_top_in[6] mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_113 vgnd vpwr scs8hd_decap_8
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XFILLER_25_91 vpwr vgnd scs8hd_fill_2
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_left_track_9.LATCH_4_.latch data_in mem_left_track_9.LATCH_4_.latch/Q _092_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ _046_/A mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_37_3 vpwr vgnd scs8hd_fill_2
XFILLER_2_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__098__A _091_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_171 vpwr vgnd scs8hd_fill_2
X_122_ _079_/A _120_/B _122_/Y vgnd vpwr scs8hd_nor2_4
X_053_ address[3] _075_/B vgnd vpwr scs8hd_inv_8
XFILLER_11_71 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
Xmem_top_track_16.LATCH_5_.latch data_in mem_top_track_16.LATCH_5_.latch/Q _119_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_274 vgnd vpwr scs8hd_decap_3
XFILLER_29_219 vpwr vgnd scs8hd_fill_2
XFILLER_32_15 vgnd vpwr scs8hd_decap_12
XFILLER_16_27 vgnd vpwr scs8hd_decap_4
Xmux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_185 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_123 vgnd vpwr scs8hd_decap_3
X_105_ address[4] address[3] address[6] _082_/X _111_/B vgnd vpwr scs8hd_or4_4
XFILLER_27_59 vpwr vgnd scs8hd_fill_2
XFILLER_27_15 vgnd vpwr scs8hd_decap_12
XANTENNA__095__B _094_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_148 vpwr vgnd scs8hd_fill_2
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_244 vgnd vpwr scs8hd_decap_4
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_269 vgnd vpwr scs8hd_decap_8
Xmux_left_track_9.INVTX1_7_.scs8hd_inv_1 left_bottom_grid_pin_13_ mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_17.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_269 vgnd vpwr scs8hd_decap_8
XFILLER_0_140 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.INVTX1_3_.scs8hd_inv_1 right_top_grid_pin_10_ mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_5_51 vgnd vpwr scs8hd_decap_3
XFILLER_5_62 vpwr vgnd scs8hd_fill_2
XFILLER_39_177 vpwr vgnd scs8hd_fill_2
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_206 vgnd vpwr scs8hd_decap_8
XFILLER_10_228 vgnd vpwr scs8hd_decap_4
Xmux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_5_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_35_15 vgnd vpwr scs8hd_decap_12
XFILLER_27_136 vgnd vpwr scs8hd_decap_3
XFILLER_27_114 vpwr vgnd scs8hd_fill_2
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XFILLER_35_59 vpwr vgnd scs8hd_fill_2
XFILLER_27_169 vpwr vgnd scs8hd_fill_2
XFILLER_2_202 vpwr vgnd scs8hd_fill_2
XFILLER_2_257 vgnd vpwr scs8hd_decap_12
XFILLER_2_246 vgnd vpwr scs8hd_decap_8
XFILLER_2_235 vgnd vpwr scs8hd_decap_8
XFILLER_2_224 vpwr vgnd scs8hd_fill_2
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XFILLER_25_70 vgnd vpwr scs8hd_fill_1
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_128 vpwr vgnd scs8hd_fill_2
XFILLER_24_106 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__098__B _103_/B vgnd vpwr scs8hd_diode_2
XFILLER_23_150 vpwr vgnd scs8hd_fill_2
X_121_ _078_/A _120_/B _121_/Y vgnd vpwr scs8hd_nor2_4
X_052_ address[4] _075_/A vgnd vpwr scs8hd_inv_8
XANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A left_bottom_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_36_80 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_253 vpwr vgnd scs8hd_fill_2
XFILLER_37_220 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.LATCH_4_.latch data_in mem_right_track_8.LATCH_4_.latch/Q _070_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_32_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_8.LATCH_3_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_28_242 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _073_/Y vgnd vpwr scs8hd_diode_2
Xmem_left_track_17.LATCH_0_.latch data_in mem_left_track_17.LATCH_0_.latch/Q _103_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_93 vpwr vgnd scs8hd_fill_2
XFILLER_7_179 vpwr vgnd scs8hd_fill_2
XFILLER_11_142 vgnd vpwr scs8hd_decap_6
Xmem_top_track_2.LATCH_0_.latch data_in _042_/A _113_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_104_ address[6] _082_/X _104_/X vgnd vpwr scs8hd_or2_4
XFILLER_14_6 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_7 vpwr vgnd scs8hd_fill_2
XFILLER_27_27 vgnd vpwr scs8hd_decap_12
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XFILLER_25_245 vgnd vpwr scs8hd_decap_12
XFILLER_25_234 vpwr vgnd scs8hd_fill_2
XFILLER_25_223 vpwr vgnd scs8hd_fill_2
XFILLER_4_127 vgnd vpwr scs8hd_decap_3
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_234 vgnd vpwr scs8hd_fill_1
XFILLER_17_82 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _127_/HI mem_left_track_9.LATCH_2_.latch/Q
+ mux_left_track_9.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB _085_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_0_152 vgnd vpwr scs8hd_fill_1
Xmux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_2_.scs8hd_inv_1/Y
+ _042_/A mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_5_96 vpwr vgnd scs8hd_fill_2
XFILLER_39_145 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB _077_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_222 vpwr vgnd scs8hd_fill_2
Xmux_right_track_16.INVTX1_4_.scs8hd_inv_1 right_bottom_grid_pin_9_ mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_left_track_17.INVTX1_5_.scs8hd_inv_1 left_bottom_grid_pin_3_ mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_35_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _132_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_269 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
XFILLER_25_60 vgnd vpwr scs8hd_fill_1
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _154_/A vgnd vpwr scs8hd_inv_1
XFILLER_32_140 vgnd vpwr scs8hd_decap_12
XFILLER_17_192 vpwr vgnd scs8hd_fill_2
XFILLER_15_107 vpwr vgnd scs8hd_fill_2
X_120_ _059_/B _120_/B _120_/Y vgnd vpwr scs8hd_nor2_4
X_051_ address[6] _090_/C vgnd vpwr scs8hd_inv_8
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _043_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _132_/HI _045_/Y mux_top_track_14.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB _101_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_232 vgnd vpwr scs8hd_decap_12
XFILLER_20_154 vpwr vgnd scs8hd_fill_2
XFILLER_28_254 vgnd vpwr scs8hd_fill_1
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
X_103_ _096_/A _103_/B _103_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_114 vpwr vgnd scs8hd_fill_2
XFILLER_11_165 vgnd vpwr scs8hd_decap_4
XFILLER_11_176 vpwr vgnd scs8hd_fill_2
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
XFILLER_19_210 vgnd vpwr scs8hd_decap_4
XFILLER_19_254 vpwr vgnd scs8hd_fill_2
XFILLER_19_276 vgnd vpwr scs8hd_fill_1
XFILLER_8_52 vpwr vgnd scs8hd_fill_2
XFILLER_8_85 vgnd vpwr scs8hd_decap_6
XFILLER_27_39 vgnd vpwr scs8hd_decap_12
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XFILLER_25_257 vgnd vpwr scs8hd_decap_12
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_172 vpwr vgnd scs8hd_fill_2
XFILLER_30_260 vgnd vpwr scs8hd_decap_12
XFILLER_13_19 vgnd vpwr scs8hd_decap_12
XFILLER_13_227 vpwr vgnd scs8hd_fill_2
XFILLER_13_238 vpwr vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ _044_/A mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_93 vgnd vpwr scs8hd_decap_3
XFILLER_12_271 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_190 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _149_/A vgnd vpwr scs8hd_inv_1
XFILLER_5_201 vpwr vgnd scs8hd_fill_2
XFILLER_14_84 vpwr vgnd scs8hd_fill_2
XFILLER_39_70 vgnd vpwr scs8hd_decap_12
XFILLER_36_105 vgnd vpwr scs8hd_decap_12
XANTENNA__101__A _079_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_35_171 vgnd vpwr scs8hd_decap_12
XFILLER_35_39 vgnd vpwr scs8hd_decap_12
XFILLER_18_138 vpwr vgnd scs8hd_fill_2
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XPHY_61 vgnd vpwr scs8hd_decap_3
XFILLER_26_182 vpwr vgnd scs8hd_fill_2
XPHY_50 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 chanx_right_in[0] mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_87 vpwr vgnd scs8hd_fill_2
XFILLER_17_182 vgnd vpwr scs8hd_fill_1
XFILLER_32_152 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_119 vgnd vpwr scs8hd_decap_3
X_050_ enable _050_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_3 vgnd vpwr scs8hd_decap_12
XFILLER_36_93 vgnd vpwr scs8hd_decap_12
XFILLER_14_196 vpwr vgnd scs8hd_fill_2
XFILLER_35_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_84 vgnd vpwr scs8hd_decap_4
X_102_ _080_/A _103_/B _102_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_34_258 vgnd vpwr scs8hd_decap_12
XFILLER_19_266 vpwr vgnd scs8hd_fill_2
XFILLER_6_192 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_40_239 vpwr vgnd scs8hd_fill_2
XFILLER_25_269 vgnd vpwr scs8hd_decap_8
XFILLER_16_225 vpwr vgnd scs8hd_fill_2
XFILLER_17_51 vgnd vpwr scs8hd_decap_8
XFILLER_17_62 vgnd vpwr scs8hd_decap_6
XFILLER_17_95 vpwr vgnd scs8hd_fill_2
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_184 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB _057_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__104__A address[6] vgnd vpwr scs8hd_diode_2
XFILLER_22_206 vgnd vpwr scs8hd_decap_6
XFILLER_30_272 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_206 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_0_187 vgnd vpwr scs8hd_decap_4
XFILLER_0_165 vpwr vgnd scs8hd_fill_2
XFILLER_8_210 vpwr vgnd scs8hd_fill_2
XFILLER_8_254 vgnd vpwr scs8hd_fill_1
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
Xmem_top_track_0.LATCH_3_.latch data_in mem_top_track_0.LATCH_3_.latch/Q _108_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_39_169 vgnd vpwr scs8hd_decap_8
XFILLER_24_19 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_5_235 vpwr vgnd scs8hd_fill_2
XFILLER_14_30 vgnd vpwr scs8hd_fill_1
XFILLER_30_84 vgnd vpwr scs8hd_decap_8
XFILLER_39_82 vgnd vpwr scs8hd_decap_12
XFILLER_36_117 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__101__B _103_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 chanx_left_in[6] mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_73 vpwr vgnd scs8hd_fill_2
XFILLER_25_62 vpwr vgnd scs8hd_fill_2
XFILLER_25_51 vgnd vpwr scs8hd_decap_6
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_37_7 vgnd vpwr scs8hd_decap_12
XFILLER_2_55 vgnd vpwr scs8hd_decap_8
XFILLER_2_44 vgnd vpwr scs8hd_decap_8
XANTENNA__112__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_17_172 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _123_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_175 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_top_track_16.LATCH_0_.latch data_in mem_top_track_16.LATCH_0_.latch/Q _124_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XANTENNA__107__A _059_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_245 vgnd vpwr scs8hd_decap_8
XFILLER_28_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A right_bottom_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
Xmux_top_track_14.INVTX1_0_.scs8hd_inv_1 chanx_left_in[2] mux_top_track_14.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_20_145 vgnd vpwr scs8hd_decap_8
XFILLER_20_189 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_212 vpwr vgnd scs8hd_fill_2
X_101_ _079_/A _103_/B _101_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_11_134 vpwr vgnd scs8hd_fill_2
XFILLER_22_74 vgnd vpwr scs8hd_fill_1
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
XFILLER_40_207 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB _108_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_4_.scs8hd_inv_1 chanx_right_in[5] mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmem_left_track_1.LATCH_4_.latch data_in mem_left_track_1.LATCH_4_.latch/Q _085_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_270 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_16_215 vgnd vpwr scs8hd_fill_1
XFILLER_16_248 vgnd vpwr scs8hd_fill_1
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_62 vgnd vpwr scs8hd_decap_12
XFILLER_33_51 vgnd vpwr scs8hd_decap_8
XANTENNA__104__B _082_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _059_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_3_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_15_270 vgnd vpwr scs8hd_decap_6
Xmem_right_track_16.LATCH_5_.latch data_in mem_right_track_16.LATCH_5_.latch/Q _076_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmux_right_track_0.INVTX1_0_.scs8hd_inv_1 chany_top_in[2] mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_240 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A chany_top_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_0_111 vpwr vgnd scs8hd_fill_2
XFILLER_0_144 vpwr vgnd scs8hd_fill_2
XFILLER_28_84 vpwr vgnd scs8hd_fill_2
XFILLER_0_177 vpwr vgnd scs8hd_fill_2
XANTENNA__115__A _075_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_66 vpwr vgnd scs8hd_fill_2
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A right_bottom_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB _091_/Y vgnd vpwr scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _135_/HI _043_/Y mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_39_94 vgnd vpwr scs8hd_decap_12
XFILLER_36_129 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _044_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_228 vgnd vpwr scs8hd_decap_4
XFILLER_2_206 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_0.INVTX1_4_.scs8hd_inv_1 chanx_left_in[3] mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_30 vgnd vpwr scs8hd_decap_3
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_67 vgnd vpwr scs8hd_decap_4
XANTENNA__112__B _075_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
XFILLER_32_121 vgnd vpwr scs8hd_decap_12
XFILLER_17_151 vpwr vgnd scs8hd_fill_2
XFILLER_17_184 vpwr vgnd scs8hd_fill_2
XFILLER_23_187 vpwr vgnd scs8hd_fill_2
XFILLER_23_154 vpwr vgnd scs8hd_fill_2
XFILLER_23_132 vgnd vpwr scs8hd_decap_3
XFILLER_11_98 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_5_.scs8hd_inv_1 right_bottom_grid_pin_13_ mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_110 vgnd vpwr scs8hd_decap_6
XFILLER_14_132 vgnd vpwr scs8hd_decap_4
XFILLER_14_154 vpwr vgnd scs8hd_fill_2
XANTENNA__107__B _111_/B vgnd vpwr scs8hd_diode_2
XANTENNA__123__A _080_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_102 vpwr vgnd scs8hd_fill_2
XFILLER_20_168 vgnd vpwr scs8hd_decap_8
X_100_ _078_/A _103_/B _100_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_128 vpwr vgnd scs8hd_fill_2
XFILLER_11_102 vpwr vgnd scs8hd_fill_2
XFILLER_22_97 vgnd vpwr scs8hd_decap_4
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A address[4] vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_10_190 vgnd vpwr scs8hd_decap_4
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_238 vpwr vgnd scs8hd_fill_2
XFILLER_25_227 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB _088_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _046_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_1.INVTX1_7_.scs8hd_inv_1 left_bottom_grid_pin_11_ mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_153 vpwr vgnd scs8hd_fill_2
XANTENNA__120__B _120_/B vgnd vpwr scs8hd_diode_2
XFILLER_38_19 vgnd vpwr scs8hd_decap_12
XFILLER_21_252 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB _080_/Y vgnd vpwr scs8hd_diode_2
XFILLER_28_74 vgnd vpwr scs8hd_fill_1
Xmem_right_track_0.LATCH_4_.latch data_in mem_right_track_0.LATCH_4_.latch/Q _059_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__115__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_5_56 vpwr vgnd scs8hd_fill_2
XFILLER_39_149 vgnd vpwr scs8hd_decap_12
XFILLER_39_127 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__041__A _041_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.INVTX1_2_.scs8hd_inv_1 chany_top_in[7] mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_43 vpwr vgnd scs8hd_fill_2
XFILLER_14_54 vgnd vpwr scs8hd_decap_12
XFILLER_5_248 vpwr vgnd scs8hd_fill_2
XFILLER_5_259 vpwr vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 _133_/HI mem_top_track_16.LATCH_5_.latch/Q
+ mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_29_182 vgnd vpwr scs8hd_fill_1
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_64 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vpwr scs8hd_diode_2
XPHY_53 vgnd vpwr scs8hd_decap_3
Xmux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_5_.latch/Q mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__112__C _104_/X vgnd vpwr scs8hd_diode_2
XFILLER_32_166 vgnd vpwr scs8hd_decap_12
XFILLER_32_133 vgnd vpwr scs8hd_decap_4
XFILLER_17_196 vpwr vgnd scs8hd_fill_2
XFILLER_23_100 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_77 vpwr vgnd scs8hd_fill_2
XANTENNA__123__B _120_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_37_258 vpwr vgnd scs8hd_fill_2
XFILLER_20_125 vgnd vpwr scs8hd_decap_4
XFILLER_20_158 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_225 vgnd vpwr scs8hd_decap_8
XFILLER_11_114 vpwr vgnd scs8hd_fill_2
XFILLER_22_32 vgnd vpwr scs8hd_decap_12
XFILLER_7_118 vpwr vgnd scs8hd_fill_2
XFILLER_0_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XFILLER_19_225 vpwr vgnd scs8hd_fill_2
XFILLER_19_236 vpwr vgnd scs8hd_fill_2
XFILLER_19_258 vgnd vpwr scs8hd_decap_4
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XFILLER_8_56 vpwr vgnd scs8hd_fill_2
XANTENNA__118__B address[3] vgnd vpwr scs8hd_diode_2
X_159_ chanx_right_in[5] chany_top_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_6_173 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_33_3 vgnd vpwr scs8hd_decap_12
XFILLER_25_206 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_5_.latch data_in mem_left_track_9.LATCH_5_.latch/Q _091_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__044__A _044_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _126_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_16_206 vpwr vgnd scs8hd_fill_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_86 vgnd vpwr scs8hd_decap_12
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_132 vpwr vgnd scs8hd_fill_2
XFILLER_3_176 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_2.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_224 vpwr vgnd scs8hd_fill_2
XFILLER_8_235 vgnd vpwr scs8hd_decap_8
XFILLER_8_246 vgnd vpwr scs8hd_decap_8
XANTENNA__115__C _104_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_79 vpwr vgnd scs8hd_fill_2
XFILLER_39_139 vpwr vgnd scs8hd_fill_2
XFILLER_39_106 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_66 vgnd vpwr scs8hd_fill_1
XFILLER_14_88 vpwr vgnd scs8hd_fill_2
XFILLER_30_32 vgnd vpwr scs8hd_decap_12
XFILLER_5_205 vpwr vgnd scs8hd_fill_2
XFILLER_39_41 vgnd vpwr scs8hd_decap_12
XFILLER_29_172 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ _046_/Y mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__142__A chanx_right_in[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__052__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_26_186 vgnd vpwr scs8hd_decap_6
XPHY_54 vgnd vpwr scs8hd_decap_3
XFILLER_25_87 vpwr vgnd scs8hd_fill_2
XPHY_43 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
XFILLER_1_263 vgnd vpwr scs8hd_decap_12
XFILLER_1_252 vpwr vgnd scs8hd_fill_2
XANTENNA__112__D _060_/C vgnd vpwr scs8hd_diode_2
XFILLER_32_178 vgnd vpwr scs8hd_decap_12
XANTENNA__137__A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_167 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _130_/HI mem_right_track_8.LATCH_2_.latch/Q
+ mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__047__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_145 vgnd vpwr scs8hd_decap_6
XFILLER_14_167 vgnd vpwr scs8hd_decap_12
XFILLER_9_193 vpwr vgnd scs8hd_fill_2
XFILLER_28_259 vgnd vpwr scs8hd_decap_12
XFILLER_28_215 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_44 vgnd vpwr scs8hd_decap_12
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
XFILLER_8_46 vpwr vgnd scs8hd_fill_2
XANTENNA__118__C _075_/C vgnd vpwr scs8hd_diode_2
X_158_ _158_/A chany_top_out[4] vgnd vpwr scs8hd_buf_2
X_089_ _096_/A _087_/B _089_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_26_3 vgnd vpwr scs8hd_decap_12
XANTENNA__150__A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_18_270 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB _063_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__060__A _060_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_229 vgnd vpwr scs8hd_decap_3
XFILLER_17_99 vpwr vgnd scs8hd_fill_2
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_98 vgnd vpwr scs8hd_decap_12
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_166 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__145__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XFILLER_21_276 vgnd vpwr scs8hd_fill_1
XFILLER_0_91 vpwr vgnd scs8hd_fill_2
XANTENNA__055__A enable vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_32 vgnd vpwr scs8hd_decap_12
Xmem_right_track_8.LATCH_5_.latch data_in mem_right_track_8.LATCH_5_.latch/Q _069_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_125 vgnd vpwr scs8hd_decap_4
XFILLER_0_169 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__115__D address[0] vgnd vpwr scs8hd_diode_2
Xmux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _041_/A mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XFILLER_39_118 vgnd vpwr scs8hd_decap_4
Xmem_top_track_2.LATCH_1_.latch data_in _041_/A _112_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_left_track_17.LATCH_1_.latch data_in mem_left_track_17.LATCH_1_.latch/Q _102_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_0.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_30_44 vgnd vpwr scs8hd_decap_12
XFILLER_5_239 vgnd vpwr scs8hd_decap_3
XFILLER_39_53 vgnd vpwr scs8hd_decap_8
XFILLER_29_184 vgnd vpwr scs8hd_decap_12
XFILLER_29_151 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _129_/HI mem_right_track_16.LATCH_2_.latch/Q
+ mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_35_110 vgnd vpwr scs8hd_decap_12
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_165 vgnd vpwr scs8hd_decap_8
XFILLER_25_77 vgnd vpwr scs8hd_fill_1
XFILLER_25_66 vgnd vpwr scs8hd_decap_4
XPHY_44 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
XFILLER_2_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A left_bottom_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_17_132 vpwr vgnd scs8hd_fill_2
XANTENNA__153__A _153_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_179 vpwr vgnd scs8hd_fill_2
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XANTENNA__063__A _067_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_32 vgnd vpwr scs8hd_decap_12
XFILLER_14_102 vpwr vgnd scs8hd_fill_2
XFILLER_14_179 vgnd vpwr scs8hd_decap_4
XANTENNA__148__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_9_172 vgnd vpwr scs8hd_decap_4
XANTENNA__058__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_138 vpwr vgnd scs8hd_fill_2
XFILLER_22_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
X_157_ chanx_left_in[5] chany_top_out[5] vgnd vpwr scs8hd_buf_2
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_6_186 vgnd vpwr scs8hd_decap_4
X_088_ _080_/A _087_/B _088_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__060__B address[2] vgnd vpwr scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_78 vpwr vgnd scs8hd_fill_2
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_274 vgnd vpwr scs8hd_fill_1
Xmem_right_track_16.LATCH_0_.latch data_in mem_right_track_16.LATCH_0_.latch/Q _081_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_3_112 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 _134_/HI _042_/Y mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_30_200 vgnd vpwr scs8hd_decap_12
XFILLER_15_241 vgnd vpwr scs8hd_fill_1
XANTENNA__161__A _161_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _043_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA__055__B address[5] vgnd vpwr scs8hd_diode_2
XANTENNA__071__A _078_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_115 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_28_88 vgnd vpwr scs8hd_decap_4
XFILLER_28_44 vgnd vpwr scs8hd_decap_12
XFILLER_0_148 vgnd vpwr scs8hd_decap_4
XFILLER_5_15 vgnd vpwr scs8hd_decap_12
XFILLER_8_259 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB _094_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__156__A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_38_141 vgnd vpwr scs8hd_decap_12
XANTENNA__066__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_14_35 vgnd vpwr scs8hd_decap_8
XFILLER_30_56 vgnd vpwr scs8hd_decap_12
XFILLER_5_218 vpwr vgnd scs8hd_fill_2
XFILLER_39_10 vgnd vpwr scs8hd_decap_12
XFILLER_29_196 vgnd vpwr scs8hd_decap_3
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_26_122 vpwr vgnd scs8hd_fill_2
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
XPHY_56 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XFILLER_2_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_232 vpwr vgnd scs8hd_fill_2
XFILLER_17_155 vpwr vgnd scs8hd_fill_2
XFILLER_17_188 vgnd vpwr scs8hd_fill_1
Xmux_right_track_8.INVTX1_2_.scs8hd_inv_1 chany_top_in[6] mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_114 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _045_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__063__B _079_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_44 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_106 vpwr vgnd scs8hd_fill_2
XFILLER_3_70 vpwr vgnd scs8hd_fill_2
XFILLER_28_206 vgnd vpwr scs8hd_decap_4
XANTENNA__058__B _054_/B vgnd vpwr scs8hd_diode_2
XANTENNA__074__A _096_/A vgnd vpwr scs8hd_diode_2
XFILLER_11_106 vgnd vpwr scs8hd_decap_3
XFILLER_22_68 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_9.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_19_206 vpwr vgnd scs8hd_fill_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
X_156_ chanx_left_in[4] chany_top_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_6_165 vgnd vpwr scs8hd_decap_8
Xmux_left_track_1.INVTX1_4_.scs8hd_inv_1 chanx_right_in[4] mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_194 vgnd vpwr scs8hd_fill_1
X_087_ _079_/A _087_/B _087_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__159__A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_33_220 vgnd vpwr scs8hd_decap_12
XFILLER_33_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__069__A _091_/A vgnd vpwr scs8hd_diode_2
XANTENNA__060__C _060_/C vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_68 vgnd vpwr scs8hd_fill_1
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ _044_/Y mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_212 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_139_ chanx_right_in[4] chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_31_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_190 vgnd vpwr scs8hd_decap_4
XFILLER_21_212 vpwr vgnd scs8hd_fill_2
XFILLER_0_71 vgnd vpwr scs8hd_decap_3
XFILLER_21_256 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _125_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__055__C _090_/C vgnd vpwr scs8hd_diode_2
XANTENNA__071__B _070_/B vgnd vpwr scs8hd_diode_2
XFILLER_28_56 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A _134_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A chany_top_in[6] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__066__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_14_69 vgnd vpwr scs8hd_fill_1
XFILLER_30_68 vgnd vpwr scs8hd_decap_12
XANTENNA__082__A _050_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_66 vpwr vgnd scs8hd_fill_2
XFILLER_39_22 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_263 vgnd vpwr scs8hd_decap_12
XFILLER_4_252 vgnd vpwr scs8hd_decap_8
XFILLER_4_241 vgnd vpwr scs8hd_decap_8
XFILLER_20_90 vpwr vgnd scs8hd_fill_2
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_26_145 vgnd vpwr scs8hd_decap_6
XFILLER_26_134 vpwr vgnd scs8hd_fill_2
XFILLER_26_112 vgnd vpwr scs8hd_fill_1
XPHY_46 vgnd vpwr scs8hd_decap_3
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XPHY_35 vgnd vpwr scs8hd_decap_3
XANTENNA__077__A _059_/B vgnd vpwr scs8hd_diode_2
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_25_57 vgnd vpwr scs8hd_fill_1
XFILLER_32_137 vgnd vpwr scs8hd_fill_1
XFILLER_15_90 vpwr vgnd scs8hd_fill_2
XFILLER_23_104 vgnd vpwr scs8hd_decap_4
Xmux_right_track_0.INVTX1_5_.scs8hd_inv_1 right_bottom_grid_pin_11_ mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_137 vpwr vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_4_.latch data_in mem_top_track_0.LATCH_4_.latch/Q _107_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_14.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_3_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_36_56 vgnd vpwr scs8hd_decap_12
XFILLER_22_192 vgnd vpwr scs8hd_fill_1
XFILLER_9_152 vgnd vpwr scs8hd_decap_4
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
XANTENNA__058__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__074__B _070_/B vgnd vpwr scs8hd_diode_2
XFILLER_11_118 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_0_.latch data_in mem_left_track_9.LATCH_0_.latch/Q _096_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__090__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_19_229 vpwr vgnd scs8hd_fill_2
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
X_155_ _155_/A chany_top_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_6_111 vgnd vpwr scs8hd_decap_4
X_086_ _078_/A _087_/B _086_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_12_80 vgnd vpwr scs8hd_fill_1
XFILLER_33_232 vgnd vpwr scs8hd_decap_12
XANTENNA__069__B _070_/B vgnd vpwr scs8hd_diode_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
Xmux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__085__A _059_/B vgnd vpwr scs8hd_diode_2
XFILLER_3_136 vpwr vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_1_.latch data_in mem_top_track_16.LATCH_1_.latch/Q _123_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_210 vpwr vgnd scs8hd_fill_2
XFILLER_30_224 vgnd vpwr scs8hd_decap_12
XFILLER_15_254 vpwr vgnd scs8hd_fill_2
XFILLER_15_276 vgnd vpwr scs8hd_fill_1
X_069_ _091_/A _070_/B _069_/Y vgnd vpwr scs8hd_nor2_4
X_138_ chanx_right_in[5] chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_0_94 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_top_track_16.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_268 vgnd vpwr scs8hd_decap_8
XFILLER_9_81 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_2_.latch/Q mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_28_68 vgnd vpwr scs8hd_decap_6
XFILLER_8_206 vpwr vgnd scs8hd_fill_2
XFILLER_8_228 vgnd vpwr scs8hd_decap_4
XFILLER_12_213 vgnd vpwr scs8hd_fill_1
XFILLER_12_224 vpwr vgnd scs8hd_fill_2
XFILLER_12_235 vgnd vpwr scs8hd_decap_12
XFILLER_5_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB _071_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[8] vgnd vpwr scs8hd_diode_2
XANTENNA__066__C address[0] vgnd vpwr scs8hd_diode_2
XANTENNA__082__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_29_176 vgnd vpwr scs8hd_decap_6
Xmem_left_track_1.LATCH_5_.latch data_in mem_left_track_1.LATCH_5_.latch/Q _084_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_35_135 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_3_.latch/Q mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_71 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _162_/A vgnd vpwr scs8hd_inv_1
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XANTENNA__077__B _079_/B vgnd vpwr scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA__093__A _078_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_105 vgnd vpwr scs8hd_decap_12
XFILLER_17_168 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_31_182 vgnd vpwr scs8hd_fill_1
XFILLER_11_27 vgnd vpwr scs8hd_decap_12
XANTENNA__088__A _080_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_68 vgnd vpwr scs8hd_decap_12
XFILLER_14_116 vgnd vpwr scs8hd_fill_1
XFILLER_22_182 vpwr vgnd scs8hd_fill_2
XFILLER_37_208 vgnd vpwr scs8hd_decap_12
XFILLER_20_119 vgnd vpwr scs8hd_decap_4
XFILLER_9_197 vpwr vgnd scs8hd_fill_2
XFILLER_3_83 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.INVTX1_7_.scs8hd_inv_1 left_bottom_grid_pin_15_ mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
Xmux_right_track_16.INVTX1_6_.scs8hd_inv_1 chanx_left_in[2] mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
XFILLER_22_15 vgnd vpwr scs8hd_decap_12
XANTENNA__090__B _075_/B vgnd vpwr scs8hd_diode_2
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_27_252 vgnd vpwr scs8hd_decap_3
XFILLER_27_241 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_17.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_152 vgnd vpwr scs8hd_fill_1
X_154_ _154_/A chany_top_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_6_134 vpwr vgnd scs8hd_fill_2
XFILLER_6_145 vpwr vgnd scs8hd_fill_2
X_085_ _059_/B _087_/B _085_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_9.LATCH_4_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vpwr scs8hd_ebufn_2
XFILLER_18_241 vgnd vpwr scs8hd_decap_4
XFILLER_18_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_211 vgnd vpwr scs8hd_fill_1
XFILLER_17_15 vgnd vpwr scs8hd_decap_12
XFILLER_17_59 vpwr vgnd scs8hd_fill_2
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A right_top_grid_pin_10_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA__085__B _087_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
Xmem_right_track_8.LATCH_0_.latch data_in mem_right_track_8.LATCH_0_.latch/Q _074_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_233 vpwr vgnd scs8hd_fill_2
XFILLER_15_266 vpwr vgnd scs8hd_fill_2
XFILLER_30_236 vgnd vpwr scs8hd_decap_12
Xmux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_137_ chanx_right_in[6] chanx_left_out[7] vgnd vpwr scs8hd_buf_2
X_068_ _075_/A address[3] _075_/C _070_/B vgnd vpwr scs8hd_or3_4
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
XFILLER_21_236 vpwr vgnd scs8hd_fill_2
XFILLER_21_225 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _114_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_71 vgnd vpwr scs8hd_decap_4
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _136_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB _099_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A right_bottom_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__096__A _096_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_203 vpwr vgnd scs8hd_fill_2
XFILLER_12_247 vgnd vpwr scs8hd_decap_12
Xmux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_18_80 vgnd vpwr scs8hd_fill_1
Xmux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_1_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_38_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_30_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_210 vpwr vgnd scs8hd_fill_2
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_147 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_14.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _046_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _140_/A vgnd vpwr scs8hd_inv_1
XFILLER_6_50 vgnd vpwr scs8hd_decap_6
XPHY_59 vgnd vpwr scs8hd_decap_3
XFILLER_25_15 vgnd vpwr scs8hd_decap_12
XPHY_48 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XANTENNA__093__B _094_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_202 vpwr vgnd scs8hd_fill_2
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_136 vpwr vgnd scs8hd_fill_2
XFILLER_40_183 vgnd vpwr scs8hd_decap_12
XFILLER_32_117 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_right_track_8.LATCH_2_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_right_track_0.LATCH_5_.latch data_in mem_right_track_0.LATCH_5_.latch/Q _057_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_39 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_left_track_1.LATCH_4_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__088__B _087_/B vgnd vpwr scs8hd_diode_2
XFILLER_14_106 vpwr vgnd scs8hd_fill_2
XFILLER_14_128 vpwr vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_9_132 vgnd vpwr scs8hd_decap_4
XFILLER_9_176 vgnd vpwr scs8hd_fill_1
XFILLER_3_62 vgnd vpwr scs8hd_fill_1
XFILLER_3_51 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_27 vgnd vpwr scs8hd_decap_4
XANTENNA__090__C _090_/C vgnd vpwr scs8hd_diode_2
XANTENNA__099__A _059_/B vgnd vpwr scs8hd_diode_2
XFILLER_6_102 vgnd vpwr scs8hd_decap_3
XFILLER_10_175 vgnd vpwr scs8hd_decap_8
XFILLER_10_186 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_2.INVTX1_0_.scs8hd_inv_1/Y
+ _042_/A mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
X_153_ _153_/A chanx_right_out[0] vgnd vpwr scs8hd_buf_2
X_084_ _091_/A _087_/B _084_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_19_7 vpwr vgnd scs8hd_fill_2
XFILLER_33_245 vgnd vpwr scs8hd_decap_8
Xmux_top_track_16.INVTX1_2_.scs8hd_inv_1 chanx_left_in[1] mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_234 vgnd vpwr scs8hd_decap_12
XFILLER_17_27 vgnd vpwr scs8hd_decap_12
XFILLER_33_59 vpwr vgnd scs8hd_fill_2
XFILLER_33_15 vgnd vpwr scs8hd_decap_12
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _129_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_149 vpwr vgnd scs8hd_fill_2
XFILLER_3_116 vgnd vpwr scs8hd_decap_4
XFILLER_30_215 vgnd vpwr scs8hd_decap_6
X_136_ _136_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XFILLER_30_248 vgnd vpwr scs8hd_decap_12
XFILLER_23_81 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_067_ _067_/A _096_/A _067_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_85 vgnd vpwr scs8hd_decap_4
XFILLER_21_248 vpwr vgnd scs8hd_fill_2
XFILLER_9_94 vgnd vpwr scs8hd_decap_4
XFILLER_28_15 vgnd vpwr scs8hd_decap_12
XFILLER_0_119 vgnd vpwr scs8hd_decap_3
XANTENNA__096__B _094_/B vgnd vpwr scs8hd_diode_2
XFILLER_12_259 vgnd vpwr scs8hd_decap_12
XFILLER_20_270 vgnd vpwr scs8hd_decap_4
XFILLER_34_80 vgnd vpwr scs8hd_decap_12
XFILLER_7_252 vpwr vgnd scs8hd_fill_2
XFILLER_7_263 vpwr vgnd scs8hd_fill_2
X_119_ _091_/A _120_/B _119_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_178 vgnd vpwr scs8hd_decap_12
XFILLER_30_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_29_134 vpwr vgnd scs8hd_fill_2
XFILLER_29_123 vpwr vgnd scs8hd_fill_2
XFILLER_29_101 vpwr vgnd scs8hd_fill_2
XFILLER_35_159 vgnd vpwr scs8hd_decap_12
XFILLER_6_84 vpwr vgnd scs8hd_fill_2
XFILLER_26_126 vgnd vpwr scs8hd_decap_6
XFILLER_26_104 vpwr vgnd scs8hd_fill_2
XFILLER_25_27 vgnd vpwr scs8hd_decap_12
XPHY_49 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_38 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XFILLER_1_236 vgnd vpwr scs8hd_decap_6
XFILLER_40_195 vgnd vpwr scs8hd_decap_12
XFILLER_23_118 vpwr vgnd scs8hd_fill_2
XFILLER_31_184 vgnd vpwr scs8hd_decap_12
XFILLER_31_162 vgnd vpwr scs8hd_decap_12
XFILLER_39_262 vgnd vpwr scs8hd_decap_12
XFILLER_39_240 vgnd vpwr scs8hd_fill_1
XFILLER_36_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _128_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _042_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_100 vpwr vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_184 vgnd vpwr scs8hd_decap_3
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__090__D _082_/X vgnd vpwr scs8hd_diode_2
XANTENNA__099__B _103_/B vgnd vpwr scs8hd_diode_2
XFILLER_10_154 vpwr vgnd scs8hd_fill_2
X_083_ address[4] address[3] _090_/C _082_/X _087_/B vgnd vpwr scs8hd_or4_4
X_152_ chanx_left_in[0] chanx_right_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_12_83 vgnd vpwr scs8hd_decap_3
XFILLER_18_210 vpwr vgnd scs8hd_fill_2
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
XFILLER_33_257 vgnd vpwr scs8hd_decap_12
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_246 vgnd vpwr scs8hd_decap_12
XFILLER_24_224 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB _121_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_39 vgnd vpwr scs8hd_decap_12
XFILLER_33_27 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_5_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_135_ _135_/HI _135_/LO vgnd vpwr scs8hd_conb_1
X_066_ address[1] address[2] address[0] _096_/A vgnd vpwr scs8hd_or3_4
XANTENNA_mem_top_track_0.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_172 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_28_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_93 vpwr vgnd scs8hd_fill_2
X_049_ address[0] _060_/C vgnd vpwr scs8hd_inv_8
XFILLER_7_275 vpwr vgnd scs8hd_fill_2
X_118_ address[4] address[3] _075_/C _120_/B vgnd vpwr scs8hd_or3_4
XFILLER_22_3 vgnd vpwr scs8hd_decap_12
XFILLER_14_18 vgnd vpwr scs8hd_decap_12
XFILLER_39_37 vpwr vgnd scs8hd_fill_2
XFILLER_29_168 vpwr vgnd scs8hd_fill_2
XFILLER_29_157 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB _106_/Y vgnd vpwr scs8hd_diode_2
Xmux_left_track_9.INVTX1_6_.scs8hd_inv_1 left_bottom_grid_pin_7_ mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XFILLER_25_39 vgnd vpwr scs8hd_decap_12
XPHY_39 vgnd vpwr scs8hd_decap_3
Xmux_right_track_0.INVTX1_2_.scs8hd_inv_1 chany_top_in[8] mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_215 vpwr vgnd scs8hd_fill_2
XFILLER_9_7 vpwr vgnd scs8hd_fill_2
XFILLER_1_259 vpwr vgnd scs8hd_fill_2
XFILLER_1_248 vpwr vgnd scs8hd_fill_2
XFILLER_40_141 vgnd vpwr scs8hd_decap_12
XFILLER_15_94 vpwr vgnd scs8hd_fill_2
XFILLER_31_174 vgnd vpwr scs8hd_decap_8
XFILLER_23_108 vgnd vpwr scs8hd_fill_1
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
XFILLER_39_274 vgnd vpwr scs8hd_decap_3
XFILLER_36_27 vgnd vpwr scs8hd_decap_4
Xmem_left_track_17.LATCH_2_.latch data_in mem_left_track_17.LATCH_2_.latch/Q _101_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_141 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_152 vpwr vgnd scs8hd_fill_2
XFILLER_9_156 vgnd vpwr scs8hd_fill_1
XFILLER_27_233 vpwr vgnd scs8hd_fill_2
XFILLER_27_222 vpwr vgnd scs8hd_fill_2
X_151_ chanx_left_in[1] chanx_right_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_10_111 vgnd vpwr scs8hd_decap_4
XFILLER_10_133 vpwr vgnd scs8hd_fill_2
XFILLER_10_144 vgnd vpwr scs8hd_decap_6
XFILLER_12_40 vgnd vpwr scs8hd_decap_4
X_082_ _050_/Y address[5] _082_/X vgnd vpwr scs8hd_or2_4
XFILLER_33_269 vgnd vpwr scs8hd_decap_8
XFILLER_33_39 vgnd vpwr scs8hd_decap_12
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_258 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _125_/HI mem_left_track_1.LATCH_2_.latch/Q
+ mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_15_214 vpwr vgnd scs8hd_fill_2
Xmux_top_track_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ _041_/Y mux_top_track_2.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_15_258 vpwr vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_7_.scs8hd_inv_1 chanx_left_in[5] mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_134_ _134_/HI _134_/LO vgnd vpwr scs8hd_conb_1
X_065_ _067_/A _080_/A _065_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_7 vgnd vpwr scs8hd_decap_12
XFILLER_0_32 vgnd vpwr scs8hd_decap_8
XFILLER_0_43 vpwr vgnd scs8hd_fill_2
XFILLER_0_54 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _074_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_41 vgnd vpwr scs8hd_fill_1
XFILLER_12_228 vgnd vpwr scs8hd_decap_4
XFILLER_34_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
X_117_ _075_/A _075_/B _104_/X address[0] _117_/Y vgnd vpwr scs8hd_nor4_4
X_048_ address[2] _054_/B vgnd vpwr scs8hd_inv_8
Xmem_left_track_1.LATCH_0_.latch data_in mem_left_track_1.LATCH_0_.latch/Q _089_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_15_3 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_29_114 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB _086_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_224 vpwr vgnd scs8hd_fill_2
XFILLER_4_202 vgnd vpwr scs8hd_decap_6
XFILLER_20_73 vpwr vgnd scs8hd_fill_2
XFILLER_20_84 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_29_93 vpwr vgnd scs8hd_fill_2
Xmem_right_track_16.LATCH_1_.latch data_in mem_right_track_16.LATCH_1_.latch/Q _080_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_15_51 vgnd vpwr scs8hd_decap_8
XFILLER_15_62 vpwr vgnd scs8hd_fill_2
XFILLER_15_73 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB _078_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__102__A _080_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_131 vgnd vpwr scs8hd_decap_4
XFILLER_31_120 vpwr vgnd scs8hd_fill_2
XFILLER_39_253 vpwr vgnd scs8hd_fill_2
XFILLER_39_220 vgnd vpwr scs8hd_decap_8
Xmux_left_track_17.INVTX1_4_.scs8hd_inv_1 chanx_right_in[6] mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_22_186 vgnd vpwr scs8hd_decap_6
Xmux_right_track_16.INVTX1_3_.scs8hd_inv_1 right_bottom_grid_pin_3_ mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_179 vpwr vgnd scs8hd_fill_2
XFILLER_3_87 vpwr vgnd scs8hd_fill_2
XFILLER_10_101 vgnd vpwr scs8hd_fill_1
X_150_ chanx_left_in[2] chanx_right_out[3] vgnd vpwr scs8hd_buf_2
X_081_ _096_/A _079_/B _081_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_149 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_12_63 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_3_108 vpwr vgnd scs8hd_fill_2
XFILLER_15_237 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB _102_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_62 vgnd vpwr scs8hd_decap_12
X_133_ _133_/HI _133_/LO vgnd vpwr scs8hd_conb_1
Xmux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_0_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
X_064_ address[1] address[2] _060_/C _080_/A vgnd vpwr scs8hd_or3_4
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_163 vgnd vpwr scs8hd_decap_3
XFILLER_2_130 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_14.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _045_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_2_196 vpwr vgnd scs8hd_fill_2
XANTENNA__110__A _080_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_229 vpwr vgnd scs8hd_fill_2
XFILLER_9_53 vpwr vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_207 vgnd vpwr scs8hd_decap_6
XFILLER_18_84 vpwr vgnd scs8hd_fill_2
X_116_ _075_/A _075_/B _104_/X _060_/C _116_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_7_211 vgnd vpwr scs8hd_decap_4
XANTENNA__105__A address[4] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_5_.latch_D data_in vgnd vpwr scs8hd_diode_2
X_047_ address[1] _060_/A vgnd vpwr scs8hd_inv_8
XFILLER_29_83 vgnd vpwr scs8hd_fill_1
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XPHY_19 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
Xmem_top_track_8.LATCH_0_.latch data_in _044_/A _115_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
Xmem_right_track_0.LATCH_0_.latch data_in mem_right_track_0.LATCH_0_.latch/Q _067_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_195 vpwr vgnd scs8hd_fill_2
XFILLER_31_62 vgnd vpwr scs8hd_decap_12
XFILLER_31_51 vgnd vpwr scs8hd_decap_8
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA__102__B _103_/B vgnd vpwr scs8hd_diode_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_243 vgnd vpwr scs8hd_fill_1
XFILLER_22_165 vgnd vpwr scs8hd_decap_8
XFILLER_26_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_3_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_4_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_9_114 vpwr vgnd scs8hd_fill_2
XFILLER_9_136 vgnd vpwr scs8hd_fill_1
XFILLER_13_121 vgnd vpwr scs8hd_fill_1
XFILLER_13_132 vgnd vpwr scs8hd_decap_4
XFILLER_13_165 vpwr vgnd scs8hd_fill_2
XFILLER_13_198 vgnd vpwr scs8hd_decap_6
XANTENNA__113__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_36_202 vgnd vpwr scs8hd_decap_12
XFILLER_3_66 vpwr vgnd scs8hd_fill_2
XFILLER_27_257 vgnd vpwr scs8hd_decap_12
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
X_080_ _080_/A _079_/B _080_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_128 vgnd vpwr scs8hd_decap_4
Xmux_right_track_0.tap_buf4_0_.scs8hd_inv_1 mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _153_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_18_202 vgnd vpwr scs8hd_fill_1
XFILLER_18_224 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__108__A _078_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_205 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_top_track_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_2.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_227 vgnd vpwr scs8hd_decap_4
XFILLER_23_85 vpwr vgnd scs8hd_fill_2
XFILLER_23_74 vgnd vpwr scs8hd_decap_4
X_132_ _132_/HI _132_/LO vgnd vpwr scs8hd_conb_1
Xmem_top_track_0.LATCH_5_.latch data_in mem_top_track_0.LATCH_5_.latch/Q _106_/Y vgnd
+ vpwr scs8hd_lpflow_inputisolatch_1
X_063_ _067_/A _079_/A _063_/Y vgnd vpwr scs8hd_nor2_4
Xmux_right_track_16.tap_buf4_0_.scs8hd_inv_1 mux_right_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _145_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_67 vpwr vgnd scs8hd_fill_2
XANTENNA__110__B _111_/B vgnd vpwr scs8hd_diode_2
XFILLER_21_208 vpwr vgnd scs8hd_fill_2
XFILLER_14_271 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_20_274 vgnd vpwr scs8hd_fill_1
XFILLER_11_230 vgnd vpwr scs8hd_decap_12
X_046_ _046_/A _046_/Y vgnd vpwr scs8hd_inv_8
X_115_ _075_/A address[3] _104_/X address[0] _115_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_7_201 vgnd vpwr scs8hd_fill_1
XFILLER_7_234 vpwr vgnd scs8hd_fill_2
XFILLER_7_267 vgnd vpwr scs8hd_decap_8
XFILLER_11_263 vgnd vpwr scs8hd_decap_12
XANTENNA__105__B address[3] vgnd vpwr scs8hd_diode_2
XFILLER_38_105 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A left_bottom_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_9.LATCH_1_.latch data_in mem_left_track_9.LATCH_1_.latch/Q _095_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__121__A _078_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_138 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB _059_/Y vgnd vpwr scs8hd_diode_2
XFILLER_37_171 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_top_track_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _041_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_62 vgnd vpwr scs8hd_decap_6
XFILLER_29_51 vgnd vpwr scs8hd_decap_8
XFILLER_29_73 vgnd vpwr scs8hd_decap_4
XANTENNA__116__A _075_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_88 vpwr vgnd scs8hd_fill_2
XFILLER_26_108 vgnd vpwr scs8hd_decap_4
Xmem_top_track_16.LATCH_2_.latch data_in mem_top_track_16.LATCH_2_.latch/Q _122_/Y
+ vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_34_141 vgnd vpwr scs8hd_decap_12
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_4_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_25_141 vpwr vgnd scs8hd_fill_2
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XFILLER_25_152 vpwr vgnd scs8hd_fill_2
XFILLER_31_74 vgnd vpwr scs8hd_decap_12
Xmux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_16_141 vpwr vgnd scs8hd_fill_2
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_right_track_0.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vpwr scs8hd_diode_2
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

