VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_0__3_
  CLASS BLOCK ;
  FOREIGN sb_0__3_ ;
  ORIGIN -0.005 0.000 ;
  SIZE 137.635 BY 140.000 ;
  PIN address[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.950 137.600 24.230 140.000 ;
    END
  END address[0]
  PIN address[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.430 137.600 41.710 140.000 ;
    END
  END address[1]
  PIN address[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.910 137.600 59.190 140.000 ;
    END
  END address[2]
  PIN address[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.390 137.600 76.670 140.000 ;
    END
  END address[3]
  PIN address[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 93.870 137.600 94.150 140.000 ;
    END
  END address[4]
  PIN address[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 111.350 137.600 111.630 140.000 ;
    END
  END address[5]
  PIN bottom_left_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.790 0.000 26.070 2.400 ;
    END
  END bottom_left_grid_pin_11_
  PIN bottom_left_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.850 0.000 31.130 2.400 ;
    END
  END bottom_left_grid_pin_13_
  PIN bottom_left_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.910 0.000 36.190 2.400 ;
    END
  END bottom_left_grid_pin_15_
  PIN bottom_left_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.030 0.000 0.310 2.400 ;
    END
  END bottom_left_grid_pin_1_
  PIN bottom_left_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.090 0.000 5.370 2.400 ;
    END
  END bottom_left_grid_pin_3_
  PIN bottom_left_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.150 0.000 10.430 2.400 ;
    END
  END bottom_left_grid_pin_5_
  PIN bottom_left_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.210 0.000 15.490 2.400 ;
    END
  END bottom_left_grid_pin_7_
  PIN bottom_left_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.730 0.000 21.010 2.400 ;
    END
  END bottom_left_grid_pin_9_
  PIN bottom_right_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 134.350 0.000 134.630 2.400 ;
    END
  END bottom_right_grid_pin_11_
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 53.760 137.640 54.360 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 58.520 137.640 59.120 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 63.960 137.640 64.560 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 69.400 137.640 70.000 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 74.160 137.640 74.760 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 79.600 137.640 80.200 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 85.040 137.640 85.640 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 89.800 137.640 90.400 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 95.240 137.640 95.840 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.240 6.840 137.640 7.440 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.240 12.280 137.640 12.880 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.240 17.040 137.640 17.640 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.240 22.480 137.640 23.080 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.240 27.920 137.640 28.520 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.240 32.680 137.640 33.280 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.240 38.120 137.640 38.720 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.240 43.560 137.640 44.160 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 135.240 48.320 137.640 48.920 ;
    END
  END chanx_right_out[8]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.430 0.000 41.710 2.400 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.490 0.000 46.770 2.400 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.550 0.000 51.830 2.400 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.610 0.000 56.890 2.400 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.130 0.000 62.410 2.400 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.190 0.000 67.470 2.400 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.250 0.000 72.530 2.400 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.310 0.000 77.590 2.400 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 82.830 0.000 83.110 2.400 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.890 0.000 88.170 2.400 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.950 0.000 93.230 2.400 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.010 0.000 98.290 2.400 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.530 0.000 103.810 2.400 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.590 0.000 108.870 2.400 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 113.650 0.000 113.930 2.400 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 118.710 0.000 118.990 2.400 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.230 0.000 124.510 2.400 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.290 0.000 129.570 2.400 ;
    END
  END chany_bottom_out[8]
  PIN data_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 128.830 137.600 129.110 140.000 ;
    END
  END data_in
  PIN enable
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.470 137.600 6.750 140.000 ;
    END
  END enable
  PIN right_bottom_grid_pin_12_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 2.080 137.640 2.680 ;
    END
  END right_bottom_grid_pin_12_
  PIN right_top_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 126.520 137.640 127.120 ;
    END
  END right_top_grid_pin_11_
  PIN right_top_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 131.280 137.640 131.880 ;
    END
  END right_top_grid_pin_13_
  PIN right_top_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 136.720 137.640 137.320 ;
    END
  END right_top_grid_pin_15_
  PIN right_top_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 100.000 137.640 100.600 ;
    END
  END right_top_grid_pin_1_
  PIN right_top_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 105.440 137.640 106.040 ;
    END
  END right_top_grid_pin_3_
  PIN right_top_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 110.880 137.640 111.480 ;
    END
  END right_top_grid_pin_5_
  PIN right_top_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 115.640 137.640 116.240 ;
    END
  END right_top_grid_pin_7_
  PIN right_top_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 135.240 121.080 137.640 121.680 ;
    END
  END right_top_grid_pin_9_
  PIN vpwr
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 25.695 10.640 27.295 128.080 ;
    END
  END vpwr
  PIN vgnd
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT 49.025 10.640 50.625 128.080 ;
    END
  END vgnd
  OBS
      LAYER li1 ;
        RECT 3.160 10.795 131.960 127.925 ;
      LAYER met1 ;
        RECT 3.160 10.640 131.960 137.320 ;
      LAYER met2 ;
        RECT 0.030 137.320 6.190 137.600 ;
        RECT 7.030 137.320 23.670 137.600 ;
        RECT 24.510 137.320 41.150 137.600 ;
        RECT 41.990 137.320 58.630 137.600 ;
        RECT 59.470 137.320 76.110 137.600 ;
        RECT 76.950 137.320 93.590 137.600 ;
        RECT 94.430 137.320 111.070 137.600 ;
        RECT 111.910 137.320 128.550 137.600 ;
        RECT 129.390 137.320 134.630 137.600 ;
        RECT 0.030 2.680 134.630 137.320 ;
        RECT 0.590 2.195 4.810 2.680 ;
        RECT 5.650 2.195 9.870 2.680 ;
        RECT 10.710 2.195 14.930 2.680 ;
        RECT 15.770 2.195 20.450 2.680 ;
        RECT 21.290 2.195 25.510 2.680 ;
        RECT 26.350 2.195 30.570 2.680 ;
        RECT 31.410 2.195 35.630 2.680 ;
        RECT 36.470 2.195 41.150 2.680 ;
        RECT 41.990 2.195 46.210 2.680 ;
        RECT 47.050 2.195 51.270 2.680 ;
        RECT 52.110 2.195 56.330 2.680 ;
        RECT 57.170 2.195 61.850 2.680 ;
        RECT 62.690 2.195 66.910 2.680 ;
        RECT 67.750 2.195 71.970 2.680 ;
        RECT 72.810 2.195 77.030 2.680 ;
        RECT 77.870 2.195 82.550 2.680 ;
        RECT 83.390 2.195 87.610 2.680 ;
        RECT 88.450 2.195 92.670 2.680 ;
        RECT 93.510 2.195 97.730 2.680 ;
        RECT 98.570 2.195 103.250 2.680 ;
        RECT 104.090 2.195 108.310 2.680 ;
        RECT 109.150 2.195 113.370 2.680 ;
        RECT 114.210 2.195 118.430 2.680 ;
        RECT 119.270 2.195 123.950 2.680 ;
        RECT 124.790 2.195 129.010 2.680 ;
        RECT 129.850 2.195 134.070 2.680 ;
      LAYER met3 ;
        RECT 0.005 136.320 134.840 137.185 ;
        RECT 0.005 132.280 135.240 136.320 ;
        RECT 0.005 130.880 134.840 132.280 ;
        RECT 0.005 127.520 135.240 130.880 ;
        RECT 0.005 126.120 134.840 127.520 ;
        RECT 0.005 122.080 135.240 126.120 ;
        RECT 0.005 120.680 134.840 122.080 ;
        RECT 0.005 116.640 135.240 120.680 ;
        RECT 0.005 115.240 134.840 116.640 ;
        RECT 0.005 111.880 135.240 115.240 ;
        RECT 0.005 110.480 134.840 111.880 ;
        RECT 0.005 106.440 135.240 110.480 ;
        RECT 0.005 105.040 134.840 106.440 ;
        RECT 0.005 101.000 135.240 105.040 ;
        RECT 0.005 99.600 134.840 101.000 ;
        RECT 0.005 96.240 135.240 99.600 ;
        RECT 0.005 94.840 134.840 96.240 ;
        RECT 0.005 90.800 135.240 94.840 ;
        RECT 0.005 89.400 134.840 90.800 ;
        RECT 0.005 86.040 135.240 89.400 ;
        RECT 0.005 84.640 134.840 86.040 ;
        RECT 0.005 80.600 135.240 84.640 ;
        RECT 0.005 79.200 134.840 80.600 ;
        RECT 0.005 75.160 135.240 79.200 ;
        RECT 0.005 73.760 134.840 75.160 ;
        RECT 0.005 70.400 135.240 73.760 ;
        RECT 0.005 69.000 134.840 70.400 ;
        RECT 0.005 64.960 135.240 69.000 ;
        RECT 0.005 63.560 134.840 64.960 ;
        RECT 0.005 59.520 135.240 63.560 ;
        RECT 0.005 58.120 134.840 59.520 ;
        RECT 0.005 54.760 135.240 58.120 ;
        RECT 0.005 53.360 134.840 54.760 ;
        RECT 0.005 49.320 135.240 53.360 ;
        RECT 0.005 47.920 134.840 49.320 ;
        RECT 0.005 44.560 135.240 47.920 ;
        RECT 0.005 43.160 134.840 44.560 ;
        RECT 0.005 39.120 135.240 43.160 ;
        RECT 0.005 37.720 134.840 39.120 ;
        RECT 0.005 33.680 135.240 37.720 ;
        RECT 0.005 32.280 134.840 33.680 ;
        RECT 0.005 28.920 135.240 32.280 ;
        RECT 0.005 27.520 134.840 28.920 ;
        RECT 0.005 23.480 135.240 27.520 ;
        RECT 0.005 22.080 134.840 23.480 ;
        RECT 0.005 18.040 135.240 22.080 ;
        RECT 0.005 16.640 134.840 18.040 ;
        RECT 0.005 13.280 135.240 16.640 ;
        RECT 0.005 11.880 134.840 13.280 ;
        RECT 0.005 7.840 135.240 11.880 ;
        RECT 0.005 6.440 134.840 7.840 ;
        RECT 0.005 3.080 135.240 6.440 ;
        RECT 0.005 2.215 134.840 3.080 ;
      LAYER met4 ;
        RECT 10.390 10.240 25.295 128.080 ;
        RECT 27.695 10.240 48.625 128.080 ;
        RECT 51.025 10.240 134.850 128.080 ;
        RECT 10.390 7.910 134.850 10.240 ;
      LAYER met5 ;
        RECT 10.180 7.700 135.060 39.900 ;
  END
END sb_0__3_
END LIBRARY

