* NGSPICE file created from sb_3__3_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor3_4 abstract view
.subckt scs8hd_nor3_4 A B C Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

.subckt sb_3__3_ address[0] address[1] address[2] address[3] address[4] address[5]
+ bottom_left_grid_pin_13_ bottom_right_grid_pin_11_ bottom_right_grid_pin_13_ bottom_right_grid_pin_15_
+ bottom_right_grid_pin_1_ bottom_right_grid_pin_3_ bottom_right_grid_pin_5_ bottom_right_grid_pin_7_
+ bottom_right_grid_pin_9_ chanx_left_in[0] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3]
+ chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8]
+ chanx_left_out[0] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4]
+ chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chany_bottom_in[0]
+ chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5]
+ chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_out[0] chany_bottom_out[1]
+ chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5]
+ chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8] data_in enable left_bottom_grid_pin_12_
+ left_top_grid_pin_11_ left_top_grid_pin_13_ left_top_grid_pin_15_ left_top_grid_pin_1_
+ left_top_grid_pin_3_ left_top_grid_pin_5_ left_top_grid_pin_7_ left_top_grid_pin_9_
+ vpwr vgnd
XFILLER_39_222 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 chanx_left_in[1] mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_27_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _225_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_6_129 vgnd vpwr scs8hd_decap_12
XFILLER_12_32 vgnd vpwr scs8hd_decap_6
XFILLER_37_73 vgnd vpwr scs8hd_decap_4
XFILLER_37_62 vpwr vgnd scs8hd_fill_2
XFILLER_37_95 vgnd vpwr scs8hd_decap_3
XANTENNA__108__B enable vgnd vpwr scs8hd_diode_2
XANTENNA__124__A _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_184 vgnd vpwr scs8hd_decap_12
XFILLER_24_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _190_/A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_3.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_3_ vgnd vpwr
+ scs8hd_diode_2
X_200_ _200_/A _200_/Y vgnd vpwr scs8hd_inv_8
X_131_ _147_/A _131_/B _131_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_53 vpwr vgnd scs8hd_fill_2
XFILLER_2_154 vgnd vpwr scs8hd_decap_12
XFILLER_0_57 vgnd vpwr scs8hd_decap_4
XANTENNA__110__C _123_/C vgnd vpwr scs8hd_diode_2
XANTENNA__119__A _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_9_55 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _239_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ _173_/Y mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_18_75 vpwr vgnd scs8hd_fill_2
XFILLER_11_220 vgnd vpwr scs8hd_decap_12
XFILLER_11_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _204_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_7_257 vgnd vpwr scs8hd_decap_12
X_114_ _113_/Y _115_/B vgnd vpwr scs8hd_buf_1
XFILLER_22_7 vgnd vpwr scs8hd_decap_3
XFILLER_37_172 vgnd vpwr scs8hd_decap_8
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XFILLER_20_21 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _223_/HI _194_/Y mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_20_87 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_11.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_6_23 vgnd vpwr scs8hd_decap_8
XANTENNA__116__B _115_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__132__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_6_67 vpwr vgnd scs8hd_fill_2
XFILLER_13_3 vpwr vgnd scs8hd_fill_2
XFILLER_34_142 vgnd vpwr scs8hd_decap_8
XFILLER_1_208 vgnd vpwr scs8hd_decap_12
XFILLER_25_175 vgnd vpwr scs8hd_decap_8
XFILLER_25_142 vpwr vgnd scs8hd_fill_2
XFILLER_25_120 vpwr vgnd scs8hd_fill_2
XFILLER_40_178 vgnd vpwr scs8hd_decap_12
XFILLER_31_53 vpwr vgnd scs8hd_fill_2
XFILLER_15_65 vgnd vpwr scs8hd_decap_4
XFILLER_31_97 vpwr vgnd scs8hd_fill_2
XFILLER_31_75 vpwr vgnd scs8hd_fill_2
XFILLER_0_230 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _187_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_31_123 vgnd vpwr scs8hd_decap_3
XFILLER_16_131 vgnd vpwr scs8hd_decap_4
XFILLER_16_142 vgnd vpwr scs8hd_decap_3
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__A _096_/X vgnd vpwr scs8hd_diode_2
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_192 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_234 vgnd vpwr scs8hd_decap_8
XFILLER_39_245 vgnd vpwr scs8hd_decap_8
XFILLER_13_112 vpwr vgnd scs8hd_fill_2
XFILLER_13_123 vgnd vpwr scs8hd_decap_4
XFILLER_13_145 vgnd vpwr scs8hd_decap_4
XFILLER_42_63 vgnd vpwr scs8hd_decap_12
XFILLER_9_138 vpwr vgnd scs8hd_fill_2
XFILLER_9_149 vgnd vpwr scs8hd_decap_4
XFILLER_36_215 vgnd vpwr scs8hd_decap_12
XFILLER_42_218 vgnd vpwr scs8hd_decap_12
XFILLER_12_88 vgnd vpwr scs8hd_decap_4
XANTENNA__230__A _230_/A vgnd vpwr scs8hd_diode_2
Xmux_left_track_13.tap_buf4_0_.scs8hd_inv_1 mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ _228_/A vgnd vpwr scs8hd_inv_1
XFILLER_18_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _206_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__124__B _124_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_196 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _173_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_15.LATCH_0_.latch_SLEEPB _136_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__140__A _115_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vpwr scs8hd_diode_2
X_130_ _126_/A _115_/B _134_/C _168_/A _131_/B vgnd vpwr scs8hd_or4_4
XFILLER_23_98 vpwr vgnd scs8hd_fill_2
XFILLER_2_166 vgnd vpwr scs8hd_decap_12
XANTENNA__110__D _171_/A vgnd vpwr scs8hd_diode_2
XANTENNA__119__B _119_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA__135__A _147_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_251 vgnd vpwr scs8hd_decap_12
XFILLER_20_210 vgnd vpwr scs8hd_decap_4
XFILLER_20_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_5.tap_buf4_0_.scs8hd_inv_1 mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ _232_/A vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _189_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_18_87 vpwr vgnd scs8hd_fill_2
XFILLER_11_232 vgnd vpwr scs8hd_decap_12
X_113_ address[2] _113_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _197_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB _145_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_269 vgnd vpwr scs8hd_decap_8
XFILLER_29_118 vpwr vgnd scs8hd_fill_2
XFILLER_37_184 vgnd vpwr scs8hd_decap_12
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XFILLER_29_97 vpwr vgnd scs8hd_fill_2
XFILLER_29_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_35 vgnd vpwr scs8hd_decap_12
Xmux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ _193_/A mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_19_184 vgnd vpwr scs8hd_decap_12
XFILLER_34_154 vgnd vpwr scs8hd_decap_12
Xmem_left_track_5.LATCH_1_.latch data_in _194_/A _150_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_13.LATCH_1_.latch_SLEEPB _131_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_102 vgnd vpwr scs8hd_decap_12
XFILLER_31_10 vpwr vgnd scs8hd_fill_2
XANTENNA__233__A _233_/A vgnd vpwr scs8hd_diode_2
XFILLER_0_242 vgnd vpwr scs8hd_decap_6
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 left_bottom_grid_pin_12_ mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_31_135 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _175_/A vgnd
+ vpwr scs8hd_diode_2
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__127__B _128_/B vgnd vpwr scs8hd_diode_2
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_193 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__A _115_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_146 vgnd vpwr scs8hd_fill_1
XFILLER_26_10 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__228__A _228_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_75 vgnd vpwr scs8hd_decap_12
XFILLER_21_190 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _235_/A vgnd vpwr scs8hd_inv_1
XFILLER_3_69 vpwr vgnd scs8hd_fill_2
XFILLER_36_227 vgnd vpwr scs8hd_decap_12
XANTENNA__138__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_8_150 vgnd vpwr scs8hd_decap_3
Xmux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ _197_/Y mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_12_67 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _199_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_6 vpwr vgnd scs8hd_fill_2
XFILLER_37_86 vpwr vgnd scs8hd_fill_2
XFILLER_37_31 vgnd vpwr scs8hd_fill_1
XFILLER_33_208 vgnd vpwr scs8hd_decap_12
XFILLER_18_227 vgnd vpwr scs8hd_decap_12
XANTENNA__140__B _123_/B vgnd vpwr scs8hd_diode_2
XFILLER_32_263 vgnd vpwr scs8hd_decap_12
XFILLER_15_208 vgnd vpwr scs8hd_decap_12
XFILLER_23_252 vgnd vpwr scs8hd_decap_3
XANTENNA__241__A _241_/A vgnd vpwr scs8hd_diode_2
XFILLER_2_101 vpwr vgnd scs8hd_fill_2
XFILLER_2_178 vgnd vpwr scs8hd_decap_12
XFILLER_14_263 vgnd vpwr scs8hd_decap_12
X_189_ _189_/A _189_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__135__B _134_/X vgnd vpwr scs8hd_diode_2
XANTENNA__151__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_11 vpwr vgnd scs8hd_fill_2
XFILLER_18_22 vpwr vgnd scs8hd_fill_2
XFILLER_34_43 vgnd vpwr scs8hd_fill_1
XANTENNA__236__A _236_/A vgnd vpwr scs8hd_diode_2
X_112_ _106_/X _110_/X _112_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__146__A address[3] vgnd vpwr scs8hd_diode_2
XFILLER_37_196 vgnd vpwr scs8hd_decap_12
XFILLER_20_78 vgnd vpwr scs8hd_decap_3
XFILLER_29_76 vpwr vgnd scs8hd_fill_2
XFILLER_29_32 vgnd vpwr scs8hd_fill_1
XFILLER_28_163 vgnd vpwr scs8hd_decap_12
XFILLER_28_141 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_47 vgnd vpwr scs8hd_decap_12
XFILLER_34_166 vgnd vpwr scs8hd_decap_12
XFILLER_19_174 vpwr vgnd scs8hd_fill_2
XFILLER_19_196 vgnd vpwr scs8hd_decap_12
XFILLER_40_114 vgnd vpwr scs8hd_decap_12
XFILLER_15_12 vpwr vgnd scs8hd_fill_2
XFILLER_15_34 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[6] vgnd vpwr scs8hd_diode_2
XFILLER_31_114 vpwr vgnd scs8hd_fill_2
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_194 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__B _123_/B vgnd vpwr scs8hd_diode_2
XFILLER_39_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_136 vgnd vpwr scs8hd_decap_4
XFILLER_7_90 vgnd vpwr scs8hd_decap_3
XFILLER_42_87 vgnd vpwr scs8hd_decap_6
XFILLER_42_32 vgnd vpwr scs8hd_decap_12
XFILLER_9_118 vpwr vgnd scs8hd_fill_2
XFILLER_13_169 vgnd vpwr scs8hd_decap_12
XFILLER_36_239 vgnd vpwr scs8hd_decap_12
XANTENNA__138__B _138_/B vgnd vpwr scs8hd_diode_2
XFILLER_12_180 vgnd vpwr scs8hd_decap_12
XANTENNA__154__A _168_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_15_ mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_128 vpwr vgnd scs8hd_fill_2
XFILLER_41_220 vgnd vpwr scs8hd_decap_12
XANTENNA__239__A _239_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_239 vgnd vpwr scs8hd_decap_12
XFILLER_5_121 vgnd vpwr scs8hd_fill_1
Xmem_left_track_15.LATCH_0_.latch data_in _205_/A _169_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__140__C _143_/C vgnd vpwr scs8hd_diode_2
XANTENNA__149__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _188_/A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_80 vpwr vgnd scs8hd_fill_2
XFILLER_23_220 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_13.LATCH_0_.latch_SLEEPB _165_/Y vgnd vpwr scs8hd_diode_2
XFILLER_23_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_1_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_69 vpwr vgnd scs8hd_fill_2
X_188_ _188_/A _188_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__151__B _149_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[3] vgnd vpwr scs8hd_diode_2
XFILLER_18_45 vgnd vpwr scs8hd_decap_4
XFILLER_34_99 vgnd vpwr scs8hd_fill_1
XFILLER_11_245 vgnd vpwr scs8hd_decap_8
X_111_ _096_/X _110_/X _111_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__146__B _115_/B vgnd vpwr scs8hd_diode_2
XANTENNA__162__A _155_/X vgnd vpwr scs8hd_diode_2
XFILLER_29_22 vpwr vgnd scs8hd_fill_2
XFILLER_29_11 vpwr vgnd scs8hd_fill_2
XFILLER_20_57 vgnd vpwr scs8hd_decap_6
XFILLER_28_175 vgnd vpwr scs8hd_decap_12
XFILLER_28_120 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_7.LATCH_0_.latch_SLEEPB _120_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_59 vgnd vpwr scs8hd_decap_8
XFILLER_6_15 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_13.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_90 vpwr vgnd scs8hd_fill_2
XFILLER_20_7 vgnd vpwr scs8hd_fill_1
XFILLER_34_178 vgnd vpwr scs8hd_decap_12
XANTENNA__157__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_19_153 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_25_123 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_40_126 vgnd vpwr scs8hd_decap_12
XFILLER_15_57 vpwr vgnd scs8hd_fill_2
XFILLER_31_23 vpwr vgnd scs8hd_fill_2
XFILLER_16_101 vpwr vgnd scs8hd_fill_2
XFILLER_16_112 vgnd vpwr scs8hd_decap_8
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_11.LATCH_1_.latch_SLEEPB _161_/Y vgnd vpwr scs8hd_diode_2
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_195 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__C _143_/C vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _222_/HI _192_/Y mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_3 vgnd vpwr scs8hd_decap_3
XFILLER_30_181 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _207_/Y vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_1.LATCH_1_.latch data_in _190_/A _144_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_26_67 vpwr vgnd scs8hd_fill_2
XFILLER_26_56 vgnd vpwr scs8hd_decap_6
XFILLER_26_23 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_11.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_11_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_42_44 vgnd vpwr scs8hd_decap_12
XFILLER_21_181 vpwr vgnd scs8hd_fill_2
XFILLER_3_16 vgnd vpwr scs8hd_decap_12
XFILLER_12_192 vgnd vpwr scs8hd_decap_12
XANTENNA__154__B _153_/X vgnd vpwr scs8hd_diode_2
XANTENNA__170__A _171_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_232 vgnd vpwr scs8hd_decap_12
XFILLER_37_77 vgnd vpwr scs8hd_fill_1
XFILLER_26_251 vgnd vpwr scs8hd_decap_12
XANTENNA__140__D _153_/D vgnd vpwr scs8hd_diode_2
XANTENNA__149__B _115_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.LATCH_1_.latch_SLEEPB _116_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_262 vgnd vpwr scs8hd_decap_12
XFILLER_32_276 vgnd vpwr scs8hd_fill_1
XANTENNA__165__A _155_/X vgnd vpwr scs8hd_diode_2
XFILLER_23_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_57 vpwr vgnd scs8hd_fill_2
XFILLER_2_125 vgnd vpwr scs8hd_decap_3
Xmux_left_track_13.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_13_ mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_15 vpwr vgnd scs8hd_fill_2
XFILLER_9_37 vpwr vgnd scs8hd_fill_2
XFILLER_9_59 vpwr vgnd scs8hd_fill_2
XFILLER_14_276 vgnd vpwr scs8hd_fill_1
X_187_ _187_/A _187_/Y vgnd vpwr scs8hd_inv_8
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[3] mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_18_79 vpwr vgnd scs8hd_fill_2
XFILLER_34_56 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _186_/Y vgnd
+ vpwr scs8hd_diode_2
X_110_ _115_/A _123_/B _123_/C _171_/A _110_/X vgnd vpwr scs8hd_or4_4
X_239_ _239_/A chany_bottom_out[4] vgnd vpwr scs8hd_buf_2
XANTENNA__146__C _143_/C vgnd vpwr scs8hd_diode_2
XFILLER_41_3 vgnd vpwr scs8hd_decap_12
XANTENNA__162__B _162_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_132 vpwr vgnd scs8hd_fill_2
XFILLER_20_25 vpwr vgnd scs8hd_fill_2
XFILLER_28_187 vgnd vpwr scs8hd_decap_12
XFILLER_3_220 vgnd vpwr scs8hd_decap_12
XFILLER_13_7 vpwr vgnd scs8hd_fill_2
XFILLER_19_132 vgnd vpwr scs8hd_decap_4
XANTENNA__157__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _218_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__173__A _173_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_146 vpwr vgnd scs8hd_fill_2
XFILLER_25_113 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB _158_/Y vgnd vpwr scs8hd_diode_2
XFILLER_40_138 vgnd vpwr scs8hd_decap_12
XFILLER_15_47 vgnd vpwr scs8hd_decap_4
XFILLER_31_79 vgnd vpwr scs8hd_decap_3
XFILLER_31_57 vpwr vgnd scs8hd_fill_2
XFILLER_0_201 vgnd vpwr scs8hd_decap_12
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_135 vgnd vpwr scs8hd_fill_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__143__D _109_/A vgnd vpwr scs8hd_diode_2
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _172_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_90 vgnd vpwr scs8hd_decap_4
XANTENNA__168__A _168_/A vgnd vpwr scs8hd_diode_2
XFILLER_22_149 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ _191_/A mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_30_193 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_26_35 vgnd vpwr scs8hd_decap_8
XFILLER_13_116 vgnd vpwr scs8hd_decap_4
XFILLER_13_127 vgnd vpwr scs8hd_fill_1
XFILLER_13_149 vgnd vpwr scs8hd_fill_1
XFILLER_42_56 vgnd vpwr scs8hd_decap_6
XFILLER_21_160 vpwr vgnd scs8hd_fill_2
XFILLER_3_28 vgnd vpwr scs8hd_decap_12
XFILLER_8_142 vgnd vpwr scs8hd_decap_8
XFILLER_8_164 vgnd vpwr scs8hd_decap_8
XFILLER_8_175 vgnd vpwr scs8hd_decap_12
XANTENNA__170__B _168_/B vgnd vpwr scs8hd_diode_2
XFILLER_27_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _188_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_37_34 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _196_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_263 vgnd vpwr scs8hd_decap_12
XFILLER_5_123 vgnd vpwr scs8hd_decap_12
XANTENNA__149__C _143_/C vgnd vpwr scs8hd_diode_2
XFILLER_17_274 vgnd vpwr scs8hd_decap_3
XANTENNA__165__B _165_/B vgnd vpwr scs8hd_diode_2
XANTENNA__181__A _181_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_93 vgnd vpwr scs8hd_decap_12
XFILLER_23_36 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ _195_/Y mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_3_6 vpwr vgnd scs8hd_fill_2
XFILLER_2_137 vgnd vpwr scs8hd_decap_12
XFILLER_14_211 vgnd vpwr scs8hd_decap_3
X_186_ _186_/A _186_/Y vgnd vpwr scs8hd_inv_8
XFILLER_36_6 vgnd vpwr scs8hd_decap_12
XANTENNA__176__A _176_/A vgnd vpwr scs8hd_diode_2
Xmem_left_track_11.LATCH_0_.latch data_in _201_/A _162_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_20_258 vgnd vpwr scs8hd_decap_12
XFILLER_18_58 vpwr vgnd scs8hd_fill_2
XFILLER_34_46 vgnd vpwr scs8hd_fill_1
XFILLER_34_35 vgnd vpwr scs8hd_decap_8
XFILLER_7_218 vpwr vgnd scs8hd_fill_2
XFILLER_11_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _174_/A vgnd
+ vpwr scs8hd_diode_2
X_238_ _238_/A chany_bottom_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_6_251 vgnd vpwr scs8hd_decap_12
Xmux_left_track_11.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_11_ mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__146__D _153_/D vgnd vpwr scs8hd_diode_2
X_169_ _168_/A _168_/B _155_/X _169_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_34_3 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_7.LATCH_0_.latch data_in _179_/A _120_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_57 vpwr vgnd scs8hd_fill_2
XFILLER_28_199 vgnd vpwr scs8hd_decap_12
Xmux_left_track_7.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[2] mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_232 vgnd vpwr scs8hd_decap_12
XFILLER_19_166 vpwr vgnd scs8hd_fill_2
XFILLER_42_180 vgnd vpwr scs8hd_decap_6
XANTENNA__157__C _143_/C vgnd vpwr scs8hd_diode_2
XFILLER_33_180 vgnd vpwr scs8hd_decap_3
XFILLER_31_36 vpwr vgnd scs8hd_fill_2
XFILLER_31_14 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _198_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_213 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_31_139 vgnd vpwr scs8hd_decap_12
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_147 vpwr vgnd scs8hd_fill_2
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__168__B _168_/B vgnd vpwr scs8hd_diode_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__184__A _184_/A vgnd vpwr scs8hd_diode_2
XFILLER_7_82 vpwr vgnd scs8hd_fill_2
XFILLER_38_272 vgnd vpwr scs8hd_decap_3
XFILLER_21_194 vgnd vpwr scs8hd_decap_12
XFILLER_8_121 vpwr vgnd scs8hd_fill_2
XFILLER_8_132 vgnd vpwr scs8hd_decap_4
XFILLER_8_154 vgnd vpwr scs8hd_decap_6
XFILLER_8_187 vgnd vpwr scs8hd_decap_12
XANTENNA__170__C _168_/C vgnd vpwr scs8hd_diode_2
XANTENNA__179__A _179_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_220 vgnd vpwr scs8hd_decap_12
XFILLER_37_46 vgnd vpwr scs8hd_decap_12
XFILLER_18_209 vgnd vpwr scs8hd_decap_4
XFILLER_41_245 vgnd vpwr scs8hd_decap_12
XFILLER_5_135 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_7.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__149__D _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_253 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_190 vgnd vpwr scs8hd_decap_12
XFILLER_2_105 vgnd vpwr scs8hd_decap_6
XFILLER_2_149 vgnd vpwr scs8hd_decap_4
X_185_ _185_/A _185_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_171 vgnd vpwr scs8hd_decap_12
XFILLER_20_215 vgnd vpwr scs8hd_decap_12
XANTENNA__192__A _192_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_26 vgnd vpwr scs8hd_decap_4
XFILLER_7_208 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _186_/A mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_237_ _237_/A chany_bottom_out[6] vgnd vpwr scs8hd_buf_2
XFILLER_6_263 vgnd vpwr scs8hd_decap_12
XFILLER_10_270 vgnd vpwr scs8hd_decap_4
XFILLER_24_91 vgnd vpwr scs8hd_fill_1
X_168_ _168_/A _168_/B _168_/C _168_/Y vgnd vpwr scs8hd_nor3_4
XFILLER_27_3 vpwr vgnd scs8hd_fill_2
X_099_ address[4] address[5] _134_/C vgnd vpwr scs8hd_or2_4
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
XANTENNA__187__A _187_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_36 vpwr vgnd scs8hd_fill_2
XFILLER_28_145 vgnd vpwr scs8hd_decap_8
XANTENNA__097__A address[3] vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_15.LATCH_0_.latch data_in _187_/A _136_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_10_82 vpwr vgnd scs8hd_fill_2
XFILLER_10_93 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_34_126 vpwr vgnd scs8hd_fill_2
XFILLER_19_101 vpwr vgnd scs8hd_fill_2
XFILLER_19_112 vpwr vgnd scs8hd_fill_2
XFILLER_19_156 vgnd vpwr scs8hd_fill_1
XFILLER_19_178 vgnd vpwr scs8hd_decap_4
XANTENNA__157__D _109_/A vgnd vpwr scs8hd_diode_2
XFILLER_25_159 vpwr vgnd scs8hd_fill_2
XFILLER_15_16 vpwr vgnd scs8hd_fill_2
XFILLER_31_118 vgnd vpwr scs8hd_decap_4
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_198 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_218 vpwr vgnd scs8hd_fill_2
Xmux_left_track_5.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[1] mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__168__C _168_/C vgnd vpwr scs8hd_diode_2
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_22_118 vgnd vpwr scs8hd_fill_1
XFILLER_30_151 vpwr vgnd scs8hd_fill_2
XFILLER_7_72 vgnd vpwr scs8hd_fill_1
XFILLER_38_240 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 chanx_left_in[0] mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mem_bottom_track_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_173 vgnd vpwr scs8hd_decap_8
XFILLER_21_184 vpwr vgnd scs8hd_fill_2
XFILLER_29_262 vpwr vgnd scs8hd_fill_2
XFILLER_32_91 vgnd vpwr scs8hd_fill_1
XFILLER_8_199 vgnd vpwr scs8hd_decap_12
XFILLER_35_232 vgnd vpwr scs8hd_decap_12
XANTENNA__195__A _195_/A vgnd vpwr scs8hd_diode_2
XFILLER_12_17 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _217_/HI _190_/Y mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_37_58 vgnd vpwr scs8hd_fill_1
XFILLER_26_276 vgnd vpwr scs8hd_fill_1
XFILLER_41_257 vgnd vpwr scs8hd_decap_12
XFILLER_5_103 vgnd vpwr scs8hd_decap_12
XFILLER_5_147 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ _241_/A vgnd vpwr scs8hd_inv_1
XFILLER_32_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_84 vgnd vpwr scs8hd_decap_8
XFILLER_23_257 vgnd vpwr scs8hd_decap_12
XFILLER_13_71 vpwr vgnd scs8hd_fill_2
X_184_ _184_/A _184_/Y vgnd vpwr scs8hd_inv_8
XFILLER_29_7 vpwr vgnd scs8hd_fill_2
XFILLER_20_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_15.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_34_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_24_70 vgnd vpwr scs8hd_fill_1
XFILLER_40_80 vgnd vpwr scs8hd_decap_12
X_236_ _236_/A chany_bottom_out[7] vgnd vpwr scs8hd_buf_2
X_098_ address[2] _123_/B vgnd vpwr scs8hd_buf_1
X_167_ _167_/A _168_/B vgnd vpwr scs8hd_buf_1
XFILLER_37_113 vgnd vpwr scs8hd_decap_3
XFILLER_1_74 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _206_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_26 vgnd vpwr scs8hd_decap_6
XFILLER_20_17 vpwr vgnd scs8hd_fill_2
XFILLER_6_19 vpwr vgnd scs8hd_fill_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
X_219_ _219_/HI _219_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__198__A _198_/A vgnd vpwr scs8hd_diode_2
XFILLER_33_160 vgnd vpwr scs8hd_decap_12
XFILLER_25_127 vgnd vpwr scs8hd_decap_4
XFILLER_31_27 vgnd vpwr scs8hd_decap_6
Xmem_bottom_track_3.LATCH_0_.latch data_in _175_/A _112_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_138 vgnd vpwr scs8hd_fill_1
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_199 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_39_208 vgnd vpwr scs8hd_decap_6
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ _189_/A mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XPHY_2 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _189_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_7_95 vgnd vpwr scs8hd_decap_12
XFILLER_7_62 vgnd vpwr scs8hd_decap_4
XFILLER_38_252 vgnd vpwr scs8hd_decap_12
XFILLER_42_15 vgnd vpwr scs8hd_decap_12
XFILLER_29_274 vgnd vpwr scs8hd_decap_3
XFILLER_16_60 vpwr vgnd scs8hd_fill_2
XFILLER_16_82 vpwr vgnd scs8hd_fill_2
XFILLER_16_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_12_141 vpwr vgnd scs8hd_fill_2
XFILLER_12_163 vgnd vpwr scs8hd_decap_8
Xmux_left_track_3.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[0] mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_9_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_12_29 vpwr vgnd scs8hd_fill_2
XFILLER_37_15 vgnd vpwr scs8hd_decap_12
XFILLER_26_211 vgnd vpwr scs8hd_decap_3
XFILLER_41_269 vgnd vpwr scs8hd_decap_8
XFILLER_5_115 vgnd vpwr scs8hd_decap_6
XFILLER_5_159 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_15.INVTX1_1_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_27_81 vgnd vpwr scs8hd_decap_4
XFILLER_17_200 vgnd vpwr scs8hd_decap_12
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _234_/A vgnd vpwr scs8hd_inv_1
XFILLER_23_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _175_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_9_ mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_9_19 vpwr vgnd scs8hd_fill_2
XFILLER_13_83 vgnd vpwr scs8hd_fill_1
X_183_ _183_/A _183_/Y vgnd vpwr scs8hd_inv_8
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XFILLER_9_262 vpwr vgnd scs8hd_fill_2
XFILLER_20_239 vgnd vpwr scs8hd_decap_12
XFILLER_34_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_6 vpwr vgnd scs8hd_fill_2
X_235_ _235_/A chany_bottom_out[8] vgnd vpwr scs8hd_buf_2
Xmux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ _193_/Y mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_6_276 vgnd vpwr scs8hd_fill_1
X_166_ address[3] address[2] address[4] _138_/B _167_/A vgnd vpwr scs8hd_or4_4
X_097_ address[3] _115_/A vgnd vpwr scs8hd_buf_1
XFILLER_37_136 vgnd vpwr scs8hd_decap_12
XFILLER_1_86 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _199_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_20_29 vpwr vgnd scs8hd_fill_2
XFILLER_3_257 vgnd vpwr scs8hd_decap_12
XFILLER_19_71 vpwr vgnd scs8hd_fill_2
XFILLER_35_92 vgnd vpwr scs8hd_fill_1
XFILLER_27_180 vgnd vpwr scs8hd_decap_3
X_149_ address[3] _115_/B _143_/C _109_/A _149_/X vgnd vpwr scs8hd_or4_4
X_218_ _218_/HI _218_/LO vgnd vpwr scs8hd_conb_1
XFILLER_32_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _219_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_117 vgnd vpwr scs8hd_fill_1
XFILLER_33_172 vgnd vpwr scs8hd_decap_8
XFILLER_15_29 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ _237_/A vgnd vpwr scs8hd_inv_1
XFILLER_0_249 vgnd vpwr scs8hd_decap_12
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_94 vgnd vpwr scs8hd_fill_1
XFILLER_11_8 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_11.LATCH_0_.latch data_in _183_/A _128_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_38_264 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _177_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_42_27 vgnd vpwr scs8hd_decap_4
XFILLER_29_253 vpwr vgnd scs8hd_fill_2
XFILLER_29_220 vgnd vpwr scs8hd_decap_12
XFILLER_8_102 vgnd vpwr scs8hd_fill_1
XFILLER_16_72 vgnd vpwr scs8hd_fill_1
XFILLER_35_245 vgnd vpwr scs8hd_decap_12
XFILLER_37_27 vgnd vpwr scs8hd_decap_4
XFILLER_17_212 vgnd vpwr scs8hd_decap_12
XFILLER_17_245 vgnd vpwr scs8hd_decap_8
XFILLER_32_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _107_/Y vgnd vpwr scs8hd_diode_2
XFILLER_4_64 vgnd vpwr scs8hd_fill_1
XFILLER_23_248 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[8] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_14_215 vgnd vpwr scs8hd_decap_12
X_182_ _182_/A _182_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_95 vpwr vgnd scs8hd_fill_2
XFILLER_38_81 vgnd vpwr scs8hd_decap_8
XFILLER_1_196 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_13.INVTX1_1_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__100__A _134_/C vgnd vpwr scs8hd_diode_2
XFILLER_9_274 vgnd vpwr scs8hd_decap_3
X_234_ _234_/A chanx_left_out[0] vgnd vpwr scs8hd_buf_2
XFILLER_10_251 vgnd vpwr scs8hd_decap_4
X_165_ _155_/X _165_/B _165_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_40_93 vgnd vpwr scs8hd_decap_6
X_096_ _129_/A _096_/X vgnd vpwr scs8hd_buf_1
XFILLER_37_148 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_7.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_7_ mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_1_10 vgnd vpwr scs8hd_decap_12
XFILLER_1_98 vgnd vpwr scs8hd_fill_1
Xmem_left_track_15.LATCH_1_.latch data_in _204_/A _168_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_28_137 vpwr vgnd scs8hd_fill_2
XFILLER_28_126 vpwr vgnd scs8hd_fill_2
XFILLER_3_269 vgnd vpwr scs8hd_decap_8
XFILLER_10_30 vgnd vpwr scs8hd_fill_1
XFILLER_10_52 vgnd vpwr scs8hd_decap_4
XFILLER_19_50 vgnd vpwr scs8hd_decap_4
XFILLER_35_71 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _184_/A mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
X_217_ _217_/HI _217_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _191_/A vgnd vpwr
+ scs8hd_diode_2
X_148_ _145_/A _147_/B _148_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_25_3 vpwr vgnd scs8hd_fill_2
XFILLER_33_184 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_5.LATCH_0_.latch_SLEEPB _151_/Y vgnd vpwr scs8hd_diode_2
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_40 vpwr vgnd scs8hd_fill_2
XFILLER_21_73 vpwr vgnd scs8hd_fill_2
XFILLER_30_121 vgnd vpwr scs8hd_decap_4
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_15_162 vpwr vgnd scs8hd_fill_2
XFILLER_15_173 vpwr vgnd scs8hd_fill_2
XFILLER_15_184 vgnd vpwr scs8hd_decap_12
XFILLER_7_86 vpwr vgnd scs8hd_fill_2
XFILLER_7_53 vgnd vpwr scs8hd_decap_6
XANTENNA_mem_left_track_9.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_276 vgnd vpwr scs8hd_fill_1
XFILLER_26_29 vpwr vgnd scs8hd_fill_2
XFILLER_21_143 vpwr vgnd scs8hd_fill_2
XFILLER_29_232 vgnd vpwr scs8hd_decap_12
XFILLER_8_125 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _141_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__103__A _153_/D vgnd vpwr scs8hd_diode_2
XFILLER_35_257 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _212_/HI _188_/Y mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[1] vgnd vpwr scs8hd_diode_2
XFILLER_32_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_224 vgnd vpwr scs8hd_decap_12
XFILLER_4_76 vpwr vgnd scs8hd_fill_2
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XFILLER_4_10 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_19 vpwr vgnd scs8hd_fill_2
XFILLER_14_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_3.LATCH_1_.latch_SLEEPB _147_/Y vgnd vpwr scs8hd_diode_2
X_181_ _181_/A _181_/Y vgnd vpwr scs8hd_inv_8
XFILLER_38_71 vgnd vpwr scs8hd_decap_6
XFILLER_9_220 vgnd vpwr scs8hd_decap_12
XFILLER_9_253 vpwr vgnd scs8hd_fill_2
XFILLER_11_208 vgnd vpwr scs8hd_decap_12
XANTENNA__201__A _201_/A vgnd vpwr scs8hd_diode_2
X_233_ _233_/A chanx_left_out[1] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_13_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_10_274 vgnd vpwr scs8hd_fill_1
X_164_ _168_/C _165_/B _164_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_84 vgnd vpwr scs8hd_decap_4
X_095_ address[0] _129_/A vgnd vpwr scs8hd_inv_8
XFILLER_1_22 vgnd vpwr scs8hd_decap_12
XANTENNA__111__A _096_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_29_18 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_11.INVTX1_1_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_10_86 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_11.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_27_160 vgnd vpwr scs8hd_decap_12
XFILLER_19_62 vpwr vgnd scs8hd_fill_2
XFILLER_19_84 vpwr vgnd scs8hd_fill_2
XFILLER_19_105 vpwr vgnd scs8hd_fill_2
XFILLER_19_116 vgnd vpwr scs8hd_decap_4
XFILLER_19_138 vpwr vgnd scs8hd_fill_2
XFILLER_19_149 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
X_147_ _147_/A _147_/B _147_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__106__A address[0] vgnd vpwr scs8hd_diode_2
X_216_ _216_/HI _216_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mem_bottom_track_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_18_3 vpwr vgnd scs8hd_fill_2
XFILLER_33_196 vgnd vpwr scs8hd_decap_12
XFILLER_31_19 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_5_ mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_0_218 vgnd vpwr scs8hd_decap_12
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_152 vgnd vpwr scs8hd_fill_1
XFILLER_24_163 vgnd vpwr scs8hd_decap_12
XFILLER_21_52 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_15_141 vpwr vgnd scs8hd_fill_2
XFILLER_7_32 vgnd vpwr scs8hd_decap_6
XFILLER_15_196 vgnd vpwr scs8hd_decap_12
XFILLER_29_266 vgnd vpwr scs8hd_decap_8
XFILLER_12_100 vpwr vgnd scs8hd_fill_2
XFILLER_12_122 vgnd vpwr scs8hd_fill_1
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _206_/A mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_35_269 vgnd vpwr scs8hd_decap_8
XFILLER_7_170 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ _187_/A mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_7_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__204__A _204_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_239 vgnd vpwr scs8hd_decap_12
XFILLER_27_73 vpwr vgnd scs8hd_fill_2
XFILLER_27_40 vpwr vgnd scs8hd_fill_2
XFILLER_17_236 vgnd vpwr scs8hd_decap_8
XFILLER_17_258 vpwr vgnd scs8hd_fill_2
XFILLER_4_44 vgnd vpwr scs8hd_decap_12
XANTENNA__114__A _113_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_239 vgnd vpwr scs8hd_decap_12
X_180_ _180_/A _180_/Y vgnd vpwr scs8hd_inv_8
XFILLER_13_31 vpwr vgnd scs8hd_fill_2
XFILLER_13_53 vpwr vgnd scs8hd_fill_2
XFILLER_13_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _208_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_1_110 vgnd vpwr scs8hd_fill_1
XFILLER_1_132 vpwr vgnd scs8hd_fill_2
XFILLER_1_143 vpwr vgnd scs8hd_fill_2
XFILLER_9_232 vgnd vpwr scs8hd_decap_12
XANTENNA__109__A _109_/A vgnd vpwr scs8hd_diode_2
X_232_ _232_/A chanx_left_out[2] vgnd vpwr scs8hd_buf_2
XFILLER_24_30 vgnd vpwr scs8hd_fill_1
XFILLER_24_63 vgnd vpwr scs8hd_decap_4
XFILLER_6_202 vgnd vpwr scs8hd_decap_12
X_163_ _122_/A _113_/Y _160_/C _109_/A _165_/B vgnd vpwr scs8hd_or4_4
XFILLER_24_96 vpwr vgnd scs8hd_fill_2
XANTENNA__111__B _110_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _188_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_1_34 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB _171_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_32 vgnd vpwr scs8hd_decap_4
XFILLER_10_65 vpwr vgnd scs8hd_fill_2
XFILLER_10_98 vpwr vgnd scs8hd_fill_2
XFILLER_34_109 vgnd vpwr scs8hd_decap_8
XFILLER_27_172 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_13.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_35_95 vpwr vgnd scs8hd_fill_2
X_215_ _215_/HI _215_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__122__A _122_/A vgnd vpwr scs8hd_diode_2
X_146_ address[3] _115_/B _143_/C _153_/D _147_/B vgnd vpwr scs8hd_or4_4
XFILLER_25_109 vpwr vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ _191_/Y mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A left_bottom_grid_pin_12_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__207__A _207_/A vgnd vpwr scs8hd_diode_2
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmem_left_track_11.LATCH_1_.latch data_in _200_/A _161_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_24_131 vpwr vgnd scs8hd_fill_2
XFILLER_24_175 vgnd vpwr scs8hd_decap_12
XFILLER_21_97 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_15.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_6 vgnd vpwr scs8hd_decap_3
XANTENNA__117__A _106_/X vgnd vpwr scs8hd_diode_2
X_129_ _129_/A _147_/A vgnd vpwr scs8hd_buf_1
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _180_/A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _174_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_101 vpwr vgnd scs8hd_fill_2
XFILLER_21_123 vgnd vpwr scs8hd_decap_3
XFILLER_21_156 vpwr vgnd scs8hd_fill_2
XFILLER_29_245 vgnd vpwr scs8hd_decap_8
Xmem_bottom_track_7.LATCH_1_.latch data_in _178_/A _119_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_64 vpwr vgnd scs8hd_fill_2
XFILLER_16_86 vgnd vpwr scs8hd_decap_4
XFILLER_8_105 vpwr vgnd scs8hd_fill_2
XFILLER_8_138 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_3_ mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_12_145 vgnd vpwr scs8hd_decap_6
XFILLER_16_97 vpwr vgnd scs8hd_fill_2
XFILLER_7_182 vgnd vpwr scs8hd_fill_1
XFILLER_34_270 vgnd vpwr scs8hd_decap_4
XFILLER_26_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_15.LATCH_1_.latch_SLEEPB _168_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _201_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_251 vgnd vpwr scs8hd_decap_12
XFILLER_27_85 vgnd vpwr scs8hd_fill_1
Xmem_left_track_7.LATCH_0_.latch data_in _197_/A _156_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_141 vgnd vpwr scs8hd_decap_12
XANTENNA__130__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_56 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _198_/Y vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_11.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_22_251 vgnd vpwr scs8hd_decap_12
XFILLER_8_3 vgnd vpwr scs8hd_decap_3
XFILLER_9_266 vgnd vpwr scs8hd_decap_8
XANTENNA__125__A _106_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _124_/Y vgnd vpwr scs8hd_diode_2
XFILLER_39_181 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_10_210 vgnd vpwr scs8hd_decap_4
X_162_ _155_/X _162_/B _162_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_24_53 vgnd vpwr scs8hd_fill_1
X_231_ _231_/A chanx_left_out[3] vgnd vpwr scs8hd_buf_2
XFILLER_10_276 vgnd vpwr scs8hd_fill_1
XFILLER_37_118 vpwr vgnd scs8hd_fill_2
XFILLER_1_46 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _176_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_10_22 vpwr vgnd scs8hd_fill_2
XFILLER_27_184 vgnd vpwr scs8hd_decap_12
XFILLER_42_187 vgnd vpwr scs8hd_decap_12
X_145_ _145_/A _145_/B _145_/Y vgnd vpwr scs8hd_nor2_4
X_214_ _214_/HI _214_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _220_/HI vgnd vpwr
+ scs8hd_diode_2
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_187 vgnd vpwr scs8hd_decap_12
XFILLER_30_102 vpwr vgnd scs8hd_fill_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_30_157 vgnd vpwr scs8hd_decap_12
XANTENNA__133__A _145_/A vgnd vpwr scs8hd_diode_2
XANTENNA__117__B _115_/X vgnd vpwr scs8hd_diode_2
X_128_ _106_/X _128_/B _128_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_202 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_3 vgnd vpwr scs8hd_decap_4
XFILLER_38_235 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _182_/A mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_16_10 vpwr vgnd scs8hd_fill_2
XFILLER_16_43 vpwr vgnd scs8hd_fill_2
XFILLER_32_64 vpwr vgnd scs8hd_fill_2
XFILLER_32_20 vgnd vpwr scs8hd_decap_8
Xmem_bottom_track_15.LATCH_1_.latch data_in _186_/A _135_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__128__A _106_/X vgnd vpwr scs8hd_diode_2
XFILLER_41_208 vgnd vpwr scs8hd_decap_12
XFILLER_26_227 vgnd vpwr scs8hd_decap_12
XFILLER_27_53 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_5.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_40_263 vgnd vpwr scs8hd_decap_12
XFILLER_27_97 vpwr vgnd scs8hd_fill_2
XANTENNA__130__B _115_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_1_ mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_23_208 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _211_/HI _186_/Y mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_22 vgnd vpwr scs8hd_decap_6
XFILLER_22_263 vgnd vpwr scs8hd_decap_12
XFILLER_13_99 vpwr vgnd scs8hd_fill_2
XANTENNA__231__A _231_/A vgnd vpwr scs8hd_diode_2
XFILLER_38_96 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _190_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__125__B _124_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_245 vgnd vpwr scs8hd_decap_8
XANTENNA__141__A _147_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
X_230_ _230_/A chanx_left_out[4] vgnd vpwr scs8hd_buf_2
X_161_ _168_/C _162_/B _161_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__226__A _226_/A vgnd vpwr scs8hd_diode_2
XFILLER_24_32 vpwr vgnd scs8hd_fill_2
XFILLER_1_58 vgnd vpwr scs8hd_decap_3
XANTENNA__136__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_141 vgnd vpwr scs8hd_decap_12
XFILLER_28_108 vgnd vpwr scs8hd_decap_8
XFILLER_19_10 vpwr vgnd scs8hd_fill_2
XFILLER_19_54 vgnd vpwr scs8hd_fill_1
XFILLER_35_75 vpwr vgnd scs8hd_fill_2
XFILLER_35_53 vgnd vpwr scs8hd_decap_6
XFILLER_35_31 vgnd vpwr scs8hd_decap_4
XFILLER_27_196 vgnd vpwr scs8hd_decap_12
XFILLER_27_152 vpwr vgnd scs8hd_fill_2
XFILLER_42_199 vgnd vpwr scs8hd_decap_12
X_144_ _147_/A _145_/B _144_/Y vgnd vpwr scs8hd_nor2_4
X_213_ _213_/HI _213_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_2_251 vgnd vpwr scs8hd_decap_12
XFILLER_25_7 vgnd vpwr scs8hd_fill_1
XFILLER_18_163 vpwr vgnd scs8hd_fill_2
XFILLER_18_174 vgnd vpwr scs8hd_decap_8
XFILLER_18_185 vgnd vpwr scs8hd_decap_12
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_100 vpwr vgnd scs8hd_fill_2
XFILLER_21_44 vpwr vgnd scs8hd_fill_2
XFILLER_24_199 vgnd vpwr scs8hd_decap_12
XFILLER_21_77 vpwr vgnd scs8hd_fill_2
XFILLER_30_169 vgnd vpwr scs8hd_decap_12
XFILLER_30_125 vgnd vpwr scs8hd_fill_1
XPHY_8 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_177 vgnd vpwr scs8hd_decap_6
XFILLER_7_68 vpwr vgnd scs8hd_fill_2
XANTENNA__133__B _131_/B vgnd vpwr scs8hd_diode_2
X_127_ _096_/X _128_/B _127_/Y vgnd vpwr scs8hd_nor2_4
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _243_/A vgnd vpwr scs8hd_inv_1
XFILLER_21_114 vpwr vgnd scs8hd_fill_2
XFILLER_29_258 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_12_125 vpwr vgnd scs8hd_fill_2
XANTENNA__234__A _234_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_43 vgnd vpwr scs8hd_fill_1
XFILLER_32_32 vgnd vpwr scs8hd_decap_4
XANTENNA__144__A _147_/A vgnd vpwr scs8hd_diode_2
XANTENNA__128__B _128_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_184 vgnd vpwr scs8hd_decap_12
XFILLER_7_162 vgnd vpwr scs8hd_decap_8
XFILLER_26_239 vgnd vpwr scs8hd_decap_12
XANTENNA__229__A _229_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_154 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_3.LATCH_1_.latch data_in _174_/A _111_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__130__C _134_/C vgnd vpwr scs8hd_diode_2
XFILLER_31_220 vgnd vpwr scs8hd_decap_12
XANTENNA__139__A _160_/C vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _204_/A mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_102 vpwr vgnd scs8hd_fill_2
XFILLER_1_113 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ _185_/A mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_13_220 vgnd vpwr scs8hd_decap_12
Xmem_left_track_3.LATCH_0_.latch data_in _193_/A _148_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__141__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_13.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_39_161 vgnd vpwr scs8hd_decap_12
XFILLER_40_32 vgnd vpwr scs8hd_decap_12
XFILLER_6_227 vgnd vpwr scs8hd_decap_12
X_160_ _122_/A _113_/Y _160_/C _153_/D _162_/B vgnd vpwr scs8hd_or4_4
XFILLER_24_88 vgnd vpwr scs8hd_fill_1
XANTENNA__242__A _242_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_109 vpwr vgnd scs8hd_fill_2
XANTENNA__136__B _134_/X vgnd vpwr scs8hd_diode_2
XANTENNA__152__A _129_/A vgnd vpwr scs8hd_diode_2
XFILLER_36_175 vgnd vpwr scs8hd_decap_12
XFILLER_3_208 vgnd vpwr scs8hd_decap_12
XFILLER_19_33 vpwr vgnd scs8hd_fill_2
XFILLER_19_88 vpwr vgnd scs8hd_fill_2
XFILLER_42_156 vgnd vpwr scs8hd_decap_12
X_212_ _212_/HI _212_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__237__A _237_/A vgnd vpwr scs8hd_diode_2
X_143_ _115_/A _123_/B _143_/C _109_/A _145_/B vgnd vpwr scs8hd_or4_4
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_32_9 vgnd vpwr scs8hd_decap_8
XFILLER_2_263 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ _189_/Y mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_33_123 vpwr vgnd scs8hd_fill_2
XFILLER_33_112 vgnd vpwr scs8hd_decap_4
XFILLER_18_7 vpwr vgnd scs8hd_fill_2
XFILLER_18_197 vgnd vpwr scs8hd_decap_12
XANTENNA__147__A _147_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_2_80 vgnd vpwr scs8hd_decap_12
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_145 vgnd vpwr scs8hd_decap_4
XFILLER_21_23 vpwr vgnd scs8hd_fill_2
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_15_101 vpwr vgnd scs8hd_fill_2
XFILLER_15_123 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_3.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_5_ vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_15_145 vpwr vgnd scs8hd_fill_2
X_126_ _126_/A _123_/B _123_/C _171_/A _128_/B vgnd vpwr scs8hd_or4_4
XFILLER_38_215 vgnd vpwr scs8hd_decap_12
XFILLER_16_23 vpwr vgnd scs8hd_fill_2
XFILLER_12_104 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_13.LATCH_0_.latch_SLEEPB _133_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__144__B _145_/B vgnd vpwr scs8hd_diode_2
XFILLER_7_174 vgnd vpwr scs8hd_decap_8
XFILLER_11_181 vpwr vgnd scs8hd_fill_2
XFILLER_7_196 vgnd vpwr scs8hd_decap_12
XANTENNA__160__A _122_/A vgnd vpwr scs8hd_diode_2
X_109_ _109_/A _171_/A vgnd vpwr scs8hd_buf_1
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[7] mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_34_251 vgnd vpwr scs8hd_decap_4
XFILLER_27_77 vpwr vgnd scs8hd_fill_2
XFILLER_25_262 vgnd vpwr scs8hd_decap_12
XFILLER_40_276 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _178_/A mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_166 vgnd vpwr scs8hd_decap_12
XANTENNA__130__D _168_/A vgnd vpwr scs8hd_diode_2
XFILLER_31_232 vgnd vpwr scs8hd_decap_12
XANTENNA__155__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_16_251 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_11.LATCH_1_.latch data_in _182_/A _127_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_210 vgnd vpwr scs8hd_decap_4
XFILLER_13_35 vpwr vgnd scs8hd_fill_2
XFILLER_13_57 vpwr vgnd scs8hd_fill_2
XFILLER_13_79 vgnd vpwr scs8hd_decap_4
XFILLER_22_276 vgnd vpwr scs8hd_fill_1
XFILLER_1_136 vgnd vpwr scs8hd_decap_4
XFILLER_1_147 vgnd vpwr scs8hd_decap_12
XFILLER_13_232 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _213_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _177_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_258 vpwr vgnd scs8hd_fill_2
XFILLER_0_180 vgnd vpwr scs8hd_decap_6
XFILLER_5_91 vgnd vpwr scs8hd_decap_12
XFILLER_39_184 vgnd vpwr scs8hd_decap_12
XFILLER_39_173 vgnd vpwr scs8hd_decap_8
XFILLER_24_45 vpwr vgnd scs8hd_fill_2
XFILLER_24_67 vgnd vpwr scs8hd_fill_1
XFILLER_40_44 vgnd vpwr scs8hd_decap_12
XFILLER_6_239 vgnd vpwr scs8hd_decap_12
XFILLER_6_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_11.LATCH_1_.latch_SLEEPB _127_/Y vgnd vpwr scs8hd_diode_2
XFILLER_36_187 vgnd vpwr scs8hd_decap_12
XFILLER_36_154 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_17.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_14 vpwr vgnd scs8hd_fill_2
XFILLER_10_36 vgnd vpwr scs8hd_fill_1
XFILLER_10_69 vpwr vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ _207_/A mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_19_67 vpwr vgnd scs8hd_fill_2
XFILLER_42_168 vgnd vpwr scs8hd_decap_12
XFILLER_35_99 vpwr vgnd scs8hd_fill_2
XFILLER_35_88 vgnd vpwr scs8hd_decap_4
X_142_ _145_/A _142_/B _142_/Y vgnd vpwr scs8hd_nor2_4
X_211_ _211_/HI _211_/LO vgnd vpwr scs8hd_conb_1
XANTENNA__147__B _147_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.tap_buf4_0_.scs8hd_inv_1 mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ _227_/A vgnd vpwr scs8hd_inv_1
XFILLER_18_132 vpwr vgnd scs8hd_fill_2
XANTENNA__163__A _122_/A vgnd vpwr scs8hd_diode_2
XFILLER_32_190 vgnd vpwr scs8hd_decap_12
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_135 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _200_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_21_57 vpwr vgnd scs8hd_fill_2
X_125_ _106_/X _124_/B _125_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_15 vpwr vgnd scs8hd_fill_2
XFILLER_30_7 vgnd vpwr scs8hd_decap_12
XFILLER_38_227 vgnd vpwr scs8hd_decap_8
XANTENNA__158__A _168_/C vgnd vpwr scs8hd_diode_2
XFILLER_16_68 vpwr vgnd scs8hd_fill_2
XFILLER_8_109 vgnd vpwr scs8hd_decap_3
XFILLER_35_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _179_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_left_track_7.tap_buf4_0_.scs8hd_inv_1 mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ _231_/A vgnd vpwr scs8hd_inv_1
XFILLER_7_131 vgnd vpwr scs8hd_decap_12
X_108_ address[1] enable _109_/A vgnd vpwr scs8hd_nand2_4
XANTENNA__160__B _113_/Y vgnd vpwr scs8hd_diode_2
XFILLER_21_3 vpwr vgnd scs8hd_fill_2
XFILLER_34_274 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _183_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_91 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _191_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_25_274 vgnd vpwr scs8hd_decap_3
XFILLER_4_178 vgnd vpwr scs8hd_decap_12
XPHY_280 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_263 vgnd vpwr scs8hd_decap_12
XANTENNA__171__A _171_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_159 vgnd vpwr scs8hd_decap_12
XFILLER_38_77 vgnd vpwr scs8hd_fill_1
Xmux_left_track_15.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[6] mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _209_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA__166__A address[3] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_196 vgnd vpwr scs8hd_decap_12
XFILLER_39_130 vpwr vgnd scs8hd_fill_2
XFILLER_40_56 vgnd vpwr scs8hd_decap_12
XFILLER_10_258 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _210_/HI _184_/Y mux_bottom_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ _181_/A mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_36_199 vgnd vpwr scs8hd_decap_12
XFILLER_36_166 vgnd vpwr scs8hd_decap_6
XFILLER_10_26 vgnd vpwr scs8hd_decap_4
XFILLER_10_48 vpwr vgnd scs8hd_fill_2
XFILLER_42_125 vgnd vpwr scs8hd_decap_12
XFILLER_19_57 vpwr vgnd scs8hd_fill_2
X_141_ _147_/A _142_/B _141_/Y vgnd vpwr scs8hd_nor2_4
X_210_ _210_/HI _210_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_276 vgnd vpwr scs8hd_fill_1
XFILLER_18_111 vgnd vpwr scs8hd_decap_3
XFILLER_33_136 vgnd vpwr scs8hd_decap_12
XANTENNA__163__B _113_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_93 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _221_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _193_/A vgnd vpwr
+ scs8hd_diode_2
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_21_14 vpwr vgnd scs8hd_fill_2
XFILLER_30_128 vpwr vgnd scs8hd_fill_2
XFILLER_30_106 vpwr vgnd scs8hd_fill_2
XFILLER_15_114 vpwr vgnd scs8hd_fill_2
XFILLER_15_158 vpwr vgnd scs8hd_fill_2
XFILLER_15_169 vpwr vgnd scs8hd_fill_2
XFILLER_30_139 vgnd vpwr scs8hd_decap_12
X_124_ _096_/X _124_/B _124_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_7_49 vpwr vgnd scs8hd_fill_2
XFILLER_23_7 vgnd vpwr scs8hd_fill_1
XFILLER_16_6 vpwr vgnd scs8hd_fill_2
XANTENNA__158__B _158_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__174__A _174_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_7.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_21_139 vpwr vgnd scs8hd_fill_2
XFILLER_16_47 vpwr vgnd scs8hd_fill_2
XFILLER_32_79 vgnd vpwr scs8hd_decap_12
XFILLER_32_46 vgnd vpwr scs8hd_fill_1
XFILLER_7_143 vgnd vpwr scs8hd_decap_12
X_107_ _106_/X _105_/B _107_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__160__C _160_/C vgnd vpwr scs8hd_diode_2
XFILLER_14_3 vpwr vgnd scs8hd_fill_2
XANTENNA__169__A _168_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_11.LATCH_0_.latch_SLEEPB _162_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_57 vpwr vgnd scs8hd_fill_2
XFILLER_27_24 vgnd vpwr scs8hd_fill_1
XFILLER_25_253 vpwr vgnd scs8hd_fill_2
XFILLER_25_220 vgnd vpwr scs8hd_decap_12
XFILLER_4_17 vgnd vpwr scs8hd_decap_12
XPHY_281 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_270 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_245 vgnd vpwr scs8hd_decap_12
XANTENNA__171__B _168_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_48 vgnd vpwr scs8hd_decap_3
XFILLER_8_8 vpwr vgnd scs8hd_fill_2
XFILLER_38_89 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[7] vgnd vpwr scs8hd_diode_2
XFILLER_13_245 vgnd vpwr scs8hd_decap_12
XFILLER_0_193 vgnd vpwr scs8hd_fill_1
XANTENNA__166__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__182__A _182_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_5.LATCH_0_.latch_SLEEPB _117_/Y vgnd vpwr scs8hd_diode_2
XFILLER_10_215 vgnd vpwr scs8hd_decap_12
Xmux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _202_/A mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_40_68 vgnd vpwr scs8hd_decap_12
XFILLER_14_91 vgnd vpwr scs8hd_fill_1
Xmux_left_track_13.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[5] mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_36_112 vgnd vpwr scs8hd_decap_4
XANTENNA__177__A _177_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ _183_/A mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_27_101 vpwr vgnd scs8hd_fill_2
XFILLER_19_25 vpwr vgnd scs8hd_fill_2
XFILLER_42_137 vgnd vpwr scs8hd_decap_12
XFILLER_35_35 vgnd vpwr scs8hd_fill_1
XFILLER_27_156 vpwr vgnd scs8hd_fill_2
XFILLER_27_123 vgnd vpwr scs8hd_fill_1
X_140_ _115_/A _123_/B _143_/C _153_/D _142_/B vgnd vpwr scs8hd_or4_4
XFILLER_18_123 vpwr vgnd scs8hd_fill_2
XFILLER_18_145 vpwr vgnd scs8hd_fill_2
XFILLER_18_167 vgnd vpwr scs8hd_decap_4
XFILLER_33_148 vgnd vpwr scs8hd_decap_12
XFILLER_33_104 vpwr vgnd scs8hd_fill_2
XFILLER_25_90 vgnd vpwr scs8hd_decap_3
XANTENNA_mem_bottom_track_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__163__C _160_/C vgnd vpwr scs8hd_diode_2
XFILLER_24_104 vgnd vpwr scs8hd_decap_4
XFILLER_24_126 vgnd vpwr scs8hd_decap_3
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _221_/HI _206_/Y mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_23_170 vgnd vpwr scs8hd_decap_12
X_123_ _126_/A _123_/B _123_/C _168_/A _124_/B vgnd vpwr scs8hd_or4_4
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_11_92 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_3_ vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_118 vpwr vgnd scs8hd_fill_2
XANTENNA__190__A _190_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ _187_/Y mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_12_118 vgnd vpwr scs8hd_decap_4
XFILLER_12_129 vgnd vpwr scs8hd_fill_1
XFILLER_32_58 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[4] vgnd vpwr scs8hd_diode_2
XFILLER_28_251 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_3.LATCH_1_.latch_SLEEPB _111_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_111 vgnd vpwr scs8hd_fill_1
XFILLER_11_151 vpwr vgnd scs8hd_fill_2
XFILLER_11_173 vgnd vpwr scs8hd_decap_8
XANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB _159_/Y vgnd vpwr scs8hd_diode_2
X_106_ address[0] _106_/X vgnd vpwr scs8hd_buf_1
XFILLER_7_155 vgnd vpwr scs8hd_decap_4
XFILLER_11_184 vgnd vpwr scs8hd_decap_12
XANTENNA__160__D _153_/D vgnd vpwr scs8hd_diode_2
XFILLER_22_91 vgnd vpwr scs8hd_fill_1
XANTENNA__169__B _168_/B vgnd vpwr scs8hd_diode_2
XFILLER_34_276 vgnd vpwr scs8hd_fill_1
XANTENNA__185__A _185_/A vgnd vpwr scs8hd_diode_2
XFILLER_27_36 vpwr vgnd scs8hd_fill_2
XFILLER_27_14 vpwr vgnd scs8hd_fill_2
XFILLER_25_232 vgnd vpwr scs8hd_decap_12
XFILLER_40_202 vgnd vpwr scs8hd_decap_12
XANTENNA__095__A address[0] vgnd vpwr scs8hd_diode_2
XFILLER_4_29 vpwr vgnd scs8hd_fill_2
XFILLER_16_276 vgnd vpwr scs8hd_fill_1
XPHY_282 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_271 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_260 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_257 vgnd vpwr scs8hd_decap_12
XANTENNA__171__C _155_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_1_106 vgnd vpwr scs8hd_decap_4
XFILLER_38_35 vgnd vpwr scs8hd_decap_12
XFILLER_1_117 vgnd vpwr scs8hd_decap_3
XFILLER_13_257 vgnd vpwr scs8hd_decap_12
XANTENNA__166__C address[4] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _176_/A mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_72 vpwr vgnd scs8hd_fill_2
XFILLER_10_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_13.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_13_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_5_220 vgnd vpwr scs8hd_decap_12
XFILLER_39_6 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_7.LATCH_1_.latch_SLEEPB _154_/Y vgnd vpwr scs8hd_diode_2
Xmem_left_track_7.LATCH_1_.latch data_in _196_/A _154_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA__193__A _193_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _201_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_135 vpwr vgnd scs8hd_fill_2
XFILLER_19_37 vpwr vgnd scs8hd_fill_2
XFILLER_42_149 vgnd vpwr scs8hd_decap_6
XFILLER_33_116 vgnd vpwr scs8hd_fill_1
XFILLER_18_102 vgnd vpwr scs8hd_decap_3
XFILLER_41_171 vgnd vpwr scs8hd_decap_12
XPHY_80 vgnd vpwr scs8hd_decap_3
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__163__D _109_/A vgnd vpwr scs8hd_diode_2
X_199_ _199_/A _199_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__188__A _188_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_3 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _216_/HI _180_/Y mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_24_149 vgnd vpwr scs8hd_fill_1
Xmux_left_track_11.INVTX1_0_.scs8hd_inv_1 chany_bottom_in[4] mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_27 vpwr vgnd scs8hd_fill_2
XANTENNA__098__A address[2] vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_13.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_23_182 vgnd vpwr scs8hd_fill_1
XFILLER_11_71 vpwr vgnd scs8hd_fill_2
X_122_ _122_/A _126_/A vgnd vpwr scs8hd_buf_1
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ _205_/A mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_29_208 vgnd vpwr scs8hd_decap_12
XFILLER_12_108 vgnd vpwr scs8hd_fill_1
XFILLER_16_27 vpwr vgnd scs8hd_fill_2
XFILLER_20_163 vgnd vpwr scs8hd_decap_8
XFILLER_20_174 vgnd vpwr scs8hd_decap_12
XFILLER_28_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _176_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_11_196 vgnd vpwr scs8hd_decap_12
X_105_ _096_/X _105_/B _105_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__169__C _155_/X vgnd vpwr scs8hd_diode_2
XFILLER_8_83 vgnd vpwr scs8hd_decap_8
XPHY_261 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_250 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_283 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_272 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _203_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__196__A _196_/A vgnd vpwr scs8hd_diode_2
XFILLER_13_28 vgnd vpwr scs8hd_fill_1
XFILLER_38_47 vgnd vpwr scs8hd_decap_12
XFILLER_13_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _214_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__166__D _138_/B vgnd vpwr scs8hd_diode_2
XFILLER_5_62 vgnd vpwr scs8hd_fill_1
XFILLER_8_251 vgnd vpwr scs8hd_decap_12
XFILLER_24_49 vgnd vpwr scs8hd_decap_4
XFILLER_40_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_5_232 vgnd vpwr scs8hd_decap_12
XFILLER_36_125 vpwr vgnd scs8hd_fill_2
XFILLER_10_18 vpwr vgnd scs8hd_fill_2
XFILLER_27_114 vpwr vgnd scs8hd_fill_2
XFILLER_42_106 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _178_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_202 vgnd vpwr scs8hd_decap_12
XPHY_81 vgnd vpwr scs8hd_decap_3
XPHY_70 vgnd vpwr scs8hd_decap_3
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_198_ _198_/A _198_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _182_/A vgnd
+ vpwr scs8hd_diode_2
Xmux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _209_/HI _182_/Y mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _190_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ _179_/A mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_15_128 vpwr vgnd scs8hd_fill_2
XFILLER_7_19 vpwr vgnd scs8hd_fill_2
X_121_ address[3] _122_/A vgnd vpwr scs8hd_inv_8
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _217_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__199__A _199_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_220 vgnd vpwr scs8hd_decap_12
XFILLER_20_186 vgnd vpwr scs8hd_decap_12
Xmem_left_track_17.LATCH_0_.latch data_in _207_/A _171_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_104_ _115_/A _123_/B _123_/C _168_/A _105_/B vgnd vpwr scs8hd_or4_4
XFILLER_22_93 vgnd vpwr scs8hd_decap_6
XFILLER_19_220 vgnd vpwr scs8hd_decap_12
XFILLER_19_253 vpwr vgnd scs8hd_fill_2
XFILLER_8_51 vgnd vpwr scs8hd_decap_4
XFILLER_6_190 vgnd vpwr scs8hd_decap_12
XFILLER_8_62 vgnd vpwr scs8hd_decap_6
XFILLER_40_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_3.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_25_245 vgnd vpwr scs8hd_decap_8
XFILLER_4_105 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_16_212 vpwr vgnd scs8hd_fill_2
XPHY_284 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_273 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_262 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_251 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_240 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_60 vgnd vpwr scs8hd_fill_1
XFILLER_3_171 vgnd vpwr scs8hd_decap_12
XFILLER_12_3 vpwr vgnd scs8hd_fill_2
XFILLER_22_215 vgnd vpwr scs8hd_decap_12
XFILLER_38_59 vgnd vpwr scs8hd_decap_12
XFILLER_38_15 vgnd vpwr scs8hd_decap_12
XFILLER_9_208 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _210_/HI vgnd
+ vpwr scs8hd_diode_2
XFILLER_8_263 vgnd vpwr scs8hd_decap_12
XFILLER_39_134 vgnd vpwr scs8hd_decap_12
XFILLER_39_123 vgnd vpwr scs8hd_decap_4
XFILLER_39_112 vpwr vgnd scs8hd_fill_2
XFILLER_39_101 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _192_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_40_27 vgnd vpwr scs8hd_decap_4
XFILLER_14_83 vpwr vgnd scs8hd_fill_2
XFILLER_30_60 vpwr vgnd scs8hd_fill_2
XFILLER_42_118 vgnd vpwr scs8hd_decap_6
XFILLER_35_38 vgnd vpwr scs8hd_decap_4
XPHY_82 vgnd vpwr scs8hd_decap_3
XPHY_71 vgnd vpwr scs8hd_decap_3
XPHY_60 vgnd vpwr scs8hd_decap_3
Xmux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _200_/A mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_41_184 vgnd vpwr scs8hd_decap_12
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
X_197_ _197_/A _197_/Y vgnd vpwr scs8hd_inv_8
XFILLER_32_140 vgnd vpwr scs8hd_decap_12
XFILLER_24_118 vgnd vpwr scs8hd_decap_8
Xmem_left_track_3.LATCH_1_.latch data_in _192_/A _147_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_21_18 vgnd vpwr scs8hd_decap_3
XFILLER_15_118 vpwr vgnd scs8hd_fill_2
X_120_ _106_/X _119_/B _120_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_184 vgnd vpwr scs8hd_decap_12
XFILLER_36_81 vgnd vpwr scs8hd_decap_8
XFILLER_14_151 vpwr vgnd scs8hd_fill_2
XFILLER_42_3 vgnd vpwr scs8hd_decap_12
XFILLER_37_232 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_32_39 vgnd vpwr scs8hd_decap_4
XFILLER_32_28 vgnd vpwr scs8hd_decap_3
XFILLER_20_132 vpwr vgnd scs8hd_fill_2
XFILLER_20_198 vgnd vpwr scs8hd_decap_12
XFILLER_28_276 vgnd vpwr scs8hd_fill_1
XFILLER_7_114 vgnd vpwr scs8hd_decap_8
X_103_ _153_/D _168_/A vgnd vpwr scs8hd_buf_1
XFILLER_22_83 vgnd vpwr scs8hd_decap_6
XFILLER_34_202 vgnd vpwr scs8hd_decap_12
Xmux_left_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _220_/HI _204_/Y mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_19_232 vgnd vpwr scs8hd_decap_12
XFILLER_8_41 vgnd vpwr scs8hd_fill_1
XFILLER_8_96 vgnd vpwr scs8hd_decap_6
XFILLER_40_227 vgnd vpwr scs8hd_decap_12
XFILLER_4_117 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ _185_/Y mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_left_track_15.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XPHY_285 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_274 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_263 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_252 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_241 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_230 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_22_227 vgnd vpwr scs8hd_decap_12
XFILLER_30_271 vgnd vpwr scs8hd_decap_4
XFILLER_38_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_120 vgnd vpwr scs8hd_decap_4
XFILLER_0_197 vpwr vgnd scs8hd_fill_2
XFILLER_28_93 vpwr vgnd scs8hd_fill_2
XFILLER_28_71 vgnd vpwr scs8hd_decap_4
XFILLER_28_60 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_11.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_5_31 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_15.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_15_ mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_39_157 vpwr vgnd scs8hd_fill_2
XFILLER_39_146 vgnd vpwr scs8hd_decap_8
XFILLER_24_18 vgnd vpwr scs8hd_decap_12
XFILLER_38_190 vgnd vpwr scs8hd_decap_12
XFILLER_30_83 vgnd vpwr scs8hd_fill_1
XFILLER_5_245 vgnd vpwr scs8hd_decap_12
XANTENNA__101__A enable vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_1_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_19_29 vpwr vgnd scs8hd_fill_2
XFILLER_35_182 vgnd vpwr scs8hd_fill_1
XFILLER_35_171 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _174_/A mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_4_6 vpwr vgnd scs8hd_fill_2
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_127 vgnd vpwr scs8hd_decap_3
XFILLER_18_149 vpwr vgnd scs8hd_fill_2
XPHY_83 vgnd vpwr scs8hd_decap_3
XPHY_72 vgnd vpwr scs8hd_decap_3
XFILLER_33_119 vgnd vpwr scs8hd_decap_3
XFILLER_33_108 vpwr vgnd scs8hd_fill_2
XPHY_61 vgnd vpwr scs8hd_decap_3
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_50 vgnd vpwr scs8hd_decap_3
XFILLER_41_196 vgnd vpwr scs8hd_decap_12
X_196_ _196_/A _196_/Y vgnd vpwr scs8hd_inv_8
Xmux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ _240_/A vgnd vpwr scs8hd_inv_1
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_24_108 vgnd vpwr scs8hd_fill_1
XFILLER_32_152 vgnd vpwr scs8hd_fill_1
XFILLER_23_196 vgnd vpwr scs8hd_decap_12
XFILLER_2_3 vpwr vgnd scs8hd_fill_2
XFILLER_36_60 vgnd vpwr scs8hd_decap_8
XFILLER_36_93 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_14_163 vgnd vpwr scs8hd_decap_12
X_179_ _179_/A _179_/Y vgnd vpwr scs8hd_inv_8
XFILLER_35_3 vpwr vgnd scs8hd_fill_2
XFILLER_20_111 vpwr vgnd scs8hd_fill_2
XFILLER_28_211 vgnd vpwr scs8hd_decap_3
Xmux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _215_/HI _178_/Y mux_bottom_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_11_111 vpwr vgnd scs8hd_fill_2
XFILLER_11_155 vpwr vgnd scs8hd_fill_2
XFILLER_7_159 vgnd vpwr scs8hd_fill_1
XFILLER_7_126 vgnd vpwr scs8hd_decap_3
X_102_ address[1] _102_/B _153_/D vgnd vpwr scs8hd_or2_4
XFILLER_22_62 vpwr vgnd scs8hd_fill_2
XFILLER_34_258 vgnd vpwr scs8hd_decap_12
XFILLER_27_18 vgnd vpwr scs8hd_decap_6
Xmux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ _203_/A mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_40_239 vgnd vpwr scs8hd_decap_12
XFILLER_25_258 vpwr vgnd scs8hd_fill_2
XFILLER_4_129 vgnd vpwr scs8hd_decap_12
XFILLER_17_73 vgnd vpwr scs8hd_fill_1
XPHY_275 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_264 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_253 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_242 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_231 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_220 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_184 vgnd vpwr scs8hd_decap_12
XANTENNA__104__A _115_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _200_/Y vgnd vpwr
+ scs8hd_diode_2
Xmem_left_track_13.LATCH_0_.latch data_in _203_/A _165_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_22_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_187 vgnd vpwr scs8hd_decap_6
XFILLER_5_10 vpwr vgnd scs8hd_fill_2
XFILLER_8_276 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_9.LATCH_0_.latch data_in _181_/A _125_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_87 vpwr vgnd scs8hd_fill_2
XFILLER_5_76 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _179_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ _207_/Y mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_left_track_11.tap_buf4_0_.scs8hd_inv_1 mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ _229_/A vgnd vpwr scs8hd_inv_1
XFILLER_14_30 vgnd vpwr scs8hd_fill_1
XFILLER_14_63 vgnd vpwr scs8hd_fill_1
XFILLER_39_60 vgnd vpwr scs8hd_fill_1
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _183_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_15.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_7.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_27_139 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_13.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_13_ mux_bottom_track_13.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
XANTENNA__202__A _202_/A vgnd vpwr scs8hd_diode_2
XPHY_84 vgnd vpwr scs8hd_decap_3
XPHY_73 vgnd vpwr scs8hd_decap_3
XPHY_62 vgnd vpwr scs8hd_decap_3
XFILLER_26_150 vgnd vpwr scs8hd_decap_3
XPHY_51 vgnd vpwr scs8hd_decap_3
XFILLER_25_95 vgnd vpwr scs8hd_decap_3
XFILLER_25_73 vpwr vgnd scs8hd_fill_2
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vpwr scs8hd_decap_3
X_195_ _195_/A _195_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XANTENNA__112__A _106_/X vgnd vpwr scs8hd_diode_2
Xmux_left_track_3.tap_buf4_0_.scs8hd_inv_1 mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ _233_/A vgnd vpwr scs8hd_inv_1
XFILLER_23_153 vgnd vpwr scs8hd_fill_1
XFILLER_11_53 vpwr vgnd scs8hd_fill_2
XFILLER_11_75 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _202_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_14_175 vgnd vpwr scs8hd_decap_12
XANTENNA__107__A _106_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
X_178_ _178_/A _178_/Y vgnd vpwr scs8hd_inv_8
XFILLER_37_245 vgnd vpwr scs8hd_decap_12
XFILLER_28_3 vpwr vgnd scs8hd_fill_2
XFILLER_20_145 vpwr vgnd scs8hd_fill_2
X_101_ enable _102_/B vgnd vpwr scs8hd_inv_8
XFILLER_11_134 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ _177_/A mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_19_245 vgnd vpwr scs8hd_decap_8
XFILLER_34_215 vgnd vpwr scs8hd_decap_12
XFILLER_8_32 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _181_/A vgnd
+ vpwr scs8hd_diode_2
XPHY_243 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_232 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_221 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_210 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _185_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_16_204 vgnd vpwr scs8hd_decap_8
XFILLER_16_215 vgnd vpwr scs8hd_decap_12
XFILLER_17_52 vpwr vgnd scs8hd_fill_2
XFILLER_17_85 vpwr vgnd scs8hd_fill_2
XFILLER_17_96 vpwr vgnd scs8hd_fill_2
XPHY_276 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_265 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_254 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_84 vgnd vpwr scs8hd_decap_3
XFILLER_33_73 vgnd vpwr scs8hd_decap_6
XFILLER_33_40 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _193_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_3_196 vgnd vpwr scs8hd_decap_12
XANTENNA__104__B _123_/B vgnd vpwr scs8hd_diode_2
XANTENNA__120__A _106_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_251 vgnd vpwr scs8hd_decap_4
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ _198_/A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _142_/Y vgnd vpwr scs8hd_diode_2
XANTENNA__205__A _205_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ _236_/A vgnd vpwr scs8hd_inv_1
XFILLER_28_84 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _215_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_8_211 vgnd vpwr scs8hd_decap_3
XFILLER_12_251 vgnd vpwr scs8hd_decap_12
XANTENNA__115__A _115_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ _181_/Y mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_10_3 vpwr vgnd scs8hd_fill_2
Xmem_bottom_track_17.LATCH_0_.latch data_in _189_/A _142_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_5_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_94 vgnd vpwr scs8hd_decap_3
XFILLER_36_129 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_3.LATCH_0_.latch_SLEEPB _148_/Y vgnd vpwr scs8hd_diode_2
XFILLER_27_118 vpwr vgnd scs8hd_fill_2
XFILLER_35_184 vgnd vpwr scs8hd_decap_12
XFILLER_35_19 vgnd vpwr scs8hd_decap_12
XFILLER_2_239 vgnd vpwr scs8hd_decap_12
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_18_107 vpwr vgnd scs8hd_fill_2
XPHY_85 vgnd vpwr scs8hd_decap_3
XFILLER_41_110 vgnd vpwr scs8hd_decap_12
XPHY_74 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_decap_3
XPHY_52 vgnd vpwr scs8hd_decap_3
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_41_62 vgnd vpwr scs8hd_decap_12
XFILLER_41_51 vgnd vpwr scs8hd_decap_8
X_194_ _194_/A _194_/Y vgnd vpwr scs8hd_inv_8
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XANTENNA__112__B _110_/X vgnd vpwr scs8hd_diode_2
XFILLER_32_154 vgnd vpwr scs8hd_decap_12
XFILLER_17_162 vpwr vgnd scs8hd_fill_2
XFILLER_17_184 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_7.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_23_132 vgnd vpwr scs8hd_decap_4
XANTENNA_mem_bottom_track_15.LATCH_1_.latch_SLEEPB _135_/Y vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_11.INVTX1_0_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _195_/A vgnd vpwr
+ scs8hd_diode_2
X_177_ _177_/A _177_/Y vgnd vpwr scs8hd_inv_8
XFILLER_14_187 vgnd vpwr scs8hd_decap_12
XANTENNA__107__B _105_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_5.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__123__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _222_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_9_180 vgnd vpwr scs8hd_decap_3
X_100_ _134_/C _123_/C vgnd vpwr scs8hd_buf_1
XFILLER_11_168 vgnd vpwr scs8hd_decap_3
XFILLER_19_257 vgnd vpwr scs8hd_decap_12
XFILLER_34_227 vgnd vpwr scs8hd_decap_12
XANTENNA__118__A _115_/A vgnd vpwr scs8hd_diode_2
XFILLER_8_55 vgnd vpwr scs8hd_fill_1
X_229_ _229_/A chanx_left_out[5] vgnd vpwr scs8hd_buf_2
XFILLER_40_3 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB _144_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_31 vpwr vgnd scs8hd_fill_2
XPHY_277 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_266 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_255 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_244 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_233 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_31_208 vgnd vpwr scs8hd_decap_12
XPHY_222 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_211 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_227 vgnd vpwr scs8hd_decap_12
XPHY_200 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_24_271 vgnd vpwr scs8hd_decap_4
XANTENNA__104__C _123_/C vgnd vpwr scs8hd_diode_2
XFILLER_12_7 vgnd vpwr scs8hd_fill_1
XANTENNA__120__B _119_/B vgnd vpwr scs8hd_diode_2
Xmux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _219_/HI _202_/Y mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_13_208 vgnd vpwr scs8hd_decap_12
XFILLER_21_230 vgnd vpwr scs8hd_decap_12
XFILLER_0_101 vgnd vpwr scs8hd_decap_12
XFILLER_0_145 vpwr vgnd scs8hd_fill_2
XFILLER_0_156 vgnd vpwr scs8hd_decap_12
XFILLER_28_30 vgnd vpwr scs8hd_fill_1
XFILLER_12_263 vgnd vpwr scs8hd_decap_12
XFILLER_5_34 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _211_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA__115__B _115_/B vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ _183_/Y mux_bottom_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_116 vgnd vpwr scs8hd_decap_6
XFILLER_39_105 vgnd vpwr scs8hd_decap_4
XANTENNA__131__A _147_/A vgnd vpwr scs8hd_diode_2
XFILLER_14_32 vpwr vgnd scs8hd_fill_2
XFILLER_14_87 vpwr vgnd scs8hd_fill_2
XFILLER_30_86 vgnd vpwr scs8hd_decap_4
XFILLER_30_64 vpwr vgnd scs8hd_fill_2
XFILLER_39_62 vgnd vpwr scs8hd_decap_12
XFILLER_36_108 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__126__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_35_196 vgnd vpwr scs8hd_decap_12
XFILLER_35_174 vgnd vpwr scs8hd_decap_8
Xmem_bottom_track_5.LATCH_0_.latch data_in _177_/A _117_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_64 vgnd vpwr scs8hd_decap_3
XPHY_53 vgnd vpwr scs8hd_decap_3
XFILLER_26_163 vgnd vpwr scs8hd_decap_12
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_42 vgnd vpwr scs8hd_decap_3
XFILLER_25_42 vgnd vpwr scs8hd_decap_3
XFILLER_25_53 vgnd vpwr scs8hd_decap_8
XFILLER_41_74 vgnd vpwr scs8hd_decap_12
XPHY_75 vgnd vpwr scs8hd_decap_3
X_193_ _193_/A _193_/Y vgnd vpwr scs8hd_inv_8
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mem_bottom_track_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[2] vgnd vpwr scs8hd_diode_2
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XFILLER_32_166 vgnd vpwr scs8hd_decap_12
XFILLER_17_141 vpwr vgnd scs8hd_fill_2
XFILLER_23_166 vpwr vgnd scs8hd_fill_2
XFILLER_11_88 vpwr vgnd scs8hd_fill_2
XFILLER_36_30 vgnd vpwr scs8hd_fill_1
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _172_/A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_14_199 vgnd vpwr scs8hd_decap_12
X_176_ _176_/A _176_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__B _123_/B vgnd vpwr scs8hd_diode_2
XFILLER_37_269 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_7_107 vgnd vpwr scs8hd_decap_4
XFILLER_22_43 vpwr vgnd scs8hd_fill_2
XFILLER_22_54 vpwr vgnd scs8hd_fill_2
XFILLER_34_239 vgnd vpwr scs8hd_decap_12
XFILLER_19_269 vgnd vpwr scs8hd_decap_8
XFILLER_42_261 vgnd vpwr scs8hd_decap_12
XFILLER_8_23 vgnd vpwr scs8hd_decap_8
XANTENNA__118__B _115_/B vgnd vpwr scs8hd_diode_2
X_228_ _228_/A chanx_left_out[6] vgnd vpwr scs8hd_buf_2
XANTENNA_mux_bottom_track_15.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_15_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA__134__A _126_/A vgnd vpwr scs8hd_diode_2
X_159_ _155_/X _158_/B _159_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_16_239 vgnd vpwr scs8hd_decap_12
XFILLER_17_65 vpwr vgnd scs8hd_fill_2
XPHY_278 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_267 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_256 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_245 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_53 vpwr vgnd scs8hd_fill_2
XPHY_234 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_223 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_212 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_201 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__104__D _168_/A vgnd vpwr scs8hd_diode_2
XANTENNA__129__A _129_/A vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _214_/HI _176_/Y mux_bottom_track_5.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_21_242 vpwr vgnd scs8hd_fill_2
XFILLER_0_168 vgnd vpwr scs8hd_decap_12
Xmux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ _201_/A mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_28_97 vpwr vgnd scs8hd_fill_2
XFILLER_28_42 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_15.LATCH_0_.latch_SLEEPB _169_/Y vgnd vpwr scs8hd_diode_2
XFILLER_5_46 vgnd vpwr scs8hd_decap_12
XANTENNA__131__B _131_/B vgnd vpwr scs8hd_diode_2
XANTENNA__115__C _123_/C vgnd vpwr scs8hd_diode_2
XFILLER_38_150 vgnd vpwr scs8hd_decap_3
XFILLER_14_22 vpwr vgnd scs8hd_fill_2
XFILLER_14_66 vpwr vgnd scs8hd_fill_2
XFILLER_30_43 vpwr vgnd scs8hd_fill_2
XFILLER_30_32 vpwr vgnd scs8hd_fill_2
XANTENNA__232__A _232_/A vgnd vpwr scs8hd_diode_2
XFILLER_39_74 vgnd vpwr scs8hd_decap_12
XFILLER_39_52 vpwr vgnd scs8hd_fill_2
XANTENNA__126__B _123_/B vgnd vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__142__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_41_123 vgnd vpwr scs8hd_decap_12
XPHY_76 vgnd vpwr scs8hd_decap_3
XPHY_65 vgnd vpwr scs8hd_decap_3
XFILLER_26_175 vgnd vpwr scs8hd_decap_12
XFILLER_26_142 vgnd vpwr scs8hd_decap_8
XANTENNA__227__A _227_/A vgnd vpwr scs8hd_diode_2
XPHY_54 vgnd vpwr scs8hd_decap_3
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _203_/Y vgnd vpwr
+ scs8hd_diode_2
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_32 vgnd vpwr scs8hd_decap_3
XPHY_43 vgnd vpwr scs8hd_decap_3
XFILLER_25_21 vgnd vpwr scs8hd_decap_6
XFILLER_25_65 vpwr vgnd scs8hd_fill_2
XFILLER_41_86 vgnd vpwr scs8hd_decap_12
X_192_ _192_/A _192_/Y vgnd vpwr scs8hd_inv_8
Xmux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ _205_/Y mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmem_bottom_track_13.LATCH_0_.latch data_in _185_/A _133_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_9_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _125_/Y vgnd vpwr scs8hd_diode_2
XFILLER_32_178 vgnd vpwr scs8hd_decap_12
XFILLER_32_123 vgnd vpwr scs8hd_decap_3
XANTENNA__137__A address[5] vgnd vpwr scs8hd_diode_2
XFILLER_17_175 vgnd vpwr scs8hd_decap_8
XFILLER_23_156 vgnd vpwr scs8hd_fill_1
XFILLER_11_23 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_11.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_2_7 vgnd vpwr scs8hd_decap_12
XFILLER_11_34 vpwr vgnd scs8hd_fill_2
XFILLER_14_123 vgnd vpwr scs8hd_decap_4
X_175_ _175_/A _175_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__C _123_/C vgnd vpwr scs8hd_diode_2
XFILLER_35_7 vgnd vpwr scs8hd_decap_12
XFILLER_9_160 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_13.LATCH_1_.latch_SLEEPB _164_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_115 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_28_215 vgnd vpwr scs8hd_decap_12
XFILLER_11_115 vgnd vpwr scs8hd_decap_4
XANTENNA__240__A _240_/A vgnd vpwr scs8hd_diode_2
XFILLER_42_273 vgnd vpwr scs8hd_decap_4
X_227_ _227_/A chanx_left_out[7] vgnd vpwr scs8hd_buf_2
XFILLER_8_79 vpwr vgnd scs8hd_fill_2
XANTENNA__118__C _123_/C vgnd vpwr scs8hd_diode_2
XFILLER_6_141 vgnd vpwr scs8hd_decap_12
XANTENNA__134__B _115_/B vgnd vpwr scs8hd_diode_2
X_158_ _168_/C _158_/B _158_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA_mux_bottom_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _178_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA__150__A _147_/A vgnd vpwr scs8hd_diode_2
XPHY_279 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_268 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__235__A _235_/A vgnd vpwr scs8hd_diode_2
XPHY_257 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_246 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_235 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_224 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_213 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _182_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_24_251 vgnd vpwr scs8hd_decap_4
XPHY_202 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_276 vgnd vpwr scs8hd_fill_1
XANTENNA__145__A _145_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_15.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_3.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_0_.scs8hd_inv_1/Y
+ _175_/A mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XANTENNA_mem_bottom_track_7.LATCH_1_.latch_SLEEPB _119_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _205_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_0_125 vgnd vpwr scs8hd_decap_12
XFILLER_12_276 vgnd vpwr scs8hd_fill_1
XANTENNA__115__D _168_/A vgnd vpwr scs8hd_diode_2
XFILLER_5_58 vgnd vpwr scs8hd_fill_1
XFILLER_5_14 vpwr vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_1_.latch data_in _206_/A _170_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
Xmux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ _196_/A mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_30_77 vgnd vpwr scs8hd_decap_6
XFILLER_39_86 vgnd vpwr scs8hd_decap_8
XFILLER_29_184 vgnd vpwr scs8hd_decap_12
XANTENNA__142__B _142_/B vgnd vpwr scs8hd_diode_2
XANTENNA__126__C _123_/C vgnd vpwr scs8hd_diode_2
Xmux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ _179_/Y mux_bottom_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_41_135 vgnd vpwr scs8hd_decap_12
XPHY_77 vgnd vpwr scs8hd_decap_3
XPHY_66 vgnd vpwr scs8hd_decap_3
XPHY_55 vgnd vpwr scs8hd_decap_3
XFILLER_26_187 vgnd vpwr scs8hd_decap_12
XPHY_11 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XPHY_44 vgnd vpwr scs8hd_decap_3
XFILLER_41_98 vgnd vpwr scs8hd_decap_12
X_191_ _191_/A _191_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__243__A _243_/A vgnd vpwr scs8hd_diode_2
XFILLER_1_220 vgnd vpwr scs8hd_decap_12
XFILLER_40_190 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _180_/A vgnd
+ vpwr scs8hd_diode_2
XANTENNA__153__A _126_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_102 vgnd vpwr scs8hd_decap_4
XFILLER_23_113 vpwr vgnd scs8hd_fill_2
XFILLER_11_57 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _184_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_36_54 vgnd vpwr scs8hd_decap_3
XFILLER_36_43 vgnd vpwr scs8hd_fill_1
XFILLER_36_32 vgnd vpwr scs8hd_decap_4
XANTENNA__238__A _238_/A vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_1.LATCH_0_.latch data_in _173_/A _107_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_102 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_left_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _192_/Y vgnd vpwr
+ scs8hd_diode_2
X_243_ _243_/A chany_bottom_out[0] vgnd vpwr scs8hd_buf_2
X_174_ _174_/A _174_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__123__D _168_/A vgnd vpwr scs8hd_diode_2
XFILLER_37_238 vgnd vpwr scs8hd_decap_6
XFILLER_28_7 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_11.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XANTENNA__148__A _145_/A vgnd vpwr scs8hd_diode_2
XFILLER_20_149 vgnd vpwr scs8hd_decap_4
XFILLER_28_227 vgnd vpwr scs8hd_decap_12
XFILLER_11_138 vpwr vgnd scs8hd_fill_2
XFILLER_22_23 vgnd vpwr scs8hd_decap_4
XFILLER_42_230 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_9_ mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_8_58 vgnd vpwr scs8hd_fill_1
XANTENNA__134__C _134_/C vgnd vpwr scs8hd_diode_2
X_157_ _126_/A address[2] _143_/C _109_/A _158_/B vgnd vpwr scs8hd_or4_4
X_226_ _226_/A chanx_left_out[8] vgnd vpwr scs8hd_buf_2
XANTENNA__118__D _171_/A vgnd vpwr scs8hd_diode_2
XANTENNA__150__B _149_/X vgnd vpwr scs8hd_diode_2
XFILLER_25_208 vgnd vpwr scs8hd_decap_12
XFILLER_33_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_1.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XPHY_225 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_214 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_203 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_12 vpwr vgnd scs8hd_fill_2
XFILLER_17_56 vpwr vgnd scs8hd_fill_2
XFILLER_17_89 vpwr vgnd scs8hd_fill_2
XPHY_269 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_258 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_247 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_11 vgnd vpwr scs8hd_decap_12
XPHY_236 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
XFILLER_15_252 vgnd vpwr scs8hd_decap_12
XANTENNA__145__B _145_/B vgnd vpwr scs8hd_diode_2
XANTENNA__161__A _168_/C vgnd vpwr scs8hd_diode_2
X_209_ _209_/HI _209_/LO vgnd vpwr scs8hd_conb_1
XFILLER_0_137 vgnd vpwr scs8hd_decap_4
XFILLER_8_215 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _216_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__156__A _155_/X vgnd vpwr scs8hd_diode_2
XFILLER_38_130 vgnd vpwr scs8hd_decap_12
XFILLER_30_23 vgnd vpwr scs8hd_decap_8
XFILLER_14_79 vpwr vgnd scs8hd_fill_2
XFILLER_39_10 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _194_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_29_196 vgnd vpwr scs8hd_decap_12
XFILLER_29_152 vpwr vgnd scs8hd_fill_2
Xmux_left_track_11.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _218_/HI _200_/Y mux_left_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA__126__D _171_/A vgnd vpwr scs8hd_diode_2
XFILLER_4_251 vgnd vpwr scs8hd_decap_12
XFILLER_6_80 vpwr vgnd scs8hd_fill_2
XFILLER_26_133 vgnd vpwr scs8hd_decap_6
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_41_147 vgnd vpwr scs8hd_decap_12
XPHY_78 vgnd vpwr scs8hd_decap_3
XPHY_67 vgnd vpwr scs8hd_decap_3
X_190_ _190_/A _190_/Y vgnd vpwr scs8hd_inv_8
XPHY_56 vgnd vpwr scs8hd_decap_3
XFILLER_26_199 vgnd vpwr scs8hd_decap_12
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_34 vgnd vpwr scs8hd_decap_3
XPHY_45 vgnd vpwr scs8hd_decap_3
XFILLER_1_232 vgnd vpwr scs8hd_decap_12
XFILLER_17_100 vgnd vpwr scs8hd_decap_3
XFILLER_17_188 vgnd vpwr scs8hd_decap_12
XANTENNA__153__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_36_77 vpwr vgnd scs8hd_fill_2
XFILLER_14_136 vgnd vpwr scs8hd_decap_12
X_173_ _173_/A _173_/Y vgnd vpwr scs8hd_inv_8
X_242_ _242_/A chany_bottom_out[1] vgnd vpwr scs8hd_buf_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ _199_/A mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XANTENNA__148__B _147_/B vgnd vpwr scs8hd_diode_2
XFILLER_20_128 vpwr vgnd scs8hd_fill_2
XFILLER_9_184 vgnd vpwr scs8hd_decap_12
XANTENNA__164__A _168_/C vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _223_/HI vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_239 vgnd vpwr scs8hd_decap_12
XFILLER_0_6 vpwr vgnd scs8hd_fill_2
XFILLER_22_79 vpwr vgnd scs8hd_fill_2
XFILLER_42_242 vgnd vpwr scs8hd_decap_6
XFILLER_6_154 vgnd vpwr scs8hd_decap_12
XANTENNA__134__D _171_/A vgnd vpwr scs8hd_diode_2
X_156_ _155_/X _153_/X _156_/Y vgnd vpwr scs8hd_nor2_4
X_225_ _225_/HI _225_/LO vgnd vpwr scs8hd_conb_1
XFILLER_33_220 vgnd vpwr scs8hd_decap_12
XANTENNA__159__A _155_/X vgnd vpwr scs8hd_diode_2
XFILLER_33_275 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_259 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_248 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_23 vpwr vgnd scs8hd_fill_2
XPHY_237 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_226 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_215 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_204 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_35 vpwr vgnd scs8hd_fill_2
XFILLER_33_89 vpwr vgnd scs8hd_fill_2
XFILLER_3_135 vgnd vpwr scs8hd_decap_12
XFILLER_15_220 vgnd vpwr scs8hd_decap_12
XFILLER_15_264 vgnd vpwr scs8hd_decap_12
X_139_ _160_/C _143_/C vgnd vpwr scs8hd_buf_1
XANTENNA__161__B _162_/B vgnd vpwr scs8hd_diode_2
X_208_ _208_/HI _208_/LO vgnd vpwr scs8hd_conb_1
XFILLER_2_190 vgnd vpwr scs8hd_decap_12
Xmux_left_track_7.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_7_ mux_left_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_21_245 vgnd vpwr scs8hd_decap_12
XFILLER_0_116 vpwr vgnd scs8hd_fill_2
XFILLER_0_149 vgnd vpwr scs8hd_decap_6
XFILLER_28_67 vpwr vgnd scs8hd_fill_2
XFILLER_28_56 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_8_227 vgnd vpwr scs8hd_decap_12
XFILLER_12_212 vpwr vgnd scs8hd_fill_2
XFILLER_5_27 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _212_/HI vgnd
+ vpwr scs8hd_diode_2
XANTENNA__172__A _172_/A vgnd vpwr scs8hd_diode_2
XANTENNA__156__B _153_/X vgnd vpwr scs8hd_diode_2
XFILLER_38_142 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_3.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _213_/HI _174_/Y mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_14_14 vpwr vgnd scs8hd_fill_2
XFILLER_14_36 vpwr vgnd scs8hd_fill_2
XFILLER_14_47 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ _242_/A vgnd vpwr scs8hd_inv_1
XFILLER_5_208 vgnd vpwr scs8hd_decap_12
XFILLER_39_22 vgnd vpwr scs8hd_decap_12
XFILLER_4_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_35_112 vgnd vpwr scs8hd_decap_4
XFILLER_35_123 vgnd vpwr scs8hd_decap_12
XANTENNA__167__A _167_/A vgnd vpwr scs8hd_diode_2
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
Xmem_left_track_13.LATCH_1_.latch data_in _202_/A _164_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_46 vgnd vpwr scs8hd_decap_3
XFILLER_41_159 vgnd vpwr scs8hd_decap_12
XPHY_79 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_decap_3
XFILLER_9_3 vgnd vpwr scs8hd_decap_3
XFILLER_32_104 vgnd vpwr scs8hd_decap_8
XFILLER_17_123 vgnd vpwr scs8hd_decap_4
XFILLER_17_145 vpwr vgnd scs8hd_fill_2
XFILLER_15_90 vpwr vgnd scs8hd_fill_2
XANTENNA__153__C _143_/C vgnd vpwr scs8hd_diode_2
Xmem_bottom_track_9.LATCH_1_.latch data_in _180_/A _124_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_36_89 vgnd vpwr scs8hd_decap_3
XFILLER_14_148 vgnd vpwr scs8hd_fill_1
XANTENNA_mem_bottom_track_11.LATCH_0_.latch_SLEEPB _128_/Y vgnd vpwr scs8hd_diode_2
X_241_ _241_/A chany_bottom_out[2] vgnd vpwr scs8hd_buf_2
X_172_ _172_/A _172_/Y vgnd vpwr scs8hd_inv_8
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA__164__B _165_/B vgnd vpwr scs8hd_diode_2
XFILLER_13_181 vpwr vgnd scs8hd_fill_2
XANTENNA__180__A _180_/A vgnd vpwr scs8hd_diode_2
XFILLER_9_196 vgnd vpwr scs8hd_decap_12
XFILLER_3_60 vgnd vpwr scs8hd_fill_1
Xmux_left_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_13.INVTX1_1_.scs8hd_inv_1/Y
+ _203_/Y mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_36_251 vgnd vpwr scs8hd_decap_12
XFILLER_11_107 vpwr vgnd scs8hd_fill_2
XFILLER_22_47 vpwr vgnd scs8hd_fill_2
XFILLER_22_58 vpwr vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_0_.latch data_in _199_/A _159_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_224_ _224_/HI _224_/LO vgnd vpwr scs8hd_conb_1
XFILLER_8_38 vgnd vpwr scs8hd_fill_1
X_155_ address[0] _155_/X vgnd vpwr scs8hd_buf_1
XFILLER_6_166 vgnd vpwr scs8hd_decap_12
XFILLER_33_7 vpwr vgnd scs8hd_fill_2
XFILLER_26_6 vpwr vgnd scs8hd_fill_2
XFILLER_33_232 vgnd vpwr scs8hd_decap_12
XANTENNA__159__B _158_/B vgnd vpwr scs8hd_diode_2
XFILLER_18_251 vgnd vpwr scs8hd_decap_12
XANTENNA__175__A _175_/A vgnd vpwr scs8hd_diode_2
XPHY_249 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_57 vpwr vgnd scs8hd_fill_2
XPHY_238 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_227 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_216 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_205 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_69 vgnd vpwr scs8hd_decap_4
XFILLER_24_276 vgnd vpwr scs8hd_fill_1
XFILLER_3_114 vgnd vpwr scs8hd_decap_8
XFILLER_3_147 vgnd vpwr scs8hd_decap_12
XFILLER_15_232 vgnd vpwr scs8hd_decap_12
X_207_ _207_/A _207_/Y vgnd vpwr scs8hd_inv_8
XFILLER_30_213 vgnd vpwr scs8hd_fill_1
XFILLER_15_276 vgnd vpwr scs8hd_fill_1
X_138_ address[4] _138_/B _160_/C vgnd vpwr scs8hd_nand2_4
XFILLER_24_3 vgnd vpwr scs8hd_decap_4
XFILLER_0_61 vgnd vpwr scs8hd_fill_1
XFILLER_21_257 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _202_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_28_46 vgnd vpwr scs8hd_fill_1
XFILLER_28_35 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_3.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[0] vgnd vpwr scs8hd_diode_2
XFILLER_8_239 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_7_ vgnd vpwr
+ scs8hd_diode_2
XFILLER_38_154 vgnd vpwr scs8hd_decap_12
XFILLER_14_26 vpwr vgnd scs8hd_fill_2
XFILLER_14_59 vgnd vpwr scs8hd_decap_4
XFILLER_30_47 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ _173_/A mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_39_56 vgnd vpwr scs8hd_decap_4
XFILLER_39_34 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_5_ mux_left_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_29_132 vgnd vpwr scs8hd_decap_4
XFILLER_29_110 vpwr vgnd scs8hd_fill_2
XFILLER_29_165 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _181_/Y vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_left_track_13.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_20_91 vgnd vpwr scs8hd_fill_1
XFILLER_35_135 vgnd vpwr scs8hd_decap_12
XANTENNA__183__A _183_/A vgnd vpwr scs8hd_diode_2
XFILLER_6_93 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_13.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _185_/Y vgnd
+ vpwr scs8hd_diode_2
XPHY_69 vgnd vpwr scs8hd_decap_3
XPHY_58 vgnd vpwr scs8hd_decap_3
XFILLER_25_69 vpwr vgnd scs8hd_fill_2
XPHY_14 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_47 vgnd vpwr scs8hd_decap_3
XFILLER_25_47 vgnd vpwr scs8hd_decap_3
XFILLER_34_190 vgnd vpwr scs8hd_decap_12
XFILLER_1_245 vgnd vpwr scs8hd_decap_12
Xmux_left_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _194_/A mux_left_track_5.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XANTENNA__153__D _153_/D vgnd vpwr scs8hd_diode_2
XANTENNA__178__A _178_/A vgnd vpwr scs8hd_diode_2
XFILLER_23_138 vpwr vgnd scs8hd_fill_2
XFILLER_23_149 vgnd vpwr scs8hd_decap_4
XFILLER_11_27 vgnd vpwr scs8hd_decap_4
XFILLER_11_38 vpwr vgnd scs8hd_fill_2
XFILLER_36_46 vgnd vpwr scs8hd_decap_8
X_240_ _240_/A chany_bottom_out[3] vgnd vpwr scs8hd_buf_2
X_171_ _171_/A _168_/B _155_/X _171_/Y vgnd vpwr scs8hd_nor3_4
Xmux_bottom_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ _177_/Y mux_bottom_track_5.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XFILLER_37_208 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_17.LATCH_1_.latch data_in _188_/A _141_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_3.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_9_153 vgnd vpwr scs8hd_fill_1
XFILLER_9_164 vpwr vgnd scs8hd_fill_2
XFILLER_36_263 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _204_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_11_119 vgnd vpwr scs8hd_fill_1
XFILLER_42_211 vgnd vpwr scs8hd_decap_6
XFILLER_19_208 vgnd vpwr scs8hd_decap_12
X_223_ _223_/HI _223_/LO vgnd vpwr scs8hd_conb_1
XFILLER_6_178 vgnd vpwr scs8hd_decap_12
XFILLER_10_163 vgnd vpwr scs8hd_decap_8
XFILLER_10_174 vgnd vpwr scs8hd_decap_12
X_154_ _168_/C _153_/X _154_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_19_6 vpwr vgnd scs8hd_fill_2
XFILLER_18_263 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _225_/HI _198_/Y mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_11.tap_buf4_0_.scs8hd_inv_1/A
+ _238_/A vgnd vpwr scs8hd_inv_1
XANTENNA__191__A _191_/A vgnd vpwr scs8hd_diode_2
XFILLER_17_48 vpwr vgnd scs8hd_fill_2
XFILLER_24_211 vgnd vpwr scs8hd_decap_3
XPHY_239 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_33_36 vpwr vgnd scs8hd_fill_2
XPHY_228 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_217 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_206 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_3_159 vgnd vpwr scs8hd_decap_12
X_137_ address[5] _138_/B vgnd vpwr scs8hd_inv_8
X_206_ _206_/A _206_/Y vgnd vpwr scs8hd_inv_8
XANTENNA__186__A _186_/A vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _187_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_269 vgnd vpwr scs8hd_decap_8
XFILLER_9_82 vgnd vpwr scs8hd_decap_8
XFILLER_9_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _195_/Y vgnd vpwr
+ scs8hd_diode_2
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 mux_left_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _226_/A vgnd vpwr scs8hd_inv_1
XANTENNA__096__A _129_/A vgnd vpwr scs8hd_diode_2
XFILLER_18_91 vgnd vpwr scs8hd_fill_1
XFILLER_38_166 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_39_46 vgnd vpwr scs8hd_decap_3
XFILLER_29_177 vgnd vpwr scs8hd_decap_6
XFILLER_4_276 vgnd vpwr scs8hd_fill_1
XFILLER_35_147 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _230_/A vgnd vpwr scs8hd_inv_1
XPHY_59 vgnd vpwr scs8hd_decap_3
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _173_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_2_19 vgnd vpwr scs8hd_decap_12
XFILLER_1_257 vgnd vpwr scs8hd_decap_12
XFILLER_17_114 vpwr vgnd scs8hd_fill_2
XFILLER_17_158 vpwr vgnd scs8hd_fill_2
XFILLER_40_150 vgnd vpwr scs8hd_decap_3
XFILLER_32_128 vgnd vpwr scs8hd_decap_3
Xmux_left_track_3.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_3_ mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__194__A _194_/A vgnd vpwr scs8hd_diode_2
XFILLER_16_180 vgnd vpwr scs8hd_decap_12
XFILLER_23_117 vgnd vpwr scs8hd_decap_3
X_170_ _171_/A _168_/B _168_/C _170_/Y vgnd vpwr scs8hd_nor3_4
XANTENNA_mem_left_track_3.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_9_132 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_13.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_13.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_161 vpwr vgnd scs8hd_fill_2
XFILLER_3_40 vgnd vpwr scs8hd_decap_12
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XANTENNA__189__A _189_/A vgnd vpwr scs8hd_diode_2
XFILLER_3_73 vgnd vpwr scs8hd_decap_12
XFILLER_3_62 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _197_/A vgnd vpwr
+ scs8hd_diode_2
XANTENNA__099__A address[4] vgnd vpwr scs8hd_diode_2
XFILLER_27_220 vgnd vpwr scs8hd_decap_12
X_222_ _222_/HI _222_/LO vgnd vpwr scs8hd_conb_1
XFILLER_10_186 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_5.LATCH_1_.latch data_in _176_/A _116_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_153_ _126_/A address[2] _143_/C _153_/D _153_/X vgnd vpwr scs8hd_or4_4
XFILLER_37_90 vgnd vpwr scs8hd_decap_3
XFILLER_33_245 vgnd vpwr scs8hd_decap_8
Xmux_left_track_7.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_7.INVTX1_0_.scs8hd_inv_1/Y
+ _197_/A mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_207 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_16 vpwr vgnd scs8hd_fill_2
XPHY_229 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_218 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_30_215 vgnd vpwr scs8hd_decap_12
XFILLER_30_259 vgnd vpwr scs8hd_decap_12
X_205_ _205_/A _205_/Y vgnd vpwr scs8hd_inv_8
Xmem_left_track_5.LATCH_0_.latch data_in _195_/A _151_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
X_136_ _145_/A _134_/X _136_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_23_81 vpwr vgnd scs8hd_fill_2
XFILLER_31_6 vpwr vgnd scs8hd_fill_2
XFILLER_0_30 vgnd vpwr scs8hd_fill_1
XFILLER_0_63 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_3.LATCH_0_.latch_SLEEPB _112_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_204 vgnd vpwr scs8hd_decap_8
XFILLER_12_215 vgnd vpwr scs8hd_decap_12
XFILLER_20_270 vgnd vpwr scs8hd_decap_4
X_119_ _096_/X _119_/B _119_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_38_178 vgnd vpwr scs8hd_decap_12
XANTENNA__197__A _197_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_80 vpwr vgnd scs8hd_fill_2
XFILLER_20_93 vpwr vgnd scs8hd_fill_2
XFILLER_35_159 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_7.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_6_84 vgnd vpwr scs8hd_decap_8
XFILLER_26_104 vpwr vgnd scs8hd_fill_2
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_decap_3
XFILLER_41_59 vpwr vgnd scs8hd_fill_2
XFILLER_41_15 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_269 vgnd vpwr scs8hd_decap_8
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _208_/HI _172_/Y mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_15_71 vpwr vgnd scs8hd_fill_2
XFILLER_31_151 vgnd vpwr scs8hd_decap_12
XFILLER_16_192 vgnd vpwr scs8hd_decap_12
XFILLER_31_184 vgnd vpwr scs8hd_decap_12
XFILLER_39_262 vgnd vpwr scs8hd_decap_12
XFILLER_14_107 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_11.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _105_/Y vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_7.LATCH_0_.latch_SLEEPB _156_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_3 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[8] vgnd vpwr scs8hd_diode_2
XFILLER_13_184 vgnd vpwr scs8hd_decap_12
XFILLER_3_52 vgnd vpwr scs8hd_decap_8
XFILLER_36_276 vgnd vpwr scs8hd_fill_1
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 left_top_grid_pin_1_ mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_3_85 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A _224_/HI vgnd vpwr
+ scs8hd_diode_2
XANTENNA__099__B address[5] vgnd vpwr scs8hd_diode_2
XFILLER_27_232 vgnd vpwr scs8hd_decap_12
XFILLER_10_132 vgnd vpwr scs8hd_decap_4
XFILLER_10_198 vgnd vpwr scs8hd_decap_12
XFILLER_12_72 vgnd vpwr scs8hd_decap_3
X_152_ _129_/A _168_/C vgnd vpwr scs8hd_buf_1
X_221_ _221_/HI _221_/LO vgnd vpwr scs8hd_conb_1
XFILLER_37_80 vpwr vgnd scs8hd_fill_2
XFILLER_18_276 vgnd vpwr scs8hd_fill_1
Xmem_bottom_track_13.LATCH_1_.latch data_in _184_/A _131_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XPHY_219 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_208 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xmux_left_track_11.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_11.INVTX1_1_.scs8hd_inv_1/Y
+ _201_/Y mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
Xmux_bottom_track_7.INVTX1_1_.scs8hd_inv_1 chanx_left_in[4] mux_bottom_track_7.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XFILLER_30_227 vgnd vpwr scs8hd_decap_12
XFILLER_30_205 vgnd vpwr scs8hd_decap_8
X_204_ _204_/A _204_/Y vgnd vpwr scs8hd_inv_8
X_135_ _147_/A _134_/X _135_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_0_53 vpwr vgnd scs8hd_fill_2
XFILLER_0_75 vgnd vpwr scs8hd_decap_12
XFILLER_0_97 vpwr vgnd scs8hd_fill_2
XFILLER_9_51 vpwr vgnd scs8hd_fill_2
XFILLER_12_227 vgnd vpwr scs8hd_decap_12
XANTENNA_mem_left_track_5.LATCH_1_.latch_SLEEPB _150_/Y vgnd vpwr scs8hd_diode_2
XFILLER_7_242 vpwr vgnd scs8hd_fill_2
X_118_ _115_/A _115_/B _123_/C _171_/A _119_/B vgnd vpwr scs8hd_or4_4
XFILLER_38_113 vgnd vpwr scs8hd_decap_8
XFILLER_38_102 vpwr vgnd scs8hd_fill_2
XFILLER_22_3 vpwr vgnd scs8hd_fill_2
XFILLER_14_18 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_5.INVTX1_0_.scs8hd_inv_1_A bottom_right_grid_pin_5_ vgnd
+ vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A chanx_left_in[5] vgnd vpwr scs8hd_diode_2
XFILLER_20_83 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_15.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_15.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_116 vpwr vgnd scs8hd_fill_2
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_28 vgnd vpwr scs8hd_decap_3
XFILLER_25_17 vpwr vgnd scs8hd_fill_2
XFILLER_41_27 vgnd vpwr scs8hd_decap_12
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_17_127 vgnd vpwr scs8hd_fill_1
XFILLER_31_71 vpwr vgnd scs8hd_fill_2
XFILLER_31_93 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _205_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_31_163 vgnd vpwr scs8hd_decap_12
XFILLER_31_196 vgnd vpwr scs8hd_decap_12
XFILLER_39_274 vgnd vpwr scs8hd_decap_3
XFILLER_14_119 vpwr vgnd scs8hd_fill_2
XFILLER_22_163 vgnd vpwr scs8hd_decap_8
XFILLER_22_174 vgnd vpwr scs8hd_decap_12
XFILLER_26_71 vpwr vgnd scs8hd_fill_2
XFILLER_9_112 vgnd vpwr scs8hd_decap_4
XFILLER_13_141 vpwr vgnd scs8hd_fill_2
XFILLER_9_156 vgnd vpwr scs8hd_fill_1
XFILLER_13_196 vgnd vpwr scs8hd_decap_12
XFILLER_3_97 vgnd vpwr scs8hd_decap_4
Xmux_left_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ _192_/A mux_left_track_3.tap_buf4_0_.scs8hd_inv_1/A vgnd vpwr scs8hd_ebufn_2
XFILLER_36_211 vgnd vpwr scs8hd_decap_3
XFILLER_22_29 vpwr vgnd scs8hd_fill_2
X_220_ _220_/HI _220_/LO vgnd vpwr scs8hd_conb_1
XANTENNA_mux_left_track_11.INVTX1_0_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vpwr scs8hd_diode_2
X_151_ _145_/A _149_/X _151_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_10_111 vgnd vpwr scs8hd_decap_8
XFILLER_12_40 vgnd vpwr scs8hd_fill_1
XFILLER_12_84 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_15.INVTX1_1_.scs8hd_inv_1_A left_top_grid_pin_15_ vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_3.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ _175_/Y mux_bottom_track_3.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vpwr scs8hd_ebufn_2
XPHY_209 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _180_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_30_239 vgnd vpwr scs8hd_decap_12
X_203_ _203_/A _203_/Y vgnd vpwr scs8hd_inv_8
X_134_ _126_/A _115_/B _134_/C _171_/A _134_/X vgnd vpwr scs8hd_or4_4
XFILLER_0_10 vgnd vpwr scs8hd_decap_12
Xmem_bottom_track_1.LATCH_1_.latch data_in _172_/A _105_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_32 vgnd vpwr scs8hd_decap_12
XFILLER_0_87 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_bottom_track_13.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _184_/Y vgnd
+ vpwr scs8hd_diode_2
XFILLER_21_206 vgnd vpwr scs8hd_decap_12
XFILLER_9_41 vgnd vpwr scs8hd_fill_1
XFILLER_28_39 vgnd vpwr scs8hd_fill_1
Xmux_left_track_7.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 _224_/HI _196_/Y mux_left_track_7.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_ebufn_2
XFILLER_12_239 vgnd vpwr scs8hd_decap_12
XFILLER_18_83 vpwr vgnd scs8hd_fill_2
XFILLER_34_93 vgnd vpwr scs8hd_decap_6
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _207_/A vgnd vpwr
+ scs8hd_diode_2
Xmux_bottom_track_5.INVTX1_1_.scs8hd_inv_1 chanx_left_in[3] mux_bottom_track_5.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
X_117_ _106_/X _115_/X _117_/Y vgnd vpwr scs8hd_nor2_4
Xmem_left_track_1.LATCH_0_.latch data_in _191_/A _145_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_29_136 vgnd vpwr scs8hd_fill_1
XFILLER_29_114 vpwr vgnd scs8hd_fill_2
XFILLER_37_180 vgnd vpwr scs8hd_decap_3
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_202 vgnd vpwr scs8hd_decap_12
XFILLER_29_93 vpwr vgnd scs8hd_fill_2
XFILLER_34_150 vgnd vpwr scs8hd_decap_3
XPHY_18 vgnd vpwr scs8hd_decap_3
XPHY_29 vgnd vpwr scs8hd_decap_3
XFILLER_25_29 vpwr vgnd scs8hd_fill_2
XFILLER_41_39 vgnd vpwr scs8hd_decap_12
XANTENNA__102__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_23_109 vpwr vgnd scs8hd_fill_2
XFILLER_31_175 vgnd vpwr scs8hd_decap_8
XFILLER_39_253 vpwr vgnd scs8hd_fill_2
XFILLER_39_242 vpwr vgnd scs8hd_fill_2
XFILLER_36_39 vgnd vpwr scs8hd_decap_4
XFILLER_22_142 vgnd vpwr scs8hd_decap_4
XFILLER_22_186 vgnd vpwr scs8hd_decap_12
XFILLER_9_102 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_bottom_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _186_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_9_168 vgnd vpwr scs8hd_decap_12
XFILLER_3_10 vgnd vpwr scs8hd_decap_4
XANTENNA_mux_left_track_5.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB _194_/Y vgnd vpwr
+ scs8hd_diode_2
XFILLER_27_245 vgnd vpwr scs8hd_decap_12
X_150_ _147_/A _149_/X _150_/Y vgnd vpwr scs8hd_nor2_4
XFILLER_6_105 vgnd vpwr scs8hd_decap_12
XFILLER_10_145 vgnd vpwr scs8hd_decap_6
XFILLER_12_52 vgnd vpwr scs8hd_decap_8
XFILLER_12_96 vpwr vgnd scs8hd_fill_2
XFILLER_33_259 vpwr vgnd scs8hd_fill_2
XFILLER_5_171 vgnd vpwr scs8hd_decap_12
XFILLER_24_215 vgnd vpwr scs8hd_decap_12
XFILLER_24_259 vgnd vpwr scs8hd_decap_12
XANTENNA__200__A _200_/A vgnd vpwr scs8hd_diode_2
XFILLER_15_248 vpwr vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB _170_/Y vgnd vpwr scs8hd_diode_2
X_133_ _145_/A _131_/B _133_/Y vgnd vpwr scs8hd_nor2_4
X_202_ _202_/A _202_/Y vgnd vpwr scs8hd_inv_8
XFILLER_23_40 vpwr vgnd scs8hd_fill_2
XFILLER_23_62 vgnd vpwr scs8hd_decap_4
XFILLER_0_22 vgnd vpwr scs8hd_decap_8
XFILLER_0_44 vgnd vpwr scs8hd_decap_6
XANTENNA__110__A _115_/A vgnd vpwr scs8hd_diode_2
XFILLER_21_218 vgnd vpwr scs8hd_decap_12
XFILLER_9_97 vgnd vpwr scs8hd_decap_3
XFILLER_28_18 vgnd vpwr scs8hd_decap_12
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _172_/A vgnd
+ vpwr scs8hd_diode_2
XFILLER_20_251 vgnd vpwr scs8hd_decap_4
Xmux_left_track_5.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_5.INVTX1_0_.scs8hd_inv_1/Y
+ _195_/A mux_left_track_5.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_18_62 vpwr vgnd scs8hd_fill_2
XFILLER_7_222 vgnd vpwr scs8hd_decap_12
XFILLER_11_262 vgnd vpwr scs8hd_decap_12
X_116_ _096_/X _115_/X _116_/Y vgnd vpwr scs8hd_nor2_4
XANTENNA__105__A _096_/X vgnd vpwr scs8hd_diode_2
XFILLER_30_19 vgnd vpwr scs8hd_fill_1
XFILLER_29_148 vpwr vgnd scs8hd_fill_2
XFILLER_29_126 vgnd vpwr scs8hd_decap_4
XFILLER_20_41 vgnd vpwr scs8hd_decap_8
XFILLER_20_74 vpwr vgnd scs8hd_fill_2
XFILLER_35_118 vgnd vpwr scs8hd_decap_4
XFILLER_29_72 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_7.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB _196_/A vgnd vpwr
+ scs8hd_diode_2
XFILLER_26_129 vpwr vgnd scs8hd_fill_2
Xmux_bottom_track_3.INVTX1_1_.scs8hd_inv_1 chanx_left_in[2] mux_bottom_track_3.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_inv_1
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_19_170 vpwr vgnd scs8hd_fill_2
XANTENNA_mux_left_track_13.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_13.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_118 vpwr vgnd scs8hd_fill_2
XFILLER_40_154 vgnd vpwr scs8hd_decap_12
XFILLER_25_184 vgnd vpwr scs8hd_decap_12
XFILLER_31_40 vpwr vgnd scs8hd_fill_2
XANTENNA__102__B _102_/B vgnd vpwr scs8hd_diode_2
XFILLER_0_261 vgnd vpwr scs8hd_decap_12
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ _199_/Y mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vpwr scs8hd_ebufn_2
XFILLER_31_110 vpwr vgnd scs8hd_fill_2
XFILLER_16_151 vpwr vgnd scs8hd_fill_2
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_36_18 vgnd vpwr scs8hd_decap_12
XFILLER_22_110 vgnd vpwr scs8hd_decap_8
XFILLER_22_121 vpwr vgnd scs8hd_fill_2
XFILLER_22_198 vgnd vpwr scs8hd_decap_12
XANTENNA__203__A _203_/A vgnd vpwr scs8hd_diode_2
XFILLER_26_84 vgnd vpwr scs8hd_decap_8
XANTENNA_mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_15.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vpwr scs8hd_diode_2
XFILLER_42_94 vgnd vpwr scs8hd_decap_12
XFILLER_13_165 vpwr vgnd scs8hd_fill_2
XANTENNA__113__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_3_66 vgnd vpwr scs8hd_fill_1
XANTENNA_mux_left_track_15.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_15.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vpwr scs8hd_diode_2
XFILLER_27_257 vgnd vpwr scs8hd_decap_12
XFILLER_42_249 vgnd vpwr scs8hd_decap_12
XFILLER_6_117 vgnd vpwr scs8hd_decap_12
XFILLER_18_213 vgnd vpwr scs8hd_fill_1
XANTENNA__108__A address[1] vgnd vpwr scs8hd_diode_2
XANTENNA_mux_left_track_11.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_11.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_D data_in vgnd vpwr scs8hd_diode_2
XFILLER_38_3 vgnd vpwr scs8hd_decap_12
XFILLER_24_227 vgnd vpwr scs8hd_decap_12
X_132_ address[0] _145_/A vgnd vpwr scs8hd_buf_1
X_201_ _201_/A _201_/Y vgnd vpwr scs8hd_inv_8
XFILLER_23_85 vpwr vgnd scs8hd_fill_2
XFILLER_2_120 vgnd vpwr scs8hd_decap_3
XANTENNA__110__B _123_/B vgnd vpwr scs8hd_diode_2
XFILLER_9_32 vgnd vpwr scs8hd_decap_3
XFILLER_9_65 vpwr vgnd scs8hd_fill_2
XFILLER_20_274 vgnd vpwr scs8hd_fill_1
XFILLER_18_30 vgnd vpwr scs8hd_fill_1
XFILLER_18_41 vpwr vgnd scs8hd_fill_2
XFILLER_34_84 vgnd vpwr scs8hd_decap_8
XFILLER_34_73 vgnd vpwr scs8hd_decap_6
XFILLER_7_245 vgnd vpwr scs8hd_decap_12
XFILLER_7_234 vgnd vpwr scs8hd_decap_8
XFILLER_11_274 vgnd vpwr scs8hd_decap_3
XANTENNA__105__B _105_/B vgnd vpwr scs8hd_diode_2
X_115_ _115_/A _115_/B _123_/C _168_/A _115_/X vgnd vpwr scs8hd_or4_4
XANTENNA__121__A address[3] vgnd vpwr scs8hd_diode_2
Xmem_left_track_9.LATCH_1_.latch data_in _198_/A _158_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_37_160 vgnd vpwr scs8hd_decap_12
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XANTENNA__206__A _206_/A vgnd vpwr scs8hd_diode_2
XFILLER_29_62 vgnd vpwr scs8hd_fill_1
XFILLER_29_40 vpwr vgnd scs8hd_fill_2
XFILLER_20_53 vpwr vgnd scs8hd_fill_2
XFILLER_20_97 vgnd vpwr scs8hd_decap_3
XANTENNA__116__A _096_/X vgnd vpwr scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vpwr scs8hd_diode_2
XFILLER_26_108 vgnd vpwr scs8hd_decap_8
XFILLER_20_3 vpwr vgnd scs8hd_fill_2
XFILLER_34_130 vgnd vpwr scs8hd_decap_12
XFILLER_19_182 vgnd vpwr scs8hd_fill_1
XFILLER_40_166 vgnd vpwr scs8hd_decap_12
XFILLER_25_196 vgnd vpwr scs8hd_decap_12
XFILLER_25_163 vgnd vpwr scs8hd_decap_12
XFILLER_15_53 vpwr vgnd scs8hd_fill_2
XFILLER_15_75 vpwr vgnd scs8hd_fill_2
XFILLER_15_86 vpwr vgnd scs8hd_fill_2
XFILLER_15_97 vpwr vgnd scs8hd_fill_2
XFILLER_0_273 vgnd vpwr scs8hd_decap_4
XFILLER_16_163 vgnd vpwr scs8hd_decap_8
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_191 vgnd vpwr scs8hd_tapvpwrvgnd_1
.ends

