VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_1__2_
  CLASS BLOCK ;
  FOREIGN sb_1__2_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 114.000 BY 114.000 ;
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END SC_IN_BOT
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END SC_OUT_BOT
  PIN bottom_left_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.010 0.000 1.290 4.000 ;
    END
  END bottom_left_grid_pin_42_
  PIN bottom_left_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END bottom_left_grid_pin_43_
  PIN bottom_left_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 4.000 ;
    END
  END bottom_left_grid_pin_44_
  PIN bottom_left_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END bottom_left_grid_pin_45_
  PIN bottom_left_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END bottom_left_grid_pin_46_
  PIN bottom_left_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END bottom_left_grid_pin_47_
  PIN bottom_left_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 4.000 ;
    END
  END bottom_left_grid_pin_48_
  PIN bottom_left_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END bottom_left_grid_pin_49_
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 110.000 28.890 114.000 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.650 110.000 85.930 114.000 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 4.000 103.320 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END chanx_left_out[9]
  PIN chanx_right_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 19.080 114.000 19.680 ;
    END
  END chanx_right_in[0]
  PIN chanx_right_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 42.200 114.000 42.800 ;
    END
  END chanx_right_in[10]
  PIN chanx_right_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 44.920 114.000 45.520 ;
    END
  END chanx_right_in[11]
  PIN chanx_right_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 46.960 114.000 47.560 ;
    END
  END chanx_right_in[12]
  PIN chanx_right_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 49.680 114.000 50.280 ;
    END
  END chanx_right_in[13]
  PIN chanx_right_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 51.720 114.000 52.320 ;
    END
  END chanx_right_in[14]
  PIN chanx_right_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 53.760 114.000 54.360 ;
    END
  END chanx_right_in[15]
  PIN chanx_right_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 56.480 114.000 57.080 ;
    END
  END chanx_right_in[16]
  PIN chanx_right_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 58.520 114.000 59.120 ;
    END
  END chanx_right_in[17]
  PIN chanx_right_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 61.240 114.000 61.840 ;
    END
  END chanx_right_in[18]
  PIN chanx_right_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 63.280 114.000 63.880 ;
    END
  END chanx_right_in[19]
  PIN chanx_right_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 21.120 114.000 21.720 ;
    END
  END chanx_right_in[1]
  PIN chanx_right_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 23.840 114.000 24.440 ;
    END
  END chanx_right_in[2]
  PIN chanx_right_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 25.880 114.000 26.480 ;
    END
  END chanx_right_in[3]
  PIN chanx_right_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 28.600 114.000 29.200 ;
    END
  END chanx_right_in[4]
  PIN chanx_right_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 30.640 114.000 31.240 ;
    END
  END chanx_right_in[5]
  PIN chanx_right_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 33.360 114.000 33.960 ;
    END
  END chanx_right_in[6]
  PIN chanx_right_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 35.400 114.000 36.000 ;
    END
  END chanx_right_in[7]
  PIN chanx_right_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 37.440 114.000 38.040 ;
    END
  END chanx_right_in[8]
  PIN chanx_right_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 40.160 114.000 40.760 ;
    END
  END chanx_right_in[9]
  PIN chanx_right_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 66.000 114.000 66.600 ;
    END
  END chanx_right_out[0]
  PIN chanx_right_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 89.120 114.000 89.720 ;
    END
  END chanx_right_out[10]
  PIN chanx_right_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 91.160 114.000 91.760 ;
    END
  END chanx_right_out[11]
  PIN chanx_right_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 93.880 114.000 94.480 ;
    END
  END chanx_right_out[12]
  PIN chanx_right_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 95.920 114.000 96.520 ;
    END
  END chanx_right_out[13]
  PIN chanx_right_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 98.640 114.000 99.240 ;
    END
  END chanx_right_out[14]
  PIN chanx_right_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 100.680 114.000 101.280 ;
    END
  END chanx_right_out[15]
  PIN chanx_right_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 102.720 114.000 103.320 ;
    END
  END chanx_right_out[16]
  PIN chanx_right_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 105.440 114.000 106.040 ;
    END
  END chanx_right_out[17]
  PIN chanx_right_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 107.480 114.000 108.080 ;
    END
  END chanx_right_out[18]
  PIN chanx_right_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 110.200 114.000 110.800 ;
    END
  END chanx_right_out[19]
  PIN chanx_right_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 68.040 114.000 68.640 ;
    END
  END chanx_right_out[1]
  PIN chanx_right_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 70.080 114.000 70.680 ;
    END
  END chanx_right_out[2]
  PIN chanx_right_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 72.800 114.000 73.400 ;
    END
  END chanx_right_out[3]
  PIN chanx_right_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 74.840 114.000 75.440 ;
    END
  END chanx_right_out[4]
  PIN chanx_right_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 77.560 114.000 78.160 ;
    END
  END chanx_right_out[5]
  PIN chanx_right_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 79.600 114.000 80.200 ;
    END
  END chanx_right_out[6]
  PIN chanx_right_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 82.320 114.000 82.920 ;
    END
  END chanx_right_out[7]
  PIN chanx_right_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 84.360 114.000 84.960 ;
    END
  END chanx_right_out[8]
  PIN chanx_right_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 110.000 86.400 114.000 87.000 ;
    END
  END chanx_right_out[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 4.000 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.070 0.000 52.350 4.000 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 4.000 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.150 0.000 97.430 4.000 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END chany_bottom_out[9]
  PIN left_bottom_grid_pin_34_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 4.000 1.320 ;
    END
  END left_bottom_grid_pin_34_
  PIN left_bottom_grid_pin_35_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END left_bottom_grid_pin_35_
  PIN left_bottom_grid_pin_36_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END left_bottom_grid_pin_36_
  PIN left_bottom_grid_pin_37_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END left_bottom_grid_pin_37_
  PIN left_bottom_grid_pin_38_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END left_bottom_grid_pin_38_
  PIN left_bottom_grid_pin_39_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END left_bottom_grid_pin_39_
  PIN left_bottom_grid_pin_40_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END left_bottom_grid_pin_40_
  PIN left_bottom_grid_pin_41_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END left_bottom_grid_pin_41_
  PIN left_top_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END left_top_grid_pin_1_
  PIN prog_clk_0_S_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END prog_clk_0_S_in
  PIN right_bottom_grid_pin_34_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 0.720 114.000 1.320 ;
    END
  END right_bottom_grid_pin_34_
  PIN right_bottom_grid_pin_35_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 2.760 114.000 3.360 ;
    END
  END right_bottom_grid_pin_35_
  PIN right_bottom_grid_pin_36_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 4.800 114.000 5.400 ;
    END
  END right_bottom_grid_pin_36_
  PIN right_bottom_grid_pin_37_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 7.520 114.000 8.120 ;
    END
  END right_bottom_grid_pin_37_
  PIN right_bottom_grid_pin_38_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 9.560 114.000 10.160 ;
    END
  END right_bottom_grid_pin_38_
  PIN right_bottom_grid_pin_39_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 12.280 114.000 12.880 ;
    END
  END right_bottom_grid_pin_39_
  PIN right_bottom_grid_pin_40_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 14.320 114.000 14.920 ;
    END
  END right_bottom_grid_pin_40_
  PIN right_bottom_grid_pin_41_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 17.040 114.000 17.640 ;
    END
  END right_bottom_grid_pin_41_
  PIN right_top_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 112.240 114.000 112.840 ;
    END
  END right_top_grid_pin_1_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.880 10.640 23.480 100.880 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.040 10.640 40.640 100.880 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 108.100 100.725 ;
      LAYER met1 ;
        RECT 0.990 5.820 113.090 100.880 ;
      LAYER met2 ;
        RECT 1.020 109.720 28.330 112.725 ;
        RECT 29.170 109.720 85.370 112.725 ;
        RECT 86.210 109.720 113.060 112.725 ;
        RECT 1.020 4.280 113.060 109.720 ;
        RECT 1.570 0.835 2.570 4.280 ;
        RECT 3.410 0.835 4.870 4.280 ;
        RECT 5.710 0.835 7.170 4.280 ;
        RECT 8.010 0.835 9.470 4.280 ;
        RECT 10.310 0.835 11.770 4.280 ;
        RECT 12.610 0.835 14.070 4.280 ;
        RECT 14.910 0.835 16.370 4.280 ;
        RECT 17.210 0.835 18.210 4.280 ;
        RECT 19.050 0.835 20.510 4.280 ;
        RECT 21.350 0.835 22.810 4.280 ;
        RECT 23.650 0.835 25.110 4.280 ;
        RECT 25.950 0.835 27.410 4.280 ;
        RECT 28.250 0.835 29.710 4.280 ;
        RECT 30.550 0.835 32.010 4.280 ;
        RECT 32.850 0.835 33.850 4.280 ;
        RECT 34.690 0.835 36.150 4.280 ;
        RECT 36.990 0.835 38.450 4.280 ;
        RECT 39.290 0.835 40.750 4.280 ;
        RECT 41.590 0.835 43.050 4.280 ;
        RECT 43.890 0.835 45.350 4.280 ;
        RECT 46.190 0.835 47.650 4.280 ;
        RECT 48.490 0.835 49.490 4.280 ;
        RECT 50.330 0.835 51.790 4.280 ;
        RECT 52.630 0.835 54.090 4.280 ;
        RECT 54.930 0.835 56.390 4.280 ;
        RECT 57.230 0.835 58.690 4.280 ;
        RECT 59.530 0.835 60.990 4.280 ;
        RECT 61.830 0.835 63.290 4.280 ;
        RECT 64.130 0.835 65.590 4.280 ;
        RECT 66.430 0.835 67.430 4.280 ;
        RECT 68.270 0.835 69.730 4.280 ;
        RECT 70.570 0.835 72.030 4.280 ;
        RECT 72.870 0.835 74.330 4.280 ;
        RECT 75.170 0.835 76.630 4.280 ;
        RECT 77.470 0.835 78.930 4.280 ;
        RECT 79.770 0.835 81.230 4.280 ;
        RECT 82.070 0.835 83.070 4.280 ;
        RECT 83.910 0.835 85.370 4.280 ;
        RECT 86.210 0.835 87.670 4.280 ;
        RECT 88.510 0.835 89.970 4.280 ;
        RECT 90.810 0.835 92.270 4.280 ;
        RECT 93.110 0.835 94.570 4.280 ;
        RECT 95.410 0.835 96.870 4.280 ;
        RECT 97.710 0.835 98.710 4.280 ;
        RECT 99.550 0.835 101.010 4.280 ;
        RECT 101.850 0.835 103.310 4.280 ;
        RECT 104.150 0.835 105.610 4.280 ;
        RECT 106.450 0.835 107.910 4.280 ;
        RECT 108.750 0.835 110.210 4.280 ;
        RECT 111.050 0.835 112.510 4.280 ;
      LAYER met3 ;
        RECT 4.400 111.840 109.600 112.705 ;
        RECT 4.000 111.200 110.000 111.840 ;
        RECT 4.400 109.800 109.600 111.200 ;
        RECT 4.000 108.480 110.000 109.800 ;
        RECT 4.400 107.080 109.600 108.480 ;
        RECT 4.000 106.440 110.000 107.080 ;
        RECT 4.400 105.040 109.600 106.440 ;
        RECT 4.000 103.720 110.000 105.040 ;
        RECT 4.400 102.320 109.600 103.720 ;
        RECT 4.000 101.680 110.000 102.320 ;
        RECT 4.400 100.280 109.600 101.680 ;
        RECT 4.000 99.640 110.000 100.280 ;
        RECT 4.400 98.240 109.600 99.640 ;
        RECT 4.000 96.920 110.000 98.240 ;
        RECT 4.400 95.520 109.600 96.920 ;
        RECT 4.000 94.880 110.000 95.520 ;
        RECT 4.400 93.480 109.600 94.880 ;
        RECT 4.000 92.160 110.000 93.480 ;
        RECT 4.400 90.760 109.600 92.160 ;
        RECT 4.000 90.120 110.000 90.760 ;
        RECT 4.400 88.720 109.600 90.120 ;
        RECT 4.000 87.400 110.000 88.720 ;
        RECT 4.400 86.000 109.600 87.400 ;
        RECT 4.000 85.360 110.000 86.000 ;
        RECT 4.400 83.960 109.600 85.360 ;
        RECT 4.000 83.320 110.000 83.960 ;
        RECT 4.400 81.920 109.600 83.320 ;
        RECT 4.000 80.600 110.000 81.920 ;
        RECT 4.400 79.200 109.600 80.600 ;
        RECT 4.000 78.560 110.000 79.200 ;
        RECT 4.400 77.160 109.600 78.560 ;
        RECT 4.000 75.840 110.000 77.160 ;
        RECT 4.400 74.440 109.600 75.840 ;
        RECT 4.000 73.800 110.000 74.440 ;
        RECT 4.400 72.400 109.600 73.800 ;
        RECT 4.000 71.080 110.000 72.400 ;
        RECT 4.400 69.680 109.600 71.080 ;
        RECT 4.000 69.040 110.000 69.680 ;
        RECT 4.400 67.640 109.600 69.040 ;
        RECT 4.000 67.000 110.000 67.640 ;
        RECT 4.400 65.600 109.600 67.000 ;
        RECT 4.000 64.280 110.000 65.600 ;
        RECT 4.400 62.880 109.600 64.280 ;
        RECT 4.000 62.240 110.000 62.880 ;
        RECT 4.400 60.840 109.600 62.240 ;
        RECT 4.000 59.520 110.000 60.840 ;
        RECT 4.400 58.120 109.600 59.520 ;
        RECT 4.000 57.480 110.000 58.120 ;
        RECT 4.400 56.080 109.600 57.480 ;
        RECT 4.000 54.760 110.000 56.080 ;
        RECT 4.400 53.360 109.600 54.760 ;
        RECT 4.000 52.720 110.000 53.360 ;
        RECT 4.400 51.320 109.600 52.720 ;
        RECT 4.000 50.680 110.000 51.320 ;
        RECT 4.400 49.280 109.600 50.680 ;
        RECT 4.000 47.960 110.000 49.280 ;
        RECT 4.400 46.560 109.600 47.960 ;
        RECT 4.000 45.920 110.000 46.560 ;
        RECT 4.400 44.520 109.600 45.920 ;
        RECT 4.000 43.200 110.000 44.520 ;
        RECT 4.400 41.800 109.600 43.200 ;
        RECT 4.000 41.160 110.000 41.800 ;
        RECT 4.400 39.760 109.600 41.160 ;
        RECT 4.000 38.440 110.000 39.760 ;
        RECT 4.400 37.040 109.600 38.440 ;
        RECT 4.000 36.400 110.000 37.040 ;
        RECT 4.400 35.000 109.600 36.400 ;
        RECT 4.000 34.360 110.000 35.000 ;
        RECT 4.400 32.960 109.600 34.360 ;
        RECT 4.000 31.640 110.000 32.960 ;
        RECT 4.400 30.240 109.600 31.640 ;
        RECT 4.000 29.600 110.000 30.240 ;
        RECT 4.400 28.200 109.600 29.600 ;
        RECT 4.000 26.880 110.000 28.200 ;
        RECT 4.400 25.480 109.600 26.880 ;
        RECT 4.000 24.840 110.000 25.480 ;
        RECT 4.400 23.440 109.600 24.840 ;
        RECT 4.000 22.120 110.000 23.440 ;
        RECT 4.400 20.720 109.600 22.120 ;
        RECT 4.000 20.080 110.000 20.720 ;
        RECT 4.400 18.680 109.600 20.080 ;
        RECT 4.000 18.040 110.000 18.680 ;
        RECT 4.400 16.640 109.600 18.040 ;
        RECT 4.000 15.320 110.000 16.640 ;
        RECT 4.400 13.920 109.600 15.320 ;
        RECT 4.000 13.280 110.000 13.920 ;
        RECT 4.400 11.880 109.600 13.280 ;
        RECT 4.000 10.560 110.000 11.880 ;
        RECT 4.400 9.160 109.600 10.560 ;
        RECT 4.000 8.520 110.000 9.160 ;
        RECT 4.400 7.120 109.600 8.520 ;
        RECT 4.000 5.800 110.000 7.120 ;
        RECT 4.400 4.400 109.600 5.800 ;
        RECT 4.000 3.760 110.000 4.400 ;
        RECT 4.400 2.360 109.600 3.760 ;
        RECT 4.000 1.720 110.000 2.360 ;
        RECT 4.400 0.855 109.600 1.720 ;
      LAYER met4 ;
        RECT 26.055 10.240 38.640 100.880 ;
        RECT 41.040 10.240 97.225 100.880 ;
        RECT 26.055 9.695 97.225 10.240 ;
  END
END sb_1__2_
END LIBRARY

