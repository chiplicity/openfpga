magic
tech sky130A
magscale 1 2
timestamp 1606473813
<< locali >>
rect 16405 17927 16439 18165
rect 17969 16839 18003 16941
rect 21741 16635 21775 17281
rect 13829 14187 13863 14425
rect 8585 12079 8619 12181
rect 15761 10923 15795 11025
rect 11161 7047 11195 7217
<< viali >>
rect 5089 19865 5123 19899
rect 17877 19865 17911 19899
rect 18613 19865 18647 19899
rect 20729 19865 20763 19899
rect 4997 19729 5031 19763
rect 17693 19729 17727 19763
rect 18429 19729 18463 19763
rect 19533 19729 19567 19763
rect 20545 19729 20579 19763
rect 5181 19661 5215 19695
rect 19809 19661 19843 19695
rect 4629 19525 4663 19559
rect 7481 19321 7515 19355
rect 9137 19321 9171 19355
rect 15853 19185 15887 19219
rect 17141 19185 17175 19219
rect 4077 19117 4111 19151
rect 4344 19117 4378 19151
rect 6101 19117 6135 19151
rect 7757 19117 7791 19151
rect 9689 19117 9723 19151
rect 12357 19117 12391 19151
rect 16865 19117 16899 19151
rect 18153 19117 18187 19151
rect 19533 19117 19567 19151
rect 19809 19117 19843 19151
rect 20269 19117 20303 19151
rect 6368 19049 6402 19083
rect 8002 19049 8036 19083
rect 9956 19049 9990 19083
rect 12624 19049 12658 19083
rect 15761 19049 15795 19083
rect 18797 19049 18831 19083
rect 5457 18981 5491 19015
rect 11069 18981 11103 19015
rect 13737 18981 13771 19015
rect 14013 18981 14047 19015
rect 15301 18981 15335 19015
rect 15669 18981 15703 19015
rect 20453 18981 20487 19015
rect 3801 18777 3835 18811
rect 5181 18777 5215 18811
rect 9689 18777 9723 18811
rect 14841 18777 14875 18811
rect 16773 18777 16807 18811
rect 20729 18777 20763 18811
rect 10968 18709 11002 18743
rect 12909 18709 12943 18743
rect 15384 18709 15418 18743
rect 17233 18709 17267 18743
rect 18337 18709 18371 18743
rect 2688 18641 2722 18675
rect 5089 18641 5123 18675
rect 5733 18641 5767 18675
rect 7757 18641 7791 18675
rect 8401 18641 8435 18675
rect 9597 18641 9631 18675
rect 10701 18641 10735 18675
rect 12817 18641 12851 18675
rect 13461 18641 13495 18675
rect 13728 18641 13762 18675
rect 15117 18641 15151 18675
rect 17141 18641 17175 18675
rect 18061 18641 18095 18675
rect 19533 18641 19567 18675
rect 20545 18641 20579 18675
rect 2421 18573 2455 18607
rect 5365 18573 5399 18607
rect 7849 18573 7883 18607
rect 8033 18573 8067 18607
rect 9873 18573 9907 18607
rect 10241 18573 10275 18607
rect 13001 18573 13035 18607
rect 17325 18573 17359 18607
rect 19717 18573 19751 18607
rect 12081 18505 12115 18539
rect 4721 18437 4755 18471
rect 7389 18437 7423 18471
rect 9229 18437 9263 18471
rect 12449 18437 12483 18471
rect 16497 18437 16531 18471
rect 13369 18233 13403 18267
rect 19809 18233 19843 18267
rect 10425 18165 10459 18199
rect 16405 18165 16439 18199
rect 8217 18097 8251 18131
rect 10885 18097 10919 18131
rect 11069 18097 11103 18131
rect 13921 18097 13955 18131
rect 5181 18029 5215 18063
rect 8125 18029 8159 18063
rect 10793 18029 10827 18063
rect 5457 17961 5491 17995
rect 13737 17961 13771 17995
rect 16589 18097 16623 18131
rect 19625 18029 19659 18063
rect 20269 18029 20303 18063
rect 7665 17893 7699 17927
rect 8033 17893 8067 17927
rect 13829 17893 13863 17927
rect 16405 17893 16439 17927
rect 20453 17893 20487 17927
rect 2973 17689 3007 17723
rect 17049 17689 17083 17723
rect 20361 17689 20395 17723
rect 20913 17689 20947 17723
rect 5172 17621 5206 17655
rect 1860 17553 1894 17587
rect 4905 17553 4939 17587
rect 16957 17553 16991 17587
rect 19349 17553 19383 17587
rect 20177 17553 20211 17587
rect 20729 17553 20763 17587
rect 1593 17485 1627 17519
rect 3341 17485 3375 17519
rect 17141 17485 17175 17519
rect 19625 17485 19659 17519
rect 6285 17349 6319 17383
rect 16589 17349 16623 17383
rect 21741 17281 21775 17315
rect 12817 17145 12851 17179
rect 18153 17145 18187 17179
rect 7941 17077 7975 17111
rect 3525 17009 3559 17043
rect 4537 17009 4571 17043
rect 4629 17009 4663 17043
rect 9137 17009 9171 17043
rect 10333 17009 10367 17043
rect 12265 17009 12299 17043
rect 12449 17009 12483 17043
rect 13369 17009 13403 17043
rect 18613 17009 18647 17043
rect 18705 17009 18739 17043
rect 20177 17009 20211 17043
rect 3341 16941 3375 16975
rect 6561 16941 6595 16975
rect 9045 16941 9079 16975
rect 16497 16941 16531 16975
rect 16764 16941 16798 16975
rect 17969 16941 18003 16975
rect 19257 16941 19291 16975
rect 19993 16941 20027 16975
rect 6828 16873 6862 16907
rect 10241 16873 10275 16907
rect 13277 16873 13311 16907
rect 19533 16873 19567 16907
rect 2973 16805 3007 16839
rect 3433 16805 3467 16839
rect 4077 16805 4111 16839
rect 4445 16805 4479 16839
rect 8585 16805 8619 16839
rect 8953 16805 8987 16839
rect 9781 16805 9815 16839
rect 10149 16805 10183 16839
rect 11805 16805 11839 16839
rect 12173 16805 12207 16839
rect 13185 16805 13219 16839
rect 17877 16805 17911 16839
rect 17969 16805 18003 16839
rect 18521 16805 18555 16839
rect 6929 16601 6963 16635
rect 10057 16601 10091 16635
rect 11713 16601 11747 16635
rect 12541 16601 12575 16635
rect 16957 16601 16991 16635
rect 18061 16601 18095 16635
rect 20177 16601 20211 16635
rect 20729 16601 20763 16635
rect 21741 16601 21775 16635
rect 4169 16533 4203 16567
rect 8944 16533 8978 16567
rect 10578 16533 10612 16567
rect 19073 16533 19107 16567
rect 3893 16465 3927 16499
rect 7297 16465 7331 16499
rect 7941 16465 7975 16499
rect 8677 16465 8711 16499
rect 13257 16465 13291 16499
rect 15025 16465 15059 16499
rect 15844 16465 15878 16499
rect 18797 16465 18831 16499
rect 19993 16465 20027 16499
rect 20545 16465 20579 16499
rect 7389 16397 7423 16431
rect 7481 16397 7515 16431
rect 10333 16397 10367 16431
rect 13001 16397 13035 16431
rect 15577 16397 15611 16431
rect 14381 16261 14415 16295
rect 3157 16057 3191 16091
rect 7021 16057 7055 16091
rect 7297 16057 7331 16091
rect 12909 16057 12943 16091
rect 15301 16057 15335 16091
rect 20453 16057 20487 16091
rect 14105 15989 14139 16023
rect 19901 15989 19935 16023
rect 5641 15921 5675 15955
rect 7757 15921 7791 15955
rect 7849 15921 7883 15955
rect 10149 15921 10183 15955
rect 14657 15921 14691 15955
rect 15761 15921 15795 15955
rect 15853 15921 15887 15955
rect 1777 15853 1811 15887
rect 5908 15853 5942 15887
rect 11529 15853 11563 15887
rect 11796 15853 11830 15887
rect 14473 15853 14507 15887
rect 15669 15853 15703 15887
rect 19717 15853 19751 15887
rect 20269 15853 20303 15887
rect 2044 15785 2078 15819
rect 14565 15785 14599 15819
rect 7665 15717 7699 15751
rect 3065 15513 3099 15547
rect 6285 15513 6319 15547
rect 20729 15513 20763 15547
rect 19165 15445 19199 15479
rect 3433 15377 3467 15411
rect 5172 15377 5206 15411
rect 7389 15377 7423 15411
rect 18889 15377 18923 15411
rect 19625 15377 19659 15411
rect 19901 15377 19935 15411
rect 20545 15377 20579 15411
rect 3525 15309 3559 15343
rect 3617 15309 3651 15343
rect 4905 15309 4939 15343
rect 7205 15173 7239 15207
rect 2973 14969 3007 15003
rect 4077 14969 4111 15003
rect 13185 14969 13219 15003
rect 14933 14969 14967 15003
rect 20453 14969 20487 15003
rect 7941 14901 7975 14935
rect 3433 14833 3467 14867
rect 4629 14833 4663 14867
rect 8401 14833 8435 14867
rect 8585 14833 8619 14867
rect 10149 14833 10183 14867
rect 10241 14833 10275 14867
rect 12541 14833 12575 14867
rect 13553 14833 13587 14867
rect 17141 14833 17175 14867
rect 19073 14833 19107 14867
rect 1593 14765 1627 14799
rect 4537 14765 4571 14799
rect 12449 14765 12483 14799
rect 13369 14765 13403 14799
rect 13820 14765 13854 14799
rect 18797 14765 18831 14799
rect 20269 14765 20303 14799
rect 1860 14697 1894 14731
rect 10057 14697 10091 14731
rect 10701 14697 10735 14731
rect 4445 14629 4479 14663
rect 8309 14629 8343 14663
rect 9689 14629 9723 14663
rect 11989 14629 12023 14663
rect 12357 14629 12391 14663
rect 16589 14629 16623 14663
rect 16957 14629 16991 14663
rect 17049 14629 17083 14663
rect 3617 14425 3651 14459
rect 9689 14425 9723 14459
rect 12909 14425 12943 14459
rect 13829 14425 13863 14459
rect 20913 14425 20947 14459
rect 2504 14357 2538 14391
rect 2237 14289 2271 14323
rect 6101 14289 6135 14323
rect 8576 14289 8610 14323
rect 12817 14289 12851 14323
rect 6193 14221 6227 14255
rect 6285 14221 6319 14255
rect 8309 14221 8343 14255
rect 13001 14221 13035 14255
rect 14188 14357 14222 14391
rect 19533 14357 19567 14391
rect 13921 14289 13955 14323
rect 15577 14289 15611 14323
rect 15844 14289 15878 14323
rect 19257 14289 19291 14323
rect 19993 14289 20027 14323
rect 20269 14289 20303 14323
rect 20729 14289 20763 14323
rect 17417 14221 17451 14255
rect 12449 14153 12483 14187
rect 13829 14153 13863 14187
rect 15301 14153 15335 14187
rect 5733 14085 5767 14119
rect 16957 14085 16991 14119
rect 6193 13881 6227 13915
rect 8677 13881 8711 13915
rect 12633 13881 12667 13915
rect 17509 13881 17543 13915
rect 18981 13881 19015 13915
rect 19901 13881 19935 13915
rect 20453 13881 20487 13915
rect 8953 13813 8987 13847
rect 12357 13813 12391 13847
rect 16497 13813 16531 13847
rect 6469 13745 6503 13779
rect 13185 13745 13219 13779
rect 17141 13745 17175 13779
rect 18061 13745 18095 13779
rect 4813 13677 4847 13711
rect 7297 13677 7331 13711
rect 7564 13677 7598 13711
rect 9137 13677 9171 13711
rect 10977 13677 11011 13711
rect 17877 13677 17911 13711
rect 18797 13677 18831 13711
rect 19717 13677 19751 13711
rect 20269 13677 20303 13711
rect 5080 13609 5114 13643
rect 11222 13609 11256 13643
rect 13001 13609 13035 13643
rect 13645 13609 13679 13643
rect 17969 13609 18003 13643
rect 13093 13541 13127 13575
rect 16865 13541 16899 13575
rect 16957 13541 16991 13575
rect 5641 13337 5675 13371
rect 11345 13337 11379 13371
rect 20177 13337 20211 13371
rect 20729 13337 20763 13371
rect 4160 13269 4194 13303
rect 10059 13269 10093 13303
rect 18613 13269 18647 13303
rect 3893 13201 3927 13235
rect 6009 13201 6043 13235
rect 18337 13201 18371 13235
rect 19441 13201 19475 13235
rect 19993 13201 20027 13235
rect 20545 13201 20579 13235
rect 6101 13133 6135 13167
rect 6193 13133 6227 13167
rect 5273 13065 5307 13099
rect 19625 13065 19659 13099
rect 11253 12793 11287 12827
rect 12449 12793 12483 12827
rect 20085 12793 20119 12827
rect 7665 12725 7699 12759
rect 12909 12725 12943 12759
rect 9873 12657 9907 12691
rect 13369 12657 13403 12691
rect 13553 12657 13587 12691
rect 14749 12657 14783 12691
rect 15577 12657 15611 12691
rect 7849 12589 7883 12623
rect 11345 12589 11379 12623
rect 12633 12589 12667 12623
rect 15301 12589 15335 12623
rect 16589 12589 16623 12623
rect 19073 12589 19107 12623
rect 19349 12589 19383 12623
rect 19901 12589 19935 12623
rect 10140 12521 10174 12555
rect 11621 12521 11655 12555
rect 14565 12521 14599 12555
rect 16856 12521 16890 12555
rect 13277 12453 13311 12487
rect 14105 12453 14139 12487
rect 14473 12453 14507 12487
rect 17969 12453 18003 12487
rect 10333 12249 10367 12283
rect 14565 12249 14599 12283
rect 16681 12249 16715 12283
rect 18061 12249 18095 12283
rect 20085 12249 20119 12283
rect 20637 12249 20671 12283
rect 7288 12181 7322 12215
rect 8585 12181 8619 12215
rect 14473 12181 14507 12215
rect 15568 12181 15602 12215
rect 7021 12113 7055 12147
rect 8933 12113 8967 12147
rect 10701 12113 10735 12147
rect 12716 12113 12750 12147
rect 18429 12113 18463 12147
rect 19901 12113 19935 12147
rect 20453 12113 20487 12147
rect 8585 12045 8619 12079
rect 8677 12045 8711 12079
rect 10793 12045 10827 12079
rect 10885 12045 10919 12079
rect 12449 12045 12483 12079
rect 14657 12045 14691 12079
rect 15301 12045 15335 12079
rect 18521 12045 18555 12079
rect 18613 12045 18647 12079
rect 10057 11977 10091 12011
rect 13829 11977 13863 12011
rect 8401 11909 8435 11943
rect 14105 11909 14139 11943
rect 7941 11705 7975 11739
rect 10333 11705 10367 11739
rect 13369 11705 13403 11739
rect 13645 11705 13679 11739
rect 18061 11705 18095 11739
rect 20453 11705 20487 11739
rect 6837 11637 6871 11671
rect 7389 11569 7423 11603
rect 8585 11569 8619 11603
rect 10885 11569 10919 11603
rect 14197 11569 14231 11603
rect 18613 11569 18647 11603
rect 7205 11501 7239 11535
rect 10793 11501 10827 11535
rect 13553 11501 13587 11535
rect 14105 11501 14139 11535
rect 20269 11501 20303 11535
rect 8401 11433 8435 11467
rect 10701 11433 10735 11467
rect 11345 11433 11379 11467
rect 18429 11433 18463 11467
rect 19073 11433 19107 11467
rect 7297 11365 7331 11399
rect 8309 11365 8343 11399
rect 14013 11365 14047 11399
rect 18521 11365 18555 11399
rect 8217 11161 8251 11195
rect 8677 11161 8711 11195
rect 13737 11161 13771 11195
rect 14197 11161 14231 11195
rect 15945 11161 15979 11195
rect 17417 11161 17451 11195
rect 18797 11161 18831 11195
rect 20729 11161 20763 11195
rect 8585 11093 8619 11127
rect 11069 11093 11103 11127
rect 10793 11025 10827 11059
rect 14105 11025 14139 11059
rect 14749 11025 14783 11059
rect 15761 11025 15795 11059
rect 16313 11025 16347 11059
rect 17325 11025 17359 11059
rect 19165 11025 19199 11059
rect 20545 11025 20579 11059
rect 8769 10957 8803 10991
rect 14289 10957 14323 10991
rect 16405 10957 16439 10991
rect 16589 10957 16623 10991
rect 17509 10957 17543 10991
rect 19257 10957 19291 10991
rect 19349 10957 19383 10991
rect 15761 10889 15795 10923
rect 16957 10889 16991 10923
rect 8585 10617 8619 10651
rect 10241 10617 10275 10651
rect 14197 10617 14231 10651
rect 16497 10617 16531 10651
rect 18705 10617 18739 10651
rect 20453 10617 20487 10651
rect 10793 10481 10827 10515
rect 11897 10481 11931 10515
rect 12817 10481 12851 10515
rect 17141 10481 17175 10515
rect 19257 10481 19291 10515
rect 7205 10413 7239 10447
rect 11621 10413 11655 10447
rect 13084 10413 13118 10447
rect 20269 10413 20303 10447
rect 7472 10345 7506 10379
rect 10609 10345 10643 10379
rect 11713 10345 11747 10379
rect 16865 10345 16899 10379
rect 19073 10345 19107 10379
rect 10701 10277 10735 10311
rect 11253 10277 11287 10311
rect 16957 10277 16991 10311
rect 19165 10277 19199 10311
rect 9505 10073 9539 10107
rect 10609 10073 10643 10107
rect 11069 10073 11103 10107
rect 17325 10073 17359 10107
rect 18061 10073 18095 10107
rect 19901 10073 19935 10107
rect 20729 10073 20763 10107
rect 16212 10005 16246 10039
rect 8392 9937 8426 9971
rect 10977 9937 11011 9971
rect 15945 9937 15979 9971
rect 18521 9937 18555 9971
rect 18788 9937 18822 9971
rect 20545 9937 20579 9971
rect 8125 9869 8159 9903
rect 11161 9869 11195 9903
rect 9321 9529 9355 9563
rect 10793 9529 10827 9563
rect 18705 9529 18739 9563
rect 15485 9461 15519 9495
rect 11345 9393 11379 9427
rect 12909 9393 12943 9427
rect 13553 9393 13587 9427
rect 19257 9393 19291 9427
rect 7941 9325 7975 9359
rect 12817 9325 12851 9359
rect 13820 9325 13854 9359
rect 15301 9325 15335 9359
rect 19073 9325 19107 9359
rect 8208 9257 8242 9291
rect 11161 9257 11195 9291
rect 11805 9257 11839 9291
rect 11253 9189 11287 9223
rect 12357 9189 12391 9223
rect 12725 9189 12759 9223
rect 14933 9189 14967 9223
rect 19165 9189 19199 9223
rect 11069 8985 11103 9019
rect 11529 8985 11563 9019
rect 13461 8985 13495 9019
rect 19717 8985 19751 9019
rect 20729 8985 20763 9019
rect 11437 8917 11471 8951
rect 15761 8917 15795 8951
rect 13277 8849 13311 8883
rect 15485 8849 15519 8883
rect 18337 8849 18371 8883
rect 18604 8849 18638 8883
rect 19993 8849 20027 8883
rect 20545 8849 20579 8883
rect 11621 8781 11655 8815
rect 20177 8713 20211 8747
rect 11437 8441 11471 8475
rect 20453 8441 20487 8475
rect 13553 8305 13587 8339
rect 11253 8237 11287 8271
rect 13369 8237 13403 8271
rect 20269 8237 20303 8271
rect 13737 7897 13771 7931
rect 16405 7897 16439 7931
rect 19441 7897 19475 7931
rect 20729 7897 20763 7931
rect 11161 7829 11195 7863
rect 9496 7761 9530 7795
rect 10885 7761 10919 7795
rect 14105 7761 14139 7795
rect 15005 7761 15039 7795
rect 16773 7761 16807 7795
rect 17417 7761 17451 7795
rect 18317 7761 18351 7795
rect 19993 7761 20027 7795
rect 20545 7761 20579 7795
rect 9229 7693 9263 7727
rect 14197 7693 14231 7727
rect 14381 7693 14415 7727
rect 14749 7693 14783 7727
rect 16865 7693 16899 7727
rect 17049 7693 17083 7727
rect 18061 7693 18095 7727
rect 10609 7557 10643 7591
rect 16129 7557 16163 7591
rect 20177 7557 20211 7591
rect 10241 7353 10275 7387
rect 14289 7353 14323 7387
rect 17601 7353 17635 7387
rect 10793 7217 10827 7251
rect 11161 7217 11195 7251
rect 11253 7217 11287 7251
rect 14565 7217 14599 7251
rect 9781 7081 9815 7115
rect 10609 7081 10643 7115
rect 12909 7149 12943 7183
rect 16221 7149 16255 7183
rect 11498 7081 11532 7115
rect 13176 7081 13210 7115
rect 16488 7081 16522 7115
rect 10701 7013 10735 7047
rect 11161 7013 11195 7047
rect 12633 7013 12667 7047
rect 10609 6809 10643 6843
rect 14105 6809 14139 6843
rect 16865 6809 16899 6843
rect 17325 6809 17359 6843
rect 10977 6741 11011 6775
rect 14473 6741 14507 6775
rect 17233 6741 17267 6775
rect 7553 6673 7587 6707
rect 20545 6673 20579 6707
rect 7297 6605 7331 6639
rect 11069 6605 11103 6639
rect 11161 6605 11195 6639
rect 14565 6605 14599 6639
rect 14657 6605 14691 6639
rect 17417 6605 17451 6639
rect 8677 6537 8711 6571
rect 20729 6469 20763 6503
rect 20729 5721 20763 5755
rect 20545 5585 20579 5619
rect 20729 4633 20763 4667
rect 20545 4497 20579 4531
<< metal1 >>
rect 1104 20010 21620 20032
rect 1104 19958 7846 20010
rect 7898 19958 7910 20010
rect 7962 19958 7974 20010
rect 8026 19958 8038 20010
rect 8090 19958 14710 20010
rect 14762 19958 14774 20010
rect 14826 19958 14838 20010
rect 14890 19958 14902 20010
rect 14954 19958 21620 20010
rect 1104 19936 21620 19958
rect 4706 19856 4712 19908
rect 4764 19896 4770 19908
rect 5077 19899 5135 19905
rect 5077 19896 5089 19899
rect 4764 19868 5089 19896
rect 4764 19856 4770 19868
rect 5077 19865 5089 19868
rect 5123 19865 5135 19899
rect 5077 19859 5135 19865
rect 17865 19899 17923 19905
rect 17865 19865 17877 19899
rect 17911 19896 17923 19899
rect 17954 19896 17960 19908
rect 17911 19868 17960 19896
rect 17911 19865 17923 19868
rect 17865 19859 17923 19865
rect 17954 19856 17960 19868
rect 18012 19856 18018 19908
rect 18601 19899 18659 19905
rect 18601 19865 18613 19899
rect 18647 19896 18659 19899
rect 18690 19896 18696 19908
rect 18647 19868 18696 19896
rect 18647 19865 18659 19868
rect 18601 19859 18659 19865
rect 18690 19856 18696 19868
rect 18748 19856 18754 19908
rect 20622 19856 20628 19908
rect 20680 19896 20686 19908
rect 20717 19899 20775 19905
rect 20717 19896 20729 19899
rect 20680 19868 20729 19896
rect 20680 19856 20686 19868
rect 20717 19865 20729 19868
rect 20763 19865 20775 19899
rect 20717 19859 20775 19865
rect 4985 19763 5043 19769
rect 4985 19729 4997 19763
rect 5031 19760 5043 19763
rect 9582 19760 9588 19772
rect 5031 19732 9588 19760
rect 5031 19729 5043 19732
rect 4985 19723 5043 19729
rect 9582 19720 9588 19732
rect 9640 19720 9646 19772
rect 17678 19760 17684 19772
rect 17639 19732 17684 19760
rect 17678 19720 17684 19732
rect 17736 19720 17742 19772
rect 18417 19763 18475 19769
rect 18417 19729 18429 19763
rect 18463 19760 18475 19763
rect 18506 19760 18512 19772
rect 18463 19732 18512 19760
rect 18463 19729 18475 19732
rect 18417 19723 18475 19729
rect 18506 19720 18512 19732
rect 18564 19720 18570 19772
rect 19334 19720 19340 19772
rect 19392 19760 19398 19772
rect 19521 19763 19579 19769
rect 19521 19760 19533 19763
rect 19392 19732 19533 19760
rect 19392 19720 19398 19732
rect 19521 19729 19533 19732
rect 19567 19729 19579 19763
rect 19521 19723 19579 19729
rect 19702 19720 19708 19772
rect 19760 19760 19766 19772
rect 20533 19763 20591 19769
rect 20533 19760 20545 19763
rect 19760 19732 20545 19760
rect 19760 19720 19766 19732
rect 20533 19729 20545 19732
rect 20579 19729 20591 19763
rect 20533 19723 20591 19729
rect 4706 19652 4712 19704
rect 4764 19692 4770 19704
rect 5169 19695 5227 19701
rect 5169 19692 5181 19695
rect 4764 19664 5181 19692
rect 4764 19652 4770 19664
rect 5169 19661 5181 19664
rect 5215 19661 5227 19695
rect 19794 19692 19800 19704
rect 19755 19664 19800 19692
rect 5169 19655 5227 19661
rect 19794 19652 19800 19664
rect 19852 19652 19858 19704
rect 4617 19559 4675 19565
rect 4617 19525 4629 19559
rect 4663 19556 4675 19559
rect 5166 19556 5172 19568
rect 4663 19528 5172 19556
rect 4663 19525 4675 19528
rect 4617 19519 4675 19525
rect 5166 19516 5172 19528
rect 5224 19516 5230 19568
rect 1104 19466 21620 19488
rect 1104 19414 4414 19466
rect 4466 19414 4478 19466
rect 4530 19414 4542 19466
rect 4594 19414 4606 19466
rect 4658 19414 11278 19466
rect 11330 19414 11342 19466
rect 11394 19414 11406 19466
rect 11458 19414 11470 19466
rect 11522 19414 18142 19466
rect 18194 19414 18206 19466
rect 18258 19414 18270 19466
rect 18322 19414 18334 19466
rect 18386 19414 21620 19466
rect 1104 19392 21620 19414
rect 7469 19355 7527 19361
rect 7469 19321 7481 19355
rect 7515 19352 7527 19355
rect 7926 19352 7932 19364
rect 7515 19324 7932 19352
rect 7515 19321 7527 19324
rect 7469 19315 7527 19321
rect 7926 19312 7932 19324
rect 7984 19312 7990 19364
rect 9125 19355 9183 19361
rect 9125 19321 9137 19355
rect 9171 19352 9183 19355
rect 9950 19352 9956 19364
rect 9171 19324 9956 19352
rect 9171 19321 9183 19324
rect 9125 19315 9183 19321
rect 9950 19312 9956 19324
rect 10008 19312 10014 19364
rect 7668 19188 7880 19216
rect 106 19108 112 19160
rect 164 19148 170 19160
rect 842 19148 848 19160
rect 164 19120 848 19148
rect 164 19108 170 19120
rect 842 19108 848 19120
rect 900 19108 906 19160
rect 2406 19108 2412 19160
rect 2464 19148 2470 19160
rect 4065 19151 4123 19157
rect 4065 19148 4077 19151
rect 2464 19120 4077 19148
rect 2464 19108 2470 19120
rect 4065 19117 4077 19120
rect 4111 19117 4123 19151
rect 4065 19111 4123 19117
rect 4332 19151 4390 19157
rect 4332 19117 4344 19151
rect 4378 19148 4390 19151
rect 4706 19148 4712 19160
rect 4378 19120 4712 19148
rect 4378 19117 4390 19120
rect 4332 19111 4390 19117
rect 4706 19108 4712 19120
rect 4764 19108 4770 19160
rect 6086 19148 6092 19160
rect 6047 19120 6092 19148
rect 6086 19108 6092 19120
rect 6144 19108 6150 19160
rect 7668 19148 7696 19188
rect 6288 19120 7696 19148
rect 7745 19151 7803 19157
rect 5810 19040 5816 19092
rect 5868 19080 5874 19092
rect 6288 19080 6316 19120
rect 7745 19117 7757 19151
rect 7791 19117 7803 19151
rect 7852 19148 7880 19188
rect 9600 19188 9812 19216
rect 9600 19148 9628 19188
rect 7852 19120 9628 19148
rect 9677 19151 9735 19157
rect 7745 19111 7803 19117
rect 9677 19117 9689 19151
rect 9723 19117 9735 19151
rect 9784 19148 9812 19188
rect 15378 19176 15384 19228
rect 15436 19216 15442 19228
rect 15841 19219 15899 19225
rect 15841 19216 15853 19219
rect 15436 19188 15853 19216
rect 15436 19176 15442 19188
rect 15841 19185 15853 19188
rect 15887 19185 15899 19219
rect 15841 19179 15899 19185
rect 17129 19219 17187 19225
rect 17129 19185 17141 19219
rect 17175 19216 17187 19219
rect 17678 19216 17684 19228
rect 17175 19188 17684 19216
rect 17175 19185 17187 19188
rect 17129 19179 17187 19185
rect 17678 19176 17684 19188
rect 17736 19176 17742 19228
rect 11146 19148 11152 19160
rect 9784 19120 11152 19148
rect 9677 19111 9735 19117
rect 5868 19052 6316 19080
rect 6356 19083 6414 19089
rect 5868 19040 5874 19052
rect 6356 19049 6368 19083
rect 6402 19080 6414 19083
rect 7558 19080 7564 19092
rect 6402 19052 7564 19080
rect 6402 19049 6414 19052
rect 6356 19043 6414 19049
rect 7558 19040 7564 19052
rect 7616 19040 7622 19092
rect 5442 19012 5448 19024
rect 5403 18984 5448 19012
rect 5442 18972 5448 18984
rect 5500 18972 5506 19024
rect 6086 18972 6092 19024
rect 6144 19012 6150 19024
rect 6546 19012 6552 19024
rect 6144 18984 6552 19012
rect 6144 18972 6150 18984
rect 6546 18972 6552 18984
rect 6604 19012 6610 19024
rect 7760 19012 7788 19111
rect 7926 19040 7932 19092
rect 7984 19089 7990 19092
rect 7984 19083 8048 19089
rect 7984 19049 8002 19083
rect 8036 19080 8048 19083
rect 8202 19080 8208 19092
rect 8036 19052 8208 19080
rect 8036 19049 8048 19052
rect 7984 19043 8048 19049
rect 7984 19040 7990 19043
rect 8202 19040 8208 19052
rect 8260 19040 8266 19092
rect 9692 19012 9720 19111
rect 11146 19108 11152 19120
rect 11204 19108 11210 19160
rect 12342 19148 12348 19160
rect 12303 19120 12348 19148
rect 12342 19108 12348 19120
rect 12400 19108 12406 19160
rect 13354 19108 13360 19160
rect 13412 19148 13418 19160
rect 13412 19120 15884 19148
rect 13412 19108 13418 19120
rect 9950 19089 9956 19092
rect 9944 19080 9956 19089
rect 9911 19052 9956 19080
rect 9944 19043 9956 19052
rect 9950 19040 9956 19043
rect 10008 19040 10014 19092
rect 12618 19089 12624 19092
rect 12612 19080 12624 19089
rect 12579 19052 12624 19080
rect 12612 19043 12624 19052
rect 12618 19040 12624 19043
rect 12676 19040 12682 19092
rect 15746 19080 15752 19092
rect 13556 19052 15608 19080
rect 15707 19052 15752 19080
rect 10686 19012 10692 19024
rect 6604 18984 10692 19012
rect 6604 18972 6610 18984
rect 10686 18972 10692 18984
rect 10744 18972 10750 19024
rect 11054 19012 11060 19024
rect 11015 18984 11060 19012
rect 11054 18972 11060 18984
rect 11112 18972 11118 19024
rect 11882 18972 11888 19024
rect 11940 19012 11946 19024
rect 13556 19012 13584 19052
rect 13722 19012 13728 19024
rect 11940 18984 13584 19012
rect 13683 18984 13728 19012
rect 11940 18972 11946 18984
rect 13722 18972 13728 18984
rect 13780 18972 13786 19024
rect 13814 18972 13820 19024
rect 13872 19012 13878 19024
rect 14001 19015 14059 19021
rect 14001 19012 14013 19015
rect 13872 18984 14013 19012
rect 13872 18972 13878 18984
rect 14001 18981 14013 18984
rect 14047 18981 14059 19015
rect 14001 18975 14059 18981
rect 15289 19015 15347 19021
rect 15289 18981 15301 19015
rect 15335 19012 15347 19015
rect 15470 19012 15476 19024
rect 15335 18984 15476 19012
rect 15335 18981 15347 18984
rect 15289 18975 15347 18981
rect 15470 18972 15476 18984
rect 15528 18972 15534 19024
rect 15580 19012 15608 19052
rect 15746 19040 15752 19052
rect 15804 19040 15810 19092
rect 15654 19012 15660 19024
rect 15580 18984 15660 19012
rect 15654 18972 15660 18984
rect 15712 19012 15718 19024
rect 15856 19012 15884 19120
rect 16758 19108 16764 19160
rect 16816 19148 16822 19160
rect 16853 19151 16911 19157
rect 16853 19148 16865 19151
rect 16816 19120 16865 19148
rect 16816 19108 16822 19120
rect 16853 19117 16865 19120
rect 16899 19117 16911 19151
rect 16853 19111 16911 19117
rect 18141 19151 18199 19157
rect 18141 19117 18153 19151
rect 18187 19148 18199 19151
rect 18874 19148 18880 19160
rect 18187 19120 18880 19148
rect 18187 19117 18199 19120
rect 18141 19111 18199 19117
rect 18874 19108 18880 19120
rect 18932 19108 18938 19160
rect 19521 19151 19579 19157
rect 19521 19117 19533 19151
rect 19567 19117 19579 19151
rect 19521 19111 19579 19117
rect 19797 19151 19855 19157
rect 19797 19117 19809 19151
rect 19843 19148 19855 19151
rect 20257 19151 20315 19157
rect 20257 19148 20269 19151
rect 19843 19120 20269 19148
rect 19843 19117 19855 19120
rect 19797 19111 19855 19117
rect 20257 19117 20269 19120
rect 20303 19117 20315 19151
rect 20257 19111 20315 19117
rect 18782 19080 18788 19092
rect 18743 19052 18788 19080
rect 18782 19040 18788 19052
rect 18840 19040 18846 19092
rect 19536 19080 19564 19111
rect 18892 19052 19564 19080
rect 18892 19012 18920 19052
rect 15712 18984 15805 19012
rect 15856 18984 18920 19012
rect 15712 18972 15718 18984
rect 19242 18972 19248 19024
rect 19300 19012 19306 19024
rect 20441 19015 20499 19021
rect 20441 19012 20453 19015
rect 19300 18984 20453 19012
rect 19300 18972 19306 18984
rect 20441 18981 20453 18984
rect 20487 18981 20499 19015
rect 20441 18975 20499 18981
rect 1104 18922 21620 18944
rect 1104 18870 7846 18922
rect 7898 18870 7910 18922
rect 7962 18870 7974 18922
rect 8026 18870 8038 18922
rect 8090 18870 14710 18922
rect 14762 18870 14774 18922
rect 14826 18870 14838 18922
rect 14890 18870 14902 18922
rect 14954 18870 21620 18922
rect 1104 18848 21620 18870
rect 3789 18811 3847 18817
rect 3789 18777 3801 18811
rect 3835 18808 3847 18811
rect 4706 18808 4712 18820
rect 3835 18780 4712 18808
rect 3835 18777 3847 18780
rect 3789 18771 3847 18777
rect 4706 18768 4712 18780
rect 4764 18768 4770 18820
rect 5166 18808 5172 18820
rect 5127 18780 5172 18808
rect 5166 18768 5172 18780
rect 5224 18768 5230 18820
rect 8294 18808 8300 18820
rect 6288 18780 8300 18808
rect 2498 18700 2504 18752
rect 2556 18740 2562 18752
rect 6288 18740 6316 18780
rect 8294 18768 8300 18780
rect 8352 18768 8358 18820
rect 9122 18768 9128 18820
rect 9180 18808 9186 18820
rect 9677 18811 9735 18817
rect 9677 18808 9689 18811
rect 9180 18780 9689 18808
rect 9180 18768 9186 18780
rect 9677 18777 9689 18780
rect 9723 18777 9735 18811
rect 9677 18771 9735 18777
rect 9858 18768 9864 18820
rect 9916 18808 9922 18820
rect 9916 18780 11192 18808
rect 9916 18768 9922 18780
rect 2556 18712 6316 18740
rect 2556 18700 2562 18712
rect 6362 18700 6368 18752
rect 6420 18740 6426 18752
rect 9398 18740 9404 18752
rect 6420 18712 9404 18740
rect 6420 18700 6426 18712
rect 9398 18700 9404 18712
rect 9456 18700 9462 18752
rect 10956 18743 11014 18749
rect 10956 18709 10968 18743
rect 11002 18740 11014 18743
rect 11054 18740 11060 18752
rect 11002 18712 11060 18740
rect 11002 18709 11014 18712
rect 10956 18703 11014 18709
rect 11054 18700 11060 18712
rect 11112 18700 11118 18752
rect 11164 18740 11192 18780
rect 12434 18768 12440 18820
rect 12492 18808 12498 18820
rect 14829 18811 14887 18817
rect 12492 18780 14596 18808
rect 12492 18768 12498 18780
rect 12897 18743 12955 18749
rect 12897 18740 12909 18743
rect 11164 18712 12909 18740
rect 12897 18709 12909 18712
rect 12943 18709 12955 18743
rect 12897 18703 12955 18709
rect 2676 18675 2734 18681
rect 2676 18641 2688 18675
rect 2722 18672 2734 18675
rect 2958 18672 2964 18684
rect 2722 18644 2964 18672
rect 2722 18641 2734 18644
rect 2676 18635 2734 18641
rect 2958 18632 2964 18644
rect 3016 18632 3022 18684
rect 5077 18675 5135 18681
rect 5077 18641 5089 18675
rect 5123 18672 5135 18675
rect 5721 18675 5779 18681
rect 5721 18672 5733 18675
rect 5123 18644 5733 18672
rect 5123 18641 5135 18644
rect 5077 18635 5135 18641
rect 5721 18641 5733 18644
rect 5767 18641 5779 18675
rect 5721 18635 5779 18641
rect 7745 18675 7803 18681
rect 7745 18641 7757 18675
rect 7791 18672 7803 18675
rect 8389 18675 8447 18681
rect 8389 18672 8401 18675
rect 7791 18644 8401 18672
rect 7791 18641 7803 18644
rect 7745 18635 7803 18641
rect 8389 18641 8401 18644
rect 8435 18641 8447 18675
rect 9582 18672 9588 18684
rect 9495 18644 9588 18672
rect 8389 18635 8447 18641
rect 9582 18632 9588 18644
rect 9640 18632 9646 18684
rect 10686 18672 10692 18684
rect 10647 18644 10692 18672
rect 10686 18632 10692 18644
rect 10744 18632 10750 18684
rect 12802 18672 12808 18684
rect 12763 18644 12808 18672
rect 12802 18632 12808 18644
rect 12860 18632 12866 18684
rect 13464 18681 13492 18780
rect 13722 18681 13728 18684
rect 13449 18675 13507 18681
rect 13449 18641 13461 18675
rect 13495 18641 13507 18675
rect 13716 18672 13728 18681
rect 13635 18644 13728 18672
rect 13449 18635 13507 18641
rect 13716 18635 13728 18644
rect 13780 18672 13786 18684
rect 13998 18672 14004 18684
rect 13780 18644 14004 18672
rect 13722 18632 13728 18635
rect 13780 18632 13786 18644
rect 13998 18632 14004 18644
rect 14056 18632 14062 18684
rect 14568 18672 14596 18780
rect 14829 18777 14841 18811
rect 14875 18777 14887 18811
rect 16758 18808 16764 18820
rect 16719 18780 16764 18808
rect 14829 18771 14887 18777
rect 14844 18740 14872 18771
rect 16758 18768 16764 18780
rect 16816 18768 16822 18820
rect 17954 18768 17960 18820
rect 18012 18808 18018 18820
rect 20070 18808 20076 18820
rect 18012 18780 20076 18808
rect 18012 18768 18018 18780
rect 20070 18768 20076 18780
rect 20128 18768 20134 18820
rect 20714 18808 20720 18820
rect 20675 18780 20720 18808
rect 20714 18768 20720 18780
rect 20772 18768 20778 18820
rect 15378 18749 15384 18752
rect 15372 18740 15384 18749
rect 14844 18712 15384 18740
rect 15372 18703 15384 18712
rect 15378 18700 15384 18703
rect 15436 18700 15442 18752
rect 15470 18700 15476 18752
rect 15528 18740 15534 18752
rect 17221 18743 17279 18749
rect 17221 18740 17233 18743
rect 15528 18712 17233 18740
rect 15528 18700 15534 18712
rect 17221 18709 17233 18712
rect 17267 18709 17279 18743
rect 17221 18703 17279 18709
rect 18325 18743 18383 18749
rect 18325 18709 18337 18743
rect 18371 18740 18383 18743
rect 18506 18740 18512 18752
rect 18371 18712 18512 18740
rect 18371 18709 18383 18712
rect 18325 18703 18383 18709
rect 18506 18700 18512 18712
rect 18564 18700 18570 18752
rect 15105 18675 15163 18681
rect 15105 18672 15117 18675
rect 14568 18644 15117 18672
rect 15105 18641 15117 18644
rect 15151 18641 15163 18675
rect 15105 18635 15163 18641
rect 16574 18632 16580 18684
rect 16632 18672 16638 18684
rect 17129 18675 17187 18681
rect 17129 18672 17141 18675
rect 16632 18644 17141 18672
rect 16632 18632 16638 18644
rect 17129 18641 17141 18644
rect 17175 18641 17187 18675
rect 17129 18635 17187 18641
rect 17954 18632 17960 18684
rect 18012 18672 18018 18684
rect 18049 18675 18107 18681
rect 18049 18672 18061 18675
rect 18012 18644 18061 18672
rect 18012 18632 18018 18644
rect 18049 18641 18061 18644
rect 18095 18641 18107 18675
rect 19518 18672 19524 18684
rect 19479 18644 19524 18672
rect 18049 18635 18107 18641
rect 19518 18632 19524 18644
rect 19576 18632 19582 18684
rect 19794 18632 19800 18684
rect 19852 18672 19858 18684
rect 20533 18675 20591 18681
rect 20533 18672 20545 18675
rect 19852 18644 20545 18672
rect 19852 18632 19858 18644
rect 20533 18641 20545 18644
rect 20579 18641 20591 18675
rect 20533 18635 20591 18641
rect 2406 18604 2412 18616
rect 2367 18576 2412 18604
rect 2406 18564 2412 18576
rect 2464 18564 2470 18616
rect 5353 18607 5411 18613
rect 5353 18573 5365 18607
rect 5399 18604 5411 18607
rect 5442 18604 5448 18616
rect 5399 18576 5448 18604
rect 5399 18573 5411 18576
rect 5353 18567 5411 18573
rect 5442 18564 5448 18576
rect 5500 18564 5506 18616
rect 7650 18564 7656 18616
rect 7708 18604 7714 18616
rect 7837 18607 7895 18613
rect 7837 18604 7849 18607
rect 7708 18576 7849 18604
rect 7708 18564 7714 18576
rect 7837 18573 7849 18576
rect 7883 18573 7895 18607
rect 7837 18567 7895 18573
rect 8021 18607 8079 18613
rect 8021 18573 8033 18607
rect 8067 18604 8079 18607
rect 8202 18604 8208 18616
rect 8067 18576 8208 18604
rect 8067 18573 8079 18576
rect 8021 18567 8079 18573
rect 8202 18564 8208 18576
rect 8260 18564 8266 18616
rect 6822 18536 6828 18548
rect 4632 18508 6828 18536
rect 290 18428 296 18480
rect 348 18468 354 18480
rect 4632 18468 4660 18508
rect 6822 18496 6828 18508
rect 6880 18496 6886 18548
rect 7466 18496 7472 18548
rect 7524 18536 7530 18548
rect 8386 18536 8392 18548
rect 7524 18508 8392 18536
rect 7524 18496 7530 18508
rect 8386 18496 8392 18508
rect 8444 18496 8450 18548
rect 9600 18536 9628 18632
rect 9861 18607 9919 18613
rect 9861 18573 9873 18607
rect 9907 18604 9919 18607
rect 9950 18604 9956 18616
rect 9907 18576 9956 18604
rect 9907 18573 9919 18576
rect 9861 18567 9919 18573
rect 9950 18564 9956 18576
rect 10008 18564 10014 18616
rect 10226 18604 10232 18616
rect 10187 18576 10232 18604
rect 10226 18564 10232 18576
rect 10284 18564 10290 18616
rect 12989 18607 13047 18613
rect 12989 18573 13001 18607
rect 13035 18573 13047 18607
rect 17313 18607 17371 18613
rect 17313 18604 17325 18607
rect 12989 18567 13047 18573
rect 16500 18576 17325 18604
rect 10686 18536 10692 18548
rect 9600 18508 10692 18536
rect 10686 18496 10692 18508
rect 10744 18496 10750 18548
rect 12069 18539 12127 18545
rect 12069 18505 12081 18539
rect 12115 18536 12127 18539
rect 12618 18536 12624 18548
rect 12115 18508 12624 18536
rect 12115 18505 12127 18508
rect 12069 18499 12127 18505
rect 12618 18496 12624 18508
rect 12676 18536 12682 18548
rect 13004 18536 13032 18567
rect 12676 18508 13032 18536
rect 12676 18496 12682 18508
rect 348 18440 4660 18468
rect 4709 18471 4767 18477
rect 348 18428 354 18440
rect 4709 18437 4721 18471
rect 4755 18468 4767 18471
rect 5166 18468 5172 18480
rect 4755 18440 5172 18468
rect 4755 18437 4767 18440
rect 4709 18431 4767 18437
rect 5166 18428 5172 18440
rect 5224 18428 5230 18480
rect 7377 18471 7435 18477
rect 7377 18437 7389 18471
rect 7423 18468 7435 18471
rect 9122 18468 9128 18480
rect 7423 18440 9128 18468
rect 7423 18437 7435 18440
rect 7377 18431 7435 18437
rect 9122 18428 9128 18440
rect 9180 18428 9186 18480
rect 9217 18471 9275 18477
rect 9217 18437 9229 18471
rect 9263 18468 9275 18471
rect 10870 18468 10876 18480
rect 9263 18440 10876 18468
rect 9263 18437 9275 18440
rect 9217 18431 9275 18437
rect 10870 18428 10876 18440
rect 10928 18428 10934 18480
rect 10962 18428 10968 18480
rect 11020 18468 11026 18480
rect 11698 18468 11704 18480
rect 11020 18440 11704 18468
rect 11020 18428 11026 18440
rect 11698 18428 11704 18440
rect 11756 18428 11762 18480
rect 12437 18471 12495 18477
rect 12437 18437 12449 18471
rect 12483 18468 12495 18471
rect 13262 18468 13268 18480
rect 12483 18440 13268 18468
rect 12483 18437 12495 18440
rect 12437 18431 12495 18437
rect 13262 18428 13268 18440
rect 13320 18428 13326 18480
rect 16390 18428 16396 18480
rect 16448 18468 16454 18480
rect 16500 18477 16528 18576
rect 17313 18573 17325 18576
rect 17359 18573 17371 18607
rect 19702 18604 19708 18616
rect 19663 18576 19708 18604
rect 17313 18567 17371 18573
rect 19702 18564 19708 18576
rect 19760 18564 19766 18616
rect 16485 18471 16543 18477
rect 16485 18468 16497 18471
rect 16448 18440 16497 18468
rect 16448 18428 16454 18440
rect 16485 18437 16497 18440
rect 16531 18437 16543 18471
rect 16485 18431 16543 18437
rect 16942 18428 16948 18480
rect 17000 18468 17006 18480
rect 21174 18468 21180 18480
rect 17000 18440 21180 18468
rect 17000 18428 17006 18440
rect 21174 18428 21180 18440
rect 21232 18428 21238 18480
rect 1104 18378 21620 18400
rect 1104 18326 4414 18378
rect 4466 18326 4478 18378
rect 4530 18326 4542 18378
rect 4594 18326 4606 18378
rect 4658 18326 11278 18378
rect 11330 18326 11342 18378
rect 11394 18326 11406 18378
rect 11458 18326 11470 18378
rect 11522 18326 18142 18378
rect 18194 18326 18206 18378
rect 18258 18326 18270 18378
rect 18322 18326 18334 18378
rect 18386 18326 21620 18378
rect 1104 18304 21620 18326
rect 1946 18224 1952 18276
rect 2004 18264 2010 18276
rect 6730 18264 6736 18276
rect 2004 18236 6736 18264
rect 2004 18224 2010 18236
rect 6730 18224 6736 18236
rect 6788 18224 6794 18276
rect 6822 18224 6828 18276
rect 6880 18264 6886 18276
rect 9030 18264 9036 18276
rect 6880 18236 9036 18264
rect 6880 18224 6886 18236
rect 9030 18224 9036 18236
rect 9088 18224 9094 18276
rect 9122 18224 9128 18276
rect 9180 18264 9186 18276
rect 13354 18264 13360 18276
rect 9180 18236 13216 18264
rect 13315 18236 13360 18264
rect 9180 18224 9186 18236
rect 6914 18156 6920 18208
rect 6972 18196 6978 18208
rect 10413 18199 10471 18205
rect 6972 18168 8340 18196
rect 6972 18156 6978 18168
rect 7558 18088 7564 18140
rect 7616 18128 7622 18140
rect 8205 18131 8263 18137
rect 8205 18128 8217 18131
rect 7616 18100 8217 18128
rect 7616 18088 7622 18100
rect 8205 18097 8217 18100
rect 8251 18097 8263 18131
rect 8312 18128 8340 18168
rect 10413 18165 10425 18199
rect 10459 18196 10471 18199
rect 13188 18196 13216 18236
rect 13354 18224 13360 18236
rect 13412 18224 13418 18276
rect 13906 18224 13912 18276
rect 13964 18264 13970 18276
rect 14550 18264 14556 18276
rect 13964 18236 14556 18264
rect 13964 18224 13970 18236
rect 14550 18224 14556 18236
rect 14608 18224 14614 18276
rect 15838 18224 15844 18276
rect 15896 18264 15902 18276
rect 19702 18264 19708 18276
rect 15896 18236 19708 18264
rect 15896 18224 15902 18236
rect 19702 18224 19708 18236
rect 19760 18224 19766 18276
rect 19797 18267 19855 18273
rect 19797 18233 19809 18267
rect 19843 18264 19855 18267
rect 19886 18264 19892 18276
rect 19843 18236 19892 18264
rect 19843 18233 19855 18236
rect 19797 18227 19855 18233
rect 19886 18224 19892 18236
rect 19944 18224 19950 18276
rect 16393 18199 16451 18205
rect 10459 18168 13124 18196
rect 13188 18168 14136 18196
rect 10459 18165 10471 18168
rect 10413 18159 10471 18165
rect 10686 18128 10692 18140
rect 8312 18100 10692 18128
rect 8205 18091 8263 18097
rect 10686 18088 10692 18100
rect 10744 18088 10750 18140
rect 10870 18128 10876 18140
rect 10831 18100 10876 18128
rect 10870 18088 10876 18100
rect 10928 18088 10934 18140
rect 11054 18128 11060 18140
rect 11015 18100 11060 18128
rect 11054 18088 11060 18100
rect 11112 18088 11118 18140
rect 11514 18088 11520 18140
rect 11572 18128 11578 18140
rect 11974 18128 11980 18140
rect 11572 18100 11980 18128
rect 11572 18088 11578 18100
rect 11974 18088 11980 18100
rect 12032 18088 12038 18140
rect 3602 18020 3608 18072
rect 3660 18060 3666 18072
rect 4246 18060 4252 18072
rect 3660 18032 4252 18060
rect 3660 18020 3666 18032
rect 4246 18020 4252 18032
rect 4304 18020 4310 18072
rect 5166 18060 5172 18072
rect 5127 18032 5172 18060
rect 5166 18020 5172 18032
rect 5224 18020 5230 18072
rect 8113 18063 8171 18069
rect 8113 18029 8125 18063
rect 8159 18060 8171 18063
rect 8570 18060 8576 18072
rect 8159 18032 8576 18060
rect 8159 18029 8171 18032
rect 8113 18023 8171 18029
rect 8570 18020 8576 18032
rect 8628 18020 8634 18072
rect 10226 18020 10232 18072
rect 10284 18060 10290 18072
rect 10781 18063 10839 18069
rect 10781 18060 10793 18063
rect 10284 18032 10793 18060
rect 10284 18020 10290 18032
rect 10781 18029 10793 18032
rect 10827 18029 10839 18063
rect 13096 18060 13124 18168
rect 13909 18131 13967 18137
rect 13909 18097 13921 18131
rect 13955 18128 13967 18131
rect 14108 18128 14136 18168
rect 16393 18165 16405 18199
rect 16439 18196 16451 18199
rect 19518 18196 19524 18208
rect 16439 18168 19524 18196
rect 16439 18165 16451 18168
rect 16393 18159 16451 18165
rect 19518 18156 19524 18168
rect 19576 18156 19582 18208
rect 16574 18128 16580 18140
rect 13955 18100 14044 18128
rect 14108 18100 16436 18128
rect 16535 18100 16580 18128
rect 13955 18097 13967 18100
rect 13909 18091 13967 18097
rect 14016 18072 14044 18100
rect 13096 18032 13952 18060
rect 10781 18023 10839 18029
rect 5445 17995 5503 18001
rect 5445 17961 5457 17995
rect 5491 17992 5503 17995
rect 10594 17992 10600 18004
rect 5491 17964 10600 17992
rect 5491 17961 5503 17964
rect 5445 17955 5503 17961
rect 10594 17952 10600 17964
rect 10652 17952 10658 18004
rect 13722 17952 13728 18004
rect 13780 17992 13786 18004
rect 13780 17964 13825 17992
rect 13780 17952 13786 17964
rect 3050 17884 3056 17936
rect 3108 17924 3114 17936
rect 5902 17924 5908 17936
rect 3108 17896 5908 17924
rect 3108 17884 3114 17896
rect 5902 17884 5908 17896
rect 5960 17884 5966 17936
rect 7650 17924 7656 17936
rect 7611 17896 7656 17924
rect 7650 17884 7656 17896
rect 7708 17884 7714 17936
rect 8021 17927 8079 17933
rect 8021 17893 8033 17927
rect 8067 17924 8079 17927
rect 8202 17924 8208 17936
rect 8067 17896 8208 17924
rect 8067 17893 8079 17896
rect 8021 17887 8079 17893
rect 8202 17884 8208 17896
rect 8260 17884 8266 17936
rect 8294 17884 8300 17936
rect 8352 17924 8358 17936
rect 9950 17924 9956 17936
rect 8352 17896 9956 17924
rect 8352 17884 8358 17896
rect 9950 17884 9956 17896
rect 10008 17884 10014 17936
rect 11606 17884 11612 17936
rect 11664 17924 11670 17936
rect 12066 17924 12072 17936
rect 11664 17896 12072 17924
rect 11664 17884 11670 17896
rect 12066 17884 12072 17896
rect 12124 17884 12130 17936
rect 12526 17884 12532 17936
rect 12584 17924 12590 17936
rect 12986 17924 12992 17936
rect 12584 17896 12992 17924
rect 12584 17884 12590 17896
rect 12986 17884 12992 17896
rect 13044 17884 13050 17936
rect 13262 17884 13268 17936
rect 13320 17924 13326 17936
rect 13817 17927 13875 17933
rect 13817 17924 13829 17927
rect 13320 17896 13829 17924
rect 13320 17884 13326 17896
rect 13817 17893 13829 17896
rect 13863 17893 13875 17927
rect 13924 17924 13952 18032
rect 13998 18020 14004 18072
rect 14056 18020 14062 18072
rect 15286 18020 15292 18072
rect 15344 18060 15350 18072
rect 16298 18060 16304 18072
rect 15344 18032 16304 18060
rect 15344 18020 15350 18032
rect 16298 18020 16304 18032
rect 16356 18020 16362 18072
rect 16408 18060 16436 18100
rect 16574 18088 16580 18100
rect 16632 18088 16638 18140
rect 19702 18088 19708 18140
rect 19760 18128 19766 18140
rect 21910 18128 21916 18140
rect 19760 18100 21916 18128
rect 19760 18088 19766 18100
rect 21910 18088 21916 18100
rect 21968 18088 21974 18140
rect 19334 18060 19340 18072
rect 16408 18032 19340 18060
rect 19334 18020 19340 18032
rect 19392 18020 19398 18072
rect 19610 18060 19616 18072
rect 19571 18032 19616 18060
rect 19610 18020 19616 18032
rect 19668 18020 19674 18072
rect 20257 18063 20315 18069
rect 20257 18029 20269 18063
rect 20303 18029 20315 18063
rect 20257 18023 20315 18029
rect 14182 17952 14188 18004
rect 14240 17992 14246 18004
rect 15102 17992 15108 18004
rect 14240 17964 15108 17992
rect 14240 17952 14246 17964
rect 15102 17952 15108 17964
rect 15160 17952 15166 18004
rect 15194 17952 15200 18004
rect 15252 17992 15258 18004
rect 20272 17992 20300 18023
rect 20622 18020 20628 18072
rect 20680 18060 20686 18072
rect 21358 18060 21364 18072
rect 20680 18032 21364 18060
rect 20680 18020 20686 18032
rect 21358 18020 21364 18032
rect 21416 18020 21422 18072
rect 15252 17964 20300 17992
rect 15252 17952 15258 17964
rect 16393 17927 16451 17933
rect 16393 17924 16405 17927
rect 13924 17896 16405 17924
rect 13817 17887 13875 17893
rect 16393 17893 16405 17896
rect 16439 17893 16451 17927
rect 16393 17887 16451 17893
rect 16482 17884 16488 17936
rect 16540 17924 16546 17936
rect 19518 17924 19524 17936
rect 16540 17896 19524 17924
rect 16540 17884 16546 17896
rect 19518 17884 19524 17896
rect 19576 17884 19582 17936
rect 19886 17884 19892 17936
rect 19944 17924 19950 17936
rect 20254 17924 20260 17936
rect 19944 17896 20260 17924
rect 19944 17884 19950 17896
rect 20254 17884 20260 17896
rect 20312 17884 20318 17936
rect 20438 17924 20444 17936
rect 20399 17896 20444 17924
rect 20438 17884 20444 17896
rect 20496 17884 20502 17936
rect 20806 17884 20812 17936
rect 20864 17924 20870 17936
rect 22462 17924 22468 17936
rect 20864 17896 22468 17924
rect 20864 17884 20870 17896
rect 22462 17884 22468 17896
rect 22520 17884 22526 17936
rect 1104 17834 21620 17856
rect 1104 17782 7846 17834
rect 7898 17782 7910 17834
rect 7962 17782 7974 17834
rect 8026 17782 8038 17834
rect 8090 17782 14710 17834
rect 14762 17782 14774 17834
rect 14826 17782 14838 17834
rect 14890 17782 14902 17834
rect 14954 17782 21620 17834
rect 1104 17760 21620 17782
rect 2958 17720 2964 17732
rect 2919 17692 2964 17720
rect 2958 17680 2964 17692
rect 3016 17680 3022 17732
rect 17034 17720 17040 17732
rect 16995 17692 17040 17720
rect 17034 17680 17040 17692
rect 17092 17680 17098 17732
rect 20346 17720 20352 17732
rect 20307 17692 20352 17720
rect 20346 17680 20352 17692
rect 20404 17680 20410 17732
rect 20898 17720 20904 17732
rect 20859 17692 20904 17720
rect 20898 17680 20904 17692
rect 20956 17680 20962 17732
rect 2406 17652 2412 17664
rect 1596 17624 2412 17652
rect 1596 17528 1624 17624
rect 2406 17612 2412 17624
rect 2464 17652 2470 17664
rect 5160 17655 5218 17661
rect 2464 17624 4936 17652
rect 2464 17612 2470 17624
rect 1848 17587 1906 17593
rect 1848 17553 1860 17587
rect 1894 17584 1906 17587
rect 3142 17584 3148 17596
rect 1894 17556 3148 17584
rect 1894 17553 1906 17556
rect 1848 17547 1906 17553
rect 3142 17544 3148 17556
rect 3200 17544 3206 17596
rect 4908 17593 4936 17624
rect 5160 17621 5172 17655
rect 5206 17652 5218 17655
rect 5442 17652 5448 17664
rect 5206 17624 5448 17652
rect 5206 17621 5218 17624
rect 5160 17615 5218 17621
rect 5442 17612 5448 17624
rect 5500 17612 5506 17664
rect 5626 17612 5632 17664
rect 5684 17652 5690 17664
rect 18874 17652 18880 17664
rect 5684 17624 18880 17652
rect 5684 17612 5690 17624
rect 18874 17612 18880 17624
rect 18932 17612 18938 17664
rect 4893 17587 4951 17593
rect 4893 17553 4905 17587
rect 4939 17553 4951 17587
rect 4893 17547 4951 17553
rect 14458 17544 14464 17596
rect 14516 17584 14522 17596
rect 16945 17587 17003 17593
rect 16945 17584 16957 17587
rect 14516 17556 16957 17584
rect 14516 17544 14522 17556
rect 16945 17553 16957 17556
rect 16991 17553 17003 17587
rect 16945 17547 17003 17553
rect 17218 17544 17224 17596
rect 17276 17584 17282 17596
rect 19337 17587 19395 17593
rect 19337 17584 19349 17587
rect 17276 17556 19349 17584
rect 17276 17544 17282 17556
rect 19337 17553 19349 17556
rect 19383 17553 19395 17587
rect 20162 17584 20168 17596
rect 20123 17556 20168 17584
rect 19337 17547 19395 17553
rect 20162 17544 20168 17556
rect 20220 17544 20226 17596
rect 20717 17587 20775 17593
rect 20717 17553 20729 17587
rect 20763 17553 20775 17587
rect 20717 17547 20775 17553
rect 1578 17516 1584 17528
rect 1539 17488 1584 17516
rect 1578 17476 1584 17488
rect 1636 17476 1642 17528
rect 3326 17516 3332 17528
rect 3287 17488 3332 17516
rect 3326 17476 3332 17488
rect 3384 17476 3390 17528
rect 10686 17476 10692 17528
rect 10744 17516 10750 17528
rect 16758 17516 16764 17528
rect 10744 17488 16764 17516
rect 10744 17476 10750 17488
rect 16758 17476 16764 17488
rect 16816 17476 16822 17528
rect 17126 17476 17132 17528
rect 17184 17516 17190 17528
rect 19613 17519 19671 17525
rect 17184 17488 17229 17516
rect 17184 17476 17190 17488
rect 19613 17485 19625 17519
rect 19659 17516 19671 17519
rect 20732 17516 20760 17547
rect 19659 17488 20760 17516
rect 19659 17485 19671 17488
rect 19613 17479 19671 17485
rect 6273 17383 6331 17389
rect 6273 17349 6285 17383
rect 6319 17380 6331 17383
rect 9122 17380 9128 17392
rect 6319 17352 9128 17380
rect 6319 17349 6331 17352
rect 6273 17343 6331 17349
rect 9122 17340 9128 17352
rect 9180 17340 9186 17392
rect 12802 17340 12808 17392
rect 12860 17380 12866 17392
rect 14274 17380 14280 17392
rect 12860 17352 14280 17380
rect 12860 17340 12866 17352
rect 14274 17340 14280 17352
rect 14332 17340 14338 17392
rect 16577 17383 16635 17389
rect 16577 17349 16589 17383
rect 16623 17380 16635 17383
rect 18598 17380 18604 17392
rect 16623 17352 18604 17380
rect 16623 17349 16635 17352
rect 16577 17343 16635 17349
rect 18598 17340 18604 17352
rect 18656 17340 18662 17392
rect 21726 17312 21732 17324
rect 1104 17290 21620 17312
rect 1104 17238 4414 17290
rect 4466 17238 4478 17290
rect 4530 17238 4542 17290
rect 4594 17238 4606 17290
rect 4658 17238 11278 17290
rect 11330 17238 11342 17290
rect 11394 17238 11406 17290
rect 11458 17238 11470 17290
rect 11522 17238 18142 17290
rect 18194 17238 18206 17290
rect 18258 17238 18270 17290
rect 18322 17238 18334 17290
rect 18386 17238 21620 17290
rect 21687 17284 21732 17312
rect 21726 17272 21732 17284
rect 21784 17272 21790 17324
rect 1104 17216 21620 17238
rect 4062 17136 4068 17188
rect 4120 17176 4126 17188
rect 4120 17148 9260 17176
rect 4120 17136 4126 17148
rect 3142 17068 3148 17120
rect 3200 17108 3206 17120
rect 3200 17080 4660 17108
rect 3200 17068 3206 17080
rect 2958 17000 2964 17052
rect 3016 17040 3022 17052
rect 3513 17043 3571 17049
rect 3513 17040 3525 17043
rect 3016 17012 3525 17040
rect 3016 17000 3022 17012
rect 3513 17009 3525 17012
rect 3559 17009 3571 17043
rect 3513 17003 3571 17009
rect 4154 17000 4160 17052
rect 4212 17040 4218 17052
rect 4632 17049 4660 17080
rect 7558 17068 7564 17120
rect 7616 17108 7622 17120
rect 7929 17111 7987 17117
rect 7929 17108 7941 17111
rect 7616 17080 7941 17108
rect 7616 17068 7622 17080
rect 7929 17077 7941 17080
rect 7975 17077 7987 17111
rect 7929 17071 7987 17077
rect 4525 17043 4583 17049
rect 4525 17040 4537 17043
rect 4212 17012 4537 17040
rect 4212 17000 4218 17012
rect 4525 17009 4537 17012
rect 4571 17009 4583 17043
rect 4525 17003 4583 17009
rect 4617 17043 4675 17049
rect 4617 17009 4629 17043
rect 4663 17009 4675 17043
rect 4617 17003 4675 17009
rect 5534 17000 5540 17052
rect 5592 17040 5598 17052
rect 9122 17040 9128 17052
rect 5592 17012 6684 17040
rect 9083 17012 9128 17040
rect 5592 17000 5598 17012
rect 3326 16972 3332 16984
rect 3287 16944 3332 16972
rect 3326 16932 3332 16944
rect 3384 16932 3390 16984
rect 5442 16932 5448 16984
rect 5500 16972 5506 16984
rect 6546 16972 6552 16984
rect 5500 16944 6552 16972
rect 5500 16932 5506 16944
rect 6546 16932 6552 16944
rect 6604 16932 6610 16984
rect 6656 16972 6684 17012
rect 9122 17000 9128 17012
rect 9180 17000 9186 17052
rect 9033 16975 9091 16981
rect 9033 16972 9045 16975
rect 6656 16944 9045 16972
rect 9033 16941 9045 16944
rect 9079 16941 9091 16975
rect 9232 16972 9260 17148
rect 11146 17136 11152 17188
rect 11204 17176 11210 17188
rect 12805 17179 12863 17185
rect 11204 17148 12296 17176
rect 11204 17136 11210 17148
rect 10318 17040 10324 17052
rect 10279 17012 10324 17040
rect 10318 17000 10324 17012
rect 10376 17000 10382 17052
rect 12268 17049 12296 17148
rect 12805 17145 12817 17179
rect 12851 17176 12863 17179
rect 17218 17176 17224 17188
rect 12851 17148 17224 17176
rect 12851 17145 12863 17148
rect 12805 17139 12863 17145
rect 17218 17136 17224 17148
rect 17276 17136 17282 17188
rect 17954 17136 17960 17188
rect 18012 17176 18018 17188
rect 18141 17179 18199 17185
rect 18141 17176 18153 17179
rect 18012 17148 18153 17176
rect 18012 17136 18018 17148
rect 18141 17145 18153 17148
rect 18187 17145 18199 17179
rect 18141 17139 18199 17145
rect 20070 17136 20076 17188
rect 20128 17176 20134 17188
rect 20346 17176 20352 17188
rect 20128 17148 20352 17176
rect 20128 17136 20134 17148
rect 20346 17136 20352 17148
rect 20404 17136 20410 17188
rect 12342 17068 12348 17120
rect 12400 17108 12406 17120
rect 12400 17080 12480 17108
rect 12400 17068 12406 17080
rect 12452 17049 12480 17080
rect 12253 17043 12311 17049
rect 11992 17012 12204 17040
rect 11992 16972 12020 17012
rect 9232 16944 12020 16972
rect 12176 16972 12204 17012
rect 12253 17009 12265 17043
rect 12299 17009 12311 17043
rect 12253 17003 12311 17009
rect 12437 17043 12495 17049
rect 12437 17009 12449 17043
rect 12483 17009 12495 17043
rect 12437 17003 12495 17009
rect 12894 17000 12900 17052
rect 12952 17040 12958 17052
rect 13357 17043 13415 17049
rect 13357 17040 13369 17043
rect 12952 17012 13369 17040
rect 12952 17000 12958 17012
rect 13357 17009 13369 17012
rect 13403 17009 13415 17043
rect 18598 17040 18604 17052
rect 18559 17012 18604 17040
rect 13357 17003 13415 17009
rect 18598 17000 18604 17012
rect 18656 17000 18662 17052
rect 18693 17043 18751 17049
rect 18693 17009 18705 17043
rect 18739 17009 18751 17043
rect 20162 17040 20168 17052
rect 20123 17012 20168 17040
rect 18693 17003 18751 17009
rect 16482 16972 16488 16984
rect 12176 16944 15424 16972
rect 16443 16944 16488 16972
rect 9033 16935 9091 16941
rect 6816 16907 6874 16913
rect 6816 16873 6828 16907
rect 6862 16904 6874 16907
rect 7006 16904 7012 16916
rect 6862 16876 7012 16904
rect 6862 16873 6874 16876
rect 6816 16867 6874 16873
rect 7006 16864 7012 16876
rect 7064 16864 7070 16916
rect 10229 16907 10287 16913
rect 10229 16904 10241 16907
rect 8588 16876 10241 16904
rect 2958 16836 2964 16848
rect 2919 16808 2964 16836
rect 2958 16796 2964 16808
rect 3016 16796 3022 16848
rect 3421 16839 3479 16845
rect 3421 16805 3433 16839
rect 3467 16836 3479 16839
rect 4065 16839 4123 16845
rect 4065 16836 4077 16839
rect 3467 16808 4077 16836
rect 3467 16805 3479 16808
rect 3421 16799 3479 16805
rect 4065 16805 4077 16808
rect 4111 16805 4123 16839
rect 4065 16799 4123 16805
rect 4433 16839 4491 16845
rect 4433 16805 4445 16839
rect 4479 16836 4491 16839
rect 8294 16836 8300 16848
rect 4479 16808 8300 16836
rect 4479 16805 4491 16808
rect 4433 16799 4491 16805
rect 8294 16796 8300 16808
rect 8352 16796 8358 16848
rect 8588 16845 8616 16876
rect 10229 16873 10241 16876
rect 10275 16873 10287 16907
rect 13265 16907 13323 16913
rect 13265 16904 13277 16907
rect 10229 16867 10287 16873
rect 11808 16876 13277 16904
rect 8573 16839 8631 16845
rect 8573 16805 8585 16839
rect 8619 16805 8631 16839
rect 8938 16836 8944 16848
rect 8899 16808 8944 16836
rect 8573 16799 8631 16805
rect 8938 16796 8944 16808
rect 8996 16796 9002 16848
rect 9766 16836 9772 16848
rect 9727 16808 9772 16836
rect 9766 16796 9772 16808
rect 9824 16796 9830 16848
rect 10134 16836 10140 16848
rect 10095 16808 10140 16836
rect 10134 16796 10140 16808
rect 10192 16796 10198 16848
rect 11808 16845 11836 16876
rect 13265 16873 13277 16876
rect 13311 16873 13323 16907
rect 13265 16867 13323 16873
rect 11793 16839 11851 16845
rect 11793 16805 11805 16839
rect 11839 16805 11851 16839
rect 11793 16799 11851 16805
rect 11882 16796 11888 16848
rect 11940 16836 11946 16848
rect 12161 16839 12219 16845
rect 12161 16836 12173 16839
rect 11940 16808 12173 16836
rect 11940 16796 11946 16808
rect 12161 16805 12173 16808
rect 12207 16805 12219 16839
rect 13170 16836 13176 16848
rect 13131 16808 13176 16836
rect 12161 16799 12219 16805
rect 13170 16796 13176 16808
rect 13228 16796 13234 16848
rect 15396 16836 15424 16944
rect 16482 16932 16488 16944
rect 16540 16932 16546 16984
rect 16752 16975 16810 16981
rect 16752 16941 16764 16975
rect 16798 16972 16810 16975
rect 17126 16972 17132 16984
rect 16798 16944 17132 16972
rect 16798 16941 16810 16944
rect 16752 16935 16810 16941
rect 17126 16932 17132 16944
rect 17184 16932 17190 16984
rect 17957 16975 18015 16981
rect 17957 16941 17969 16975
rect 18003 16972 18015 16975
rect 18708 16972 18736 17003
rect 20162 17000 20168 17012
rect 20220 17000 20226 17052
rect 19242 16972 19248 16984
rect 18003 16944 18736 16972
rect 19203 16944 19248 16972
rect 18003 16941 18015 16944
rect 17957 16935 18015 16941
rect 19242 16932 19248 16944
rect 19300 16932 19306 16984
rect 19334 16932 19340 16984
rect 19392 16972 19398 16984
rect 19981 16975 20039 16981
rect 19981 16972 19993 16975
rect 19392 16944 19993 16972
rect 19392 16932 19398 16944
rect 19981 16941 19993 16944
rect 20027 16941 20039 16975
rect 19981 16935 20039 16941
rect 19521 16907 19579 16913
rect 19521 16873 19533 16907
rect 19567 16873 19579 16907
rect 19521 16867 19579 16873
rect 17865 16839 17923 16845
rect 17865 16836 17877 16839
rect 15396 16808 17877 16836
rect 17865 16805 17877 16808
rect 17911 16836 17923 16839
rect 17957 16839 18015 16845
rect 17957 16836 17969 16839
rect 17911 16808 17969 16836
rect 17911 16805 17923 16808
rect 17865 16799 17923 16805
rect 17957 16805 17969 16808
rect 18003 16805 18015 16839
rect 17957 16799 18015 16805
rect 18046 16796 18052 16848
rect 18104 16836 18110 16848
rect 18509 16839 18567 16845
rect 18509 16836 18521 16839
rect 18104 16808 18521 16836
rect 18104 16796 18110 16808
rect 18509 16805 18521 16808
rect 18555 16805 18567 16839
rect 19536 16836 19564 16867
rect 20438 16836 20444 16848
rect 19536 16808 20444 16836
rect 18509 16799 18567 16805
rect 20438 16796 20444 16808
rect 20496 16796 20502 16848
rect 1104 16746 21620 16768
rect 1104 16694 7846 16746
rect 7898 16694 7910 16746
rect 7962 16694 7974 16746
rect 8026 16694 8038 16746
rect 8090 16694 14710 16746
rect 14762 16694 14774 16746
rect 14826 16694 14838 16746
rect 14890 16694 14902 16746
rect 14954 16694 21620 16746
rect 1104 16672 21620 16694
rect 6917 16635 6975 16641
rect 6917 16601 6929 16635
rect 6963 16632 6975 16635
rect 10045 16635 10103 16641
rect 6963 16604 9996 16632
rect 6963 16601 6975 16604
rect 6917 16595 6975 16601
rect 4157 16567 4215 16573
rect 4157 16533 4169 16567
rect 4203 16564 4215 16567
rect 5626 16564 5632 16576
rect 4203 16536 5632 16564
rect 4203 16533 4215 16536
rect 4157 16527 4215 16533
rect 5626 16524 5632 16536
rect 5684 16524 5690 16576
rect 8932 16567 8990 16573
rect 8932 16533 8944 16567
rect 8978 16564 8990 16567
rect 9122 16564 9128 16576
rect 8978 16536 9128 16564
rect 8978 16533 8990 16536
rect 8932 16527 8990 16533
rect 9122 16524 9128 16536
rect 9180 16524 9186 16576
rect 2958 16456 2964 16508
rect 3016 16496 3022 16508
rect 3881 16499 3939 16505
rect 3881 16496 3893 16499
rect 3016 16468 3893 16496
rect 3016 16456 3022 16468
rect 3881 16465 3893 16468
rect 3927 16465 3939 16499
rect 3881 16459 3939 16465
rect 7285 16499 7343 16505
rect 7285 16465 7297 16499
rect 7331 16496 7343 16499
rect 7929 16499 7987 16505
rect 7929 16496 7941 16499
rect 7331 16468 7941 16496
rect 7331 16465 7343 16468
rect 7285 16459 7343 16465
rect 7929 16465 7941 16468
rect 7975 16465 7987 16499
rect 8665 16499 8723 16505
rect 8665 16496 8677 16499
rect 7929 16459 7987 16465
rect 8220 16468 8677 16496
rect 7374 16428 7380 16440
rect 7335 16400 7380 16428
rect 7374 16388 7380 16400
rect 7432 16388 7438 16440
rect 7469 16431 7527 16437
rect 7469 16397 7481 16431
rect 7515 16397 7527 16431
rect 7469 16391 7527 16397
rect 7006 16320 7012 16372
rect 7064 16360 7070 16372
rect 7484 16360 7512 16391
rect 7558 16388 7564 16440
rect 7616 16428 7622 16440
rect 8220 16428 8248 16468
rect 8665 16465 8677 16468
rect 8711 16496 8723 16499
rect 9968 16496 9996 16604
rect 10045 16601 10057 16635
rect 10091 16601 10103 16635
rect 10045 16595 10103 16601
rect 11701 16635 11759 16641
rect 11701 16601 11713 16635
rect 11747 16632 11759 16635
rect 11790 16632 11796 16644
rect 11747 16604 11796 16632
rect 11747 16601 11759 16604
rect 11701 16595 11759 16601
rect 10060 16564 10088 16595
rect 11790 16592 11796 16604
rect 11848 16632 11854 16644
rect 12342 16632 12348 16644
rect 11848 16604 12348 16632
rect 11848 16592 11854 16604
rect 12342 16592 12348 16604
rect 12400 16592 12406 16644
rect 12529 16635 12587 16641
rect 12529 16601 12541 16635
rect 12575 16632 12587 16635
rect 13170 16632 13176 16644
rect 12575 16604 13176 16632
rect 12575 16601 12587 16604
rect 12529 16595 12587 16601
rect 13170 16592 13176 16604
rect 13228 16592 13234 16644
rect 15562 16592 15568 16644
rect 15620 16632 15626 16644
rect 16482 16632 16488 16644
rect 15620 16604 16488 16632
rect 15620 16592 15626 16604
rect 16482 16592 16488 16604
rect 16540 16592 16546 16644
rect 16945 16635 17003 16641
rect 16945 16601 16957 16635
rect 16991 16632 17003 16635
rect 17126 16632 17132 16644
rect 16991 16604 17132 16632
rect 16991 16601 17003 16604
rect 16945 16595 17003 16601
rect 17126 16592 17132 16604
rect 17184 16592 17190 16644
rect 18046 16632 18052 16644
rect 18007 16604 18052 16632
rect 18046 16592 18052 16604
rect 18104 16592 18110 16644
rect 20162 16632 20168 16644
rect 20123 16604 20168 16632
rect 20162 16592 20168 16604
rect 20220 16592 20226 16644
rect 20717 16635 20775 16641
rect 20717 16601 20729 16635
rect 20763 16632 20775 16635
rect 21729 16635 21787 16641
rect 21729 16632 21741 16635
rect 20763 16604 21741 16632
rect 20763 16601 20775 16604
rect 20717 16595 20775 16601
rect 21729 16601 21741 16604
rect 21775 16601 21787 16635
rect 21729 16595 21787 16601
rect 10318 16564 10324 16576
rect 10060 16536 10324 16564
rect 10318 16524 10324 16536
rect 10376 16564 10382 16576
rect 10566 16567 10624 16573
rect 10566 16564 10578 16567
rect 10376 16536 10578 16564
rect 10376 16524 10382 16536
rect 10566 16533 10578 16536
rect 10612 16533 10624 16567
rect 19061 16567 19119 16573
rect 10566 16527 10624 16533
rect 10704 16536 18828 16564
rect 10704 16496 10732 16536
rect 8711 16468 9904 16496
rect 9968 16468 10732 16496
rect 8711 16465 8723 16468
rect 8665 16459 8723 16465
rect 7616 16400 8248 16428
rect 9876 16428 9904 16468
rect 12894 16456 12900 16508
rect 12952 16496 12958 16508
rect 13245 16499 13303 16505
rect 13245 16496 13257 16499
rect 12952 16468 13257 16496
rect 12952 16456 12958 16468
rect 13245 16465 13257 16468
rect 13291 16465 13303 16499
rect 13245 16459 13303 16465
rect 13722 16456 13728 16508
rect 13780 16496 13786 16508
rect 15013 16499 15071 16505
rect 13780 16468 14964 16496
rect 13780 16456 13786 16468
rect 10321 16431 10379 16437
rect 10321 16428 10333 16431
rect 9876 16400 10333 16428
rect 7616 16388 7622 16400
rect 10321 16397 10333 16400
rect 10367 16397 10379 16431
rect 10321 16391 10379 16397
rect 12434 16388 12440 16440
rect 12492 16428 12498 16440
rect 12989 16431 13047 16437
rect 12989 16428 13001 16431
rect 12492 16400 13001 16428
rect 12492 16388 12498 16400
rect 12989 16397 13001 16400
rect 13035 16397 13047 16431
rect 14936 16428 14964 16468
rect 15013 16465 15025 16499
rect 15059 16496 15071 16499
rect 15654 16496 15660 16508
rect 15059 16468 15660 16496
rect 15059 16465 15071 16468
rect 15013 16459 15071 16465
rect 15654 16456 15660 16468
rect 15712 16456 15718 16508
rect 15832 16499 15890 16505
rect 15832 16465 15844 16499
rect 15878 16496 15890 16499
rect 16390 16496 16396 16508
rect 15878 16468 16396 16496
rect 15878 16465 15890 16468
rect 15832 16459 15890 16465
rect 16390 16456 16396 16468
rect 16448 16456 16454 16508
rect 18800 16505 18828 16536
rect 19061 16533 19073 16567
rect 19107 16564 19119 16567
rect 19610 16564 19616 16576
rect 19107 16536 19616 16564
rect 19107 16533 19119 16536
rect 19061 16527 19119 16533
rect 19610 16524 19616 16536
rect 19668 16524 19674 16576
rect 18785 16499 18843 16505
rect 18785 16465 18797 16499
rect 18831 16465 18843 16499
rect 18785 16459 18843 16465
rect 18874 16456 18880 16508
rect 18932 16496 18938 16508
rect 19981 16499 20039 16505
rect 19981 16496 19993 16499
rect 18932 16468 19993 16496
rect 18932 16456 18938 16468
rect 19981 16465 19993 16468
rect 20027 16465 20039 16499
rect 19981 16459 20039 16465
rect 20438 16456 20444 16508
rect 20496 16496 20502 16508
rect 20533 16499 20591 16505
rect 20533 16496 20545 16499
rect 20496 16468 20545 16496
rect 20496 16456 20502 16468
rect 20533 16465 20545 16468
rect 20579 16465 20591 16499
rect 20533 16459 20591 16465
rect 15562 16428 15568 16440
rect 14936 16400 15568 16428
rect 12989 16391 13047 16397
rect 7064 16332 7512 16360
rect 7064 16320 7070 16332
rect 13004 16292 13032 16391
rect 15562 16388 15568 16400
rect 15620 16388 15626 16440
rect 13722 16292 13728 16304
rect 13004 16264 13728 16292
rect 13722 16252 13728 16264
rect 13780 16252 13786 16304
rect 14366 16292 14372 16304
rect 14327 16264 14372 16292
rect 14366 16252 14372 16264
rect 14424 16252 14430 16304
rect 1104 16202 21620 16224
rect 1104 16150 4414 16202
rect 4466 16150 4478 16202
rect 4530 16150 4542 16202
rect 4594 16150 4606 16202
rect 4658 16150 11278 16202
rect 11330 16150 11342 16202
rect 11394 16150 11406 16202
rect 11458 16150 11470 16202
rect 11522 16150 18142 16202
rect 18194 16150 18206 16202
rect 18258 16150 18270 16202
rect 18322 16150 18334 16202
rect 18386 16150 21620 16202
rect 1104 16128 21620 16150
rect 3142 16088 3148 16100
rect 3103 16060 3148 16088
rect 3142 16048 3148 16060
rect 3200 16048 3206 16100
rect 7006 16088 7012 16100
rect 6967 16060 7012 16088
rect 7006 16048 7012 16060
rect 7064 16048 7070 16100
rect 7285 16091 7343 16097
rect 7285 16057 7297 16091
rect 7331 16088 7343 16091
rect 7374 16088 7380 16100
rect 7331 16060 7380 16088
rect 7331 16057 7343 16060
rect 7285 16051 7343 16057
rect 7374 16048 7380 16060
rect 7432 16048 7438 16100
rect 12894 16088 12900 16100
rect 12855 16060 12900 16088
rect 12894 16048 12900 16060
rect 12952 16048 12958 16100
rect 15289 16091 15347 16097
rect 15289 16057 15301 16091
rect 15335 16088 15347 16091
rect 15335 16060 17632 16088
rect 15335 16057 15347 16060
rect 15289 16051 15347 16057
rect 14093 16023 14151 16029
rect 14093 15989 14105 16023
rect 14139 16020 14151 16023
rect 17604 16020 17632 16060
rect 19058 16048 19064 16100
rect 19116 16088 19122 16100
rect 20441 16091 20499 16097
rect 20441 16088 20453 16091
rect 19116 16060 20453 16088
rect 19116 16048 19122 16060
rect 20441 16057 20453 16060
rect 20487 16057 20499 16091
rect 20441 16051 20499 16057
rect 19334 16020 19340 16032
rect 14139 15992 15792 16020
rect 17604 15992 19340 16020
rect 14139 15989 14151 15992
rect 14093 15983 14151 15989
rect 4890 15912 4896 15964
rect 4948 15952 4954 15964
rect 5442 15952 5448 15964
rect 4948 15924 5448 15952
rect 4948 15912 4954 15924
rect 5442 15912 5448 15924
rect 5500 15952 5506 15964
rect 5629 15955 5687 15961
rect 5629 15952 5641 15955
rect 5500 15924 5641 15952
rect 5500 15912 5506 15924
rect 5629 15921 5641 15924
rect 5675 15921 5687 15955
rect 7742 15952 7748 15964
rect 7703 15924 7748 15952
rect 5629 15915 5687 15921
rect 7742 15912 7748 15924
rect 7800 15912 7806 15964
rect 7837 15955 7895 15961
rect 7837 15921 7849 15955
rect 7883 15921 7895 15955
rect 10134 15952 10140 15964
rect 10095 15924 10140 15952
rect 7837 15915 7895 15921
rect 1578 15844 1584 15896
rect 1636 15884 1642 15896
rect 1765 15887 1823 15893
rect 1765 15884 1777 15887
rect 1636 15856 1777 15884
rect 1636 15844 1642 15856
rect 1765 15853 1777 15856
rect 1811 15853 1823 15887
rect 1765 15847 1823 15853
rect 5896 15887 5954 15893
rect 5896 15853 5908 15887
rect 5942 15884 5954 15887
rect 6270 15884 6276 15896
rect 5942 15856 6276 15884
rect 5942 15853 5954 15856
rect 5896 15847 5954 15853
rect 6270 15844 6276 15856
rect 6328 15884 6334 15896
rect 7852 15884 7880 15915
rect 10134 15912 10140 15924
rect 10192 15912 10198 15964
rect 14366 15912 14372 15964
rect 14424 15952 14430 15964
rect 15764 15961 15792 15992
rect 19334 15980 19340 15992
rect 19392 15980 19398 16032
rect 19889 16023 19947 16029
rect 19889 15989 19901 16023
rect 19935 16020 19947 16023
rect 20070 16020 20076 16032
rect 19935 15992 20076 16020
rect 19935 15989 19947 15992
rect 19889 15983 19947 15989
rect 20070 15980 20076 15992
rect 20128 15980 20134 16032
rect 14645 15955 14703 15961
rect 14645 15952 14657 15955
rect 14424 15924 14657 15952
rect 14424 15912 14430 15924
rect 14645 15921 14657 15924
rect 14691 15921 14703 15955
rect 14645 15915 14703 15921
rect 15749 15955 15807 15961
rect 15749 15921 15761 15955
rect 15795 15921 15807 15955
rect 15749 15915 15807 15921
rect 15838 15912 15844 15964
rect 15896 15952 15902 15964
rect 15896 15924 15941 15952
rect 15896 15912 15902 15924
rect 6328 15856 7880 15884
rect 6328 15844 6334 15856
rect 11054 15844 11060 15896
rect 11112 15884 11118 15896
rect 11790 15893 11796 15896
rect 11517 15887 11575 15893
rect 11517 15884 11529 15887
rect 11112 15856 11529 15884
rect 11112 15844 11118 15856
rect 11517 15853 11529 15856
rect 11563 15853 11575 15887
rect 11784 15884 11796 15893
rect 11751 15856 11796 15884
rect 11517 15847 11575 15853
rect 11784 15847 11796 15856
rect 11790 15844 11796 15847
rect 11848 15844 11854 15896
rect 14458 15884 14464 15896
rect 14419 15856 14464 15884
rect 14458 15844 14464 15856
rect 14516 15844 14522 15896
rect 15654 15884 15660 15896
rect 15615 15856 15660 15884
rect 15654 15844 15660 15856
rect 15712 15844 15718 15896
rect 19150 15844 19156 15896
rect 19208 15884 19214 15896
rect 19705 15887 19763 15893
rect 19705 15884 19717 15887
rect 19208 15856 19717 15884
rect 19208 15844 19214 15856
rect 19705 15853 19717 15856
rect 19751 15853 19763 15887
rect 19705 15847 19763 15853
rect 19794 15844 19800 15896
rect 19852 15884 19858 15896
rect 20257 15887 20315 15893
rect 20257 15884 20269 15887
rect 19852 15856 20269 15884
rect 19852 15844 19858 15856
rect 20257 15853 20269 15856
rect 20303 15853 20315 15887
rect 20257 15847 20315 15853
rect 2032 15819 2090 15825
rect 2032 15785 2044 15819
rect 2078 15816 2090 15819
rect 2958 15816 2964 15828
rect 2078 15788 2964 15816
rect 2078 15785 2090 15788
rect 2032 15779 2090 15785
rect 2958 15776 2964 15788
rect 3016 15776 3022 15828
rect 9398 15776 9404 15828
rect 9456 15816 9462 15828
rect 14553 15819 14611 15825
rect 14553 15816 14565 15819
rect 9456 15788 14565 15816
rect 9456 15776 9462 15788
rect 14553 15785 14565 15788
rect 14599 15785 14611 15819
rect 14553 15779 14611 15785
rect 7650 15748 7656 15760
rect 7611 15720 7656 15748
rect 7650 15708 7656 15720
rect 7708 15708 7714 15760
rect 1104 15658 21620 15680
rect 1104 15606 7846 15658
rect 7898 15606 7910 15658
rect 7962 15606 7974 15658
rect 8026 15606 8038 15658
rect 8090 15606 14710 15658
rect 14762 15606 14774 15658
rect 14826 15606 14838 15658
rect 14890 15606 14902 15658
rect 14954 15606 21620 15658
rect 1104 15584 21620 15606
rect 3053 15547 3111 15553
rect 3053 15513 3065 15547
rect 3099 15513 3111 15547
rect 6270 15544 6276 15556
rect 6231 15516 6276 15544
rect 3053 15507 3111 15513
rect 3068 15476 3096 15507
rect 6270 15504 6276 15516
rect 6328 15504 6334 15556
rect 20717 15547 20775 15553
rect 20717 15513 20729 15547
rect 20763 15544 20775 15547
rect 20990 15544 20996 15556
rect 20763 15516 20996 15544
rect 20763 15513 20775 15516
rect 20717 15507 20775 15513
rect 20990 15504 20996 15516
rect 21048 15504 21054 15556
rect 19150 15476 19156 15488
rect 3068 15448 18920 15476
rect 19111 15448 19156 15476
rect 3418 15408 3424 15420
rect 3379 15380 3424 15408
rect 3418 15368 3424 15380
rect 3476 15368 3482 15420
rect 5160 15411 5218 15417
rect 5160 15377 5172 15411
rect 5206 15408 5218 15411
rect 6822 15408 6828 15420
rect 5206 15380 6828 15408
rect 5206 15377 5218 15380
rect 5160 15371 5218 15377
rect 6822 15368 6828 15380
rect 6880 15368 6886 15420
rect 7377 15411 7435 15417
rect 7377 15377 7389 15411
rect 7423 15408 7435 15411
rect 8202 15408 8208 15420
rect 7423 15380 8208 15408
rect 7423 15377 7435 15380
rect 7377 15371 7435 15377
rect 8202 15368 8208 15380
rect 8260 15368 8266 15420
rect 18892 15417 18920 15448
rect 19150 15436 19156 15448
rect 19208 15436 19214 15488
rect 18877 15411 18935 15417
rect 18877 15377 18889 15411
rect 18923 15377 18935 15411
rect 18877 15371 18935 15377
rect 19334 15368 19340 15420
rect 19392 15408 19398 15420
rect 19613 15411 19671 15417
rect 19613 15408 19625 15411
rect 19392 15380 19625 15408
rect 19392 15368 19398 15380
rect 19613 15377 19625 15380
rect 19659 15377 19671 15411
rect 19613 15371 19671 15377
rect 19889 15411 19947 15417
rect 19889 15377 19901 15411
rect 19935 15408 19947 15411
rect 20533 15411 20591 15417
rect 20533 15408 20545 15411
rect 19935 15380 20545 15408
rect 19935 15377 19947 15380
rect 19889 15371 19947 15377
rect 20533 15377 20545 15380
rect 20579 15377 20591 15411
rect 20533 15371 20591 15377
rect 3510 15340 3516 15352
rect 3471 15312 3516 15340
rect 3510 15300 3516 15312
rect 3568 15300 3574 15352
rect 3605 15343 3663 15349
rect 3605 15309 3617 15343
rect 3651 15309 3663 15343
rect 4890 15340 4896 15352
rect 4803 15312 4896 15340
rect 3605 15303 3663 15309
rect 2958 15232 2964 15284
rect 3016 15272 3022 15284
rect 3620 15272 3648 15303
rect 4890 15300 4896 15312
rect 4948 15300 4954 15352
rect 3016 15244 3648 15272
rect 3016 15232 3022 15244
rect 2222 15164 2228 15216
rect 2280 15204 2286 15216
rect 4908 15204 4936 15300
rect 7193 15207 7251 15213
rect 7193 15204 7205 15207
rect 2280 15176 7205 15204
rect 2280 15164 2286 15176
rect 7193 15173 7205 15176
rect 7239 15204 7251 15207
rect 7558 15204 7564 15216
rect 7239 15176 7564 15204
rect 7239 15173 7251 15176
rect 7193 15167 7251 15173
rect 7558 15164 7564 15176
rect 7616 15164 7622 15216
rect 10042 15164 10048 15216
rect 10100 15204 10106 15216
rect 18782 15204 18788 15216
rect 10100 15176 18788 15204
rect 10100 15164 10106 15176
rect 18782 15164 18788 15176
rect 18840 15164 18846 15216
rect 1104 15114 21620 15136
rect 1104 15062 4414 15114
rect 4466 15062 4478 15114
rect 4530 15062 4542 15114
rect 4594 15062 4606 15114
rect 4658 15062 11278 15114
rect 11330 15062 11342 15114
rect 11394 15062 11406 15114
rect 11458 15062 11470 15114
rect 11522 15062 18142 15114
rect 18194 15062 18206 15114
rect 18258 15062 18270 15114
rect 18322 15062 18334 15114
rect 18386 15062 21620 15114
rect 1104 15040 21620 15062
rect 2958 15000 2964 15012
rect 2919 14972 2964 15000
rect 2958 14960 2964 14972
rect 3016 14960 3022 15012
rect 3510 14960 3516 15012
rect 3568 15000 3574 15012
rect 4065 15003 4123 15009
rect 4065 15000 4077 15003
rect 3568 14972 4077 15000
rect 3568 14960 3574 14972
rect 4065 14969 4077 14972
rect 4111 14969 4123 15003
rect 4065 14963 4123 14969
rect 10962 14960 10968 15012
rect 11020 15000 11026 15012
rect 12434 15000 12440 15012
rect 11020 14972 12440 15000
rect 11020 14960 11026 14972
rect 12434 14960 12440 14972
rect 12492 15000 12498 15012
rect 13173 15003 13231 15009
rect 13173 15000 13185 15003
rect 12492 14972 13185 15000
rect 12492 14960 12498 14972
rect 13173 14969 13185 14972
rect 13219 14969 13231 15003
rect 13173 14963 13231 14969
rect 14921 15003 14979 15009
rect 14921 14969 14933 15003
rect 14967 15000 14979 15003
rect 15194 15000 15200 15012
rect 14967 14972 15200 15000
rect 14967 14969 14979 14972
rect 14921 14963 14979 14969
rect 7929 14935 7987 14941
rect 7929 14901 7941 14935
rect 7975 14932 7987 14935
rect 7975 14904 10180 14932
rect 7975 14901 7987 14904
rect 7929 14895 7987 14901
rect 3418 14864 3424 14876
rect 3379 14836 3424 14864
rect 3418 14824 3424 14836
rect 3476 14824 3482 14876
rect 3602 14824 3608 14876
rect 3660 14864 3666 14876
rect 4617 14867 4675 14873
rect 4617 14864 4629 14867
rect 3660 14836 4629 14864
rect 3660 14824 3666 14836
rect 4617 14833 4629 14836
rect 4663 14833 4675 14867
rect 8386 14864 8392 14876
rect 8347 14836 8392 14864
rect 4617 14827 4675 14833
rect 8386 14824 8392 14836
rect 8444 14824 8450 14876
rect 8570 14864 8576 14876
rect 8531 14836 8576 14864
rect 8570 14824 8576 14836
rect 8628 14824 8634 14876
rect 10152 14873 10180 14904
rect 10137 14867 10195 14873
rect 10137 14833 10149 14867
rect 10183 14833 10195 14867
rect 10137 14827 10195 14833
rect 10226 14824 10232 14876
rect 10284 14864 10290 14876
rect 12526 14864 12532 14876
rect 10284 14836 10329 14864
rect 12487 14836 12532 14864
rect 10284 14824 10290 14836
rect 12526 14824 12532 14836
rect 12584 14824 12590 14876
rect 13188 14864 13216 14963
rect 15194 14960 15200 14972
rect 15252 15000 15258 15012
rect 15838 15000 15844 15012
rect 15252 14972 15844 15000
rect 15252 14960 15258 14972
rect 15838 14960 15844 14972
rect 15896 14960 15902 15012
rect 20438 15000 20444 15012
rect 20399 14972 20444 15000
rect 20438 14960 20444 14972
rect 20496 14960 20502 15012
rect 19334 14932 19340 14944
rect 16040 14904 19340 14932
rect 13538 14864 13544 14876
rect 13188 14836 13544 14864
rect 13538 14824 13544 14836
rect 13596 14824 13602 14876
rect 1578 14796 1584 14808
rect 1491 14768 1584 14796
rect 1578 14756 1584 14768
rect 1636 14796 1642 14808
rect 2222 14796 2228 14808
rect 1636 14768 2228 14796
rect 1636 14756 1642 14768
rect 2222 14756 2228 14768
rect 2280 14756 2286 14808
rect 4246 14756 4252 14808
rect 4304 14796 4310 14808
rect 4525 14799 4583 14805
rect 4525 14796 4537 14799
rect 4304 14768 4537 14796
rect 4304 14756 4310 14768
rect 4525 14765 4537 14768
rect 4571 14765 4583 14799
rect 4525 14759 4583 14765
rect 9950 14756 9956 14808
rect 10008 14796 10014 14808
rect 12437 14799 12495 14805
rect 12437 14796 12449 14799
rect 10008 14768 12449 14796
rect 10008 14756 10014 14768
rect 12437 14765 12449 14768
rect 12483 14765 12495 14799
rect 12437 14759 12495 14765
rect 12710 14756 12716 14808
rect 12768 14796 12774 14808
rect 13357 14799 13415 14805
rect 13357 14796 13369 14799
rect 12768 14768 13369 14796
rect 12768 14756 12774 14768
rect 13357 14765 13369 14768
rect 13403 14765 13415 14799
rect 13357 14759 13415 14765
rect 13808 14799 13866 14805
rect 13808 14765 13820 14799
rect 13854 14796 13866 14799
rect 14366 14796 14372 14808
rect 13854 14768 14372 14796
rect 13854 14765 13866 14768
rect 13808 14759 13866 14765
rect 14366 14756 14372 14768
rect 14424 14756 14430 14808
rect 1848 14731 1906 14737
rect 1848 14697 1860 14731
rect 1894 14728 1906 14731
rect 3602 14728 3608 14740
rect 1894 14700 3608 14728
rect 1894 14697 1906 14700
rect 1848 14691 1906 14697
rect 3602 14688 3608 14700
rect 3660 14688 3666 14740
rect 10045 14731 10103 14737
rect 10045 14697 10057 14731
rect 10091 14728 10103 14731
rect 10689 14731 10747 14737
rect 10689 14728 10701 14731
rect 10091 14700 10701 14728
rect 10091 14697 10103 14700
rect 10045 14691 10103 14697
rect 10689 14697 10701 14700
rect 10735 14697 10747 14731
rect 16040 14728 16068 14904
rect 19334 14892 19340 14904
rect 19392 14892 19398 14944
rect 16850 14824 16856 14876
rect 16908 14864 16914 14876
rect 17129 14867 17187 14873
rect 17129 14864 17141 14867
rect 16908 14836 17141 14864
rect 16908 14824 16914 14836
rect 17129 14833 17141 14836
rect 17175 14833 17187 14867
rect 17129 14827 17187 14833
rect 19061 14867 19119 14873
rect 19061 14833 19073 14867
rect 19107 14864 19119 14867
rect 19794 14864 19800 14876
rect 19107 14836 19800 14864
rect 19107 14833 19119 14836
rect 19061 14827 19119 14833
rect 19794 14824 19800 14836
rect 19852 14824 19858 14876
rect 18785 14799 18843 14805
rect 18785 14796 18797 14799
rect 10689 14691 10747 14697
rect 11072 14700 16068 14728
rect 16592 14768 18797 14796
rect 4433 14663 4491 14669
rect 4433 14629 4445 14663
rect 4479 14660 4491 14663
rect 7650 14660 7656 14672
rect 4479 14632 7656 14660
rect 4479 14629 4491 14632
rect 4433 14623 4491 14629
rect 7650 14620 7656 14632
rect 7708 14620 7714 14672
rect 8297 14663 8355 14669
rect 8297 14629 8309 14663
rect 8343 14660 8355 14663
rect 8478 14660 8484 14672
rect 8343 14632 8484 14660
rect 8343 14629 8355 14632
rect 8297 14623 8355 14629
rect 8478 14620 8484 14632
rect 8536 14620 8542 14672
rect 9677 14663 9735 14669
rect 9677 14629 9689 14663
rect 9723 14660 9735 14663
rect 11072 14660 11100 14700
rect 11974 14660 11980 14672
rect 9723 14632 11100 14660
rect 11935 14632 11980 14660
rect 9723 14629 9735 14632
rect 9677 14623 9735 14629
rect 11974 14620 11980 14632
rect 12032 14620 12038 14672
rect 12066 14620 12072 14672
rect 12124 14660 12130 14672
rect 16592 14669 16620 14768
rect 18785 14765 18797 14768
rect 18831 14765 18843 14799
rect 18785 14759 18843 14765
rect 19518 14756 19524 14808
rect 19576 14796 19582 14808
rect 20257 14799 20315 14805
rect 20257 14796 20269 14799
rect 19576 14768 20269 14796
rect 19576 14756 19582 14768
rect 20257 14765 20269 14768
rect 20303 14765 20315 14799
rect 20257 14759 20315 14765
rect 12345 14663 12403 14669
rect 12345 14660 12357 14663
rect 12124 14632 12357 14660
rect 12124 14620 12130 14632
rect 12345 14629 12357 14632
rect 12391 14629 12403 14663
rect 12345 14623 12403 14629
rect 16577 14663 16635 14669
rect 16577 14629 16589 14663
rect 16623 14629 16635 14663
rect 16942 14660 16948 14672
rect 16903 14632 16948 14660
rect 16577 14623 16635 14629
rect 16942 14620 16948 14632
rect 17000 14620 17006 14672
rect 17034 14620 17040 14672
rect 17092 14660 17098 14672
rect 17092 14632 17137 14660
rect 17092 14620 17098 14632
rect 1104 14570 21620 14592
rect 1104 14518 7846 14570
rect 7898 14518 7910 14570
rect 7962 14518 7974 14570
rect 8026 14518 8038 14570
rect 8090 14518 14710 14570
rect 14762 14518 14774 14570
rect 14826 14518 14838 14570
rect 14890 14518 14902 14570
rect 14954 14518 21620 14570
rect 1104 14496 21620 14518
rect 3602 14456 3608 14468
rect 3563 14428 3608 14456
rect 3602 14416 3608 14428
rect 3660 14416 3666 14468
rect 6822 14416 6828 14468
rect 6880 14456 6886 14468
rect 9677 14459 9735 14465
rect 9677 14456 9689 14459
rect 6880 14428 9689 14456
rect 6880 14416 6886 14428
rect 9677 14425 9689 14428
rect 9723 14456 9735 14459
rect 10226 14456 10232 14468
rect 9723 14428 10232 14456
rect 9723 14425 9735 14428
rect 9677 14419 9735 14425
rect 10226 14416 10232 14428
rect 10284 14416 10290 14468
rect 11974 14416 11980 14468
rect 12032 14456 12038 14468
rect 12897 14459 12955 14465
rect 12897 14456 12909 14459
rect 12032 14428 12909 14456
rect 12032 14416 12038 14428
rect 12897 14425 12909 14428
rect 12943 14425 12955 14459
rect 12897 14419 12955 14425
rect 13817 14459 13875 14465
rect 13817 14425 13829 14459
rect 13863 14456 13875 14459
rect 20898 14456 20904 14468
rect 13863 14428 20024 14456
rect 20859 14428 20904 14456
rect 13863 14425 13875 14428
rect 13817 14419 13875 14425
rect 2492 14391 2550 14397
rect 2492 14357 2504 14391
rect 2538 14388 2550 14391
rect 2538 14360 6224 14388
rect 2538 14357 2550 14360
rect 2492 14351 2550 14357
rect 2222 14320 2228 14332
rect 2183 14292 2228 14320
rect 2222 14280 2228 14292
rect 2280 14280 2286 14332
rect 6086 14320 6092 14332
rect 6047 14292 6092 14320
rect 6086 14280 6092 14292
rect 6144 14280 6150 14332
rect 6196 14320 6224 14360
rect 7650 14348 7656 14400
rect 7708 14388 7714 14400
rect 14176 14391 14234 14397
rect 7708 14360 12020 14388
rect 7708 14348 7714 14360
rect 11992 14332 12020 14360
rect 14176 14357 14188 14391
rect 14222 14388 14234 14391
rect 15194 14388 15200 14400
rect 14222 14360 15200 14388
rect 14222 14357 14234 14360
rect 14176 14351 14234 14357
rect 15194 14348 15200 14360
rect 15252 14348 15258 14400
rect 16390 14348 16396 14400
rect 16448 14388 16454 14400
rect 18506 14388 18512 14400
rect 16448 14360 18512 14388
rect 16448 14348 16454 14360
rect 18506 14348 18512 14360
rect 18564 14348 18570 14400
rect 19518 14388 19524 14400
rect 19479 14360 19524 14388
rect 19518 14348 19524 14360
rect 19576 14348 19582 14400
rect 8570 14329 8576 14332
rect 8564 14320 8576 14329
rect 6196 14292 6316 14320
rect 8531 14292 8576 14320
rect 6288 14264 6316 14292
rect 8564 14283 8576 14292
rect 8570 14280 8576 14283
rect 8628 14280 8634 14332
rect 11974 14280 11980 14332
rect 12032 14280 12038 14332
rect 12618 14280 12624 14332
rect 12676 14320 12682 14332
rect 12805 14323 12863 14329
rect 12805 14320 12817 14323
rect 12676 14292 12817 14320
rect 12676 14280 12682 14292
rect 12805 14289 12817 14292
rect 12851 14289 12863 14323
rect 12805 14283 12863 14289
rect 13538 14280 13544 14332
rect 13596 14320 13602 14332
rect 13909 14323 13967 14329
rect 13909 14320 13921 14323
rect 13596 14292 13921 14320
rect 13596 14280 13602 14292
rect 13909 14289 13921 14292
rect 13955 14320 13967 14323
rect 15565 14323 15623 14329
rect 15565 14320 15577 14323
rect 13955 14292 15577 14320
rect 13955 14289 13967 14292
rect 13909 14283 13967 14289
rect 15565 14289 15577 14292
rect 15611 14289 15623 14323
rect 15832 14323 15890 14329
rect 15832 14320 15844 14323
rect 15565 14283 15623 14289
rect 15672 14292 15844 14320
rect 6178 14252 6184 14264
rect 6139 14224 6184 14252
rect 6178 14212 6184 14224
rect 6236 14212 6242 14264
rect 6270 14212 6276 14264
rect 6328 14252 6334 14264
rect 6328 14224 6421 14252
rect 6328 14212 6334 14224
rect 7742 14212 7748 14264
rect 7800 14252 7806 14264
rect 8297 14255 8355 14261
rect 8297 14252 8309 14255
rect 7800 14224 8309 14252
rect 7800 14212 7806 14224
rect 8297 14221 8309 14224
rect 8343 14221 8355 14255
rect 8297 14215 8355 14221
rect 12250 14212 12256 14264
rect 12308 14252 12314 14264
rect 12989 14255 13047 14261
rect 12989 14252 13001 14255
rect 12308 14224 13001 14252
rect 12308 14212 12314 14224
rect 12989 14221 13001 14224
rect 13035 14221 13047 14255
rect 15672 14252 15700 14292
rect 15832 14289 15844 14292
rect 15878 14320 15890 14323
rect 17126 14320 17132 14332
rect 15878 14292 17132 14320
rect 15878 14289 15890 14292
rect 15832 14283 15890 14289
rect 17126 14280 17132 14292
rect 17184 14280 17190 14332
rect 19996 14329 20024 14428
rect 20898 14416 20904 14428
rect 20956 14416 20962 14468
rect 19245 14323 19303 14329
rect 19245 14289 19257 14323
rect 19291 14289 19303 14323
rect 19245 14283 19303 14289
rect 19981 14323 20039 14329
rect 19981 14289 19993 14323
rect 20027 14289 20039 14323
rect 19981 14283 20039 14289
rect 20257 14323 20315 14329
rect 20257 14289 20269 14323
rect 20303 14320 20315 14323
rect 20717 14323 20775 14329
rect 20717 14320 20729 14323
rect 20303 14292 20729 14320
rect 20303 14289 20315 14292
rect 20257 14283 20315 14289
rect 20717 14289 20729 14292
rect 20763 14289 20775 14323
rect 20717 14283 20775 14289
rect 17402 14252 17408 14264
rect 12989 14215 13047 14221
rect 15304 14224 15700 14252
rect 17363 14224 17408 14252
rect 15304 14193 15332 14224
rect 17402 14212 17408 14224
rect 17460 14212 17466 14264
rect 12437 14187 12495 14193
rect 9600 14156 9812 14184
rect 5721 14119 5779 14125
rect 5721 14085 5733 14119
rect 5767 14116 5779 14119
rect 9600 14116 9628 14156
rect 5767 14088 9628 14116
rect 9784 14116 9812 14156
rect 12437 14153 12449 14187
rect 12483 14184 12495 14187
rect 13817 14187 13875 14193
rect 13817 14184 13829 14187
rect 12483 14156 13829 14184
rect 12483 14153 12495 14156
rect 12437 14147 12495 14153
rect 13817 14153 13829 14156
rect 13863 14153 13875 14187
rect 13817 14147 13875 14153
rect 15289 14187 15347 14193
rect 15289 14153 15301 14187
rect 15335 14153 15347 14187
rect 19260 14184 19288 14283
rect 15289 14147 15347 14153
rect 16500 14156 19288 14184
rect 16500 14116 16528 14156
rect 9784 14088 16528 14116
rect 5767 14085 5779 14088
rect 5721 14079 5779 14085
rect 16850 14076 16856 14128
rect 16908 14116 16914 14128
rect 16945 14119 17003 14125
rect 16945 14116 16957 14119
rect 16908 14088 16957 14116
rect 16908 14076 16914 14088
rect 16945 14085 16957 14088
rect 16991 14085 17003 14119
rect 16945 14079 17003 14085
rect 1104 14026 21620 14048
rect 1104 13974 4414 14026
rect 4466 13974 4478 14026
rect 4530 13974 4542 14026
rect 4594 13974 4606 14026
rect 4658 13974 11278 14026
rect 11330 13974 11342 14026
rect 11394 13974 11406 14026
rect 11458 13974 11470 14026
rect 11522 13974 18142 14026
rect 18194 13974 18206 14026
rect 18258 13974 18270 14026
rect 18322 13974 18334 14026
rect 18386 13974 21620 14026
rect 1104 13952 21620 13974
rect 6181 13915 6239 13921
rect 6181 13881 6193 13915
rect 6227 13912 6239 13915
rect 6270 13912 6276 13924
rect 6227 13884 6276 13912
rect 6227 13881 6239 13884
rect 6181 13875 6239 13881
rect 6270 13872 6276 13884
rect 6328 13872 6334 13924
rect 8202 13872 8208 13924
rect 8260 13872 8266 13924
rect 8570 13872 8576 13924
rect 8628 13912 8634 13924
rect 8665 13915 8723 13921
rect 8665 13912 8677 13915
rect 8628 13884 8677 13912
rect 8628 13872 8634 13884
rect 8665 13881 8677 13884
rect 8711 13881 8723 13915
rect 12618 13912 12624 13924
rect 8665 13875 8723 13881
rect 9048 13884 12480 13912
rect 12579 13884 12624 13912
rect 8220 13844 8248 13872
rect 8941 13847 8999 13853
rect 8941 13844 8953 13847
rect 8220 13816 8953 13844
rect 8941 13813 8953 13816
rect 8987 13813 8999 13847
rect 8941 13807 8999 13813
rect 6086 13736 6092 13788
rect 6144 13776 6150 13788
rect 6457 13779 6515 13785
rect 6457 13776 6469 13779
rect 6144 13748 6469 13776
rect 6144 13736 6150 13748
rect 6457 13745 6469 13748
rect 6503 13745 6515 13779
rect 6457 13739 6515 13745
rect 4430 13668 4436 13720
rect 4488 13708 4494 13720
rect 4801 13711 4859 13717
rect 4801 13708 4813 13711
rect 4488 13680 4813 13708
rect 4488 13668 4494 13680
rect 4801 13677 4813 13680
rect 4847 13708 4859 13711
rect 7285 13711 7343 13717
rect 7285 13708 7297 13711
rect 4847 13680 7297 13708
rect 4847 13677 4859 13680
rect 4801 13671 4859 13677
rect 7285 13677 7297 13680
rect 7331 13677 7343 13711
rect 7285 13671 7343 13677
rect 7552 13711 7610 13717
rect 7552 13677 7564 13711
rect 7598 13708 7610 13711
rect 9048 13708 9076 13884
rect 12250 13844 12256 13856
rect 11992 13816 12256 13844
rect 9582 13736 9588 13788
rect 9640 13776 9646 13788
rect 9640 13748 11100 13776
rect 9640 13736 9646 13748
rect 7598 13680 9076 13708
rect 9125 13711 9183 13717
rect 7598 13677 7610 13680
rect 7552 13671 7610 13677
rect 9125 13677 9137 13711
rect 9171 13708 9183 13711
rect 10778 13708 10784 13720
rect 9171 13680 10784 13708
rect 9171 13677 9183 13680
rect 9125 13671 9183 13677
rect 5068 13643 5126 13649
rect 5068 13609 5080 13643
rect 5114 13640 5126 13643
rect 5258 13640 5264 13652
rect 5114 13612 5264 13640
rect 5114 13609 5126 13612
rect 5068 13603 5126 13609
rect 5258 13600 5264 13612
rect 5316 13600 5322 13652
rect 7300 13640 7328 13671
rect 10778 13668 10784 13680
rect 10836 13668 10842 13720
rect 10962 13708 10968 13720
rect 10923 13680 10968 13708
rect 10962 13668 10968 13680
rect 11020 13668 11026 13720
rect 11072 13708 11100 13748
rect 11992 13708 12020 13816
rect 12250 13804 12256 13816
rect 12308 13844 12314 13856
rect 12345 13847 12403 13853
rect 12345 13844 12357 13847
rect 12308 13816 12357 13844
rect 12308 13804 12314 13816
rect 12345 13813 12357 13816
rect 12391 13813 12403 13847
rect 12452 13844 12480 13884
rect 12618 13872 12624 13884
rect 12676 13872 12682 13924
rect 16850 13912 16856 13924
rect 15764 13884 16856 13912
rect 15764 13844 15792 13884
rect 16850 13872 16856 13884
rect 16908 13872 16914 13924
rect 16942 13872 16948 13924
rect 17000 13912 17006 13924
rect 17497 13915 17555 13921
rect 17497 13912 17509 13915
rect 17000 13884 17509 13912
rect 17000 13872 17006 13884
rect 17497 13881 17509 13884
rect 17543 13881 17555 13915
rect 17497 13875 17555 13881
rect 18690 13872 18696 13924
rect 18748 13912 18754 13924
rect 18969 13915 19027 13921
rect 18969 13912 18981 13915
rect 18748 13884 18981 13912
rect 18748 13872 18754 13884
rect 18969 13881 18981 13884
rect 19015 13881 19027 13915
rect 18969 13875 19027 13881
rect 19702 13872 19708 13924
rect 19760 13912 19766 13924
rect 19889 13915 19947 13921
rect 19889 13912 19901 13915
rect 19760 13884 19901 13912
rect 19760 13872 19766 13884
rect 19889 13881 19901 13884
rect 19935 13881 19947 13915
rect 20438 13912 20444 13924
rect 20399 13884 20444 13912
rect 19889 13875 19947 13881
rect 20438 13872 20444 13884
rect 20496 13872 20502 13924
rect 12452 13816 15792 13844
rect 16485 13847 16543 13853
rect 12345 13807 12403 13813
rect 16485 13813 16497 13847
rect 16531 13844 16543 13847
rect 17034 13844 17040 13856
rect 16531 13816 17040 13844
rect 16531 13813 16543 13816
rect 16485 13807 16543 13813
rect 17034 13804 17040 13816
rect 17092 13804 17098 13856
rect 12434 13736 12440 13788
rect 12492 13776 12498 13788
rect 13173 13779 13231 13785
rect 13173 13776 13185 13779
rect 12492 13748 13185 13776
rect 12492 13736 12498 13748
rect 13173 13745 13185 13748
rect 13219 13745 13231 13779
rect 17126 13776 17132 13788
rect 17039 13748 17132 13776
rect 13173 13739 13231 13745
rect 17126 13736 17132 13748
rect 17184 13776 17190 13788
rect 18049 13779 18107 13785
rect 18049 13776 18061 13779
rect 17184 13748 18061 13776
rect 17184 13736 17190 13748
rect 18049 13745 18061 13748
rect 18095 13745 18107 13779
rect 18049 13739 18107 13745
rect 18506 13736 18512 13788
rect 18564 13776 18570 13788
rect 18564 13748 20300 13776
rect 18564 13736 18570 13748
rect 11072 13680 12020 13708
rect 13740 13680 17356 13708
rect 7742 13640 7748 13652
rect 7300 13612 7748 13640
rect 7742 13600 7748 13612
rect 7800 13600 7806 13652
rect 11146 13600 11152 13652
rect 11204 13649 11210 13652
rect 11204 13643 11268 13649
rect 11204 13609 11222 13643
rect 11256 13640 11268 13643
rect 12342 13640 12348 13652
rect 11256 13612 12348 13640
rect 11256 13609 11268 13612
rect 11204 13603 11268 13609
rect 11204 13600 11210 13603
rect 12342 13600 12348 13612
rect 12400 13600 12406 13652
rect 12989 13643 13047 13649
rect 12989 13609 13001 13643
rect 13035 13640 13047 13643
rect 13633 13643 13691 13649
rect 13633 13640 13645 13643
rect 13035 13612 13645 13640
rect 13035 13609 13047 13612
rect 12989 13603 13047 13609
rect 13633 13609 13645 13612
rect 13679 13609 13691 13643
rect 13633 13603 13691 13609
rect 106 13532 112 13584
rect 164 13572 170 13584
rect 7558 13572 7564 13584
rect 164 13544 7564 13572
rect 164 13532 170 13544
rect 7558 13532 7564 13544
rect 7616 13532 7622 13584
rect 13081 13575 13139 13581
rect 13081 13541 13093 13575
rect 13127 13572 13139 13575
rect 13740 13572 13768 13680
rect 17328 13640 17356 13680
rect 17402 13668 17408 13720
rect 17460 13708 17466 13720
rect 17865 13711 17923 13717
rect 17865 13708 17877 13711
rect 17460 13680 17877 13708
rect 17460 13668 17466 13680
rect 17865 13677 17877 13680
rect 17911 13677 17923 13711
rect 18782 13708 18788 13720
rect 18743 13680 18788 13708
rect 17865 13671 17923 13677
rect 18782 13668 18788 13680
rect 18840 13668 18846 13720
rect 19702 13708 19708 13720
rect 19663 13680 19708 13708
rect 19702 13668 19708 13680
rect 19760 13668 19766 13720
rect 20272 13717 20300 13748
rect 20257 13711 20315 13717
rect 20257 13677 20269 13711
rect 20303 13677 20315 13711
rect 20257 13671 20315 13677
rect 17957 13643 18015 13649
rect 17957 13640 17969 13643
rect 17328 13612 17969 13640
rect 17880 13584 17908 13612
rect 17957 13609 17969 13612
rect 18003 13609 18015 13643
rect 17957 13603 18015 13609
rect 16850 13572 16856 13584
rect 13127 13544 13768 13572
rect 16811 13544 16856 13572
rect 13127 13541 13139 13544
rect 13081 13535 13139 13541
rect 16850 13532 16856 13544
rect 16908 13532 16914 13584
rect 16942 13532 16948 13584
rect 17000 13572 17006 13584
rect 17000 13544 17045 13572
rect 17000 13532 17006 13544
rect 17862 13532 17868 13584
rect 17920 13532 17926 13584
rect 1104 13482 21620 13504
rect 1104 13430 7846 13482
rect 7898 13430 7910 13482
rect 7962 13430 7974 13482
rect 8026 13430 8038 13482
rect 8090 13430 14710 13482
rect 14762 13430 14774 13482
rect 14826 13430 14838 13482
rect 14890 13430 14902 13482
rect 14954 13430 21620 13482
rect 1104 13408 21620 13430
rect 5629 13371 5687 13377
rect 5629 13337 5641 13371
rect 5675 13368 5687 13371
rect 6178 13368 6184 13380
rect 5675 13340 6184 13368
rect 5675 13337 5687 13340
rect 5629 13331 5687 13337
rect 6178 13328 6184 13340
rect 6236 13328 6242 13380
rect 10778 13328 10784 13380
rect 10836 13368 10842 13380
rect 11333 13371 11391 13377
rect 11333 13368 11345 13371
rect 10836 13340 11345 13368
rect 10836 13328 10842 13340
rect 11333 13337 11345 13340
rect 11379 13337 11391 13371
rect 11333 13331 11391 13337
rect 20165 13371 20223 13377
rect 20165 13337 20177 13371
rect 20211 13368 20223 13371
rect 20530 13368 20536 13380
rect 20211 13340 20536 13368
rect 20211 13337 20223 13340
rect 20165 13331 20223 13337
rect 20530 13328 20536 13340
rect 20588 13328 20594 13380
rect 20714 13368 20720 13380
rect 20675 13340 20720 13368
rect 20714 13328 20720 13340
rect 20772 13328 20778 13380
rect 4148 13303 4206 13309
rect 4148 13269 4160 13303
rect 4194 13300 4206 13303
rect 9582 13300 9588 13312
rect 4194 13272 9588 13300
rect 4194 13269 4206 13272
rect 4148 13263 4206 13269
rect 9582 13260 9588 13272
rect 9640 13260 9646 13312
rect 10042 13300 10048 13312
rect 10005 13272 10048 13300
rect 10042 13260 10048 13272
rect 10100 13260 10106 13312
rect 18601 13303 18659 13309
rect 18601 13269 18613 13303
rect 18647 13300 18659 13303
rect 18782 13300 18788 13312
rect 18647 13272 18788 13300
rect 18647 13269 18659 13272
rect 18601 13263 18659 13269
rect 18782 13260 18788 13272
rect 18840 13260 18846 13312
rect 3881 13235 3939 13241
rect 3881 13201 3893 13235
rect 3927 13232 3939 13235
rect 4430 13232 4436 13244
rect 3927 13204 4436 13232
rect 3927 13201 3939 13204
rect 3881 13195 3939 13201
rect 4430 13192 4436 13204
rect 4488 13192 4494 13244
rect 5997 13235 6055 13241
rect 5997 13201 6009 13235
rect 6043 13232 6055 13235
rect 8570 13232 8576 13244
rect 6043 13204 8576 13232
rect 6043 13201 6055 13204
rect 5997 13195 6055 13201
rect 8570 13192 8576 13204
rect 8628 13232 8634 13244
rect 13722 13232 13728 13244
rect 8628 13204 13728 13232
rect 8628 13192 8634 13204
rect 13722 13192 13728 13204
rect 13780 13192 13786 13244
rect 18325 13235 18383 13241
rect 18325 13201 18337 13235
rect 18371 13232 18383 13235
rect 18690 13232 18696 13244
rect 18371 13204 18696 13232
rect 18371 13201 18383 13204
rect 18325 13195 18383 13201
rect 18690 13192 18696 13204
rect 18748 13192 18754 13244
rect 19242 13192 19248 13244
rect 19300 13232 19306 13244
rect 19429 13235 19487 13241
rect 19429 13232 19441 13235
rect 19300 13204 19441 13232
rect 19300 13192 19306 13204
rect 19429 13201 19441 13204
rect 19475 13201 19487 13235
rect 19429 13195 19487 13201
rect 19981 13235 20039 13241
rect 19981 13201 19993 13235
rect 20027 13232 20039 13235
rect 20162 13232 20168 13244
rect 20027 13204 20168 13232
rect 20027 13201 20039 13204
rect 19981 13195 20039 13201
rect 20162 13192 20168 13204
rect 20220 13192 20226 13244
rect 20533 13235 20591 13241
rect 20533 13201 20545 13235
rect 20579 13201 20591 13235
rect 20533 13195 20591 13201
rect 5902 13124 5908 13176
rect 5960 13164 5966 13176
rect 6089 13167 6147 13173
rect 6089 13164 6101 13167
rect 5960 13136 6101 13164
rect 5960 13124 5966 13136
rect 6089 13133 6101 13136
rect 6135 13133 6147 13167
rect 6089 13127 6147 13133
rect 6181 13167 6239 13173
rect 6181 13133 6193 13167
rect 6227 13133 6239 13167
rect 6181 13127 6239 13133
rect 5258 13096 5264 13108
rect 5171 13068 5264 13096
rect 5258 13056 5264 13068
rect 5316 13096 5322 13108
rect 6196 13096 6224 13127
rect 7558 13124 7564 13176
rect 7616 13164 7622 13176
rect 13354 13164 13360 13176
rect 7616 13136 13360 13164
rect 7616 13124 7622 13136
rect 13354 13124 13360 13136
rect 13412 13124 13418 13176
rect 15562 13124 15568 13176
rect 15620 13164 15626 13176
rect 20548 13164 20576 13195
rect 15620 13136 20576 13164
rect 15620 13124 15626 13136
rect 5316 13068 6224 13096
rect 19613 13099 19671 13105
rect 5316 13056 5322 13068
rect 19613 13065 19625 13099
rect 19659 13096 19671 13099
rect 20622 13096 20628 13108
rect 19659 13068 20628 13096
rect 19659 13065 19671 13068
rect 19613 13059 19671 13065
rect 20622 13056 20628 13068
rect 20680 13056 20686 13108
rect 1104 12938 21620 12960
rect 1104 12886 4414 12938
rect 4466 12886 4478 12938
rect 4530 12886 4542 12938
rect 4594 12886 4606 12938
rect 4658 12886 11278 12938
rect 11330 12886 11342 12938
rect 11394 12886 11406 12938
rect 11458 12886 11470 12938
rect 11522 12886 18142 12938
rect 18194 12886 18206 12938
rect 18258 12886 18270 12938
rect 18322 12886 18334 12938
rect 18386 12886 21620 12938
rect 1104 12864 21620 12886
rect 11146 12784 11152 12836
rect 11204 12824 11210 12836
rect 11241 12827 11299 12833
rect 11241 12824 11253 12827
rect 11204 12796 11253 12824
rect 11204 12784 11210 12796
rect 11241 12793 11253 12796
rect 11287 12793 11299 12827
rect 11241 12787 11299 12793
rect 12437 12827 12495 12833
rect 12437 12793 12449 12827
rect 12483 12824 12495 12827
rect 12710 12824 12716 12836
rect 12483 12796 12716 12824
rect 12483 12793 12495 12796
rect 12437 12787 12495 12793
rect 12710 12784 12716 12796
rect 12768 12784 12774 12836
rect 13722 12784 13728 12836
rect 13780 12824 13786 12836
rect 18874 12824 18880 12836
rect 13780 12796 18880 12824
rect 13780 12784 13786 12796
rect 18874 12784 18880 12796
rect 18932 12784 18938 12836
rect 20070 12824 20076 12836
rect 20031 12796 20076 12824
rect 20070 12784 20076 12796
rect 20128 12784 20134 12836
rect 7653 12759 7711 12765
rect 7653 12725 7665 12759
rect 7699 12725 7711 12759
rect 7653 12719 7711 12725
rect 12897 12759 12955 12765
rect 12897 12725 12909 12759
rect 12943 12756 12955 12759
rect 14550 12756 14556 12768
rect 12943 12728 14556 12756
rect 12943 12725 12955 12728
rect 12897 12719 12955 12725
rect 7668 12688 7696 12719
rect 14550 12716 14556 12728
rect 14608 12716 14614 12768
rect 19886 12716 19892 12768
rect 19944 12756 19950 12768
rect 20622 12756 20628 12768
rect 19944 12728 20628 12756
rect 19944 12716 19950 12728
rect 20622 12716 20628 12728
rect 20680 12716 20686 12768
rect 7742 12688 7748 12700
rect 7655 12660 7748 12688
rect 7742 12648 7748 12660
rect 7800 12688 7806 12700
rect 9861 12691 9919 12697
rect 9861 12688 9873 12691
rect 7800 12660 9873 12688
rect 7800 12648 7806 12660
rect 9861 12657 9873 12660
rect 9907 12657 9919 12691
rect 13354 12688 13360 12700
rect 13315 12660 13360 12688
rect 9861 12651 9919 12657
rect 13354 12648 13360 12660
rect 13412 12648 13418 12700
rect 13538 12688 13544 12700
rect 13499 12660 13544 12688
rect 13538 12648 13544 12660
rect 13596 12648 13602 12700
rect 14737 12691 14795 12697
rect 14737 12657 14749 12691
rect 14783 12688 14795 12691
rect 15010 12688 15016 12700
rect 14783 12660 15016 12688
rect 14783 12657 14795 12660
rect 14737 12651 14795 12657
rect 15010 12648 15016 12660
rect 15068 12648 15074 12700
rect 15562 12688 15568 12700
rect 15523 12660 15568 12688
rect 15562 12648 15568 12660
rect 15620 12648 15626 12700
rect 7837 12623 7895 12629
rect 7837 12589 7849 12623
rect 7883 12620 7895 12623
rect 8202 12620 8208 12632
rect 7883 12592 8208 12620
rect 7883 12589 7895 12592
rect 7837 12583 7895 12589
rect 8202 12580 8208 12592
rect 8260 12580 8266 12632
rect 11330 12620 11336 12632
rect 11291 12592 11336 12620
rect 11330 12580 11336 12592
rect 11388 12580 11394 12632
rect 12621 12623 12679 12629
rect 12621 12620 12633 12623
rect 11440 12592 12633 12620
rect 10134 12561 10140 12564
rect 10128 12515 10140 12561
rect 10192 12552 10198 12564
rect 10192 12524 10228 12552
rect 10134 12512 10140 12515
rect 10192 12512 10198 12524
rect 10778 12512 10784 12564
rect 10836 12552 10842 12564
rect 11440 12552 11468 12592
rect 12621 12589 12633 12592
rect 12667 12589 12679 12623
rect 12621 12583 12679 12589
rect 13096 12592 14688 12620
rect 10836 12524 11468 12552
rect 11609 12555 11667 12561
rect 10836 12512 10842 12524
rect 11609 12521 11621 12555
rect 11655 12552 11667 12555
rect 13096 12552 13124 12592
rect 13814 12552 13820 12564
rect 11655 12524 13124 12552
rect 13188 12524 13820 12552
rect 11655 12521 11667 12524
rect 11609 12515 11667 12521
rect 8294 12444 8300 12496
rect 8352 12484 8358 12496
rect 8662 12484 8668 12496
rect 8352 12456 8668 12484
rect 8352 12444 8358 12456
rect 8662 12444 8668 12456
rect 8720 12484 8726 12496
rect 13188 12484 13216 12524
rect 13814 12512 13820 12524
rect 13872 12552 13878 12564
rect 14553 12555 14611 12561
rect 14553 12552 14565 12555
rect 13872 12524 14565 12552
rect 13872 12512 13878 12524
rect 14553 12521 14565 12524
rect 14599 12521 14611 12555
rect 14660 12552 14688 12592
rect 15194 12580 15200 12632
rect 15252 12620 15258 12632
rect 15289 12623 15347 12629
rect 15289 12620 15301 12623
rect 15252 12592 15301 12620
rect 15252 12580 15258 12592
rect 15289 12589 15301 12592
rect 15335 12589 15347 12623
rect 15289 12583 15347 12589
rect 15838 12580 15844 12632
rect 15896 12620 15902 12632
rect 16577 12623 16635 12629
rect 16577 12620 16589 12623
rect 15896 12592 16589 12620
rect 15896 12580 15902 12592
rect 16577 12589 16589 12592
rect 16623 12589 16635 12623
rect 19058 12620 19064 12632
rect 19019 12592 19064 12620
rect 16577 12583 16635 12589
rect 19058 12580 19064 12592
rect 19116 12580 19122 12632
rect 19337 12623 19395 12629
rect 19337 12589 19349 12623
rect 19383 12620 19395 12623
rect 19889 12623 19947 12629
rect 19889 12620 19901 12623
rect 19383 12592 19901 12620
rect 19383 12589 19395 12592
rect 19337 12583 19395 12589
rect 19889 12589 19901 12592
rect 19935 12589 19947 12623
rect 19889 12583 19947 12589
rect 16390 12552 16396 12564
rect 14660 12524 16396 12552
rect 14553 12515 14611 12521
rect 16390 12512 16396 12524
rect 16448 12512 16454 12564
rect 16844 12555 16902 12561
rect 16844 12521 16856 12555
rect 16890 12552 16902 12555
rect 17494 12552 17500 12564
rect 16890 12524 17500 12552
rect 16890 12521 16902 12524
rect 16844 12515 16902 12521
rect 17494 12512 17500 12524
rect 17552 12512 17558 12564
rect 8720 12456 13216 12484
rect 13265 12487 13323 12493
rect 8720 12444 8726 12456
rect 13265 12453 13277 12487
rect 13311 12484 13323 12487
rect 13722 12484 13728 12496
rect 13311 12456 13728 12484
rect 13311 12453 13323 12456
rect 13265 12447 13323 12453
rect 13722 12444 13728 12456
rect 13780 12444 13786 12496
rect 14090 12484 14096 12496
rect 14051 12456 14096 12484
rect 14090 12444 14096 12456
rect 14148 12444 14154 12496
rect 14274 12444 14280 12496
rect 14332 12484 14338 12496
rect 14461 12487 14519 12493
rect 14461 12484 14473 12487
rect 14332 12456 14473 12484
rect 14332 12444 14338 12456
rect 14461 12453 14473 12456
rect 14507 12453 14519 12487
rect 17954 12484 17960 12496
rect 17915 12456 17960 12484
rect 14461 12447 14519 12453
rect 17954 12444 17960 12456
rect 18012 12444 18018 12496
rect 1104 12394 21620 12416
rect 1104 12342 7846 12394
rect 7898 12342 7910 12394
rect 7962 12342 7974 12394
rect 8026 12342 8038 12394
rect 8090 12342 14710 12394
rect 14762 12342 14774 12394
rect 14826 12342 14838 12394
rect 14890 12342 14902 12394
rect 14954 12342 21620 12394
rect 1104 12320 21620 12342
rect 8938 12240 8944 12292
rect 8996 12240 9002 12292
rect 10321 12283 10379 12289
rect 10321 12249 10333 12283
rect 10367 12280 10379 12283
rect 11330 12280 11336 12292
rect 10367 12252 11336 12280
rect 10367 12249 10379 12252
rect 10321 12243 10379 12249
rect 11330 12240 11336 12252
rect 11388 12240 11394 12292
rect 14550 12280 14556 12292
rect 14511 12252 14556 12280
rect 14550 12240 14556 12252
rect 14608 12240 14614 12292
rect 15010 12240 15016 12292
rect 15068 12280 15074 12292
rect 16669 12283 16727 12289
rect 16669 12280 16681 12283
rect 15068 12252 16681 12280
rect 15068 12240 15074 12252
rect 16669 12249 16681 12252
rect 16715 12249 16727 12283
rect 16669 12243 16727 12249
rect 17954 12240 17960 12292
rect 18012 12240 18018 12292
rect 18049 12283 18107 12289
rect 18049 12249 18061 12283
rect 18095 12280 18107 12283
rect 19058 12280 19064 12292
rect 18095 12252 19064 12280
rect 18095 12249 18107 12252
rect 18049 12243 18107 12249
rect 19058 12240 19064 12252
rect 19116 12240 19122 12292
rect 19978 12240 19984 12292
rect 20036 12280 20042 12292
rect 20073 12283 20131 12289
rect 20073 12280 20085 12283
rect 20036 12252 20085 12280
rect 20036 12240 20042 12252
rect 20073 12249 20085 12252
rect 20119 12249 20131 12283
rect 20073 12243 20131 12249
rect 20254 12240 20260 12292
rect 20312 12280 20318 12292
rect 20625 12283 20683 12289
rect 20625 12280 20637 12283
rect 20312 12252 20637 12280
rect 20312 12240 20318 12252
rect 20625 12249 20637 12252
rect 20671 12249 20683 12283
rect 20625 12243 20683 12249
rect 7276 12215 7334 12221
rect 7276 12181 7288 12215
rect 7322 12212 7334 12215
rect 7374 12212 7380 12224
rect 7322 12184 7380 12212
rect 7322 12181 7334 12184
rect 7276 12175 7334 12181
rect 7374 12172 7380 12184
rect 7432 12172 7438 12224
rect 7742 12172 7748 12224
rect 7800 12212 7806 12224
rect 8573 12215 8631 12221
rect 8573 12212 8585 12215
rect 7800 12184 8585 12212
rect 7800 12172 7806 12184
rect 8573 12181 8585 12184
rect 8619 12181 8631 12215
rect 8956 12212 8984 12240
rect 13998 12212 14004 12224
rect 8956 12184 14004 12212
rect 8573 12175 8631 12181
rect 13998 12172 14004 12184
rect 14056 12172 14062 12224
rect 14090 12172 14096 12224
rect 14148 12212 14154 12224
rect 14461 12215 14519 12221
rect 14461 12212 14473 12215
rect 14148 12184 14473 12212
rect 14148 12172 14154 12184
rect 14461 12181 14473 12184
rect 14507 12181 14519 12215
rect 14461 12175 14519 12181
rect 7009 12147 7067 12153
rect 7009 12113 7021 12147
rect 7055 12144 7067 12147
rect 7760 12144 7788 12172
rect 8921 12147 8979 12153
rect 8921 12144 8933 12147
rect 7055 12116 7788 12144
rect 8404 12116 8933 12144
rect 7055 12113 7067 12116
rect 7009 12107 7067 12113
rect 8404 11952 8432 12116
rect 8921 12113 8933 12116
rect 8967 12113 8979 12147
rect 8921 12107 8979 12113
rect 10318 12104 10324 12156
rect 10376 12144 10382 12156
rect 10689 12147 10747 12153
rect 10689 12144 10701 12147
rect 10376 12116 10701 12144
rect 10376 12104 10382 12116
rect 10689 12113 10701 12116
rect 10735 12113 10747 12147
rect 10689 12107 10747 12113
rect 12704 12147 12762 12153
rect 12704 12113 12716 12147
rect 12750 12144 12762 12147
rect 13538 12144 13544 12156
rect 12750 12116 13544 12144
rect 12750 12113 12762 12116
rect 12704 12107 12762 12113
rect 13538 12104 13544 12116
rect 13596 12144 13602 12156
rect 15028 12144 15056 12240
rect 15556 12215 15614 12221
rect 15556 12181 15568 12215
rect 15602 12212 15614 12215
rect 17972 12212 18000 12240
rect 15602 12184 18552 12212
rect 15602 12181 15614 12184
rect 15556 12175 15614 12181
rect 15838 12144 15844 12156
rect 13596 12116 15056 12144
rect 15304 12116 15844 12144
rect 13596 12104 13602 12116
rect 15304 12088 15332 12116
rect 15838 12104 15844 12116
rect 15896 12104 15902 12156
rect 17954 12104 17960 12156
rect 18012 12144 18018 12156
rect 18417 12147 18475 12153
rect 18417 12144 18429 12147
rect 18012 12116 18429 12144
rect 18012 12104 18018 12116
rect 18417 12113 18429 12116
rect 18463 12113 18475 12147
rect 18524 12144 18552 12184
rect 19886 12144 19892 12156
rect 18524 12116 18644 12144
rect 19847 12116 19892 12144
rect 18417 12107 18475 12113
rect 8573 12079 8631 12085
rect 8573 12045 8585 12079
rect 8619 12076 8631 12079
rect 8665 12079 8723 12085
rect 8665 12076 8677 12079
rect 8619 12048 8677 12076
rect 8619 12045 8631 12048
rect 8573 12039 8631 12045
rect 8665 12045 8677 12048
rect 8711 12045 8723 12079
rect 8665 12039 8723 12045
rect 9674 12036 9680 12088
rect 9732 12076 9738 12088
rect 10781 12079 10839 12085
rect 10781 12076 10793 12079
rect 9732 12048 10793 12076
rect 9732 12036 9738 12048
rect 10781 12045 10793 12048
rect 10827 12045 10839 12079
rect 10781 12039 10839 12045
rect 10873 12079 10931 12085
rect 10873 12045 10885 12079
rect 10919 12045 10931 12079
rect 10873 12039 10931 12045
rect 10045 12011 10103 12017
rect 10045 11977 10057 12011
rect 10091 12008 10103 12011
rect 10134 12008 10140 12020
rect 10091 11980 10140 12008
rect 10091 11977 10103 11980
rect 10045 11971 10103 11977
rect 10134 11968 10140 11980
rect 10192 12008 10198 12020
rect 10888 12008 10916 12039
rect 12434 12036 12440 12088
rect 12492 12076 12498 12088
rect 14645 12079 14703 12085
rect 14645 12076 14657 12079
rect 12492 12048 12537 12076
rect 14292 12048 14657 12076
rect 12492 12036 12498 12048
rect 14292 12020 14320 12048
rect 14645 12045 14657 12048
rect 14691 12045 14703 12079
rect 15286 12076 15292 12088
rect 15247 12048 15292 12076
rect 14645 12039 14703 12045
rect 15286 12036 15292 12048
rect 15344 12036 15350 12088
rect 16942 12036 16948 12088
rect 17000 12076 17006 12088
rect 18616 12085 18644 12116
rect 19886 12104 19892 12116
rect 19944 12104 19950 12156
rect 20438 12144 20444 12156
rect 20399 12116 20444 12144
rect 20438 12104 20444 12116
rect 20496 12104 20502 12156
rect 18509 12079 18567 12085
rect 18509 12076 18521 12079
rect 17000 12048 18521 12076
rect 17000 12036 17006 12048
rect 18509 12045 18521 12048
rect 18555 12045 18567 12079
rect 18509 12039 18567 12045
rect 18601 12079 18659 12085
rect 18601 12045 18613 12079
rect 18647 12045 18659 12079
rect 18601 12039 18659 12045
rect 10192 11980 10916 12008
rect 13817 12011 13875 12017
rect 10192 11968 10198 11980
rect 13817 11977 13829 12011
rect 13863 12008 13875 12011
rect 14274 12008 14280 12020
rect 13863 11980 14280 12008
rect 13863 11977 13875 11980
rect 13817 11971 13875 11977
rect 14274 11968 14280 11980
rect 14332 11968 14338 12020
rect 8386 11940 8392 11952
rect 8347 11912 8392 11940
rect 8386 11900 8392 11912
rect 8444 11900 8450 11952
rect 14090 11940 14096 11952
rect 14051 11912 14096 11940
rect 14090 11900 14096 11912
rect 14148 11900 14154 11952
rect 14182 11900 14188 11952
rect 14240 11940 14246 11952
rect 18966 11940 18972 11952
rect 14240 11912 18972 11940
rect 14240 11900 14246 11912
rect 18966 11900 18972 11912
rect 19024 11900 19030 11952
rect 1104 11850 21620 11872
rect 1104 11798 4414 11850
rect 4466 11798 4478 11850
rect 4530 11798 4542 11850
rect 4594 11798 4606 11850
rect 4658 11798 11278 11850
rect 11330 11798 11342 11850
rect 11394 11798 11406 11850
rect 11458 11798 11470 11850
rect 11522 11798 18142 11850
rect 18194 11798 18206 11850
rect 18258 11798 18270 11850
rect 18322 11798 18334 11850
rect 18386 11798 21620 11850
rect 1104 11776 21620 11798
rect 7929 11739 7987 11745
rect 7929 11705 7941 11739
rect 7975 11736 7987 11739
rect 9674 11736 9680 11748
rect 7975 11708 9680 11736
rect 7975 11705 7987 11708
rect 7929 11699 7987 11705
rect 9674 11696 9680 11708
rect 9732 11696 9738 11748
rect 10318 11736 10324 11748
rect 10279 11708 10324 11736
rect 10318 11696 10324 11708
rect 10376 11696 10382 11748
rect 12434 11696 12440 11748
rect 12492 11736 12498 11748
rect 12802 11736 12808 11748
rect 12492 11708 12808 11736
rect 12492 11696 12498 11708
rect 12802 11696 12808 11708
rect 12860 11736 12866 11748
rect 13357 11739 13415 11745
rect 13357 11736 13369 11739
rect 12860 11708 13369 11736
rect 12860 11696 12866 11708
rect 13357 11705 13369 11708
rect 13403 11705 13415 11739
rect 13357 11699 13415 11705
rect 13633 11739 13691 11745
rect 13633 11705 13645 11739
rect 13679 11736 13691 11739
rect 15194 11736 15200 11748
rect 13679 11708 15200 11736
rect 13679 11705 13691 11708
rect 13633 11699 13691 11705
rect 15194 11696 15200 11708
rect 15252 11696 15258 11748
rect 15746 11696 15752 11748
rect 15804 11736 15810 11748
rect 16390 11736 16396 11748
rect 15804 11708 16396 11736
rect 15804 11696 15810 11708
rect 16390 11696 16396 11708
rect 16448 11696 16454 11748
rect 17954 11696 17960 11748
rect 18012 11736 18018 11748
rect 18049 11739 18107 11745
rect 18049 11736 18061 11739
rect 18012 11708 18061 11736
rect 18012 11696 18018 11708
rect 18049 11705 18061 11708
rect 18095 11705 18107 11739
rect 18049 11699 18107 11705
rect 19150 11696 19156 11748
rect 19208 11736 19214 11748
rect 20441 11739 20499 11745
rect 20441 11736 20453 11739
rect 19208 11708 20453 11736
rect 19208 11696 19214 11708
rect 20441 11705 20453 11708
rect 20487 11705 20499 11739
rect 20441 11699 20499 11705
rect 6825 11671 6883 11677
rect 6825 11637 6837 11671
rect 6871 11637 6883 11671
rect 6825 11631 6883 11637
rect 6840 11600 6868 11631
rect 12158 11628 12164 11680
rect 12216 11668 12222 11680
rect 14550 11668 14556 11680
rect 12216 11640 14556 11668
rect 12216 11628 12222 11640
rect 14550 11628 14556 11640
rect 14608 11628 14614 11680
rect 7374 11600 7380 11612
rect 6840 11572 7144 11600
rect 7335 11572 7380 11600
rect 6730 11492 6736 11544
rect 6788 11532 6794 11544
rect 6788 11504 7052 11532
rect 6788 11492 6794 11504
rect 7024 11396 7052 11504
rect 7116 11464 7144 11572
rect 7374 11560 7380 11572
rect 7432 11600 7438 11612
rect 8294 11600 8300 11612
rect 7432 11572 8300 11600
rect 7432 11560 7438 11572
rect 8294 11560 8300 11572
rect 8352 11560 8358 11612
rect 8386 11560 8392 11612
rect 8444 11600 8450 11612
rect 8573 11603 8631 11609
rect 8573 11600 8585 11603
rect 8444 11572 8585 11600
rect 8444 11560 8450 11572
rect 8573 11569 8585 11572
rect 8619 11600 8631 11603
rect 10873 11603 10931 11609
rect 10873 11600 10885 11603
rect 8619 11572 10885 11600
rect 8619 11569 8631 11572
rect 8573 11563 8631 11569
rect 10873 11569 10885 11572
rect 10919 11569 10931 11603
rect 14182 11600 14188 11612
rect 14143 11572 14188 11600
rect 10873 11563 10931 11569
rect 14182 11560 14188 11572
rect 14240 11560 14246 11612
rect 17494 11560 17500 11612
rect 17552 11600 17558 11612
rect 18601 11603 18659 11609
rect 18601 11600 18613 11603
rect 17552 11572 18613 11600
rect 17552 11560 17558 11572
rect 18601 11569 18613 11572
rect 18647 11569 18659 11603
rect 18601 11563 18659 11569
rect 7193 11535 7251 11541
rect 7193 11501 7205 11535
rect 7239 11532 7251 11535
rect 8478 11532 8484 11544
rect 7239 11504 8484 11532
rect 7239 11501 7251 11504
rect 7193 11495 7251 11501
rect 8478 11492 8484 11504
rect 8536 11492 8542 11544
rect 10781 11535 10839 11541
rect 10781 11501 10793 11535
rect 10827 11532 10839 11535
rect 10827 11504 12664 11532
rect 10827 11501 10839 11504
rect 10781 11495 10839 11501
rect 8389 11467 8447 11473
rect 8389 11464 8401 11467
rect 7116 11436 8401 11464
rect 8389 11433 8401 11436
rect 8435 11433 8447 11467
rect 8389 11427 8447 11433
rect 10689 11467 10747 11473
rect 10689 11433 10701 11467
rect 10735 11464 10747 11467
rect 11333 11467 11391 11473
rect 11333 11464 11345 11467
rect 10735 11436 11345 11464
rect 10735 11433 10747 11436
rect 10689 11427 10747 11433
rect 11333 11433 11345 11436
rect 11379 11433 11391 11467
rect 12636 11464 12664 11504
rect 12710 11492 12716 11544
rect 12768 11532 12774 11544
rect 13541 11535 13599 11541
rect 13541 11532 13553 11535
rect 12768 11504 13553 11532
rect 12768 11492 12774 11504
rect 13541 11501 13553 11504
rect 13587 11501 13599 11535
rect 14090 11532 14096 11544
rect 14051 11504 14096 11532
rect 13541 11495 13599 11501
rect 14090 11492 14096 11504
rect 14148 11492 14154 11544
rect 20254 11532 20260 11544
rect 20215 11504 20260 11532
rect 20254 11492 20260 11504
rect 20312 11492 20318 11544
rect 14458 11464 14464 11476
rect 12636 11436 14464 11464
rect 11333 11427 11391 11433
rect 14458 11424 14464 11436
rect 14516 11424 14522 11476
rect 18417 11467 18475 11473
rect 18417 11433 18429 11467
rect 18463 11464 18475 11467
rect 19061 11467 19119 11473
rect 19061 11464 19073 11467
rect 18463 11436 19073 11464
rect 18463 11433 18475 11436
rect 18417 11427 18475 11433
rect 19061 11433 19073 11436
rect 19107 11433 19119 11467
rect 19061 11427 19119 11433
rect 7285 11399 7343 11405
rect 7285 11396 7297 11399
rect 7024 11368 7297 11396
rect 7285 11365 7297 11368
rect 7331 11365 7343 11399
rect 7285 11359 7343 11365
rect 8202 11356 8208 11408
rect 8260 11396 8266 11408
rect 8297 11399 8355 11405
rect 8297 11396 8309 11399
rect 8260 11368 8309 11396
rect 8260 11356 8266 11368
rect 8297 11365 8309 11368
rect 8343 11365 8355 11399
rect 8297 11359 8355 11365
rect 13722 11356 13728 11408
rect 13780 11396 13786 11408
rect 14001 11399 14059 11405
rect 14001 11396 14013 11399
rect 13780 11368 14013 11396
rect 13780 11356 13786 11368
rect 14001 11365 14013 11368
rect 14047 11365 14059 11399
rect 14001 11359 14059 11365
rect 18509 11399 18567 11405
rect 18509 11365 18521 11399
rect 18555 11396 18567 11399
rect 18782 11396 18788 11408
rect 18555 11368 18788 11396
rect 18555 11365 18567 11368
rect 18509 11359 18567 11365
rect 18782 11356 18788 11368
rect 18840 11356 18846 11408
rect 1104 11306 21620 11328
rect 1104 11254 7846 11306
rect 7898 11254 7910 11306
rect 7962 11254 7974 11306
rect 8026 11254 8038 11306
rect 8090 11254 14710 11306
rect 14762 11254 14774 11306
rect 14826 11254 14838 11306
rect 14890 11254 14902 11306
rect 14954 11254 21620 11306
rect 1104 11232 21620 11254
rect 8202 11192 8208 11204
rect 8163 11164 8208 11192
rect 8202 11152 8208 11164
rect 8260 11152 8266 11204
rect 8662 11192 8668 11204
rect 8623 11164 8668 11192
rect 8662 11152 8668 11164
rect 8720 11152 8726 11204
rect 13722 11192 13728 11204
rect 13683 11164 13728 11192
rect 13722 11152 13728 11164
rect 13780 11152 13786 11204
rect 14185 11195 14243 11201
rect 14185 11161 14197 11195
rect 14231 11192 14243 11195
rect 14458 11192 14464 11204
rect 14231 11164 14464 11192
rect 14231 11161 14243 11164
rect 14185 11155 14243 11161
rect 14458 11152 14464 11164
rect 14516 11152 14522 11204
rect 15933 11195 15991 11201
rect 15933 11161 15945 11195
rect 15979 11192 15991 11195
rect 17405 11195 17463 11201
rect 17405 11192 17417 11195
rect 15979 11164 17417 11192
rect 15979 11161 15991 11164
rect 15933 11155 15991 11161
rect 17405 11161 17417 11164
rect 17451 11161 17463 11195
rect 18782 11192 18788 11204
rect 18743 11164 18788 11192
rect 17405 11155 17463 11161
rect 18782 11152 18788 11164
rect 18840 11152 18846 11204
rect 19426 11152 19432 11204
rect 19484 11192 19490 11204
rect 20717 11195 20775 11201
rect 20717 11192 20729 11195
rect 19484 11164 20729 11192
rect 19484 11152 19490 11164
rect 20717 11161 20729 11164
rect 20763 11161 20775 11195
rect 20717 11155 20775 11161
rect 8573 11127 8631 11133
rect 8573 11093 8585 11127
rect 8619 11124 8631 11127
rect 8938 11124 8944 11136
rect 8619 11096 8944 11124
rect 8619 11093 8631 11096
rect 8573 11087 8631 11093
rect 8938 11084 8944 11096
rect 8996 11084 9002 11136
rect 11057 11127 11115 11133
rect 11057 11093 11069 11127
rect 11103 11124 11115 11127
rect 20254 11124 20260 11136
rect 11103 11096 20260 11124
rect 11103 11093 11115 11096
rect 11057 11087 11115 11093
rect 20254 11084 20260 11096
rect 20312 11084 20318 11136
rect 10778 11056 10784 11068
rect 10739 11028 10784 11056
rect 10778 11016 10784 11028
rect 10836 11016 10842 11068
rect 14093 11059 14151 11065
rect 14093 11025 14105 11059
rect 14139 11056 14151 11059
rect 14737 11059 14795 11065
rect 14737 11056 14749 11059
rect 14139 11028 14749 11056
rect 14139 11025 14151 11028
rect 14093 11019 14151 11025
rect 14737 11025 14749 11028
rect 14783 11025 14795 11059
rect 14737 11019 14795 11025
rect 15749 11059 15807 11065
rect 15749 11025 15761 11059
rect 15795 11056 15807 11059
rect 16301 11059 16359 11065
rect 16301 11056 16313 11059
rect 15795 11028 16313 11056
rect 15795 11025 15807 11028
rect 15749 11019 15807 11025
rect 16301 11025 16313 11028
rect 16347 11056 16359 11059
rect 17310 11056 17316 11068
rect 16347 11028 16712 11056
rect 17271 11028 17316 11056
rect 16347 11025 16359 11028
rect 16301 11019 16359 11025
rect 8294 10948 8300 11000
rect 8352 10988 8358 11000
rect 8757 10991 8815 10997
rect 8757 10988 8769 10991
rect 8352 10960 8769 10988
rect 8352 10948 8358 10960
rect 8757 10957 8769 10960
rect 8803 10957 8815 10991
rect 8757 10951 8815 10957
rect 14274 10948 14280 11000
rect 14332 10988 14338 11000
rect 14332 10960 14377 10988
rect 14332 10948 14338 10960
rect 14550 10948 14556 11000
rect 14608 10988 14614 11000
rect 16393 10991 16451 10997
rect 16393 10988 16405 10991
rect 14608 10960 16405 10988
rect 14608 10948 14614 10960
rect 16393 10957 16405 10960
rect 16439 10957 16451 10991
rect 16393 10951 16451 10957
rect 16577 10991 16635 10997
rect 16577 10957 16589 10991
rect 16623 10957 16635 10991
rect 16684 10988 16712 11028
rect 17310 11016 17316 11028
rect 17368 11016 17374 11068
rect 17862 11016 17868 11068
rect 17920 11056 17926 11068
rect 19153 11059 19211 11065
rect 19153 11056 19165 11059
rect 17920 11028 19165 11056
rect 17920 11016 17926 11028
rect 19153 11025 19165 11028
rect 19199 11025 19211 11059
rect 20530 11056 20536 11068
rect 20491 11028 20536 11056
rect 19153 11019 19211 11025
rect 20530 11016 20536 11028
rect 20588 11016 20594 11068
rect 16850 10988 16856 11000
rect 16684 10960 16856 10988
rect 16577 10951 16635 10957
rect 11974 10880 11980 10932
rect 12032 10920 12038 10932
rect 12250 10920 12256 10932
rect 12032 10892 12256 10920
rect 12032 10880 12038 10892
rect 12250 10880 12256 10892
rect 12308 10920 12314 10932
rect 15749 10923 15807 10929
rect 15749 10920 15761 10923
rect 12308 10892 15761 10920
rect 12308 10880 12314 10892
rect 15749 10889 15761 10892
rect 15795 10889 15807 10923
rect 15749 10883 15807 10889
rect 16482 10880 16488 10932
rect 16540 10920 16546 10932
rect 16592 10920 16620 10951
rect 16850 10948 16856 10960
rect 16908 10988 16914 11000
rect 17218 10988 17224 11000
rect 16908 10960 17224 10988
rect 16908 10948 16914 10960
rect 17218 10948 17224 10960
rect 17276 10948 17282 11000
rect 17494 10988 17500 11000
rect 17455 10960 17500 10988
rect 17494 10948 17500 10960
rect 17552 10948 17558 11000
rect 19245 10991 19303 10997
rect 19245 10988 19257 10991
rect 17604 10960 19257 10988
rect 16942 10920 16948 10932
rect 16540 10892 16620 10920
rect 16903 10892 16948 10920
rect 16540 10880 16546 10892
rect 16942 10880 16948 10892
rect 17000 10880 17006 10932
rect 12802 10812 12808 10864
rect 12860 10852 12866 10864
rect 15286 10852 15292 10864
rect 12860 10824 15292 10852
rect 12860 10812 12866 10824
rect 15286 10812 15292 10824
rect 15344 10812 15350 10864
rect 16390 10812 16396 10864
rect 16448 10852 16454 10864
rect 17604 10852 17632 10960
rect 19245 10957 19257 10960
rect 19291 10957 19303 10991
rect 19245 10951 19303 10957
rect 19337 10991 19395 10997
rect 19337 10957 19349 10991
rect 19383 10957 19395 10991
rect 19337 10951 19395 10957
rect 16448 10824 17632 10852
rect 16448 10812 16454 10824
rect 19242 10812 19248 10864
rect 19300 10852 19306 10864
rect 19352 10852 19380 10951
rect 19300 10824 19380 10852
rect 19300 10812 19306 10824
rect 1104 10762 21620 10784
rect 1104 10710 4414 10762
rect 4466 10710 4478 10762
rect 4530 10710 4542 10762
rect 4594 10710 4606 10762
rect 4658 10710 11278 10762
rect 11330 10710 11342 10762
rect 11394 10710 11406 10762
rect 11458 10710 11470 10762
rect 11522 10710 18142 10762
rect 18194 10710 18206 10762
rect 18258 10710 18270 10762
rect 18322 10710 18334 10762
rect 18386 10710 21620 10762
rect 1104 10688 21620 10710
rect 1670 10608 1676 10660
rect 1728 10648 1734 10660
rect 1728 10620 8156 10648
rect 1728 10608 1734 10620
rect 8128 10580 8156 10620
rect 8294 10608 8300 10660
rect 8352 10648 8358 10660
rect 8573 10651 8631 10657
rect 8573 10648 8585 10651
rect 8352 10620 8585 10648
rect 8352 10608 8358 10620
rect 8573 10617 8585 10620
rect 8619 10617 8631 10651
rect 8573 10611 8631 10617
rect 10229 10651 10287 10657
rect 10229 10617 10241 10651
rect 10275 10648 10287 10651
rect 10778 10648 10784 10660
rect 10275 10620 10784 10648
rect 10275 10617 10287 10620
rect 10229 10611 10287 10617
rect 10778 10608 10784 10620
rect 10836 10608 10842 10660
rect 14182 10648 14188 10660
rect 14143 10620 14188 10648
rect 14182 10608 14188 10620
rect 14240 10608 14246 10660
rect 16485 10651 16543 10657
rect 16485 10617 16497 10651
rect 16531 10648 16543 10651
rect 17310 10648 17316 10660
rect 16531 10620 17316 10648
rect 16531 10617 16543 10620
rect 16485 10611 16543 10617
rect 17310 10608 17316 10620
rect 17368 10608 17374 10660
rect 18690 10648 18696 10660
rect 18651 10620 18696 10648
rect 18690 10608 18696 10620
rect 18748 10608 18754 10660
rect 20346 10608 20352 10660
rect 20404 10648 20410 10660
rect 20441 10651 20499 10657
rect 20441 10648 20453 10651
rect 20404 10620 20453 10648
rect 20404 10608 20410 10620
rect 20441 10617 20453 10620
rect 20487 10617 20499 10651
rect 20441 10611 20499 10617
rect 8128 10552 10916 10580
rect 10781 10515 10839 10521
rect 10781 10512 10793 10515
rect 9508 10484 10793 10512
rect 7193 10447 7251 10453
rect 7193 10413 7205 10447
rect 7239 10444 7251 10447
rect 7742 10444 7748 10456
rect 7239 10416 7748 10444
rect 7239 10413 7251 10416
rect 7193 10407 7251 10413
rect 7742 10404 7748 10416
rect 7800 10404 7806 10456
rect 9508 10388 9536 10484
rect 10781 10481 10793 10484
rect 10827 10481 10839 10515
rect 10781 10475 10839 10481
rect 7460 10379 7518 10385
rect 7460 10345 7472 10379
rect 7506 10376 7518 10379
rect 9490 10376 9496 10388
rect 7506 10348 9496 10376
rect 7506 10345 7518 10348
rect 7460 10339 7518 10345
rect 9490 10336 9496 10348
rect 9548 10336 9554 10388
rect 10594 10376 10600 10388
rect 10555 10348 10600 10376
rect 10594 10336 10600 10348
rect 10652 10336 10658 10388
rect 10888 10376 10916 10552
rect 11885 10515 11943 10521
rect 11885 10481 11897 10515
rect 11931 10512 11943 10515
rect 12250 10512 12256 10524
rect 11931 10484 12256 10512
rect 11931 10481 11943 10484
rect 11885 10475 11943 10481
rect 12250 10472 12256 10484
rect 12308 10472 12314 10524
rect 12802 10512 12808 10524
rect 12763 10484 12808 10512
rect 12802 10472 12808 10484
rect 12860 10472 12866 10524
rect 16206 10472 16212 10524
rect 16264 10512 16270 10524
rect 16482 10512 16488 10524
rect 16264 10484 16488 10512
rect 16264 10472 16270 10484
rect 16482 10472 16488 10484
rect 16540 10512 16546 10524
rect 17129 10515 17187 10521
rect 17129 10512 17141 10515
rect 16540 10484 17141 10512
rect 16540 10472 16546 10484
rect 17129 10481 17141 10484
rect 17175 10512 17187 10515
rect 19150 10512 19156 10524
rect 17175 10484 19156 10512
rect 17175 10481 17187 10484
rect 17129 10475 17187 10481
rect 19150 10472 19156 10484
rect 19208 10472 19214 10524
rect 19245 10515 19303 10521
rect 19245 10481 19257 10515
rect 19291 10512 19303 10515
rect 19702 10512 19708 10524
rect 19291 10484 19708 10512
rect 19291 10481 19303 10484
rect 19245 10475 19303 10481
rect 19702 10472 19708 10484
rect 19760 10472 19766 10524
rect 11609 10447 11667 10453
rect 11609 10413 11621 10447
rect 11655 10444 11667 10447
rect 11974 10444 11980 10456
rect 11655 10416 11980 10444
rect 11655 10413 11667 10416
rect 11609 10407 11667 10413
rect 11974 10404 11980 10416
rect 12032 10404 12038 10456
rect 13072 10447 13130 10453
rect 13072 10413 13084 10447
rect 13118 10444 13130 10447
rect 14274 10444 14280 10456
rect 13118 10416 14280 10444
rect 13118 10413 13130 10416
rect 13072 10407 13130 10413
rect 14274 10404 14280 10416
rect 14332 10404 14338 10456
rect 20254 10444 20260 10456
rect 20215 10416 20260 10444
rect 20254 10404 20260 10416
rect 20312 10404 20318 10456
rect 11701 10379 11759 10385
rect 11701 10376 11713 10379
rect 10888 10348 11713 10376
rect 11701 10345 11713 10348
rect 11747 10345 11759 10379
rect 16850 10376 16856 10388
rect 16811 10348 16856 10376
rect 11701 10339 11759 10345
rect 16850 10336 16856 10348
rect 16908 10336 16914 10388
rect 18046 10336 18052 10388
rect 18104 10376 18110 10388
rect 19061 10379 19119 10385
rect 19061 10376 19073 10379
rect 18104 10348 19073 10376
rect 18104 10336 18110 10348
rect 19061 10345 19073 10348
rect 19107 10345 19119 10379
rect 19061 10339 19119 10345
rect 10686 10308 10692 10320
rect 10647 10280 10692 10308
rect 10686 10268 10692 10280
rect 10744 10268 10750 10320
rect 11054 10268 11060 10320
rect 11112 10308 11118 10320
rect 11241 10311 11299 10317
rect 11241 10308 11253 10311
rect 11112 10280 11253 10308
rect 11112 10268 11118 10280
rect 11241 10277 11253 10280
rect 11287 10277 11299 10311
rect 16942 10308 16948 10320
rect 16903 10280 16948 10308
rect 11241 10271 11299 10277
rect 16942 10268 16948 10280
rect 17000 10268 17006 10320
rect 19150 10308 19156 10320
rect 19111 10280 19156 10308
rect 19150 10268 19156 10280
rect 19208 10268 19214 10320
rect 1104 10218 21620 10240
rect 1104 10166 7846 10218
rect 7898 10166 7910 10218
rect 7962 10166 7974 10218
rect 8026 10166 8038 10218
rect 8090 10166 14710 10218
rect 14762 10166 14774 10218
rect 14826 10166 14838 10218
rect 14890 10166 14902 10218
rect 14954 10166 21620 10218
rect 1104 10144 21620 10166
rect 9490 10104 9496 10116
rect 9451 10076 9496 10104
rect 9490 10064 9496 10076
rect 9548 10064 9554 10116
rect 10597 10107 10655 10113
rect 10597 10073 10609 10107
rect 10643 10104 10655 10107
rect 10686 10104 10692 10116
rect 10643 10076 10692 10104
rect 10643 10073 10655 10076
rect 10597 10067 10655 10073
rect 10686 10064 10692 10076
rect 10744 10064 10750 10116
rect 11054 10104 11060 10116
rect 11015 10076 11060 10104
rect 11054 10064 11060 10076
rect 11112 10064 11118 10116
rect 17313 10107 17371 10113
rect 17313 10073 17325 10107
rect 17359 10104 17371 10107
rect 17494 10104 17500 10116
rect 17359 10076 17500 10104
rect 17359 10073 17371 10076
rect 17313 10067 17371 10073
rect 17494 10064 17500 10076
rect 17552 10064 17558 10116
rect 18046 10104 18052 10116
rect 18007 10076 18052 10104
rect 18046 10064 18052 10076
rect 18104 10064 18110 10116
rect 19242 10064 19248 10116
rect 19300 10104 19306 10116
rect 19889 10107 19947 10113
rect 19889 10104 19901 10107
rect 19300 10076 19901 10104
rect 19300 10064 19306 10076
rect 19889 10073 19901 10076
rect 19935 10073 19947 10107
rect 19889 10067 19947 10073
rect 20717 10107 20775 10113
rect 20717 10073 20729 10107
rect 20763 10073 20775 10107
rect 20717 10067 20775 10073
rect 16206 10045 16212 10048
rect 16200 10036 16212 10045
rect 16167 10008 16212 10036
rect 16200 9999 16212 10008
rect 16206 9996 16212 9999
rect 16264 9996 16270 10048
rect 17770 9996 17776 10048
rect 17828 10036 17834 10048
rect 20732 10036 20760 10067
rect 17828 10008 20760 10036
rect 17828 9996 17834 10008
rect 8380 9971 8438 9977
rect 8380 9937 8392 9971
rect 8426 9968 8438 9971
rect 9306 9968 9312 9980
rect 8426 9940 9312 9968
rect 8426 9937 8438 9940
rect 8380 9931 8438 9937
rect 9306 9928 9312 9940
rect 9364 9928 9370 9980
rect 10965 9971 11023 9977
rect 10965 9937 10977 9971
rect 11011 9968 11023 9971
rect 11054 9968 11060 9980
rect 11011 9940 11060 9968
rect 11011 9937 11023 9940
rect 10965 9931 11023 9937
rect 11054 9928 11060 9940
rect 11112 9928 11118 9980
rect 15286 9928 15292 9980
rect 15344 9968 15350 9980
rect 15933 9971 15991 9977
rect 15933 9968 15945 9971
rect 15344 9940 15945 9968
rect 15344 9928 15350 9940
rect 15933 9937 15945 9940
rect 15979 9968 15991 9971
rect 18506 9968 18512 9980
rect 15979 9940 18512 9968
rect 15979 9937 15991 9940
rect 15933 9931 15991 9937
rect 18506 9928 18512 9940
rect 18564 9928 18570 9980
rect 18776 9971 18834 9977
rect 18776 9937 18788 9971
rect 18822 9968 18834 9971
rect 19702 9968 19708 9980
rect 18822 9940 19708 9968
rect 18822 9937 18834 9940
rect 18776 9931 18834 9937
rect 19702 9928 19708 9940
rect 19760 9928 19766 9980
rect 20530 9968 20536 9980
rect 20491 9940 20536 9968
rect 20530 9928 20536 9940
rect 20588 9928 20594 9980
rect 7742 9860 7748 9912
rect 7800 9900 7806 9912
rect 8113 9903 8171 9909
rect 8113 9900 8125 9903
rect 7800 9872 8125 9900
rect 7800 9860 7806 9872
rect 8113 9869 8125 9872
rect 8159 9869 8171 9903
rect 9324 9900 9352 9928
rect 11146 9900 11152 9912
rect 9324 9872 11152 9900
rect 8113 9863 8171 9869
rect 11146 9860 11152 9872
rect 11204 9860 11210 9912
rect 12158 9724 12164 9776
rect 12216 9764 12222 9776
rect 16942 9764 16948 9776
rect 12216 9736 16948 9764
rect 12216 9724 12222 9736
rect 16942 9724 16948 9736
rect 17000 9724 17006 9776
rect 1104 9674 21620 9696
rect 1104 9622 4414 9674
rect 4466 9622 4478 9674
rect 4530 9622 4542 9674
rect 4594 9622 4606 9674
rect 4658 9622 11278 9674
rect 11330 9622 11342 9674
rect 11394 9622 11406 9674
rect 11458 9622 11470 9674
rect 11522 9622 18142 9674
rect 18194 9622 18206 9674
rect 18258 9622 18270 9674
rect 18322 9622 18334 9674
rect 18386 9622 21620 9674
rect 1104 9600 21620 9622
rect 9306 9560 9312 9572
rect 9267 9532 9312 9560
rect 9306 9520 9312 9532
rect 9364 9520 9370 9572
rect 10594 9520 10600 9572
rect 10652 9560 10658 9572
rect 10781 9563 10839 9569
rect 10781 9560 10793 9563
rect 10652 9532 10793 9560
rect 10652 9520 10658 9532
rect 10781 9529 10793 9532
rect 10827 9529 10839 9563
rect 10781 9523 10839 9529
rect 18693 9563 18751 9569
rect 18693 9529 18705 9563
rect 18739 9560 18751 9563
rect 19150 9560 19156 9572
rect 18739 9532 19156 9560
rect 18739 9529 18751 9532
rect 18693 9523 18751 9529
rect 19150 9520 19156 9532
rect 19208 9520 19214 9572
rect 12802 9452 12808 9504
rect 12860 9492 12866 9504
rect 12860 9464 13584 9492
rect 12860 9452 12866 9464
rect 11146 9384 11152 9436
rect 11204 9424 11210 9436
rect 11333 9427 11391 9433
rect 11333 9424 11345 9427
rect 11204 9396 11345 9424
rect 11204 9384 11210 9396
rect 11333 9393 11345 9396
rect 11379 9393 11391 9427
rect 11333 9387 11391 9393
rect 12250 9384 12256 9436
rect 12308 9424 12314 9436
rect 13556 9433 13584 9464
rect 15102 9452 15108 9504
rect 15160 9492 15166 9504
rect 15473 9495 15531 9501
rect 15473 9492 15485 9495
rect 15160 9464 15485 9492
rect 15160 9452 15166 9464
rect 15473 9461 15485 9464
rect 15519 9461 15531 9495
rect 15473 9455 15531 9461
rect 12897 9427 12955 9433
rect 12897 9424 12909 9427
rect 12308 9396 12909 9424
rect 12308 9384 12314 9396
rect 7742 9316 7748 9368
rect 7800 9356 7806 9368
rect 7929 9359 7987 9365
rect 7929 9356 7941 9359
rect 7800 9328 7941 9356
rect 7800 9316 7806 9328
rect 7929 9325 7941 9328
rect 7975 9325 7987 9359
rect 7929 9319 7987 9325
rect 8196 9291 8254 9297
rect 8196 9257 8208 9291
rect 8242 9288 8254 9291
rect 10962 9288 10968 9300
rect 8242 9260 10968 9288
rect 8242 9257 8254 9260
rect 8196 9251 8254 9257
rect 10962 9248 10968 9260
rect 11020 9248 11026 9300
rect 11149 9291 11207 9297
rect 11149 9257 11161 9291
rect 11195 9288 11207 9291
rect 11793 9291 11851 9297
rect 11793 9288 11805 9291
rect 11195 9260 11805 9288
rect 11195 9257 11207 9260
rect 11149 9251 11207 9257
rect 11793 9257 11805 9260
rect 11839 9257 11851 9291
rect 12728 9288 12756 9396
rect 12897 9393 12909 9396
rect 12943 9393 12955 9427
rect 12897 9387 12955 9393
rect 13541 9427 13599 9433
rect 13541 9393 13553 9427
rect 13587 9393 13599 9427
rect 13541 9387 13599 9393
rect 12805 9359 12863 9365
rect 12805 9325 12817 9359
rect 12851 9356 12863 9359
rect 13556 9356 13584 9387
rect 16850 9384 16856 9436
rect 16908 9424 16914 9436
rect 18690 9424 18696 9436
rect 16908 9396 18696 9424
rect 16908 9384 16914 9396
rect 18690 9384 18696 9396
rect 18748 9384 18754 9436
rect 19245 9427 19303 9433
rect 19245 9393 19257 9427
rect 19291 9424 19303 9427
rect 19426 9424 19432 9436
rect 19291 9396 19432 9424
rect 19291 9393 19303 9396
rect 19245 9387 19303 9393
rect 19426 9384 19432 9396
rect 19484 9384 19490 9436
rect 13630 9356 13636 9368
rect 12851 9328 13308 9356
rect 13556 9328 13636 9356
rect 12851 9325 12863 9328
rect 12805 9319 12863 9325
rect 13280 9288 13308 9328
rect 13630 9316 13636 9328
rect 13688 9316 13694 9368
rect 13808 9359 13866 9365
rect 13808 9325 13820 9359
rect 13854 9356 13866 9359
rect 14182 9356 14188 9368
rect 13854 9328 14188 9356
rect 13854 9325 13866 9328
rect 13808 9319 13866 9325
rect 14182 9316 14188 9328
rect 14240 9316 14246 9368
rect 15286 9356 15292 9368
rect 15247 9328 15292 9356
rect 15286 9316 15292 9328
rect 15344 9316 15350 9368
rect 19058 9356 19064 9368
rect 19019 9328 19064 9356
rect 19058 9316 19064 9328
rect 19116 9316 19122 9368
rect 16390 9288 16396 9300
rect 12728 9260 12848 9288
rect 13280 9260 16396 9288
rect 11793 9251 11851 9257
rect 11241 9223 11299 9229
rect 11241 9189 11253 9223
rect 11287 9220 11299 9223
rect 12345 9223 12403 9229
rect 12345 9220 12357 9223
rect 11287 9192 12357 9220
rect 11287 9189 11299 9192
rect 11241 9183 11299 9189
rect 12345 9189 12357 9192
rect 12391 9189 12403 9223
rect 12710 9220 12716 9232
rect 12671 9192 12716 9220
rect 12345 9183 12403 9189
rect 12710 9180 12716 9192
rect 12768 9180 12774 9232
rect 12820 9220 12848 9260
rect 16390 9248 16396 9260
rect 16448 9248 16454 9300
rect 14921 9223 14979 9229
rect 14921 9220 14933 9223
rect 12820 9192 14933 9220
rect 14921 9189 14933 9192
rect 14967 9189 14979 9223
rect 14921 9183 14979 9189
rect 17954 9180 17960 9232
rect 18012 9220 18018 9232
rect 19153 9223 19211 9229
rect 19153 9220 19165 9223
rect 18012 9192 19165 9220
rect 18012 9180 18018 9192
rect 19153 9189 19165 9192
rect 19199 9189 19211 9223
rect 19153 9183 19211 9189
rect 1104 9130 21620 9152
rect 1104 9078 7846 9130
rect 7898 9078 7910 9130
rect 7962 9078 7974 9130
rect 8026 9078 8038 9130
rect 8090 9078 14710 9130
rect 14762 9078 14774 9130
rect 14826 9078 14838 9130
rect 14890 9078 14902 9130
rect 14954 9078 21620 9130
rect 1104 9056 21620 9078
rect 11054 9016 11060 9028
rect 11015 8988 11060 9016
rect 11054 8976 11060 8988
rect 11112 8976 11118 9028
rect 11517 9019 11575 9025
rect 11517 8985 11529 9019
rect 11563 9016 11575 9019
rect 12158 9016 12164 9028
rect 11563 8988 12164 9016
rect 11563 8985 11575 8988
rect 11517 8979 11575 8985
rect 12158 8976 12164 8988
rect 12216 8976 12222 9028
rect 13446 9016 13452 9028
rect 13407 8988 13452 9016
rect 13446 8976 13452 8988
rect 13504 8976 13510 9028
rect 17862 9016 17868 9028
rect 13556 8988 17868 9016
rect 11425 8951 11483 8957
rect 11425 8917 11437 8951
rect 11471 8948 11483 8951
rect 11698 8948 11704 8960
rect 11471 8920 11704 8948
rect 11471 8917 11483 8920
rect 11425 8911 11483 8917
rect 11698 8908 11704 8920
rect 11756 8908 11762 8960
rect 12710 8908 12716 8960
rect 12768 8948 12774 8960
rect 13556 8948 13584 8988
rect 17862 8976 17868 8988
rect 17920 8976 17926 9028
rect 19702 9016 19708 9028
rect 19663 8988 19708 9016
rect 19702 8976 19708 8988
rect 19760 8976 19766 9028
rect 20717 9019 20775 9025
rect 20717 8985 20729 9019
rect 20763 9016 20775 9019
rect 21174 9016 21180 9028
rect 20763 8988 21180 9016
rect 20763 8985 20775 8988
rect 20717 8979 20775 8985
rect 21174 8976 21180 8988
rect 21232 8976 21238 9028
rect 12768 8920 13584 8948
rect 12768 8908 12774 8920
rect 15286 8908 15292 8960
rect 15344 8948 15350 8960
rect 15749 8951 15807 8957
rect 15749 8948 15761 8951
rect 15344 8920 15761 8948
rect 15344 8908 15350 8920
rect 15749 8917 15761 8920
rect 15795 8917 15807 8951
rect 15749 8911 15807 8917
rect 18506 8908 18512 8960
rect 18564 8908 18570 8960
rect 13265 8883 13323 8889
rect 13265 8849 13277 8883
rect 13311 8880 13323 8883
rect 13538 8880 13544 8892
rect 13311 8852 13544 8880
rect 13311 8849 13323 8852
rect 13265 8843 13323 8849
rect 13538 8840 13544 8852
rect 13596 8840 13602 8892
rect 15470 8880 15476 8892
rect 15431 8852 15476 8880
rect 15470 8840 15476 8852
rect 15528 8840 15534 8892
rect 18325 8883 18383 8889
rect 18325 8849 18337 8883
rect 18371 8880 18383 8883
rect 18524 8880 18552 8908
rect 18371 8852 18552 8880
rect 18592 8883 18650 8889
rect 18371 8849 18383 8852
rect 18325 8843 18383 8849
rect 18592 8849 18604 8883
rect 18638 8880 18650 8883
rect 19426 8880 19432 8892
rect 18638 8852 19432 8880
rect 18638 8849 18650 8852
rect 18592 8843 18650 8849
rect 19426 8840 19432 8852
rect 19484 8840 19490 8892
rect 19978 8880 19984 8892
rect 19939 8852 19984 8880
rect 19978 8840 19984 8852
rect 20036 8840 20042 8892
rect 20530 8880 20536 8892
rect 20491 8852 20536 8880
rect 20530 8840 20536 8852
rect 20588 8840 20594 8892
rect 10962 8772 10968 8824
rect 11020 8812 11026 8824
rect 11609 8815 11667 8821
rect 11609 8812 11621 8815
rect 11020 8784 11621 8812
rect 11020 8772 11026 8784
rect 11609 8781 11621 8784
rect 11655 8812 11667 8815
rect 12250 8812 12256 8824
rect 11655 8784 12256 8812
rect 11655 8781 11667 8784
rect 11609 8775 11667 8781
rect 12250 8772 12256 8784
rect 12308 8772 12314 8824
rect 11698 8704 11704 8756
rect 11756 8744 11762 8756
rect 16850 8744 16856 8756
rect 11756 8716 16856 8744
rect 11756 8704 11762 8716
rect 16850 8704 16856 8716
rect 16908 8704 16914 8756
rect 19610 8704 19616 8756
rect 19668 8744 19674 8756
rect 20165 8747 20223 8753
rect 20165 8744 20177 8747
rect 19668 8716 20177 8744
rect 19668 8704 19674 8716
rect 20165 8713 20177 8716
rect 20211 8713 20223 8747
rect 20165 8707 20223 8713
rect 1104 8586 21620 8608
rect 1104 8534 4414 8586
rect 4466 8534 4478 8586
rect 4530 8534 4542 8586
rect 4594 8534 4606 8586
rect 4658 8534 11278 8586
rect 11330 8534 11342 8586
rect 11394 8534 11406 8586
rect 11458 8534 11470 8586
rect 11522 8534 18142 8586
rect 18194 8534 18206 8586
rect 18258 8534 18270 8586
rect 18322 8534 18334 8586
rect 18386 8534 21620 8586
rect 1104 8512 21620 8534
rect 11425 8475 11483 8481
rect 11425 8441 11437 8475
rect 11471 8472 11483 8475
rect 11606 8472 11612 8484
rect 11471 8444 11612 8472
rect 11471 8441 11483 8444
rect 11425 8435 11483 8441
rect 11606 8432 11612 8444
rect 11664 8432 11670 8484
rect 20441 8475 20499 8481
rect 20441 8441 20453 8475
rect 20487 8472 20499 8475
rect 20622 8472 20628 8484
rect 20487 8444 20628 8472
rect 20487 8441 20499 8444
rect 20441 8435 20499 8441
rect 20622 8432 20628 8444
rect 20680 8432 20686 8484
rect 13538 8336 13544 8348
rect 13499 8308 13544 8336
rect 13538 8296 13544 8308
rect 13596 8296 13602 8348
rect 11238 8268 11244 8280
rect 11199 8240 11244 8268
rect 11238 8228 11244 8240
rect 11296 8228 11302 8280
rect 13354 8268 13360 8280
rect 13315 8240 13360 8268
rect 13354 8228 13360 8240
rect 13412 8228 13418 8280
rect 20254 8268 20260 8280
rect 20215 8240 20260 8268
rect 20254 8228 20260 8240
rect 20312 8228 20318 8280
rect 1104 8042 21620 8064
rect 1104 7990 7846 8042
rect 7898 7990 7910 8042
rect 7962 7990 7974 8042
rect 8026 7990 8038 8042
rect 8090 7990 14710 8042
rect 14762 7990 14774 8042
rect 14826 7990 14838 8042
rect 14890 7990 14902 8042
rect 14954 7990 21620 8042
rect 1104 7968 21620 7990
rect 13354 7888 13360 7940
rect 13412 7928 13418 7940
rect 13725 7931 13783 7937
rect 13725 7928 13737 7931
rect 13412 7900 13737 7928
rect 13412 7888 13418 7900
rect 13725 7897 13737 7900
rect 13771 7897 13783 7931
rect 13725 7891 13783 7897
rect 15470 7888 15476 7940
rect 15528 7928 15534 7940
rect 16393 7931 16451 7937
rect 16393 7928 16405 7931
rect 15528 7900 16405 7928
rect 15528 7888 15534 7900
rect 16393 7897 16405 7900
rect 16439 7897 16451 7931
rect 16393 7891 16451 7897
rect 18046 7888 18052 7940
rect 18104 7928 18110 7940
rect 18506 7928 18512 7940
rect 18104 7900 18512 7928
rect 18104 7888 18110 7900
rect 18506 7888 18512 7900
rect 18564 7888 18570 7940
rect 19426 7928 19432 7940
rect 19387 7900 19432 7928
rect 19426 7888 19432 7900
rect 19484 7888 19490 7940
rect 20717 7931 20775 7937
rect 20717 7897 20729 7931
rect 20763 7897 20775 7931
rect 20717 7891 20775 7897
rect 11149 7863 11207 7869
rect 11149 7829 11161 7863
rect 11195 7860 11207 7863
rect 11238 7860 11244 7872
rect 11195 7832 11244 7860
rect 11195 7829 11207 7832
rect 11149 7823 11207 7829
rect 11238 7820 11244 7832
rect 11296 7820 11302 7872
rect 16298 7820 16304 7872
rect 16356 7860 16362 7872
rect 20732 7860 20760 7891
rect 16356 7832 20760 7860
rect 16356 7820 16362 7832
rect 9490 7801 9496 7804
rect 9484 7792 9496 7801
rect 9451 7764 9496 7792
rect 9484 7755 9496 7764
rect 9490 7752 9496 7755
rect 9548 7752 9554 7804
rect 10226 7752 10232 7804
rect 10284 7792 10290 7804
rect 10873 7795 10931 7801
rect 10873 7792 10885 7795
rect 10284 7764 10885 7792
rect 10284 7752 10290 7764
rect 10873 7761 10885 7764
rect 10919 7761 10931 7795
rect 10873 7755 10931 7761
rect 14093 7795 14151 7801
rect 14093 7761 14105 7795
rect 14139 7792 14151 7795
rect 14550 7792 14556 7804
rect 14139 7764 14556 7792
rect 14139 7761 14151 7764
rect 14093 7755 14151 7761
rect 14550 7752 14556 7764
rect 14608 7752 14614 7804
rect 14993 7795 15051 7801
rect 14993 7792 15005 7795
rect 14660 7764 15005 7792
rect 7282 7684 7288 7736
rect 7340 7724 7346 7736
rect 7742 7724 7748 7736
rect 7340 7696 7748 7724
rect 7340 7684 7346 7696
rect 7742 7684 7748 7696
rect 7800 7724 7806 7736
rect 9217 7727 9275 7733
rect 9217 7724 9229 7727
rect 7800 7696 9229 7724
rect 7800 7684 7806 7696
rect 9217 7693 9229 7696
rect 9263 7693 9275 7727
rect 14182 7724 14188 7736
rect 14143 7696 14188 7724
rect 9217 7687 9275 7693
rect 14182 7684 14188 7696
rect 14240 7684 14246 7736
rect 14274 7684 14280 7736
rect 14332 7724 14338 7736
rect 14369 7727 14427 7733
rect 14369 7724 14381 7727
rect 14332 7696 14381 7724
rect 14332 7684 14338 7696
rect 14369 7693 14381 7696
rect 14415 7724 14427 7727
rect 14660 7724 14688 7764
rect 14993 7761 15005 7764
rect 15039 7761 15051 7795
rect 14993 7755 15051 7761
rect 16761 7795 16819 7801
rect 16761 7761 16773 7795
rect 16807 7792 16819 7795
rect 17405 7795 17463 7801
rect 17405 7792 17417 7795
rect 16807 7764 17417 7792
rect 16807 7761 16819 7764
rect 16761 7755 16819 7761
rect 17405 7761 17417 7764
rect 17451 7761 17463 7795
rect 18305 7795 18363 7801
rect 18305 7792 18317 7795
rect 17405 7755 17463 7761
rect 17512 7764 18317 7792
rect 14415 7696 14688 7724
rect 14737 7727 14795 7733
rect 14415 7693 14427 7696
rect 14369 7687 14427 7693
rect 14737 7693 14749 7727
rect 14783 7693 14795 7727
rect 16850 7724 16856 7736
rect 16811 7696 16856 7724
rect 14737 7687 14795 7693
rect 13630 7616 13636 7668
rect 13688 7656 13694 7668
rect 14752 7656 14780 7687
rect 16850 7684 16856 7696
rect 16908 7684 16914 7736
rect 17037 7727 17095 7733
rect 17037 7693 17049 7727
rect 17083 7724 17095 7727
rect 17512 7724 17540 7764
rect 18305 7761 18317 7764
rect 18351 7761 18363 7795
rect 19978 7792 19984 7804
rect 19939 7764 19984 7792
rect 18305 7755 18363 7761
rect 19978 7752 19984 7764
rect 20036 7752 20042 7804
rect 20530 7792 20536 7804
rect 20491 7764 20536 7792
rect 20530 7752 20536 7764
rect 20588 7752 20594 7804
rect 17586 7724 17592 7736
rect 17083 7696 17592 7724
rect 17083 7693 17095 7696
rect 17037 7687 17095 7693
rect 17586 7684 17592 7696
rect 17644 7684 17650 7736
rect 18046 7724 18052 7736
rect 18007 7696 18052 7724
rect 18046 7684 18052 7696
rect 18104 7684 18110 7736
rect 13688 7628 14780 7656
rect 16040 7628 17080 7656
rect 13688 7616 13694 7628
rect 10597 7591 10655 7597
rect 10597 7557 10609 7591
rect 10643 7588 10655 7591
rect 10778 7588 10784 7600
rect 10643 7560 10784 7588
rect 10643 7557 10655 7560
rect 10597 7551 10655 7557
rect 10778 7548 10784 7560
rect 10836 7548 10842 7600
rect 13906 7548 13912 7600
rect 13964 7588 13970 7600
rect 16040 7588 16068 7628
rect 13964 7560 16068 7588
rect 16117 7591 16175 7597
rect 13964 7548 13970 7560
rect 16117 7557 16129 7591
rect 16163 7588 16175 7591
rect 16574 7588 16580 7600
rect 16163 7560 16580 7588
rect 16163 7557 16175 7560
rect 16117 7551 16175 7557
rect 16574 7548 16580 7560
rect 16632 7548 16638 7600
rect 17052 7588 17080 7628
rect 20165 7591 20223 7597
rect 20165 7588 20177 7591
rect 17052 7560 20177 7588
rect 20165 7557 20177 7560
rect 20211 7557 20223 7591
rect 20165 7551 20223 7557
rect 1104 7498 21620 7520
rect 1104 7446 4414 7498
rect 4466 7446 4478 7498
rect 4530 7446 4542 7498
rect 4594 7446 4606 7498
rect 4658 7446 11278 7498
rect 11330 7446 11342 7498
rect 11394 7446 11406 7498
rect 11458 7446 11470 7498
rect 11522 7446 18142 7498
rect 18194 7446 18206 7498
rect 18258 7446 18270 7498
rect 18322 7446 18334 7498
rect 18386 7446 21620 7498
rect 1104 7424 21620 7446
rect 10226 7384 10232 7396
rect 10187 7356 10232 7384
rect 10226 7344 10232 7356
rect 10284 7344 10290 7396
rect 14274 7384 14280 7396
rect 14235 7356 14280 7384
rect 14274 7344 14280 7356
rect 14332 7344 14338 7396
rect 17586 7384 17592 7396
rect 17547 7356 17592 7384
rect 17586 7344 17592 7356
rect 17644 7344 17650 7396
rect 10778 7248 10784 7260
rect 10739 7220 10784 7248
rect 10778 7208 10784 7220
rect 10836 7208 10842 7260
rect 11149 7251 11207 7257
rect 11149 7217 11161 7251
rect 11195 7248 11207 7251
rect 11241 7251 11299 7257
rect 11241 7248 11253 7251
rect 11195 7220 11253 7248
rect 11195 7217 11207 7220
rect 11149 7211 11207 7217
rect 11241 7217 11253 7220
rect 11287 7217 11299 7251
rect 14550 7248 14556 7260
rect 14511 7220 14556 7248
rect 11241 7211 11299 7217
rect 14550 7208 14556 7220
rect 14608 7208 14614 7260
rect 9769 7115 9827 7121
rect 9769 7081 9781 7115
rect 9815 7112 9827 7115
rect 10597 7115 10655 7121
rect 10597 7112 10609 7115
rect 9815 7084 10609 7112
rect 9815 7081 9827 7084
rect 9769 7075 9827 7081
rect 10597 7081 10609 7084
rect 10643 7081 10655 7115
rect 10796 7112 10824 7208
rect 12897 7183 12955 7189
rect 12897 7180 12909 7183
rect 12544 7152 12909 7180
rect 11486 7115 11544 7121
rect 11486 7112 11498 7115
rect 10796 7084 11498 7112
rect 10597 7075 10655 7081
rect 11486 7081 11498 7084
rect 11532 7081 11544 7115
rect 12544 7112 12572 7152
rect 12897 7149 12909 7152
rect 12943 7180 12955 7183
rect 13630 7180 13636 7192
rect 12943 7152 13636 7180
rect 12943 7149 12955 7152
rect 12897 7143 12955 7149
rect 13630 7140 13636 7152
rect 13688 7180 13694 7192
rect 16209 7183 16267 7189
rect 16209 7180 16221 7183
rect 13688 7152 16221 7180
rect 13688 7140 13694 7152
rect 16209 7149 16221 7152
rect 16255 7149 16267 7183
rect 16209 7143 16267 7149
rect 13164 7115 13222 7121
rect 13164 7112 13176 7115
rect 11486 7075 11544 7081
rect 12360 7084 12572 7112
rect 12636 7084 13176 7112
rect 10686 7044 10692 7056
rect 10647 7016 10692 7044
rect 10686 7004 10692 7016
rect 10744 7004 10750 7056
rect 11149 7047 11207 7053
rect 11149 7013 11161 7047
rect 11195 7044 11207 7047
rect 12360 7044 12388 7084
rect 12636 7053 12664 7084
rect 13164 7081 13176 7084
rect 13210 7112 13222 7115
rect 14550 7112 14556 7124
rect 13210 7084 14556 7112
rect 13210 7081 13222 7084
rect 13164 7075 13222 7081
rect 14550 7072 14556 7084
rect 14608 7072 14614 7124
rect 16476 7115 16534 7121
rect 16476 7081 16488 7115
rect 16522 7112 16534 7115
rect 16574 7112 16580 7124
rect 16522 7084 16580 7112
rect 16522 7081 16534 7084
rect 16476 7075 16534 7081
rect 16574 7072 16580 7084
rect 16632 7072 16638 7124
rect 11195 7016 12388 7044
rect 12621 7047 12679 7053
rect 11195 7013 11207 7016
rect 11149 7007 11207 7013
rect 12621 7013 12633 7047
rect 12667 7013 12679 7047
rect 12621 7007 12679 7013
rect 1104 6954 21620 6976
rect 1104 6902 7846 6954
rect 7898 6902 7910 6954
rect 7962 6902 7974 6954
rect 8026 6902 8038 6954
rect 8090 6902 14710 6954
rect 14762 6902 14774 6954
rect 14826 6902 14838 6954
rect 14890 6902 14902 6954
rect 14954 6902 21620 6954
rect 1104 6880 21620 6902
rect 10597 6843 10655 6849
rect 10597 6809 10609 6843
rect 10643 6840 10655 6843
rect 10686 6840 10692 6852
rect 10643 6812 10692 6840
rect 10643 6809 10655 6812
rect 10597 6803 10655 6809
rect 10686 6800 10692 6812
rect 10744 6800 10750 6852
rect 14093 6843 14151 6849
rect 14093 6809 14105 6843
rect 14139 6840 14151 6843
rect 14182 6840 14188 6852
rect 14139 6812 14188 6840
rect 14139 6809 14151 6812
rect 14093 6803 14151 6809
rect 14182 6800 14188 6812
rect 14240 6800 14246 6852
rect 16482 6840 16488 6852
rect 14384 6812 16488 6840
rect 10965 6775 11023 6781
rect 10965 6741 10977 6775
rect 11011 6772 11023 6775
rect 14384 6772 14412 6812
rect 16482 6800 16488 6812
rect 16540 6800 16546 6852
rect 16850 6840 16856 6852
rect 16811 6812 16856 6840
rect 16850 6800 16856 6812
rect 16908 6800 16914 6852
rect 17313 6843 17371 6849
rect 17313 6809 17325 6843
rect 17359 6840 17371 6843
rect 17954 6840 17960 6852
rect 17359 6812 17960 6840
rect 17359 6809 17371 6812
rect 17313 6803 17371 6809
rect 17954 6800 17960 6812
rect 18012 6800 18018 6852
rect 11011 6744 14412 6772
rect 14461 6775 14519 6781
rect 11011 6741 11023 6744
rect 10965 6735 11023 6741
rect 14461 6741 14473 6775
rect 14507 6772 14519 6775
rect 17221 6775 17279 6781
rect 14507 6744 16528 6772
rect 14507 6741 14519 6744
rect 14461 6735 14519 6741
rect 4062 6664 4068 6716
rect 4120 6704 4126 6716
rect 7541 6707 7599 6713
rect 7541 6704 7553 6707
rect 4120 6676 7553 6704
rect 4120 6664 4126 6676
rect 7541 6673 7553 6676
rect 7587 6673 7599 6707
rect 9490 6704 9496 6716
rect 7541 6667 7599 6673
rect 8680 6676 9496 6704
rect 7282 6636 7288 6648
rect 7243 6608 7288 6636
rect 7282 6596 7288 6608
rect 7340 6596 7346 6648
rect 8680 6577 8708 6676
rect 9490 6664 9496 6676
rect 9548 6704 9554 6716
rect 9548 6676 11192 6704
rect 9548 6664 9554 6676
rect 10410 6596 10416 6648
rect 10468 6636 10474 6648
rect 11164 6645 11192 6676
rect 11057 6639 11115 6645
rect 11057 6636 11069 6639
rect 10468 6608 11069 6636
rect 10468 6596 10474 6608
rect 11057 6605 11069 6608
rect 11103 6605 11115 6639
rect 11057 6599 11115 6605
rect 11149 6639 11207 6645
rect 11149 6605 11161 6639
rect 11195 6605 11207 6639
rect 11149 6599 11207 6605
rect 14553 6639 14611 6645
rect 14553 6605 14565 6639
rect 14599 6605 14611 6639
rect 14553 6599 14611 6605
rect 8665 6571 8723 6577
rect 8665 6537 8677 6571
rect 8711 6537 8723 6571
rect 8665 6531 8723 6537
rect 11072 6500 11100 6599
rect 14568 6568 14596 6599
rect 14642 6596 14648 6648
rect 14700 6636 14706 6648
rect 14700 6608 14745 6636
rect 14700 6596 14706 6608
rect 12360 6540 14596 6568
rect 16500 6568 16528 6744
rect 17221 6741 17233 6775
rect 17267 6772 17279 6775
rect 18506 6772 18512 6784
rect 17267 6744 18512 6772
rect 17267 6741 17279 6744
rect 17221 6735 17279 6741
rect 18506 6732 18512 6744
rect 18564 6732 18570 6784
rect 16574 6664 16580 6716
rect 16632 6704 16638 6716
rect 20530 6704 20536 6716
rect 16632 6676 17448 6704
rect 20491 6676 20536 6704
rect 16632 6664 16638 6676
rect 17420 6645 17448 6676
rect 20530 6664 20536 6676
rect 20588 6664 20594 6716
rect 17405 6639 17463 6645
rect 17405 6605 17417 6639
rect 17451 6605 17463 6639
rect 17405 6599 17463 6605
rect 18598 6568 18604 6580
rect 16500 6540 18604 6568
rect 12360 6500 12388 6540
rect 11072 6472 12388 6500
rect 14568 6500 14596 6540
rect 18598 6528 18604 6540
rect 18656 6528 18662 6580
rect 17954 6500 17960 6512
rect 14568 6472 17960 6500
rect 17954 6460 17960 6472
rect 18012 6460 18018 6512
rect 20714 6500 20720 6512
rect 20675 6472 20720 6500
rect 20714 6460 20720 6472
rect 20772 6460 20778 6512
rect 1104 6410 21620 6432
rect 1104 6358 4414 6410
rect 4466 6358 4478 6410
rect 4530 6358 4542 6410
rect 4594 6358 4606 6410
rect 4658 6358 11278 6410
rect 11330 6358 11342 6410
rect 11394 6358 11406 6410
rect 11458 6358 11470 6410
rect 11522 6358 18142 6410
rect 18194 6358 18206 6410
rect 18258 6358 18270 6410
rect 18322 6358 18334 6410
rect 18386 6358 21620 6410
rect 1104 6336 21620 6358
rect 13722 6256 13728 6308
rect 13780 6296 13786 6308
rect 20714 6296 20720 6308
rect 13780 6268 20720 6296
rect 13780 6256 13786 6268
rect 20714 6256 20720 6268
rect 20772 6256 20778 6308
rect 1104 5866 21620 5888
rect 1104 5814 7846 5866
rect 7898 5814 7910 5866
rect 7962 5814 7974 5866
rect 8026 5814 8038 5866
rect 8090 5814 14710 5866
rect 14762 5814 14774 5866
rect 14826 5814 14838 5866
rect 14890 5814 14902 5866
rect 14954 5814 21620 5866
rect 1104 5792 21620 5814
rect 13262 5712 13268 5764
rect 13320 5752 13326 5764
rect 20717 5755 20775 5761
rect 20717 5752 20729 5755
rect 13320 5724 20729 5752
rect 13320 5712 13326 5724
rect 20717 5721 20729 5724
rect 20763 5721 20775 5755
rect 20717 5715 20775 5721
rect 20530 5616 20536 5628
rect 20491 5588 20536 5616
rect 20530 5576 20536 5588
rect 20588 5576 20594 5628
rect 1104 5322 21620 5344
rect 1104 5270 4414 5322
rect 4466 5270 4478 5322
rect 4530 5270 4542 5322
rect 4594 5270 4606 5322
rect 4658 5270 11278 5322
rect 11330 5270 11342 5322
rect 11394 5270 11406 5322
rect 11458 5270 11470 5322
rect 11522 5270 18142 5322
rect 18194 5270 18206 5322
rect 18258 5270 18270 5322
rect 18322 5270 18334 5322
rect 18386 5270 21620 5322
rect 1104 5248 21620 5270
rect 16482 5168 16488 5220
rect 16540 5208 16546 5220
rect 17954 5208 17960 5220
rect 16540 5180 17960 5208
rect 16540 5168 16546 5180
rect 17954 5168 17960 5180
rect 18012 5168 18018 5220
rect 1104 4778 21620 4800
rect 1104 4726 7846 4778
rect 7898 4726 7910 4778
rect 7962 4726 7974 4778
rect 8026 4726 8038 4778
rect 8090 4726 14710 4778
rect 14762 4726 14774 4778
rect 14826 4726 14838 4778
rect 14890 4726 14902 4778
rect 14954 4726 21620 4778
rect 1104 4704 21620 4726
rect 20717 4667 20775 4673
rect 20717 4633 20729 4667
rect 20763 4664 20775 4667
rect 20806 4664 20812 4676
rect 20763 4636 20812 4664
rect 20763 4633 20775 4636
rect 20717 4627 20775 4633
rect 20806 4624 20812 4636
rect 20864 4624 20870 4676
rect 20530 4528 20536 4540
rect 20491 4500 20536 4528
rect 20530 4488 20536 4500
rect 20588 4488 20594 4540
rect 1104 4234 21620 4256
rect 1104 4182 4414 4234
rect 4466 4182 4478 4234
rect 4530 4182 4542 4234
rect 4594 4182 4606 4234
rect 4658 4182 11278 4234
rect 11330 4182 11342 4234
rect 11394 4182 11406 4234
rect 11458 4182 11470 4234
rect 11522 4182 18142 4234
rect 18194 4182 18206 4234
rect 18258 4182 18270 4234
rect 18322 4182 18334 4234
rect 18386 4182 21620 4234
rect 1104 4160 21620 4182
rect 16390 3944 16396 3996
rect 16448 3984 16454 3996
rect 19058 3984 19064 3996
rect 16448 3956 19064 3984
rect 16448 3944 16454 3956
rect 19058 3944 19064 3956
rect 19116 3944 19122 3996
rect 1104 3690 21620 3712
rect 1104 3638 7846 3690
rect 7898 3638 7910 3690
rect 7962 3638 7974 3690
rect 8026 3638 8038 3690
rect 8090 3638 14710 3690
rect 14762 3638 14774 3690
rect 14826 3638 14838 3690
rect 14890 3638 14902 3690
rect 14954 3638 21620 3690
rect 1104 3616 21620 3638
rect 1104 3146 21620 3168
rect 1104 3094 4414 3146
rect 4466 3094 4478 3146
rect 4530 3094 4542 3146
rect 4594 3094 4606 3146
rect 4658 3094 11278 3146
rect 11330 3094 11342 3146
rect 11394 3094 11406 3146
rect 11458 3094 11470 3146
rect 11522 3094 18142 3146
rect 18194 3094 18206 3146
rect 18258 3094 18270 3146
rect 18322 3094 18334 3146
rect 18386 3094 21620 3146
rect 1104 3072 21620 3094
rect 1104 2602 21620 2624
rect 1104 2550 7846 2602
rect 7898 2550 7910 2602
rect 7962 2550 7974 2602
rect 8026 2550 8038 2602
rect 8090 2550 14710 2602
rect 14762 2550 14774 2602
rect 14826 2550 14838 2602
rect 14890 2550 14902 2602
rect 14954 2550 21620 2602
rect 1104 2528 21620 2550
rect 1104 2058 21620 2080
rect 1104 2006 4414 2058
rect 4466 2006 4478 2058
rect 4530 2006 4542 2058
rect 4594 2006 4606 2058
rect 4658 2006 11278 2058
rect 11330 2006 11342 2058
rect 11394 2006 11406 2058
rect 11458 2006 11470 2058
rect 11522 2006 18142 2058
rect 18194 2006 18206 2058
rect 18258 2006 18270 2058
rect 18322 2006 18334 2058
rect 18386 2006 21620 2058
rect 1104 1984 21620 2006
rect 13906 1904 13912 1956
rect 13964 1944 13970 1956
rect 17954 1944 17960 1956
rect 13964 1916 17960 1944
rect 13964 1904 13970 1916
rect 17954 1904 17960 1916
rect 18012 1904 18018 1956
rect 16942 1156 16948 1208
rect 17000 1196 17006 1208
rect 17954 1196 17960 1208
rect 17000 1168 17960 1196
rect 17000 1156 17006 1168
rect 17954 1156 17960 1168
rect 18012 1156 18018 1208
<< via1 >>
rect 7846 19958 7898 20010
rect 7910 19958 7962 20010
rect 7974 19958 8026 20010
rect 8038 19958 8090 20010
rect 14710 19958 14762 20010
rect 14774 19958 14826 20010
rect 14838 19958 14890 20010
rect 14902 19958 14954 20010
rect 4712 19856 4764 19908
rect 17960 19856 18012 19908
rect 18696 19856 18748 19908
rect 20628 19856 20680 19908
rect 9588 19720 9640 19772
rect 17684 19763 17736 19772
rect 17684 19729 17693 19763
rect 17693 19729 17727 19763
rect 17727 19729 17736 19763
rect 17684 19720 17736 19729
rect 18512 19720 18564 19772
rect 19340 19720 19392 19772
rect 19708 19720 19760 19772
rect 4712 19652 4764 19704
rect 19800 19695 19852 19704
rect 19800 19661 19809 19695
rect 19809 19661 19843 19695
rect 19843 19661 19852 19695
rect 19800 19652 19852 19661
rect 5172 19516 5224 19568
rect 4414 19414 4466 19466
rect 4478 19414 4530 19466
rect 4542 19414 4594 19466
rect 4606 19414 4658 19466
rect 11278 19414 11330 19466
rect 11342 19414 11394 19466
rect 11406 19414 11458 19466
rect 11470 19414 11522 19466
rect 18142 19414 18194 19466
rect 18206 19414 18258 19466
rect 18270 19414 18322 19466
rect 18334 19414 18386 19466
rect 7932 19312 7984 19364
rect 9956 19312 10008 19364
rect 112 19108 164 19160
rect 848 19108 900 19160
rect 2412 19108 2464 19160
rect 4712 19108 4764 19160
rect 6092 19151 6144 19160
rect 6092 19117 6101 19151
rect 6101 19117 6135 19151
rect 6135 19117 6144 19151
rect 6092 19108 6144 19117
rect 5816 19040 5868 19092
rect 15384 19176 15436 19228
rect 17684 19176 17736 19228
rect 7564 19040 7616 19092
rect 5448 19015 5500 19024
rect 5448 18981 5457 19015
rect 5457 18981 5491 19015
rect 5491 18981 5500 19015
rect 5448 18972 5500 18981
rect 6092 18972 6144 19024
rect 6552 18972 6604 19024
rect 7932 19040 7984 19092
rect 8208 19040 8260 19092
rect 11152 19108 11204 19160
rect 12348 19151 12400 19160
rect 12348 19117 12357 19151
rect 12357 19117 12391 19151
rect 12391 19117 12400 19151
rect 12348 19108 12400 19117
rect 13360 19108 13412 19160
rect 9956 19083 10008 19092
rect 9956 19049 9990 19083
rect 9990 19049 10008 19083
rect 9956 19040 10008 19049
rect 12624 19083 12676 19092
rect 12624 19049 12658 19083
rect 12658 19049 12676 19083
rect 12624 19040 12676 19049
rect 15752 19083 15804 19092
rect 10692 18972 10744 19024
rect 11060 19015 11112 19024
rect 11060 18981 11069 19015
rect 11069 18981 11103 19015
rect 11103 18981 11112 19015
rect 11060 18972 11112 18981
rect 11888 18972 11940 19024
rect 13728 19015 13780 19024
rect 13728 18981 13737 19015
rect 13737 18981 13771 19015
rect 13771 18981 13780 19015
rect 13728 18972 13780 18981
rect 13820 18972 13872 19024
rect 15476 18972 15528 19024
rect 15752 19049 15761 19083
rect 15761 19049 15795 19083
rect 15795 19049 15804 19083
rect 15752 19040 15804 19049
rect 15660 19015 15712 19024
rect 15660 18981 15669 19015
rect 15669 18981 15703 19015
rect 15703 18981 15712 19015
rect 16764 19108 16816 19160
rect 18880 19108 18932 19160
rect 18788 19083 18840 19092
rect 18788 19049 18797 19083
rect 18797 19049 18831 19083
rect 18831 19049 18840 19083
rect 18788 19040 18840 19049
rect 15660 18972 15712 18981
rect 19248 18972 19300 19024
rect 7846 18870 7898 18922
rect 7910 18870 7962 18922
rect 7974 18870 8026 18922
rect 8038 18870 8090 18922
rect 14710 18870 14762 18922
rect 14774 18870 14826 18922
rect 14838 18870 14890 18922
rect 14902 18870 14954 18922
rect 4712 18768 4764 18820
rect 5172 18811 5224 18820
rect 5172 18777 5181 18811
rect 5181 18777 5215 18811
rect 5215 18777 5224 18811
rect 5172 18768 5224 18777
rect 2504 18700 2556 18752
rect 8300 18768 8352 18820
rect 9128 18768 9180 18820
rect 9864 18768 9916 18820
rect 6368 18700 6420 18752
rect 9404 18700 9456 18752
rect 11060 18700 11112 18752
rect 12440 18768 12492 18820
rect 2964 18632 3016 18684
rect 9588 18675 9640 18684
rect 9588 18641 9597 18675
rect 9597 18641 9631 18675
rect 9631 18641 9640 18675
rect 9588 18632 9640 18641
rect 10692 18675 10744 18684
rect 10692 18641 10701 18675
rect 10701 18641 10735 18675
rect 10735 18641 10744 18675
rect 10692 18632 10744 18641
rect 12808 18675 12860 18684
rect 12808 18641 12817 18675
rect 12817 18641 12851 18675
rect 12851 18641 12860 18675
rect 12808 18632 12860 18641
rect 13728 18675 13780 18684
rect 13728 18641 13762 18675
rect 13762 18641 13780 18675
rect 13728 18632 13780 18641
rect 14004 18632 14056 18684
rect 16764 18811 16816 18820
rect 16764 18777 16773 18811
rect 16773 18777 16807 18811
rect 16807 18777 16816 18811
rect 16764 18768 16816 18777
rect 17960 18768 18012 18820
rect 20076 18768 20128 18820
rect 20720 18811 20772 18820
rect 20720 18777 20729 18811
rect 20729 18777 20763 18811
rect 20763 18777 20772 18811
rect 20720 18768 20772 18777
rect 15384 18743 15436 18752
rect 15384 18709 15418 18743
rect 15418 18709 15436 18743
rect 15384 18700 15436 18709
rect 15476 18700 15528 18752
rect 18512 18700 18564 18752
rect 16580 18632 16632 18684
rect 17960 18632 18012 18684
rect 19524 18675 19576 18684
rect 19524 18641 19533 18675
rect 19533 18641 19567 18675
rect 19567 18641 19576 18675
rect 19524 18632 19576 18641
rect 19800 18632 19852 18684
rect 2412 18607 2464 18616
rect 2412 18573 2421 18607
rect 2421 18573 2455 18607
rect 2455 18573 2464 18607
rect 2412 18564 2464 18573
rect 5448 18564 5500 18616
rect 7656 18564 7708 18616
rect 8208 18564 8260 18616
rect 296 18428 348 18480
rect 6828 18496 6880 18548
rect 7472 18496 7524 18548
rect 8392 18496 8444 18548
rect 9956 18564 10008 18616
rect 10232 18607 10284 18616
rect 10232 18573 10241 18607
rect 10241 18573 10275 18607
rect 10275 18573 10284 18607
rect 10232 18564 10284 18573
rect 10692 18496 10744 18548
rect 12624 18496 12676 18548
rect 5172 18428 5224 18480
rect 9128 18428 9180 18480
rect 10876 18428 10928 18480
rect 10968 18428 11020 18480
rect 11704 18428 11756 18480
rect 13268 18428 13320 18480
rect 16396 18428 16448 18480
rect 19708 18607 19760 18616
rect 19708 18573 19717 18607
rect 19717 18573 19751 18607
rect 19751 18573 19760 18607
rect 19708 18564 19760 18573
rect 16948 18428 17000 18480
rect 21180 18428 21232 18480
rect 4414 18326 4466 18378
rect 4478 18326 4530 18378
rect 4542 18326 4594 18378
rect 4606 18326 4658 18378
rect 11278 18326 11330 18378
rect 11342 18326 11394 18378
rect 11406 18326 11458 18378
rect 11470 18326 11522 18378
rect 18142 18326 18194 18378
rect 18206 18326 18258 18378
rect 18270 18326 18322 18378
rect 18334 18326 18386 18378
rect 1952 18224 2004 18276
rect 6736 18224 6788 18276
rect 6828 18224 6880 18276
rect 9036 18224 9088 18276
rect 9128 18224 9180 18276
rect 13360 18267 13412 18276
rect 6920 18156 6972 18208
rect 7564 18088 7616 18140
rect 13360 18233 13369 18267
rect 13369 18233 13403 18267
rect 13403 18233 13412 18267
rect 13360 18224 13412 18233
rect 13912 18224 13964 18276
rect 14556 18224 14608 18276
rect 15844 18224 15896 18276
rect 19708 18224 19760 18276
rect 19892 18224 19944 18276
rect 10692 18088 10744 18140
rect 10876 18131 10928 18140
rect 10876 18097 10885 18131
rect 10885 18097 10919 18131
rect 10919 18097 10928 18131
rect 10876 18088 10928 18097
rect 11060 18131 11112 18140
rect 11060 18097 11069 18131
rect 11069 18097 11103 18131
rect 11103 18097 11112 18131
rect 11060 18088 11112 18097
rect 11520 18088 11572 18140
rect 11980 18088 12032 18140
rect 3608 18020 3660 18072
rect 4252 18020 4304 18072
rect 5172 18063 5224 18072
rect 5172 18029 5181 18063
rect 5181 18029 5215 18063
rect 5215 18029 5224 18063
rect 5172 18020 5224 18029
rect 8576 18020 8628 18072
rect 10232 18020 10284 18072
rect 19524 18156 19576 18208
rect 16580 18131 16632 18140
rect 10600 17952 10652 18004
rect 13728 17995 13780 18004
rect 13728 17961 13737 17995
rect 13737 17961 13771 17995
rect 13771 17961 13780 17995
rect 13728 17952 13780 17961
rect 3056 17884 3108 17936
rect 5908 17884 5960 17936
rect 7656 17927 7708 17936
rect 7656 17893 7665 17927
rect 7665 17893 7699 17927
rect 7699 17893 7708 17927
rect 7656 17884 7708 17893
rect 8208 17884 8260 17936
rect 8300 17884 8352 17936
rect 9956 17884 10008 17936
rect 11612 17884 11664 17936
rect 12072 17884 12124 17936
rect 12532 17884 12584 17936
rect 12992 17884 13044 17936
rect 13268 17884 13320 17936
rect 14004 18020 14056 18072
rect 15292 18020 15344 18072
rect 16304 18020 16356 18072
rect 16580 18097 16589 18131
rect 16589 18097 16623 18131
rect 16623 18097 16632 18131
rect 16580 18088 16632 18097
rect 19708 18088 19760 18140
rect 21916 18088 21968 18140
rect 19340 18020 19392 18072
rect 19616 18063 19668 18072
rect 19616 18029 19625 18063
rect 19625 18029 19659 18063
rect 19659 18029 19668 18063
rect 19616 18020 19668 18029
rect 14188 17952 14240 18004
rect 15108 17952 15160 18004
rect 15200 17952 15252 18004
rect 20628 18020 20680 18072
rect 21364 18020 21416 18072
rect 16488 17884 16540 17936
rect 19524 17884 19576 17936
rect 19892 17884 19944 17936
rect 20260 17884 20312 17936
rect 20444 17927 20496 17936
rect 20444 17893 20453 17927
rect 20453 17893 20487 17927
rect 20487 17893 20496 17927
rect 20444 17884 20496 17893
rect 20812 17884 20864 17936
rect 22468 17884 22520 17936
rect 7846 17782 7898 17834
rect 7910 17782 7962 17834
rect 7974 17782 8026 17834
rect 8038 17782 8090 17834
rect 14710 17782 14762 17834
rect 14774 17782 14826 17834
rect 14838 17782 14890 17834
rect 14902 17782 14954 17834
rect 2964 17723 3016 17732
rect 2964 17689 2973 17723
rect 2973 17689 3007 17723
rect 3007 17689 3016 17723
rect 2964 17680 3016 17689
rect 17040 17723 17092 17732
rect 17040 17689 17049 17723
rect 17049 17689 17083 17723
rect 17083 17689 17092 17723
rect 17040 17680 17092 17689
rect 20352 17723 20404 17732
rect 20352 17689 20361 17723
rect 20361 17689 20395 17723
rect 20395 17689 20404 17723
rect 20352 17680 20404 17689
rect 20904 17723 20956 17732
rect 20904 17689 20913 17723
rect 20913 17689 20947 17723
rect 20947 17689 20956 17723
rect 20904 17680 20956 17689
rect 2412 17612 2464 17664
rect 3148 17544 3200 17596
rect 5448 17612 5500 17664
rect 5632 17612 5684 17664
rect 18880 17612 18932 17664
rect 14464 17544 14516 17596
rect 17224 17544 17276 17596
rect 20168 17587 20220 17596
rect 20168 17553 20177 17587
rect 20177 17553 20211 17587
rect 20211 17553 20220 17587
rect 20168 17544 20220 17553
rect 1584 17519 1636 17528
rect 1584 17485 1593 17519
rect 1593 17485 1627 17519
rect 1627 17485 1636 17519
rect 1584 17476 1636 17485
rect 3332 17519 3384 17528
rect 3332 17485 3341 17519
rect 3341 17485 3375 17519
rect 3375 17485 3384 17519
rect 3332 17476 3384 17485
rect 10692 17476 10744 17528
rect 16764 17476 16816 17528
rect 17132 17519 17184 17528
rect 17132 17485 17141 17519
rect 17141 17485 17175 17519
rect 17175 17485 17184 17519
rect 17132 17476 17184 17485
rect 9128 17340 9180 17392
rect 12808 17340 12860 17392
rect 14280 17340 14332 17392
rect 18604 17340 18656 17392
rect 21732 17315 21784 17324
rect 4414 17238 4466 17290
rect 4478 17238 4530 17290
rect 4542 17238 4594 17290
rect 4606 17238 4658 17290
rect 11278 17238 11330 17290
rect 11342 17238 11394 17290
rect 11406 17238 11458 17290
rect 11470 17238 11522 17290
rect 18142 17238 18194 17290
rect 18206 17238 18258 17290
rect 18270 17238 18322 17290
rect 18334 17238 18386 17290
rect 21732 17281 21741 17315
rect 21741 17281 21775 17315
rect 21775 17281 21784 17315
rect 21732 17272 21784 17281
rect 4068 17136 4120 17188
rect 3148 17068 3200 17120
rect 2964 17000 3016 17052
rect 4160 17000 4212 17052
rect 7564 17068 7616 17120
rect 5540 17000 5592 17052
rect 9128 17043 9180 17052
rect 3332 16975 3384 16984
rect 3332 16941 3341 16975
rect 3341 16941 3375 16975
rect 3375 16941 3384 16975
rect 3332 16932 3384 16941
rect 5448 16932 5500 16984
rect 6552 16975 6604 16984
rect 6552 16941 6561 16975
rect 6561 16941 6595 16975
rect 6595 16941 6604 16975
rect 6552 16932 6604 16941
rect 9128 17009 9137 17043
rect 9137 17009 9171 17043
rect 9171 17009 9180 17043
rect 9128 17000 9180 17009
rect 11152 17136 11204 17188
rect 10324 17043 10376 17052
rect 10324 17009 10333 17043
rect 10333 17009 10367 17043
rect 10367 17009 10376 17043
rect 10324 17000 10376 17009
rect 17224 17136 17276 17188
rect 17960 17136 18012 17188
rect 20076 17136 20128 17188
rect 20352 17136 20404 17188
rect 12348 17068 12400 17120
rect 12900 17000 12952 17052
rect 18604 17043 18656 17052
rect 18604 17009 18613 17043
rect 18613 17009 18647 17043
rect 18647 17009 18656 17043
rect 18604 17000 18656 17009
rect 20168 17043 20220 17052
rect 16488 16975 16540 16984
rect 7012 16864 7064 16916
rect 2964 16839 3016 16848
rect 2964 16805 2973 16839
rect 2973 16805 3007 16839
rect 3007 16805 3016 16839
rect 2964 16796 3016 16805
rect 8300 16796 8352 16848
rect 8944 16839 8996 16848
rect 8944 16805 8953 16839
rect 8953 16805 8987 16839
rect 8987 16805 8996 16839
rect 8944 16796 8996 16805
rect 9772 16839 9824 16848
rect 9772 16805 9781 16839
rect 9781 16805 9815 16839
rect 9815 16805 9824 16839
rect 9772 16796 9824 16805
rect 10140 16839 10192 16848
rect 10140 16805 10149 16839
rect 10149 16805 10183 16839
rect 10183 16805 10192 16839
rect 10140 16796 10192 16805
rect 11888 16796 11940 16848
rect 13176 16839 13228 16848
rect 13176 16805 13185 16839
rect 13185 16805 13219 16839
rect 13219 16805 13228 16839
rect 13176 16796 13228 16805
rect 16488 16941 16497 16975
rect 16497 16941 16531 16975
rect 16531 16941 16540 16975
rect 16488 16932 16540 16941
rect 17132 16932 17184 16984
rect 20168 17009 20177 17043
rect 20177 17009 20211 17043
rect 20211 17009 20220 17043
rect 20168 17000 20220 17009
rect 19248 16975 19300 16984
rect 19248 16941 19257 16975
rect 19257 16941 19291 16975
rect 19291 16941 19300 16975
rect 19248 16932 19300 16941
rect 19340 16932 19392 16984
rect 18052 16796 18104 16848
rect 20444 16796 20496 16848
rect 7846 16694 7898 16746
rect 7910 16694 7962 16746
rect 7974 16694 8026 16746
rect 8038 16694 8090 16746
rect 14710 16694 14762 16746
rect 14774 16694 14826 16746
rect 14838 16694 14890 16746
rect 14902 16694 14954 16746
rect 5632 16524 5684 16576
rect 9128 16524 9180 16576
rect 2964 16456 3016 16508
rect 7380 16431 7432 16440
rect 7380 16397 7389 16431
rect 7389 16397 7423 16431
rect 7423 16397 7432 16431
rect 7380 16388 7432 16397
rect 7012 16320 7064 16372
rect 7564 16388 7616 16440
rect 11796 16592 11848 16644
rect 12348 16592 12400 16644
rect 13176 16592 13228 16644
rect 15568 16592 15620 16644
rect 16488 16592 16540 16644
rect 17132 16592 17184 16644
rect 18052 16635 18104 16644
rect 18052 16601 18061 16635
rect 18061 16601 18095 16635
rect 18095 16601 18104 16635
rect 18052 16592 18104 16601
rect 20168 16635 20220 16644
rect 20168 16601 20177 16635
rect 20177 16601 20211 16635
rect 20211 16601 20220 16635
rect 20168 16592 20220 16601
rect 10324 16524 10376 16576
rect 12900 16456 12952 16508
rect 13728 16456 13780 16508
rect 12440 16388 12492 16440
rect 15660 16456 15712 16508
rect 16396 16456 16448 16508
rect 19616 16524 19668 16576
rect 18880 16456 18932 16508
rect 20444 16456 20496 16508
rect 15568 16431 15620 16440
rect 15568 16397 15577 16431
rect 15577 16397 15611 16431
rect 15611 16397 15620 16431
rect 15568 16388 15620 16397
rect 13728 16252 13780 16304
rect 14372 16295 14424 16304
rect 14372 16261 14381 16295
rect 14381 16261 14415 16295
rect 14415 16261 14424 16295
rect 14372 16252 14424 16261
rect 4414 16150 4466 16202
rect 4478 16150 4530 16202
rect 4542 16150 4594 16202
rect 4606 16150 4658 16202
rect 11278 16150 11330 16202
rect 11342 16150 11394 16202
rect 11406 16150 11458 16202
rect 11470 16150 11522 16202
rect 18142 16150 18194 16202
rect 18206 16150 18258 16202
rect 18270 16150 18322 16202
rect 18334 16150 18386 16202
rect 3148 16091 3200 16100
rect 3148 16057 3157 16091
rect 3157 16057 3191 16091
rect 3191 16057 3200 16091
rect 3148 16048 3200 16057
rect 7012 16091 7064 16100
rect 7012 16057 7021 16091
rect 7021 16057 7055 16091
rect 7055 16057 7064 16091
rect 7012 16048 7064 16057
rect 7380 16048 7432 16100
rect 12900 16091 12952 16100
rect 12900 16057 12909 16091
rect 12909 16057 12943 16091
rect 12943 16057 12952 16091
rect 12900 16048 12952 16057
rect 19064 16048 19116 16100
rect 4896 15912 4948 15964
rect 5448 15912 5500 15964
rect 7748 15955 7800 15964
rect 7748 15921 7757 15955
rect 7757 15921 7791 15955
rect 7791 15921 7800 15955
rect 7748 15912 7800 15921
rect 10140 15955 10192 15964
rect 1584 15844 1636 15896
rect 6276 15844 6328 15896
rect 10140 15921 10149 15955
rect 10149 15921 10183 15955
rect 10183 15921 10192 15955
rect 10140 15912 10192 15921
rect 14372 15912 14424 15964
rect 19340 15980 19392 16032
rect 20076 15980 20128 16032
rect 15844 15955 15896 15964
rect 15844 15921 15853 15955
rect 15853 15921 15887 15955
rect 15887 15921 15896 15955
rect 15844 15912 15896 15921
rect 11060 15844 11112 15896
rect 11796 15887 11848 15896
rect 11796 15853 11830 15887
rect 11830 15853 11848 15887
rect 11796 15844 11848 15853
rect 14464 15887 14516 15896
rect 14464 15853 14473 15887
rect 14473 15853 14507 15887
rect 14507 15853 14516 15887
rect 14464 15844 14516 15853
rect 15660 15887 15712 15896
rect 15660 15853 15669 15887
rect 15669 15853 15703 15887
rect 15703 15853 15712 15887
rect 15660 15844 15712 15853
rect 19156 15844 19208 15896
rect 19800 15844 19852 15896
rect 2964 15776 3016 15828
rect 9404 15776 9456 15828
rect 7656 15751 7708 15760
rect 7656 15717 7665 15751
rect 7665 15717 7699 15751
rect 7699 15717 7708 15751
rect 7656 15708 7708 15717
rect 7846 15606 7898 15658
rect 7910 15606 7962 15658
rect 7974 15606 8026 15658
rect 8038 15606 8090 15658
rect 14710 15606 14762 15658
rect 14774 15606 14826 15658
rect 14838 15606 14890 15658
rect 14902 15606 14954 15658
rect 6276 15547 6328 15556
rect 6276 15513 6285 15547
rect 6285 15513 6319 15547
rect 6319 15513 6328 15547
rect 6276 15504 6328 15513
rect 20996 15504 21048 15556
rect 19156 15479 19208 15488
rect 3424 15411 3476 15420
rect 3424 15377 3433 15411
rect 3433 15377 3467 15411
rect 3467 15377 3476 15411
rect 3424 15368 3476 15377
rect 6828 15368 6880 15420
rect 8208 15368 8260 15420
rect 19156 15445 19165 15479
rect 19165 15445 19199 15479
rect 19199 15445 19208 15479
rect 19156 15436 19208 15445
rect 19340 15368 19392 15420
rect 3516 15343 3568 15352
rect 3516 15309 3525 15343
rect 3525 15309 3559 15343
rect 3559 15309 3568 15343
rect 3516 15300 3568 15309
rect 4896 15343 4948 15352
rect 2964 15232 3016 15284
rect 4896 15309 4905 15343
rect 4905 15309 4939 15343
rect 4939 15309 4948 15343
rect 4896 15300 4948 15309
rect 2228 15164 2280 15216
rect 7564 15164 7616 15216
rect 10048 15164 10100 15216
rect 18788 15164 18840 15216
rect 4414 15062 4466 15114
rect 4478 15062 4530 15114
rect 4542 15062 4594 15114
rect 4606 15062 4658 15114
rect 11278 15062 11330 15114
rect 11342 15062 11394 15114
rect 11406 15062 11458 15114
rect 11470 15062 11522 15114
rect 18142 15062 18194 15114
rect 18206 15062 18258 15114
rect 18270 15062 18322 15114
rect 18334 15062 18386 15114
rect 2964 15003 3016 15012
rect 2964 14969 2973 15003
rect 2973 14969 3007 15003
rect 3007 14969 3016 15003
rect 2964 14960 3016 14969
rect 3516 14960 3568 15012
rect 10968 14960 11020 15012
rect 12440 14960 12492 15012
rect 3424 14867 3476 14876
rect 3424 14833 3433 14867
rect 3433 14833 3467 14867
rect 3467 14833 3476 14867
rect 3424 14824 3476 14833
rect 3608 14824 3660 14876
rect 8392 14867 8444 14876
rect 8392 14833 8401 14867
rect 8401 14833 8435 14867
rect 8435 14833 8444 14867
rect 8392 14824 8444 14833
rect 8576 14867 8628 14876
rect 8576 14833 8585 14867
rect 8585 14833 8619 14867
rect 8619 14833 8628 14867
rect 8576 14824 8628 14833
rect 10232 14867 10284 14876
rect 10232 14833 10241 14867
rect 10241 14833 10275 14867
rect 10275 14833 10284 14867
rect 12532 14867 12584 14876
rect 10232 14824 10284 14833
rect 12532 14833 12541 14867
rect 12541 14833 12575 14867
rect 12575 14833 12584 14867
rect 12532 14824 12584 14833
rect 15200 14960 15252 15012
rect 15844 14960 15896 15012
rect 20444 15003 20496 15012
rect 20444 14969 20453 15003
rect 20453 14969 20487 15003
rect 20487 14969 20496 15003
rect 20444 14960 20496 14969
rect 13544 14867 13596 14876
rect 13544 14833 13553 14867
rect 13553 14833 13587 14867
rect 13587 14833 13596 14867
rect 13544 14824 13596 14833
rect 1584 14799 1636 14808
rect 1584 14765 1593 14799
rect 1593 14765 1627 14799
rect 1627 14765 1636 14799
rect 1584 14756 1636 14765
rect 2228 14756 2280 14808
rect 4252 14756 4304 14808
rect 9956 14756 10008 14808
rect 12716 14756 12768 14808
rect 14372 14756 14424 14808
rect 3608 14688 3660 14740
rect 19340 14892 19392 14944
rect 16856 14824 16908 14876
rect 19800 14824 19852 14876
rect 7656 14620 7708 14672
rect 8484 14620 8536 14672
rect 11980 14663 12032 14672
rect 11980 14629 11989 14663
rect 11989 14629 12023 14663
rect 12023 14629 12032 14663
rect 11980 14620 12032 14629
rect 12072 14620 12124 14672
rect 19524 14756 19576 14808
rect 16948 14663 17000 14672
rect 16948 14629 16957 14663
rect 16957 14629 16991 14663
rect 16991 14629 17000 14663
rect 16948 14620 17000 14629
rect 17040 14663 17092 14672
rect 17040 14629 17049 14663
rect 17049 14629 17083 14663
rect 17083 14629 17092 14663
rect 17040 14620 17092 14629
rect 7846 14518 7898 14570
rect 7910 14518 7962 14570
rect 7974 14518 8026 14570
rect 8038 14518 8090 14570
rect 14710 14518 14762 14570
rect 14774 14518 14826 14570
rect 14838 14518 14890 14570
rect 14902 14518 14954 14570
rect 3608 14459 3660 14468
rect 3608 14425 3617 14459
rect 3617 14425 3651 14459
rect 3651 14425 3660 14459
rect 3608 14416 3660 14425
rect 6828 14416 6880 14468
rect 10232 14416 10284 14468
rect 11980 14416 12032 14468
rect 20904 14459 20956 14468
rect 2228 14323 2280 14332
rect 2228 14289 2237 14323
rect 2237 14289 2271 14323
rect 2271 14289 2280 14323
rect 2228 14280 2280 14289
rect 6092 14323 6144 14332
rect 6092 14289 6101 14323
rect 6101 14289 6135 14323
rect 6135 14289 6144 14323
rect 6092 14280 6144 14289
rect 7656 14348 7708 14400
rect 15200 14348 15252 14400
rect 16396 14348 16448 14400
rect 18512 14348 18564 14400
rect 19524 14391 19576 14400
rect 19524 14357 19533 14391
rect 19533 14357 19567 14391
rect 19567 14357 19576 14391
rect 19524 14348 19576 14357
rect 8576 14323 8628 14332
rect 8576 14289 8610 14323
rect 8610 14289 8628 14323
rect 8576 14280 8628 14289
rect 11980 14280 12032 14332
rect 12624 14280 12676 14332
rect 13544 14280 13596 14332
rect 6184 14255 6236 14264
rect 6184 14221 6193 14255
rect 6193 14221 6227 14255
rect 6227 14221 6236 14255
rect 6184 14212 6236 14221
rect 6276 14255 6328 14264
rect 6276 14221 6285 14255
rect 6285 14221 6319 14255
rect 6319 14221 6328 14255
rect 6276 14212 6328 14221
rect 7748 14212 7800 14264
rect 12256 14212 12308 14264
rect 17132 14280 17184 14332
rect 20904 14425 20913 14459
rect 20913 14425 20947 14459
rect 20947 14425 20956 14459
rect 20904 14416 20956 14425
rect 17408 14255 17460 14264
rect 17408 14221 17417 14255
rect 17417 14221 17451 14255
rect 17451 14221 17460 14255
rect 17408 14212 17460 14221
rect 16856 14076 16908 14128
rect 4414 13974 4466 14026
rect 4478 13974 4530 14026
rect 4542 13974 4594 14026
rect 4606 13974 4658 14026
rect 11278 13974 11330 14026
rect 11342 13974 11394 14026
rect 11406 13974 11458 14026
rect 11470 13974 11522 14026
rect 18142 13974 18194 14026
rect 18206 13974 18258 14026
rect 18270 13974 18322 14026
rect 18334 13974 18386 14026
rect 6276 13872 6328 13924
rect 8208 13872 8260 13924
rect 8576 13872 8628 13924
rect 12624 13915 12676 13924
rect 6092 13736 6144 13788
rect 4436 13668 4488 13720
rect 9588 13736 9640 13788
rect 5264 13600 5316 13652
rect 10784 13668 10836 13720
rect 10968 13711 11020 13720
rect 10968 13677 10977 13711
rect 10977 13677 11011 13711
rect 11011 13677 11020 13711
rect 10968 13668 11020 13677
rect 12256 13804 12308 13856
rect 12624 13881 12633 13915
rect 12633 13881 12667 13915
rect 12667 13881 12676 13915
rect 12624 13872 12676 13881
rect 16856 13872 16908 13924
rect 16948 13872 17000 13924
rect 18696 13872 18748 13924
rect 19708 13872 19760 13924
rect 20444 13915 20496 13924
rect 20444 13881 20453 13915
rect 20453 13881 20487 13915
rect 20487 13881 20496 13915
rect 20444 13872 20496 13881
rect 17040 13804 17092 13856
rect 12440 13736 12492 13788
rect 17132 13779 17184 13788
rect 17132 13745 17141 13779
rect 17141 13745 17175 13779
rect 17175 13745 17184 13779
rect 17132 13736 17184 13745
rect 18512 13736 18564 13788
rect 7748 13600 7800 13652
rect 11152 13600 11204 13652
rect 12348 13600 12400 13652
rect 112 13532 164 13584
rect 7564 13532 7616 13584
rect 17408 13668 17460 13720
rect 18788 13711 18840 13720
rect 18788 13677 18797 13711
rect 18797 13677 18831 13711
rect 18831 13677 18840 13711
rect 18788 13668 18840 13677
rect 19708 13711 19760 13720
rect 19708 13677 19717 13711
rect 19717 13677 19751 13711
rect 19751 13677 19760 13711
rect 19708 13668 19760 13677
rect 16856 13575 16908 13584
rect 16856 13541 16865 13575
rect 16865 13541 16899 13575
rect 16899 13541 16908 13575
rect 16856 13532 16908 13541
rect 16948 13575 17000 13584
rect 16948 13541 16957 13575
rect 16957 13541 16991 13575
rect 16991 13541 17000 13575
rect 16948 13532 17000 13541
rect 17868 13532 17920 13584
rect 7846 13430 7898 13482
rect 7910 13430 7962 13482
rect 7974 13430 8026 13482
rect 8038 13430 8090 13482
rect 14710 13430 14762 13482
rect 14774 13430 14826 13482
rect 14838 13430 14890 13482
rect 14902 13430 14954 13482
rect 6184 13328 6236 13380
rect 10784 13328 10836 13380
rect 20536 13328 20588 13380
rect 20720 13371 20772 13380
rect 20720 13337 20729 13371
rect 20729 13337 20763 13371
rect 20763 13337 20772 13371
rect 20720 13328 20772 13337
rect 9588 13260 9640 13312
rect 10048 13303 10100 13312
rect 10048 13269 10059 13303
rect 10059 13269 10093 13303
rect 10093 13269 10100 13303
rect 10048 13260 10100 13269
rect 18788 13260 18840 13312
rect 4436 13192 4488 13244
rect 8576 13192 8628 13244
rect 13728 13192 13780 13244
rect 18696 13192 18748 13244
rect 19248 13192 19300 13244
rect 20168 13192 20220 13244
rect 5908 13124 5960 13176
rect 5264 13099 5316 13108
rect 5264 13065 5273 13099
rect 5273 13065 5307 13099
rect 5307 13065 5316 13099
rect 7564 13124 7616 13176
rect 13360 13124 13412 13176
rect 15568 13124 15620 13176
rect 5264 13056 5316 13065
rect 20628 13056 20680 13108
rect 4414 12886 4466 12938
rect 4478 12886 4530 12938
rect 4542 12886 4594 12938
rect 4606 12886 4658 12938
rect 11278 12886 11330 12938
rect 11342 12886 11394 12938
rect 11406 12886 11458 12938
rect 11470 12886 11522 12938
rect 18142 12886 18194 12938
rect 18206 12886 18258 12938
rect 18270 12886 18322 12938
rect 18334 12886 18386 12938
rect 11152 12784 11204 12836
rect 12716 12784 12768 12836
rect 13728 12784 13780 12836
rect 18880 12784 18932 12836
rect 20076 12827 20128 12836
rect 20076 12793 20085 12827
rect 20085 12793 20119 12827
rect 20119 12793 20128 12827
rect 20076 12784 20128 12793
rect 14556 12716 14608 12768
rect 19892 12716 19944 12768
rect 20628 12716 20680 12768
rect 7748 12648 7800 12700
rect 13360 12691 13412 12700
rect 13360 12657 13369 12691
rect 13369 12657 13403 12691
rect 13403 12657 13412 12691
rect 13360 12648 13412 12657
rect 13544 12691 13596 12700
rect 13544 12657 13553 12691
rect 13553 12657 13587 12691
rect 13587 12657 13596 12691
rect 13544 12648 13596 12657
rect 15016 12648 15068 12700
rect 15568 12691 15620 12700
rect 15568 12657 15577 12691
rect 15577 12657 15611 12691
rect 15611 12657 15620 12691
rect 15568 12648 15620 12657
rect 8208 12580 8260 12632
rect 11336 12623 11388 12632
rect 11336 12589 11345 12623
rect 11345 12589 11379 12623
rect 11379 12589 11388 12623
rect 11336 12580 11388 12589
rect 10140 12555 10192 12564
rect 10140 12521 10174 12555
rect 10174 12521 10192 12555
rect 10140 12512 10192 12521
rect 10784 12512 10836 12564
rect 8300 12444 8352 12496
rect 8668 12444 8720 12496
rect 13820 12512 13872 12564
rect 15200 12580 15252 12632
rect 15844 12580 15896 12632
rect 19064 12623 19116 12632
rect 19064 12589 19073 12623
rect 19073 12589 19107 12623
rect 19107 12589 19116 12623
rect 19064 12580 19116 12589
rect 16396 12512 16448 12564
rect 17500 12512 17552 12564
rect 13728 12444 13780 12496
rect 14096 12487 14148 12496
rect 14096 12453 14105 12487
rect 14105 12453 14139 12487
rect 14139 12453 14148 12487
rect 14096 12444 14148 12453
rect 14280 12444 14332 12496
rect 17960 12487 18012 12496
rect 17960 12453 17969 12487
rect 17969 12453 18003 12487
rect 18003 12453 18012 12487
rect 17960 12444 18012 12453
rect 7846 12342 7898 12394
rect 7910 12342 7962 12394
rect 7974 12342 8026 12394
rect 8038 12342 8090 12394
rect 14710 12342 14762 12394
rect 14774 12342 14826 12394
rect 14838 12342 14890 12394
rect 14902 12342 14954 12394
rect 8944 12240 8996 12292
rect 11336 12240 11388 12292
rect 14556 12283 14608 12292
rect 14556 12249 14565 12283
rect 14565 12249 14599 12283
rect 14599 12249 14608 12283
rect 14556 12240 14608 12249
rect 15016 12240 15068 12292
rect 17960 12240 18012 12292
rect 19064 12240 19116 12292
rect 19984 12240 20036 12292
rect 20260 12240 20312 12292
rect 7380 12172 7432 12224
rect 7748 12172 7800 12224
rect 14004 12172 14056 12224
rect 14096 12172 14148 12224
rect 10324 12104 10376 12156
rect 13544 12104 13596 12156
rect 15844 12104 15896 12156
rect 17960 12104 18012 12156
rect 19892 12147 19944 12156
rect 9680 12036 9732 12088
rect 10140 11968 10192 12020
rect 12440 12079 12492 12088
rect 12440 12045 12449 12079
rect 12449 12045 12483 12079
rect 12483 12045 12492 12079
rect 12440 12036 12492 12045
rect 15292 12079 15344 12088
rect 15292 12045 15301 12079
rect 15301 12045 15335 12079
rect 15335 12045 15344 12079
rect 15292 12036 15344 12045
rect 16948 12036 17000 12088
rect 19892 12113 19901 12147
rect 19901 12113 19935 12147
rect 19935 12113 19944 12147
rect 19892 12104 19944 12113
rect 20444 12147 20496 12156
rect 20444 12113 20453 12147
rect 20453 12113 20487 12147
rect 20487 12113 20496 12147
rect 20444 12104 20496 12113
rect 14280 11968 14332 12020
rect 8392 11943 8444 11952
rect 8392 11909 8401 11943
rect 8401 11909 8435 11943
rect 8435 11909 8444 11943
rect 8392 11900 8444 11909
rect 14096 11943 14148 11952
rect 14096 11909 14105 11943
rect 14105 11909 14139 11943
rect 14139 11909 14148 11943
rect 14096 11900 14148 11909
rect 14188 11900 14240 11952
rect 18972 11900 19024 11952
rect 4414 11798 4466 11850
rect 4478 11798 4530 11850
rect 4542 11798 4594 11850
rect 4606 11798 4658 11850
rect 11278 11798 11330 11850
rect 11342 11798 11394 11850
rect 11406 11798 11458 11850
rect 11470 11798 11522 11850
rect 18142 11798 18194 11850
rect 18206 11798 18258 11850
rect 18270 11798 18322 11850
rect 18334 11798 18386 11850
rect 9680 11696 9732 11748
rect 10324 11739 10376 11748
rect 10324 11705 10333 11739
rect 10333 11705 10367 11739
rect 10367 11705 10376 11739
rect 10324 11696 10376 11705
rect 12440 11696 12492 11748
rect 12808 11696 12860 11748
rect 15200 11696 15252 11748
rect 15752 11696 15804 11748
rect 16396 11696 16448 11748
rect 17960 11696 18012 11748
rect 19156 11696 19208 11748
rect 12164 11628 12216 11680
rect 14556 11628 14608 11680
rect 7380 11603 7432 11612
rect 6736 11492 6788 11544
rect 7380 11569 7389 11603
rect 7389 11569 7423 11603
rect 7423 11569 7432 11603
rect 7380 11560 7432 11569
rect 8300 11560 8352 11612
rect 8392 11560 8444 11612
rect 14188 11603 14240 11612
rect 14188 11569 14197 11603
rect 14197 11569 14231 11603
rect 14231 11569 14240 11603
rect 14188 11560 14240 11569
rect 17500 11560 17552 11612
rect 8484 11492 8536 11544
rect 12716 11492 12768 11544
rect 14096 11535 14148 11544
rect 14096 11501 14105 11535
rect 14105 11501 14139 11535
rect 14139 11501 14148 11535
rect 14096 11492 14148 11501
rect 20260 11535 20312 11544
rect 20260 11501 20269 11535
rect 20269 11501 20303 11535
rect 20303 11501 20312 11535
rect 20260 11492 20312 11501
rect 14464 11424 14516 11476
rect 8208 11356 8260 11408
rect 13728 11356 13780 11408
rect 18788 11356 18840 11408
rect 7846 11254 7898 11306
rect 7910 11254 7962 11306
rect 7974 11254 8026 11306
rect 8038 11254 8090 11306
rect 14710 11254 14762 11306
rect 14774 11254 14826 11306
rect 14838 11254 14890 11306
rect 14902 11254 14954 11306
rect 8208 11195 8260 11204
rect 8208 11161 8217 11195
rect 8217 11161 8251 11195
rect 8251 11161 8260 11195
rect 8208 11152 8260 11161
rect 8668 11195 8720 11204
rect 8668 11161 8677 11195
rect 8677 11161 8711 11195
rect 8711 11161 8720 11195
rect 8668 11152 8720 11161
rect 13728 11195 13780 11204
rect 13728 11161 13737 11195
rect 13737 11161 13771 11195
rect 13771 11161 13780 11195
rect 13728 11152 13780 11161
rect 14464 11152 14516 11204
rect 18788 11195 18840 11204
rect 18788 11161 18797 11195
rect 18797 11161 18831 11195
rect 18831 11161 18840 11195
rect 18788 11152 18840 11161
rect 19432 11152 19484 11204
rect 8944 11084 8996 11136
rect 20260 11084 20312 11136
rect 10784 11059 10836 11068
rect 10784 11025 10793 11059
rect 10793 11025 10827 11059
rect 10827 11025 10836 11059
rect 10784 11016 10836 11025
rect 17316 11059 17368 11068
rect 8300 10948 8352 11000
rect 14280 10991 14332 11000
rect 14280 10957 14289 10991
rect 14289 10957 14323 10991
rect 14323 10957 14332 10991
rect 14280 10948 14332 10957
rect 14556 10948 14608 11000
rect 17316 11025 17325 11059
rect 17325 11025 17359 11059
rect 17359 11025 17368 11059
rect 17316 11016 17368 11025
rect 17868 11016 17920 11068
rect 20536 11059 20588 11068
rect 20536 11025 20545 11059
rect 20545 11025 20579 11059
rect 20579 11025 20588 11059
rect 20536 11016 20588 11025
rect 11980 10880 12032 10932
rect 12256 10880 12308 10932
rect 16488 10880 16540 10932
rect 16856 10948 16908 11000
rect 17224 10948 17276 11000
rect 17500 10991 17552 11000
rect 17500 10957 17509 10991
rect 17509 10957 17543 10991
rect 17543 10957 17552 10991
rect 17500 10948 17552 10957
rect 16948 10923 17000 10932
rect 16948 10889 16957 10923
rect 16957 10889 16991 10923
rect 16991 10889 17000 10923
rect 16948 10880 17000 10889
rect 12808 10812 12860 10864
rect 15292 10812 15344 10864
rect 16396 10812 16448 10864
rect 19248 10812 19300 10864
rect 4414 10710 4466 10762
rect 4478 10710 4530 10762
rect 4542 10710 4594 10762
rect 4606 10710 4658 10762
rect 11278 10710 11330 10762
rect 11342 10710 11394 10762
rect 11406 10710 11458 10762
rect 11470 10710 11522 10762
rect 18142 10710 18194 10762
rect 18206 10710 18258 10762
rect 18270 10710 18322 10762
rect 18334 10710 18386 10762
rect 1676 10608 1728 10660
rect 8300 10608 8352 10660
rect 10784 10608 10836 10660
rect 14188 10651 14240 10660
rect 14188 10617 14197 10651
rect 14197 10617 14231 10651
rect 14231 10617 14240 10651
rect 14188 10608 14240 10617
rect 17316 10608 17368 10660
rect 18696 10651 18748 10660
rect 18696 10617 18705 10651
rect 18705 10617 18739 10651
rect 18739 10617 18748 10651
rect 18696 10608 18748 10617
rect 20352 10608 20404 10660
rect 7748 10404 7800 10456
rect 9496 10336 9548 10388
rect 10600 10379 10652 10388
rect 10600 10345 10609 10379
rect 10609 10345 10643 10379
rect 10643 10345 10652 10379
rect 10600 10336 10652 10345
rect 12256 10472 12308 10524
rect 12808 10515 12860 10524
rect 12808 10481 12817 10515
rect 12817 10481 12851 10515
rect 12851 10481 12860 10515
rect 12808 10472 12860 10481
rect 16212 10472 16264 10524
rect 16488 10472 16540 10524
rect 19156 10472 19208 10524
rect 19708 10472 19760 10524
rect 11980 10404 12032 10456
rect 14280 10404 14332 10456
rect 20260 10447 20312 10456
rect 20260 10413 20269 10447
rect 20269 10413 20303 10447
rect 20303 10413 20312 10447
rect 20260 10404 20312 10413
rect 16856 10379 16908 10388
rect 16856 10345 16865 10379
rect 16865 10345 16899 10379
rect 16899 10345 16908 10379
rect 16856 10336 16908 10345
rect 18052 10336 18104 10388
rect 10692 10311 10744 10320
rect 10692 10277 10701 10311
rect 10701 10277 10735 10311
rect 10735 10277 10744 10311
rect 10692 10268 10744 10277
rect 11060 10268 11112 10320
rect 16948 10311 17000 10320
rect 16948 10277 16957 10311
rect 16957 10277 16991 10311
rect 16991 10277 17000 10311
rect 16948 10268 17000 10277
rect 19156 10311 19208 10320
rect 19156 10277 19165 10311
rect 19165 10277 19199 10311
rect 19199 10277 19208 10311
rect 19156 10268 19208 10277
rect 7846 10166 7898 10218
rect 7910 10166 7962 10218
rect 7974 10166 8026 10218
rect 8038 10166 8090 10218
rect 14710 10166 14762 10218
rect 14774 10166 14826 10218
rect 14838 10166 14890 10218
rect 14902 10166 14954 10218
rect 9496 10107 9548 10116
rect 9496 10073 9505 10107
rect 9505 10073 9539 10107
rect 9539 10073 9548 10107
rect 9496 10064 9548 10073
rect 10692 10064 10744 10116
rect 11060 10107 11112 10116
rect 11060 10073 11069 10107
rect 11069 10073 11103 10107
rect 11103 10073 11112 10107
rect 11060 10064 11112 10073
rect 17500 10064 17552 10116
rect 18052 10107 18104 10116
rect 18052 10073 18061 10107
rect 18061 10073 18095 10107
rect 18095 10073 18104 10107
rect 18052 10064 18104 10073
rect 19248 10064 19300 10116
rect 16212 10039 16264 10048
rect 16212 10005 16246 10039
rect 16246 10005 16264 10039
rect 16212 9996 16264 10005
rect 17776 9996 17828 10048
rect 9312 9928 9364 9980
rect 11060 9928 11112 9980
rect 15292 9928 15344 9980
rect 18512 9971 18564 9980
rect 18512 9937 18521 9971
rect 18521 9937 18555 9971
rect 18555 9937 18564 9971
rect 18512 9928 18564 9937
rect 19708 9928 19760 9980
rect 20536 9971 20588 9980
rect 20536 9937 20545 9971
rect 20545 9937 20579 9971
rect 20579 9937 20588 9971
rect 20536 9928 20588 9937
rect 7748 9860 7800 9912
rect 11152 9903 11204 9912
rect 11152 9869 11161 9903
rect 11161 9869 11195 9903
rect 11195 9869 11204 9903
rect 11152 9860 11204 9869
rect 12164 9724 12216 9776
rect 16948 9724 17000 9776
rect 4414 9622 4466 9674
rect 4478 9622 4530 9674
rect 4542 9622 4594 9674
rect 4606 9622 4658 9674
rect 11278 9622 11330 9674
rect 11342 9622 11394 9674
rect 11406 9622 11458 9674
rect 11470 9622 11522 9674
rect 18142 9622 18194 9674
rect 18206 9622 18258 9674
rect 18270 9622 18322 9674
rect 18334 9622 18386 9674
rect 9312 9563 9364 9572
rect 9312 9529 9321 9563
rect 9321 9529 9355 9563
rect 9355 9529 9364 9563
rect 9312 9520 9364 9529
rect 10600 9520 10652 9572
rect 19156 9520 19208 9572
rect 12808 9452 12860 9504
rect 11152 9384 11204 9436
rect 12256 9384 12308 9436
rect 15108 9452 15160 9504
rect 7748 9316 7800 9368
rect 10968 9248 11020 9300
rect 16856 9384 16908 9436
rect 18696 9384 18748 9436
rect 19432 9384 19484 9436
rect 13636 9316 13688 9368
rect 14188 9316 14240 9368
rect 15292 9359 15344 9368
rect 15292 9325 15301 9359
rect 15301 9325 15335 9359
rect 15335 9325 15344 9359
rect 15292 9316 15344 9325
rect 19064 9359 19116 9368
rect 19064 9325 19073 9359
rect 19073 9325 19107 9359
rect 19107 9325 19116 9359
rect 19064 9316 19116 9325
rect 12716 9223 12768 9232
rect 12716 9189 12725 9223
rect 12725 9189 12759 9223
rect 12759 9189 12768 9223
rect 12716 9180 12768 9189
rect 16396 9248 16448 9300
rect 17960 9180 18012 9232
rect 7846 9078 7898 9130
rect 7910 9078 7962 9130
rect 7974 9078 8026 9130
rect 8038 9078 8090 9130
rect 14710 9078 14762 9130
rect 14774 9078 14826 9130
rect 14838 9078 14890 9130
rect 14902 9078 14954 9130
rect 11060 9019 11112 9028
rect 11060 8985 11069 9019
rect 11069 8985 11103 9019
rect 11103 8985 11112 9019
rect 11060 8976 11112 8985
rect 12164 8976 12216 9028
rect 13452 9019 13504 9028
rect 13452 8985 13461 9019
rect 13461 8985 13495 9019
rect 13495 8985 13504 9019
rect 13452 8976 13504 8985
rect 11704 8908 11756 8960
rect 12716 8908 12768 8960
rect 17868 8976 17920 9028
rect 19708 9019 19760 9028
rect 19708 8985 19717 9019
rect 19717 8985 19751 9019
rect 19751 8985 19760 9019
rect 19708 8976 19760 8985
rect 21180 8976 21232 9028
rect 15292 8908 15344 8960
rect 18512 8908 18564 8960
rect 13544 8840 13596 8892
rect 15476 8883 15528 8892
rect 15476 8849 15485 8883
rect 15485 8849 15519 8883
rect 15519 8849 15528 8883
rect 15476 8840 15528 8849
rect 19432 8840 19484 8892
rect 19984 8883 20036 8892
rect 19984 8849 19993 8883
rect 19993 8849 20027 8883
rect 20027 8849 20036 8883
rect 19984 8840 20036 8849
rect 20536 8883 20588 8892
rect 20536 8849 20545 8883
rect 20545 8849 20579 8883
rect 20579 8849 20588 8883
rect 20536 8840 20588 8849
rect 10968 8772 11020 8824
rect 12256 8772 12308 8824
rect 11704 8704 11756 8756
rect 16856 8704 16908 8756
rect 19616 8704 19668 8756
rect 4414 8534 4466 8586
rect 4478 8534 4530 8586
rect 4542 8534 4594 8586
rect 4606 8534 4658 8586
rect 11278 8534 11330 8586
rect 11342 8534 11394 8586
rect 11406 8534 11458 8586
rect 11470 8534 11522 8586
rect 18142 8534 18194 8586
rect 18206 8534 18258 8586
rect 18270 8534 18322 8586
rect 18334 8534 18386 8586
rect 11612 8432 11664 8484
rect 20628 8432 20680 8484
rect 13544 8339 13596 8348
rect 13544 8305 13553 8339
rect 13553 8305 13587 8339
rect 13587 8305 13596 8339
rect 13544 8296 13596 8305
rect 11244 8271 11296 8280
rect 11244 8237 11253 8271
rect 11253 8237 11287 8271
rect 11287 8237 11296 8271
rect 11244 8228 11296 8237
rect 13360 8271 13412 8280
rect 13360 8237 13369 8271
rect 13369 8237 13403 8271
rect 13403 8237 13412 8271
rect 13360 8228 13412 8237
rect 20260 8271 20312 8280
rect 20260 8237 20269 8271
rect 20269 8237 20303 8271
rect 20303 8237 20312 8271
rect 20260 8228 20312 8237
rect 7846 7990 7898 8042
rect 7910 7990 7962 8042
rect 7974 7990 8026 8042
rect 8038 7990 8090 8042
rect 14710 7990 14762 8042
rect 14774 7990 14826 8042
rect 14838 7990 14890 8042
rect 14902 7990 14954 8042
rect 13360 7888 13412 7940
rect 15476 7888 15528 7940
rect 18052 7888 18104 7940
rect 18512 7888 18564 7940
rect 19432 7931 19484 7940
rect 19432 7897 19441 7931
rect 19441 7897 19475 7931
rect 19475 7897 19484 7931
rect 19432 7888 19484 7897
rect 11244 7820 11296 7872
rect 16304 7820 16356 7872
rect 9496 7795 9548 7804
rect 9496 7761 9530 7795
rect 9530 7761 9548 7795
rect 9496 7752 9548 7761
rect 10232 7752 10284 7804
rect 14556 7752 14608 7804
rect 7288 7684 7340 7736
rect 7748 7684 7800 7736
rect 14188 7727 14240 7736
rect 14188 7693 14197 7727
rect 14197 7693 14231 7727
rect 14231 7693 14240 7727
rect 14188 7684 14240 7693
rect 14280 7684 14332 7736
rect 16856 7727 16908 7736
rect 13636 7616 13688 7668
rect 16856 7693 16865 7727
rect 16865 7693 16899 7727
rect 16899 7693 16908 7727
rect 16856 7684 16908 7693
rect 19984 7795 20036 7804
rect 19984 7761 19993 7795
rect 19993 7761 20027 7795
rect 20027 7761 20036 7795
rect 19984 7752 20036 7761
rect 20536 7795 20588 7804
rect 20536 7761 20545 7795
rect 20545 7761 20579 7795
rect 20579 7761 20588 7795
rect 20536 7752 20588 7761
rect 17592 7684 17644 7736
rect 18052 7727 18104 7736
rect 18052 7693 18061 7727
rect 18061 7693 18095 7727
rect 18095 7693 18104 7727
rect 18052 7684 18104 7693
rect 10784 7548 10836 7600
rect 13912 7548 13964 7600
rect 16580 7548 16632 7600
rect 4414 7446 4466 7498
rect 4478 7446 4530 7498
rect 4542 7446 4594 7498
rect 4606 7446 4658 7498
rect 11278 7446 11330 7498
rect 11342 7446 11394 7498
rect 11406 7446 11458 7498
rect 11470 7446 11522 7498
rect 18142 7446 18194 7498
rect 18206 7446 18258 7498
rect 18270 7446 18322 7498
rect 18334 7446 18386 7498
rect 10232 7387 10284 7396
rect 10232 7353 10241 7387
rect 10241 7353 10275 7387
rect 10275 7353 10284 7387
rect 10232 7344 10284 7353
rect 14280 7387 14332 7396
rect 14280 7353 14289 7387
rect 14289 7353 14323 7387
rect 14323 7353 14332 7387
rect 14280 7344 14332 7353
rect 17592 7387 17644 7396
rect 17592 7353 17601 7387
rect 17601 7353 17635 7387
rect 17635 7353 17644 7387
rect 17592 7344 17644 7353
rect 10784 7251 10836 7260
rect 10784 7217 10793 7251
rect 10793 7217 10827 7251
rect 10827 7217 10836 7251
rect 10784 7208 10836 7217
rect 14556 7251 14608 7260
rect 14556 7217 14565 7251
rect 14565 7217 14599 7251
rect 14599 7217 14608 7251
rect 14556 7208 14608 7217
rect 13636 7140 13688 7192
rect 10692 7047 10744 7056
rect 10692 7013 10701 7047
rect 10701 7013 10735 7047
rect 10735 7013 10744 7047
rect 10692 7004 10744 7013
rect 14556 7072 14608 7124
rect 16580 7072 16632 7124
rect 7846 6902 7898 6954
rect 7910 6902 7962 6954
rect 7974 6902 8026 6954
rect 8038 6902 8090 6954
rect 14710 6902 14762 6954
rect 14774 6902 14826 6954
rect 14838 6902 14890 6954
rect 14902 6902 14954 6954
rect 10692 6800 10744 6852
rect 14188 6800 14240 6852
rect 16488 6800 16540 6852
rect 16856 6843 16908 6852
rect 16856 6809 16865 6843
rect 16865 6809 16899 6843
rect 16899 6809 16908 6843
rect 16856 6800 16908 6809
rect 17960 6800 18012 6852
rect 4068 6664 4120 6716
rect 7288 6639 7340 6648
rect 7288 6605 7297 6639
rect 7297 6605 7331 6639
rect 7331 6605 7340 6639
rect 7288 6596 7340 6605
rect 9496 6664 9548 6716
rect 10416 6596 10468 6648
rect 14648 6639 14700 6648
rect 14648 6605 14657 6639
rect 14657 6605 14691 6639
rect 14691 6605 14700 6639
rect 14648 6596 14700 6605
rect 18512 6732 18564 6784
rect 16580 6664 16632 6716
rect 20536 6707 20588 6716
rect 20536 6673 20545 6707
rect 20545 6673 20579 6707
rect 20579 6673 20588 6707
rect 20536 6664 20588 6673
rect 18604 6528 18656 6580
rect 17960 6460 18012 6512
rect 20720 6503 20772 6512
rect 20720 6469 20729 6503
rect 20729 6469 20763 6503
rect 20763 6469 20772 6503
rect 20720 6460 20772 6469
rect 4414 6358 4466 6410
rect 4478 6358 4530 6410
rect 4542 6358 4594 6410
rect 4606 6358 4658 6410
rect 11278 6358 11330 6410
rect 11342 6358 11394 6410
rect 11406 6358 11458 6410
rect 11470 6358 11522 6410
rect 18142 6358 18194 6410
rect 18206 6358 18258 6410
rect 18270 6358 18322 6410
rect 18334 6358 18386 6410
rect 13728 6256 13780 6308
rect 20720 6256 20772 6308
rect 7846 5814 7898 5866
rect 7910 5814 7962 5866
rect 7974 5814 8026 5866
rect 8038 5814 8090 5866
rect 14710 5814 14762 5866
rect 14774 5814 14826 5866
rect 14838 5814 14890 5866
rect 14902 5814 14954 5866
rect 13268 5712 13320 5764
rect 20536 5619 20588 5628
rect 20536 5585 20545 5619
rect 20545 5585 20579 5619
rect 20579 5585 20588 5619
rect 20536 5576 20588 5585
rect 4414 5270 4466 5322
rect 4478 5270 4530 5322
rect 4542 5270 4594 5322
rect 4606 5270 4658 5322
rect 11278 5270 11330 5322
rect 11342 5270 11394 5322
rect 11406 5270 11458 5322
rect 11470 5270 11522 5322
rect 18142 5270 18194 5322
rect 18206 5270 18258 5322
rect 18270 5270 18322 5322
rect 18334 5270 18386 5322
rect 16488 5168 16540 5220
rect 17960 5168 18012 5220
rect 7846 4726 7898 4778
rect 7910 4726 7962 4778
rect 7974 4726 8026 4778
rect 8038 4726 8090 4778
rect 14710 4726 14762 4778
rect 14774 4726 14826 4778
rect 14838 4726 14890 4778
rect 14902 4726 14954 4778
rect 20812 4624 20864 4676
rect 20536 4531 20588 4540
rect 20536 4497 20545 4531
rect 20545 4497 20579 4531
rect 20579 4497 20588 4531
rect 20536 4488 20588 4497
rect 4414 4182 4466 4234
rect 4478 4182 4530 4234
rect 4542 4182 4594 4234
rect 4606 4182 4658 4234
rect 11278 4182 11330 4234
rect 11342 4182 11394 4234
rect 11406 4182 11458 4234
rect 11470 4182 11522 4234
rect 18142 4182 18194 4234
rect 18206 4182 18258 4234
rect 18270 4182 18322 4234
rect 18334 4182 18386 4234
rect 16396 3944 16448 3996
rect 19064 3944 19116 3996
rect 7846 3638 7898 3690
rect 7910 3638 7962 3690
rect 7974 3638 8026 3690
rect 8038 3638 8090 3690
rect 14710 3638 14762 3690
rect 14774 3638 14826 3690
rect 14838 3638 14890 3690
rect 14902 3638 14954 3690
rect 4414 3094 4466 3146
rect 4478 3094 4530 3146
rect 4542 3094 4594 3146
rect 4606 3094 4658 3146
rect 11278 3094 11330 3146
rect 11342 3094 11394 3146
rect 11406 3094 11458 3146
rect 11470 3094 11522 3146
rect 18142 3094 18194 3146
rect 18206 3094 18258 3146
rect 18270 3094 18322 3146
rect 18334 3094 18386 3146
rect 7846 2550 7898 2602
rect 7910 2550 7962 2602
rect 7974 2550 8026 2602
rect 8038 2550 8090 2602
rect 14710 2550 14762 2602
rect 14774 2550 14826 2602
rect 14838 2550 14890 2602
rect 14902 2550 14954 2602
rect 4414 2006 4466 2058
rect 4478 2006 4530 2058
rect 4542 2006 4594 2058
rect 4606 2006 4658 2058
rect 11278 2006 11330 2058
rect 11342 2006 11394 2058
rect 11406 2006 11458 2058
rect 11470 2006 11522 2058
rect 18142 2006 18194 2058
rect 18206 2006 18258 2058
rect 18270 2006 18322 2058
rect 18334 2006 18386 2058
rect 13912 1904 13964 1956
rect 17960 1904 18012 1956
rect 16948 1156 17000 1208
rect 17960 1156 18012 1208
<< metal2 >>
rect 294 22176 350 22656
rect 846 22176 902 22656
rect 1398 22176 1454 22656
rect 1950 22176 2006 22656
rect 2502 22176 2558 22656
rect 3054 22176 3110 22656
rect 3606 22176 3662 22656
rect 4158 22176 4214 22656
rect 4710 22176 4766 22656
rect 5262 22176 5318 22656
rect 5814 22176 5870 22656
rect 6366 22176 6422 22656
rect 6918 22176 6974 22656
rect 7470 22176 7526 22656
rect 8022 22176 8078 22656
rect 8574 22176 8630 22656
rect 9126 22176 9182 22656
rect 9678 22176 9734 22656
rect 10230 22176 10286 22656
rect 10782 22176 10838 22656
rect 11334 22176 11390 22656
rect 11978 22176 12034 22656
rect 12530 22176 12586 22656
rect 13082 22176 13138 22656
rect 13634 22176 13690 22656
rect 14186 22176 14242 22656
rect 14738 22176 14794 22656
rect 15290 22176 15346 22656
rect 15842 22176 15898 22656
rect 16394 22176 16450 22656
rect 16946 22176 17002 22656
rect 17498 22176 17554 22656
rect 18050 22176 18106 22656
rect 18602 22176 18658 22656
rect 18878 22392 18934 22401
rect 18878 22327 18934 22336
rect 112 19160 164 19166
rect 112 19102 164 19108
rect 124 13590 152 19102
rect 308 18486 336 22176
rect 860 19166 888 22176
rect 1412 22106 1440 22176
rect 1412 22078 1716 22106
rect 848 19160 900 19166
rect 848 19102 900 19108
rect 296 18480 348 18486
rect 296 18422 348 18428
rect 1584 17528 1636 17534
rect 1584 17470 1636 17476
rect 1596 15902 1624 17470
rect 1584 15896 1636 15902
rect 1584 15838 1636 15844
rect 1596 14814 1624 15838
rect 1584 14808 1636 14814
rect 1584 14750 1636 14756
rect 112 13584 164 13590
rect 112 13526 164 13532
rect 1688 10666 1716 22078
rect 1964 18282 1992 22176
rect 2412 19160 2464 19166
rect 2412 19102 2464 19108
rect 2424 18622 2452 19102
rect 2516 18758 2544 22176
rect 2504 18752 2556 18758
rect 2504 18694 2556 18700
rect 2964 18684 3016 18690
rect 2964 18626 3016 18632
rect 2412 18616 2464 18622
rect 2412 18558 2464 18564
rect 1952 18276 2004 18282
rect 1952 18218 2004 18224
rect 2424 17670 2452 18558
rect 2976 17738 3004 18626
rect 3068 17942 3096 22176
rect 3620 18078 3648 22176
rect 3608 18072 3660 18078
rect 3608 18014 3660 18020
rect 3056 17936 3108 17942
rect 3056 17878 3108 17884
rect 2964 17732 3016 17738
rect 2964 17674 3016 17680
rect 2412 17664 2464 17670
rect 2412 17606 2464 17612
rect 2976 17058 3004 17674
rect 3148 17596 3200 17602
rect 3148 17538 3200 17544
rect 3160 17126 3188 17538
rect 3332 17528 3384 17534
rect 3332 17470 3384 17476
rect 3148 17120 3200 17126
rect 3148 17062 3200 17068
rect 2964 17052 3016 17058
rect 2964 16994 3016 17000
rect 2964 16848 3016 16854
rect 2964 16790 3016 16796
rect 2976 16514 3004 16790
rect 2964 16508 3016 16514
rect 2964 16450 3016 16456
rect 3160 16106 3188 17062
rect 3344 16990 3372 17470
rect 4068 17188 4120 17194
rect 4068 17130 4120 17136
rect 4080 17097 4108 17130
rect 4066 17088 4122 17097
rect 4172 17058 4200 22176
rect 4724 19914 4752 22176
rect 4712 19908 4764 19914
rect 4712 19850 4764 19856
rect 4712 19704 4764 19710
rect 4712 19646 4764 19652
rect 4388 19468 4684 19488
rect 4444 19466 4468 19468
rect 4524 19466 4548 19468
rect 4604 19466 4628 19468
rect 4466 19414 4468 19466
rect 4530 19414 4542 19466
rect 4604 19414 4606 19466
rect 4444 19412 4468 19414
rect 4524 19412 4548 19414
rect 4604 19412 4628 19414
rect 4388 19392 4684 19412
rect 4724 19166 4752 19646
rect 5172 19568 5224 19574
rect 5172 19510 5224 19516
rect 4712 19160 4764 19166
rect 4712 19102 4764 19108
rect 4724 18826 4752 19102
rect 5184 18826 5212 19510
rect 5276 19114 5304 22176
rect 5276 19086 5580 19114
rect 5828 19098 5856 22176
rect 6092 19160 6144 19166
rect 6092 19102 6144 19108
rect 5448 19024 5500 19030
rect 5448 18966 5500 18972
rect 4712 18820 4764 18826
rect 4712 18762 4764 18768
rect 5172 18820 5224 18826
rect 5172 18762 5224 18768
rect 5460 18622 5488 18966
rect 5448 18616 5500 18622
rect 5448 18558 5500 18564
rect 5172 18480 5224 18486
rect 5172 18422 5224 18428
rect 4388 18380 4684 18400
rect 4444 18378 4468 18380
rect 4524 18378 4548 18380
rect 4604 18378 4628 18380
rect 4466 18326 4468 18378
rect 4530 18326 4542 18378
rect 4604 18326 4606 18378
rect 4444 18324 4468 18326
rect 4524 18324 4548 18326
rect 4604 18324 4628 18326
rect 4388 18304 4684 18324
rect 5184 18078 5212 18422
rect 4252 18072 4304 18078
rect 4252 18014 4304 18020
rect 5172 18072 5224 18078
rect 5172 18014 5224 18020
rect 4066 17023 4122 17032
rect 4160 17052 4212 17058
rect 4160 16994 4212 17000
rect 3332 16984 3384 16990
rect 3332 16926 3384 16932
rect 3148 16100 3200 16106
rect 3148 16042 3200 16048
rect 2964 15828 3016 15834
rect 2964 15770 3016 15776
rect 2976 15290 3004 15770
rect 3424 15420 3476 15426
rect 3424 15362 3476 15368
rect 2964 15284 3016 15290
rect 2964 15226 3016 15232
rect 2228 15216 2280 15222
rect 2228 15158 2280 15164
rect 2240 14814 2268 15158
rect 2976 15018 3004 15226
rect 2964 15012 3016 15018
rect 2964 14954 3016 14960
rect 3436 14882 3464 15362
rect 3516 15352 3568 15358
rect 3516 15294 3568 15300
rect 3528 15018 3556 15294
rect 3516 15012 3568 15018
rect 3516 14954 3568 14960
rect 3424 14876 3476 14882
rect 3424 14818 3476 14824
rect 3608 14876 3660 14882
rect 3608 14818 3660 14824
rect 2228 14808 2280 14814
rect 2228 14750 2280 14756
rect 2240 14338 2268 14750
rect 3620 14746 3648 14818
rect 4264 14814 4292 18014
rect 5460 17670 5488 18558
rect 5448 17664 5500 17670
rect 5448 17606 5500 17612
rect 4388 17292 4684 17312
rect 4444 17290 4468 17292
rect 4524 17290 4548 17292
rect 4604 17290 4628 17292
rect 4466 17238 4468 17290
rect 4530 17238 4542 17290
rect 4604 17238 4606 17290
rect 4444 17236 4468 17238
rect 4524 17236 4548 17238
rect 4604 17236 4628 17238
rect 4388 17216 4684 17236
rect 5552 17058 5580 19086
rect 5816 19092 5868 19098
rect 5816 19034 5868 19040
rect 6104 19030 6132 19102
rect 6092 19024 6144 19030
rect 6092 18966 6144 18972
rect 6380 18758 6408 22176
rect 6552 19024 6604 19030
rect 6552 18966 6604 18972
rect 6368 18752 6420 18758
rect 6368 18694 6420 18700
rect 5908 17936 5960 17942
rect 5908 17878 5960 17884
rect 5632 17664 5684 17670
rect 5632 17606 5684 17612
rect 5540 17052 5592 17058
rect 5540 16994 5592 17000
rect 5448 16984 5500 16990
rect 5448 16926 5500 16932
rect 4388 16204 4684 16224
rect 4444 16202 4468 16204
rect 4524 16202 4548 16204
rect 4604 16202 4628 16204
rect 4466 16150 4468 16202
rect 4530 16150 4542 16202
rect 4604 16150 4606 16202
rect 4444 16148 4468 16150
rect 4524 16148 4548 16150
rect 4604 16148 4628 16150
rect 4388 16128 4684 16148
rect 5460 15970 5488 16926
rect 5644 16582 5672 17606
rect 5632 16576 5684 16582
rect 5632 16518 5684 16524
rect 4896 15964 4948 15970
rect 4896 15906 4948 15912
rect 5448 15964 5500 15970
rect 5448 15906 5500 15912
rect 4908 15358 4936 15906
rect 4896 15352 4948 15358
rect 4896 15294 4948 15300
rect 4388 15116 4684 15136
rect 4444 15114 4468 15116
rect 4524 15114 4548 15116
rect 4604 15114 4628 15116
rect 4466 15062 4468 15114
rect 4530 15062 4542 15114
rect 4604 15062 4606 15114
rect 4444 15060 4468 15062
rect 4524 15060 4548 15062
rect 4604 15060 4628 15062
rect 4388 15040 4684 15060
rect 4252 14808 4304 14814
rect 4252 14750 4304 14756
rect 3608 14740 3660 14746
rect 3608 14682 3660 14688
rect 3620 14474 3648 14682
rect 3608 14468 3660 14474
rect 3608 14410 3660 14416
rect 2228 14332 2280 14338
rect 2228 14274 2280 14280
rect 4388 14028 4684 14048
rect 4444 14026 4468 14028
rect 4524 14026 4548 14028
rect 4604 14026 4628 14028
rect 4466 13974 4468 14026
rect 4530 13974 4542 14026
rect 4604 13974 4606 14026
rect 4444 13972 4468 13974
rect 4524 13972 4548 13974
rect 4604 13972 4628 13974
rect 4388 13952 4684 13972
rect 4436 13720 4488 13726
rect 4436 13662 4488 13668
rect 4448 13250 4476 13662
rect 5264 13652 5316 13658
rect 5264 13594 5316 13600
rect 4436 13244 4488 13250
rect 4436 13186 4488 13192
rect 5276 13114 5304 13594
rect 5920 13182 5948 17878
rect 6564 16990 6592 18966
rect 6828 18548 6880 18554
rect 6828 18490 6880 18496
rect 6840 18282 6868 18490
rect 6736 18276 6788 18282
rect 6736 18218 6788 18224
rect 6828 18276 6880 18282
rect 6828 18218 6880 18224
rect 6552 16984 6604 16990
rect 6552 16926 6604 16932
rect 6276 15896 6328 15902
rect 6276 15838 6328 15844
rect 6288 15562 6316 15838
rect 6276 15556 6328 15562
rect 6276 15498 6328 15504
rect 6092 14332 6144 14338
rect 6092 14274 6144 14280
rect 6104 13794 6132 14274
rect 6184 14264 6236 14270
rect 6184 14206 6236 14212
rect 6276 14264 6328 14270
rect 6276 14206 6328 14212
rect 6092 13788 6144 13794
rect 6092 13730 6144 13736
rect 6196 13386 6224 14206
rect 6288 13930 6316 14206
rect 6276 13924 6328 13930
rect 6276 13866 6328 13872
rect 6184 13380 6236 13386
rect 6184 13322 6236 13328
rect 5908 13176 5960 13182
rect 5908 13118 5960 13124
rect 5264 13108 5316 13114
rect 5264 13050 5316 13056
rect 4388 12940 4684 12960
rect 4444 12938 4468 12940
rect 4524 12938 4548 12940
rect 4604 12938 4628 12940
rect 4466 12886 4468 12938
rect 4530 12886 4542 12938
rect 4604 12886 4606 12938
rect 4444 12884 4468 12886
rect 4524 12884 4548 12886
rect 4604 12884 4628 12886
rect 4388 12864 4684 12884
rect 4388 11852 4684 11872
rect 4444 11850 4468 11852
rect 4524 11850 4548 11852
rect 4604 11850 4628 11852
rect 4466 11798 4468 11850
rect 4530 11798 4542 11850
rect 4604 11798 4606 11850
rect 4444 11796 4468 11798
rect 4524 11796 4548 11798
rect 4604 11796 4628 11798
rect 4388 11776 4684 11796
rect 6748 11550 6776 18218
rect 6932 18214 6960 22176
rect 7484 18554 7512 22176
rect 8036 20202 8064 22176
rect 7760 20174 8064 20202
rect 7564 19092 7616 19098
rect 7564 19034 7616 19040
rect 7472 18548 7524 18554
rect 7472 18490 7524 18496
rect 6920 18208 6972 18214
rect 6920 18150 6972 18156
rect 7576 18146 7604 19034
rect 7656 18616 7708 18622
rect 7656 18558 7708 18564
rect 7564 18140 7616 18146
rect 7564 18082 7616 18088
rect 7576 17126 7604 18082
rect 7668 17942 7696 18558
rect 7656 17936 7708 17942
rect 7656 17878 7708 17884
rect 7564 17120 7616 17126
rect 7564 17062 7616 17068
rect 7012 16916 7064 16922
rect 7012 16858 7064 16864
rect 7024 16378 7052 16858
rect 7380 16440 7432 16446
rect 7380 16382 7432 16388
rect 7564 16440 7616 16446
rect 7564 16382 7616 16388
rect 7012 16372 7064 16378
rect 7012 16314 7064 16320
rect 7024 16106 7052 16314
rect 7392 16106 7420 16382
rect 7012 16100 7064 16106
rect 7012 16042 7064 16048
rect 7380 16100 7432 16106
rect 7380 16042 7432 16048
rect 6828 15420 6880 15426
rect 6828 15362 6880 15368
rect 6840 14474 6868 15362
rect 7576 15222 7604 16382
rect 7760 15970 7788 20174
rect 7820 20012 8116 20032
rect 7876 20010 7900 20012
rect 7956 20010 7980 20012
rect 8036 20010 8060 20012
rect 7898 19958 7900 20010
rect 7962 19958 7974 20010
rect 8036 19958 8038 20010
rect 7876 19956 7900 19958
rect 7956 19956 7980 19958
rect 8036 19956 8060 19958
rect 7820 19936 8116 19956
rect 7932 19364 7984 19370
rect 7932 19306 7984 19312
rect 7944 19098 7972 19306
rect 7932 19092 7984 19098
rect 7932 19034 7984 19040
rect 8208 19092 8260 19098
rect 8208 19034 8260 19040
rect 7820 18924 8116 18944
rect 7876 18922 7900 18924
rect 7956 18922 7980 18924
rect 8036 18922 8060 18924
rect 7898 18870 7900 18922
rect 7962 18870 7974 18922
rect 8036 18870 8038 18922
rect 7876 18868 7900 18870
rect 7956 18868 7980 18870
rect 8036 18868 8060 18870
rect 7820 18848 8116 18868
rect 8220 18622 8248 19034
rect 8300 18820 8352 18826
rect 8300 18762 8352 18768
rect 8208 18616 8260 18622
rect 8208 18558 8260 18564
rect 8312 17942 8340 18762
rect 8392 18548 8444 18554
rect 8392 18490 8444 18496
rect 8208 17936 8260 17942
rect 8208 17878 8260 17884
rect 8300 17936 8352 17942
rect 8300 17878 8352 17884
rect 7820 17836 8116 17856
rect 7876 17834 7900 17836
rect 7956 17834 7980 17836
rect 8036 17834 8060 17836
rect 7898 17782 7900 17834
rect 7962 17782 7974 17834
rect 8036 17782 8038 17834
rect 7876 17780 7900 17782
rect 7956 17780 7980 17782
rect 8036 17780 8060 17782
rect 7820 17760 8116 17780
rect 8220 17754 8248 17878
rect 8220 17726 8340 17754
rect 8312 16854 8340 17726
rect 8300 16848 8352 16854
rect 8300 16790 8352 16796
rect 7820 16748 8116 16768
rect 7876 16746 7900 16748
rect 7956 16746 7980 16748
rect 8036 16746 8060 16748
rect 7898 16694 7900 16746
rect 7962 16694 7974 16746
rect 8036 16694 8038 16746
rect 7876 16692 7900 16694
rect 7956 16692 7980 16694
rect 8036 16692 8060 16694
rect 7820 16672 8116 16692
rect 7748 15964 7800 15970
rect 7748 15906 7800 15912
rect 7656 15760 7708 15766
rect 7656 15702 7708 15708
rect 7564 15216 7616 15222
rect 7564 15158 7616 15164
rect 7668 14678 7696 15702
rect 7820 15660 8116 15680
rect 7876 15658 7900 15660
rect 7956 15658 7980 15660
rect 8036 15658 8060 15660
rect 7898 15606 7900 15658
rect 7962 15606 7974 15658
rect 8036 15606 8038 15658
rect 7876 15604 7900 15606
rect 7956 15604 7980 15606
rect 8036 15604 8060 15606
rect 7820 15584 8116 15604
rect 8208 15420 8260 15426
rect 8208 15362 8260 15368
rect 7656 14672 7708 14678
rect 7656 14614 7708 14620
rect 6828 14468 6880 14474
rect 6828 14410 6880 14416
rect 7668 14406 7696 14614
rect 7820 14572 8116 14592
rect 7876 14570 7900 14572
rect 7956 14570 7980 14572
rect 8036 14570 8060 14572
rect 7898 14518 7900 14570
rect 7962 14518 7974 14570
rect 8036 14518 8038 14570
rect 7876 14516 7900 14518
rect 7956 14516 7980 14518
rect 8036 14516 8060 14518
rect 7820 14496 8116 14516
rect 7656 14400 7708 14406
rect 7656 14342 7708 14348
rect 7748 14264 7800 14270
rect 7748 14206 7800 14212
rect 7760 13658 7788 14206
rect 8220 13930 8248 15362
rect 8208 13924 8260 13930
rect 8208 13866 8260 13872
rect 7748 13652 7800 13658
rect 7748 13594 7800 13600
rect 7564 13584 7616 13590
rect 7564 13526 7616 13532
rect 7576 13182 7604 13526
rect 7564 13176 7616 13182
rect 7564 13118 7616 13124
rect 7760 12706 7788 13594
rect 7820 13484 8116 13504
rect 7876 13482 7900 13484
rect 7956 13482 7980 13484
rect 8036 13482 8060 13484
rect 7898 13430 7900 13482
rect 7962 13430 7974 13482
rect 8036 13430 8038 13482
rect 7876 13428 7900 13430
rect 7956 13428 7980 13430
rect 8036 13428 8060 13430
rect 7820 13408 8116 13428
rect 7748 12700 7800 12706
rect 7748 12642 7800 12648
rect 7760 12230 7788 12642
rect 8220 12638 8248 13866
rect 8208 12632 8260 12638
rect 8208 12574 8260 12580
rect 8312 12502 8340 16790
rect 8404 14882 8432 18490
rect 8588 18078 8616 22176
rect 9140 18826 9168 22176
rect 9588 19772 9640 19778
rect 9588 19714 9640 19720
rect 9128 18820 9180 18826
rect 9128 18762 9180 18768
rect 9404 18752 9456 18758
rect 9404 18694 9456 18700
rect 9128 18480 9180 18486
rect 9128 18422 9180 18428
rect 9140 18282 9168 18422
rect 9036 18276 9088 18282
rect 9036 18218 9088 18224
rect 9128 18276 9180 18282
rect 9128 18218 9180 18224
rect 9048 18185 9076 18218
rect 9034 18176 9090 18185
rect 9034 18111 9090 18120
rect 8576 18072 8628 18078
rect 8576 18014 8628 18020
rect 9128 17392 9180 17398
rect 9128 17334 9180 17340
rect 9140 17058 9168 17334
rect 9128 17052 9180 17058
rect 9128 16994 9180 17000
rect 8944 16848 8996 16854
rect 8944 16790 8996 16796
rect 8392 14876 8444 14882
rect 8392 14818 8444 14824
rect 8576 14876 8628 14882
rect 8576 14818 8628 14824
rect 8484 14672 8536 14678
rect 8484 14614 8536 14620
rect 8496 13810 8524 14614
rect 8588 14338 8616 14818
rect 8576 14332 8628 14338
rect 8576 14274 8628 14280
rect 8588 13930 8616 14274
rect 8576 13924 8628 13930
rect 8576 13866 8628 13872
rect 8496 13782 8616 13810
rect 8588 13250 8616 13782
rect 8576 13244 8628 13250
rect 8576 13186 8628 13192
rect 8300 12496 8352 12502
rect 8300 12438 8352 12444
rect 7820 12396 8116 12416
rect 7876 12394 7900 12396
rect 7956 12394 7980 12396
rect 8036 12394 8060 12396
rect 7898 12342 7900 12394
rect 7962 12342 7974 12394
rect 8036 12342 8038 12394
rect 7876 12340 7900 12342
rect 7956 12340 7980 12342
rect 8036 12340 8060 12342
rect 7820 12320 8116 12340
rect 7380 12224 7432 12230
rect 7380 12166 7432 12172
rect 7748 12224 7800 12230
rect 7748 12166 7800 12172
rect 7392 11618 7420 12166
rect 7380 11612 7432 11618
rect 7380 11554 7432 11560
rect 6736 11544 6788 11550
rect 6736 11486 6788 11492
rect 4388 10764 4684 10784
rect 4444 10762 4468 10764
rect 4524 10762 4548 10764
rect 4604 10762 4628 10764
rect 4466 10710 4468 10762
rect 4530 10710 4542 10762
rect 4604 10710 4606 10762
rect 4444 10708 4468 10710
rect 4524 10708 4548 10710
rect 4604 10708 4628 10710
rect 4388 10688 4684 10708
rect 1676 10660 1728 10666
rect 1676 10602 1728 10608
rect 7760 10462 7788 12166
rect 8392 11952 8444 11958
rect 8392 11894 8444 11900
rect 8404 11618 8432 11894
rect 8300 11612 8352 11618
rect 8300 11554 8352 11560
rect 8392 11612 8444 11618
rect 8392 11554 8444 11560
rect 8208 11408 8260 11414
rect 8208 11350 8260 11356
rect 7820 11308 8116 11328
rect 7876 11306 7900 11308
rect 7956 11306 7980 11308
rect 8036 11306 8060 11308
rect 7898 11254 7900 11306
rect 7962 11254 7974 11306
rect 8036 11254 8038 11306
rect 7876 11252 7900 11254
rect 7956 11252 7980 11254
rect 8036 11252 8060 11254
rect 7820 11232 8116 11252
rect 8220 11210 8248 11350
rect 8208 11204 8260 11210
rect 8208 11146 8260 11152
rect 8312 11006 8340 11554
rect 8484 11544 8536 11550
rect 8588 11532 8616 13186
rect 8668 12496 8720 12502
rect 8668 12438 8720 12444
rect 8536 11504 8616 11532
rect 8484 11486 8536 11492
rect 8680 11210 8708 12438
rect 8956 12298 8984 16790
rect 9140 16582 9168 16994
rect 9128 16576 9180 16582
rect 9128 16518 9180 16524
rect 9416 15834 9444 18694
rect 9600 18690 9628 19714
rect 9692 19250 9720 22176
rect 9956 19364 10008 19370
rect 9956 19306 10008 19312
rect 9692 19222 9904 19250
rect 9876 18826 9904 19222
rect 9968 19098 9996 19306
rect 10244 19137 10272 22176
rect 10230 19128 10286 19137
rect 9956 19092 10008 19098
rect 10230 19063 10286 19072
rect 9956 19034 10008 19040
rect 9864 18820 9916 18826
rect 9864 18762 9916 18768
rect 9588 18684 9640 18690
rect 9588 18626 9640 18632
rect 9968 18622 9996 19034
rect 10692 19024 10744 19030
rect 10692 18966 10744 18972
rect 10704 18690 10732 18966
rect 10796 18729 10824 22176
rect 11348 19658 11376 22176
rect 11348 19630 11652 19658
rect 11252 19468 11548 19488
rect 11308 19466 11332 19468
rect 11388 19466 11412 19468
rect 11468 19466 11492 19468
rect 11330 19414 11332 19466
rect 11394 19414 11406 19466
rect 11468 19414 11470 19466
rect 11308 19412 11332 19414
rect 11388 19412 11412 19414
rect 11468 19412 11492 19414
rect 11252 19392 11548 19412
rect 11152 19160 11204 19166
rect 11152 19102 11204 19108
rect 11060 19024 11112 19030
rect 11060 18966 11112 18972
rect 11072 18758 11100 18966
rect 11060 18752 11112 18758
rect 10782 18720 10838 18729
rect 10692 18684 10744 18690
rect 11060 18694 11112 18700
rect 10782 18655 10838 18664
rect 10692 18626 10744 18632
rect 9956 18616 10008 18622
rect 9956 18558 10008 18564
rect 10232 18616 10284 18622
rect 10232 18558 10284 18564
rect 10244 18078 10272 18558
rect 10704 18554 11008 18570
rect 10692 18548 11008 18554
rect 10744 18542 11008 18548
rect 10692 18490 10744 18496
rect 10980 18486 11008 18542
rect 10876 18480 10928 18486
rect 10876 18422 10928 18428
rect 10968 18480 11020 18486
rect 10968 18422 11020 18428
rect 10414 18176 10470 18185
rect 10888 18146 10916 18422
rect 11072 18146 11100 18694
rect 10414 18111 10470 18120
rect 10692 18140 10744 18146
rect 10232 18072 10284 18078
rect 10232 18014 10284 18020
rect 9956 17936 10008 17942
rect 9956 17878 10008 17884
rect 9770 16952 9826 16961
rect 9770 16887 9826 16896
rect 9784 16854 9812 16887
rect 9772 16848 9824 16854
rect 9772 16790 9824 16796
rect 9404 15828 9456 15834
rect 9404 15770 9456 15776
rect 9968 14814 9996 17878
rect 10324 17052 10376 17058
rect 10324 16994 10376 17000
rect 10140 16848 10192 16854
rect 10140 16790 10192 16796
rect 10152 15970 10180 16790
rect 10336 16582 10364 16994
rect 10324 16576 10376 16582
rect 10324 16518 10376 16524
rect 10140 15964 10192 15970
rect 10140 15906 10192 15912
rect 10048 15216 10100 15222
rect 10048 15158 10100 15164
rect 9956 14808 10008 14814
rect 9956 14750 10008 14756
rect 9588 13788 9640 13794
rect 9588 13730 9640 13736
rect 9600 13318 9628 13730
rect 10060 13318 10088 15158
rect 10232 14876 10284 14882
rect 10232 14818 10284 14824
rect 10244 14474 10272 14818
rect 10232 14468 10284 14474
rect 10232 14410 10284 14416
rect 9588 13312 9640 13318
rect 9588 13254 9640 13260
rect 10048 13312 10100 13318
rect 10048 13254 10100 13260
rect 10140 12564 10192 12570
rect 10140 12506 10192 12512
rect 8944 12292 8996 12298
rect 8944 12234 8996 12240
rect 8668 11204 8720 11210
rect 8668 11146 8720 11152
rect 8956 11142 8984 12234
rect 9680 12088 9732 12094
rect 9680 12030 9732 12036
rect 9692 11754 9720 12030
rect 10152 12026 10180 12506
rect 10324 12156 10376 12162
rect 10324 12098 10376 12104
rect 10140 12020 10192 12026
rect 10140 11962 10192 11968
rect 10336 11754 10364 12098
rect 9680 11748 9732 11754
rect 9680 11690 9732 11696
rect 10324 11748 10376 11754
rect 10324 11690 10376 11696
rect 8944 11136 8996 11142
rect 8944 11078 8996 11084
rect 8300 11000 8352 11006
rect 8300 10942 8352 10948
rect 8312 10666 8340 10942
rect 8300 10660 8352 10666
rect 8300 10602 8352 10608
rect 7748 10456 7800 10462
rect 7748 10398 7800 10404
rect 7760 9918 7788 10398
rect 9496 10388 9548 10394
rect 9496 10330 9548 10336
rect 7820 10220 8116 10240
rect 7876 10218 7900 10220
rect 7956 10218 7980 10220
rect 8036 10218 8060 10220
rect 7898 10166 7900 10218
rect 7962 10166 7974 10218
rect 8036 10166 8038 10218
rect 7876 10164 7900 10166
rect 7956 10164 7980 10166
rect 8036 10164 8060 10166
rect 7820 10144 8116 10164
rect 9508 10122 9536 10330
rect 9496 10116 9548 10122
rect 9496 10058 9548 10064
rect 9312 9980 9364 9986
rect 9312 9922 9364 9928
rect 7748 9912 7800 9918
rect 7748 9854 7800 9860
rect 4388 9676 4684 9696
rect 4444 9674 4468 9676
rect 4524 9674 4548 9676
rect 4604 9674 4628 9676
rect 4466 9622 4468 9674
rect 4530 9622 4542 9674
rect 4604 9622 4606 9674
rect 4444 9620 4468 9622
rect 4524 9620 4548 9622
rect 4604 9620 4628 9622
rect 4388 9600 4684 9620
rect 7760 9374 7788 9854
rect 9324 9578 9352 9922
rect 9312 9572 9364 9578
rect 9312 9514 9364 9520
rect 7748 9368 7800 9374
rect 7748 9310 7800 9316
rect 4388 8588 4684 8608
rect 4444 8586 4468 8588
rect 4524 8586 4548 8588
rect 4604 8586 4628 8588
rect 4466 8534 4468 8586
rect 4530 8534 4542 8586
rect 4604 8534 4606 8586
rect 4444 8532 4468 8534
rect 4524 8532 4548 8534
rect 4604 8532 4628 8534
rect 4388 8512 4684 8532
rect 7760 7742 7788 9310
rect 7820 9132 8116 9152
rect 7876 9130 7900 9132
rect 7956 9130 7980 9132
rect 8036 9130 8060 9132
rect 7898 9078 7900 9130
rect 7962 9078 7974 9130
rect 8036 9078 8038 9130
rect 7876 9076 7900 9078
rect 7956 9076 7980 9078
rect 8036 9076 8060 9078
rect 7820 9056 8116 9076
rect 7820 8044 8116 8064
rect 7876 8042 7900 8044
rect 7956 8042 7980 8044
rect 8036 8042 8060 8044
rect 7898 7990 7900 8042
rect 7962 7990 7974 8042
rect 8036 7990 8038 8042
rect 7876 7988 7900 7990
rect 7956 7988 7980 7990
rect 8036 7988 8060 7990
rect 7820 7968 8116 7988
rect 9496 7804 9548 7810
rect 9496 7746 9548 7752
rect 10232 7804 10284 7810
rect 10232 7746 10284 7752
rect 7288 7736 7340 7742
rect 7288 7678 7340 7684
rect 7748 7736 7800 7742
rect 7748 7678 7800 7684
rect 4388 7500 4684 7520
rect 4444 7498 4468 7500
rect 4524 7498 4548 7500
rect 4604 7498 4628 7500
rect 4466 7446 4468 7498
rect 4530 7446 4542 7498
rect 4604 7446 4606 7498
rect 4444 7444 4468 7446
rect 4524 7444 4548 7446
rect 4604 7444 4628 7446
rect 4388 7424 4684 7444
rect 4068 6716 4120 6722
rect 4068 6658 4120 6664
rect 4080 5673 4108 6658
rect 7300 6654 7328 7678
rect 7820 6956 8116 6976
rect 7876 6954 7900 6956
rect 7956 6954 7980 6956
rect 8036 6954 8060 6956
rect 7898 6902 7900 6954
rect 7962 6902 7974 6954
rect 8036 6902 8038 6954
rect 7876 6900 7900 6902
rect 7956 6900 7980 6902
rect 8036 6900 8060 6902
rect 7820 6880 8116 6900
rect 9508 6722 9536 7746
rect 10244 7402 10272 7746
rect 10232 7396 10284 7402
rect 10232 7338 10284 7344
rect 9496 6716 9548 6722
rect 9496 6658 9548 6664
rect 10428 6654 10456 18111
rect 10692 18082 10744 18088
rect 10876 18140 10928 18146
rect 10876 18082 10928 18088
rect 11060 18140 11112 18146
rect 11060 18082 11112 18088
rect 10598 18040 10654 18049
rect 10598 17975 10600 17984
rect 10652 17975 10654 17984
rect 10600 17946 10652 17952
rect 10704 17534 10732 18082
rect 10692 17528 10744 17534
rect 10692 17470 10744 17476
rect 11164 17194 11192 19102
rect 11252 18380 11548 18400
rect 11308 18378 11332 18380
rect 11388 18378 11412 18380
rect 11468 18378 11492 18380
rect 11330 18326 11332 18378
rect 11394 18326 11406 18378
rect 11468 18326 11470 18378
rect 11308 18324 11332 18326
rect 11388 18324 11412 18326
rect 11468 18324 11492 18326
rect 11252 18304 11548 18324
rect 11520 18140 11572 18146
rect 11520 18082 11572 18088
rect 11532 17482 11560 18082
rect 11624 17942 11652 19630
rect 11888 19024 11940 19030
rect 11888 18966 11940 18972
rect 11704 18480 11756 18486
rect 11704 18422 11756 18428
rect 11612 17936 11664 17942
rect 11612 17878 11664 17884
rect 11532 17454 11652 17482
rect 11252 17292 11548 17312
rect 11308 17290 11332 17292
rect 11388 17290 11412 17292
rect 11468 17290 11492 17292
rect 11330 17238 11332 17290
rect 11394 17238 11406 17290
rect 11468 17238 11470 17290
rect 11308 17236 11332 17238
rect 11388 17236 11412 17238
rect 11468 17236 11492 17238
rect 11252 17216 11548 17236
rect 11152 17188 11204 17194
rect 11152 17130 11204 17136
rect 11252 16204 11548 16224
rect 11308 16202 11332 16204
rect 11388 16202 11412 16204
rect 11468 16202 11492 16204
rect 11330 16150 11332 16202
rect 11394 16150 11406 16202
rect 11468 16150 11470 16202
rect 11308 16148 11332 16150
rect 11388 16148 11412 16150
rect 11468 16148 11492 16150
rect 11252 16128 11548 16148
rect 11060 15896 11112 15902
rect 10980 15856 11060 15884
rect 10980 15018 11008 15856
rect 11060 15838 11112 15844
rect 11252 15116 11548 15136
rect 11308 15114 11332 15116
rect 11388 15114 11412 15116
rect 11468 15114 11492 15116
rect 11330 15062 11332 15114
rect 11394 15062 11406 15114
rect 11468 15062 11470 15114
rect 11308 15060 11332 15062
rect 11388 15060 11412 15062
rect 11468 15060 11492 15062
rect 11252 15040 11548 15060
rect 10968 15012 11020 15018
rect 10968 14954 11020 14960
rect 10980 13726 11008 14954
rect 11252 14028 11548 14048
rect 11308 14026 11332 14028
rect 11388 14026 11412 14028
rect 11468 14026 11492 14028
rect 11330 13974 11332 14026
rect 11394 13974 11406 14026
rect 11468 13974 11470 14026
rect 11308 13972 11332 13974
rect 11388 13972 11412 13974
rect 11468 13972 11492 13974
rect 11252 13952 11548 13972
rect 10784 13720 10836 13726
rect 10784 13662 10836 13668
rect 10968 13720 11020 13726
rect 10968 13662 11020 13668
rect 10796 13386 10824 13662
rect 11152 13652 11204 13658
rect 11152 13594 11204 13600
rect 10784 13380 10836 13386
rect 10784 13322 10836 13328
rect 10796 12570 10824 13322
rect 11164 12842 11192 13594
rect 11252 12940 11548 12960
rect 11308 12938 11332 12940
rect 11388 12938 11412 12940
rect 11468 12938 11492 12940
rect 11330 12886 11332 12938
rect 11394 12886 11406 12938
rect 11468 12886 11470 12938
rect 11308 12884 11332 12886
rect 11388 12884 11412 12886
rect 11468 12884 11492 12886
rect 11252 12864 11548 12884
rect 11152 12836 11204 12842
rect 11152 12778 11204 12784
rect 11336 12632 11388 12638
rect 11336 12574 11388 12580
rect 10784 12564 10836 12570
rect 10784 12506 10836 12512
rect 11348 12298 11376 12574
rect 11336 12292 11388 12298
rect 11336 12234 11388 12240
rect 11252 11852 11548 11872
rect 11308 11850 11332 11852
rect 11388 11850 11412 11852
rect 11468 11850 11492 11852
rect 11330 11798 11332 11850
rect 11394 11798 11406 11850
rect 11468 11798 11470 11850
rect 11308 11796 11332 11798
rect 11388 11796 11412 11798
rect 11468 11796 11492 11798
rect 11252 11776 11548 11796
rect 10784 11068 10836 11074
rect 10784 11010 10836 11016
rect 10796 10666 10824 11010
rect 11252 10764 11548 10784
rect 11308 10762 11332 10764
rect 11388 10762 11412 10764
rect 11468 10762 11492 10764
rect 11330 10710 11332 10762
rect 11394 10710 11406 10762
rect 11468 10710 11470 10762
rect 11308 10708 11332 10710
rect 11388 10708 11412 10710
rect 11468 10708 11492 10710
rect 11252 10688 11548 10708
rect 10784 10660 10836 10666
rect 10784 10602 10836 10608
rect 10600 10388 10652 10394
rect 10600 10330 10652 10336
rect 10612 9578 10640 10330
rect 10692 10320 10744 10326
rect 10692 10262 10744 10268
rect 11060 10320 11112 10326
rect 11060 10262 11112 10268
rect 10704 10122 10732 10262
rect 11072 10122 11100 10262
rect 10692 10116 10744 10122
rect 10692 10058 10744 10064
rect 11060 10116 11112 10122
rect 11060 10058 11112 10064
rect 11060 9980 11112 9986
rect 11060 9922 11112 9928
rect 10600 9572 10652 9578
rect 10600 9514 10652 9520
rect 10968 9300 11020 9306
rect 10968 9242 11020 9248
rect 10980 8830 11008 9242
rect 11072 9034 11100 9922
rect 11152 9912 11204 9918
rect 11152 9854 11204 9860
rect 11164 9442 11192 9854
rect 11252 9676 11548 9696
rect 11308 9674 11332 9676
rect 11388 9674 11412 9676
rect 11468 9674 11492 9676
rect 11330 9622 11332 9674
rect 11394 9622 11406 9674
rect 11468 9622 11470 9674
rect 11308 9620 11332 9622
rect 11388 9620 11412 9622
rect 11468 9620 11492 9622
rect 11252 9600 11548 9620
rect 11152 9436 11204 9442
rect 11152 9378 11204 9384
rect 11060 9028 11112 9034
rect 11060 8970 11112 8976
rect 10968 8824 11020 8830
rect 10968 8766 11020 8772
rect 11252 8588 11548 8608
rect 11308 8586 11332 8588
rect 11388 8586 11412 8588
rect 11468 8586 11492 8588
rect 11330 8534 11332 8586
rect 11394 8534 11406 8586
rect 11468 8534 11470 8586
rect 11308 8532 11332 8534
rect 11388 8532 11412 8534
rect 11468 8532 11492 8534
rect 11252 8512 11548 8532
rect 11624 8490 11652 17454
rect 11716 8966 11744 18422
rect 11900 16854 11928 18966
rect 11992 18146 12020 22176
rect 12348 19160 12400 19166
rect 12400 19120 12480 19148
rect 12348 19102 12400 19108
rect 12452 18826 12480 19120
rect 12440 18820 12492 18826
rect 12440 18762 12492 18768
rect 11980 18140 12032 18146
rect 11980 18082 12032 18088
rect 12072 17936 12124 17942
rect 12072 17878 12124 17884
rect 11888 16848 11940 16854
rect 11888 16790 11940 16796
rect 12084 16802 12112 17878
rect 12348 17120 12400 17126
rect 12348 17062 12400 17068
rect 12084 16774 12204 16802
rect 11796 16644 11848 16650
rect 11796 16586 11848 16592
rect 11808 15902 11836 16586
rect 11796 15896 11848 15902
rect 11796 15838 11848 15844
rect 11980 14672 12032 14678
rect 11980 14614 12032 14620
rect 12072 14672 12124 14678
rect 12072 14614 12124 14620
rect 11992 14474 12020 14614
rect 11980 14468 12032 14474
rect 11980 14410 12032 14416
rect 11980 14332 12032 14338
rect 11980 14274 12032 14280
rect 11992 11362 12020 14274
rect 12084 11498 12112 14614
rect 12176 11686 12204 16774
rect 12360 16650 12388 17062
rect 12348 16644 12400 16650
rect 12348 16586 12400 16592
rect 12452 16446 12480 18762
rect 12544 17942 12572 22176
rect 12624 19092 12676 19098
rect 12624 19034 12676 19040
rect 12636 18554 12664 19034
rect 12808 18684 12860 18690
rect 12808 18626 12860 18632
rect 12624 18548 12676 18554
rect 12624 18490 12676 18496
rect 12532 17936 12584 17942
rect 12532 17878 12584 17884
rect 12820 17398 12848 18626
rect 12992 17936 13044 17942
rect 12992 17878 13044 17884
rect 12808 17392 12860 17398
rect 12808 17334 12860 17340
rect 13004 17210 13032 17878
rect 13096 17346 13124 22176
rect 13360 19160 13412 19166
rect 13360 19102 13412 19108
rect 13268 18480 13320 18486
rect 13268 18422 13320 18428
rect 13280 17942 13308 18422
rect 13372 18282 13400 19102
rect 13360 18276 13412 18282
rect 13360 18218 13412 18224
rect 13268 17936 13320 17942
rect 13268 17878 13320 17884
rect 13096 17318 13492 17346
rect 13004 17182 13308 17210
rect 12900 17052 12952 17058
rect 12900 16994 12952 17000
rect 12912 16514 12940 16994
rect 13176 16848 13228 16854
rect 13176 16790 13228 16796
rect 13188 16650 13216 16790
rect 13176 16644 13228 16650
rect 13176 16586 13228 16592
rect 12900 16508 12952 16514
rect 12900 16450 12952 16456
rect 12440 16440 12492 16446
rect 12440 16382 12492 16388
rect 12452 15018 12480 16382
rect 12912 16106 12940 16450
rect 12900 16100 12952 16106
rect 12900 16042 12952 16048
rect 12440 15012 12492 15018
rect 12440 14954 12492 14960
rect 12532 14876 12584 14882
rect 12452 14836 12532 14864
rect 12256 14264 12308 14270
rect 12256 14206 12308 14212
rect 12268 13862 12296 14206
rect 12256 13856 12308 13862
rect 12256 13798 12308 13804
rect 12452 13794 12480 14836
rect 12532 14818 12584 14824
rect 12716 14808 12768 14814
rect 12716 14750 12768 14756
rect 12624 14332 12676 14338
rect 12624 14274 12676 14280
rect 12636 13930 12664 14274
rect 12624 13924 12676 13930
rect 12624 13866 12676 13872
rect 12440 13788 12492 13794
rect 12360 13748 12440 13776
rect 12360 13658 12388 13748
rect 12440 13730 12492 13736
rect 12348 13652 12400 13658
rect 12348 13594 12400 13600
rect 12728 12842 12756 14750
rect 12716 12836 12768 12842
rect 12716 12778 12768 12784
rect 12440 12088 12492 12094
rect 12440 12030 12492 12036
rect 12452 11754 12480 12030
rect 12440 11748 12492 11754
rect 12440 11690 12492 11696
rect 12164 11680 12216 11686
rect 12164 11622 12216 11628
rect 12728 11550 12756 12778
rect 12808 11748 12860 11754
rect 12808 11690 12860 11696
rect 12716 11544 12768 11550
rect 12084 11470 12296 11498
rect 12716 11486 12768 11492
rect 11992 11334 12204 11362
rect 11980 10932 12032 10938
rect 11980 10874 12032 10880
rect 11992 10462 12020 10874
rect 11980 10456 12032 10462
rect 11980 10398 12032 10404
rect 12176 9782 12204 11334
rect 12268 10938 12296 11470
rect 12256 10932 12308 10938
rect 12256 10874 12308 10880
rect 12820 10870 12848 11690
rect 12808 10864 12860 10870
rect 12808 10806 12860 10812
rect 12820 10530 12848 10806
rect 12256 10524 12308 10530
rect 12256 10466 12308 10472
rect 12808 10524 12860 10530
rect 12808 10466 12860 10472
rect 12164 9776 12216 9782
rect 12164 9718 12216 9724
rect 12176 9034 12204 9718
rect 12268 9442 12296 10466
rect 12820 9510 12848 10466
rect 12808 9504 12860 9510
rect 12808 9446 12860 9452
rect 12256 9436 12308 9442
rect 12256 9378 12308 9384
rect 12164 9028 12216 9034
rect 12164 8970 12216 8976
rect 11704 8960 11756 8966
rect 11704 8902 11756 8908
rect 11716 8762 11744 8902
rect 12268 8830 12296 9378
rect 12716 9232 12768 9238
rect 12716 9174 12768 9180
rect 12728 8966 12756 9174
rect 12716 8960 12768 8966
rect 12716 8902 12768 8908
rect 12256 8824 12308 8830
rect 12256 8766 12308 8772
rect 11704 8756 11756 8762
rect 11704 8698 11756 8704
rect 11612 8484 11664 8490
rect 11612 8426 11664 8432
rect 11244 8280 11296 8286
rect 11244 8222 11296 8228
rect 11256 7878 11284 8222
rect 11244 7872 11296 7878
rect 11244 7814 11296 7820
rect 10784 7600 10836 7606
rect 10784 7542 10836 7548
rect 10796 7266 10824 7542
rect 11252 7500 11548 7520
rect 11308 7498 11332 7500
rect 11388 7498 11412 7500
rect 11468 7498 11492 7500
rect 11330 7446 11332 7498
rect 11394 7446 11406 7498
rect 11468 7446 11470 7498
rect 11308 7444 11332 7446
rect 11388 7444 11412 7446
rect 11468 7444 11492 7446
rect 11252 7424 11548 7444
rect 10784 7260 10836 7266
rect 10784 7202 10836 7208
rect 10692 7056 10744 7062
rect 10692 6998 10744 7004
rect 10704 6858 10732 6998
rect 10692 6852 10744 6858
rect 10692 6794 10744 6800
rect 7288 6648 7340 6654
rect 7288 6590 7340 6596
rect 10416 6648 10468 6654
rect 10416 6590 10468 6596
rect 4388 6412 4684 6432
rect 4444 6410 4468 6412
rect 4524 6410 4548 6412
rect 4604 6410 4628 6412
rect 4466 6358 4468 6410
rect 4530 6358 4542 6410
rect 4604 6358 4606 6410
rect 4444 6356 4468 6358
rect 4524 6356 4548 6358
rect 4604 6356 4628 6358
rect 4388 6336 4684 6356
rect 11252 6412 11548 6432
rect 11308 6410 11332 6412
rect 11388 6410 11412 6412
rect 11468 6410 11492 6412
rect 11330 6358 11332 6410
rect 11394 6358 11406 6410
rect 11468 6358 11470 6410
rect 11308 6356 11332 6358
rect 11388 6356 11412 6358
rect 11468 6356 11492 6358
rect 11252 6336 11548 6356
rect 7820 5868 8116 5888
rect 7876 5866 7900 5868
rect 7956 5866 7980 5868
rect 8036 5866 8060 5868
rect 7898 5814 7900 5866
rect 7962 5814 7974 5866
rect 8036 5814 8038 5866
rect 7876 5812 7900 5814
rect 7956 5812 7980 5814
rect 8036 5812 8060 5814
rect 7820 5792 8116 5812
rect 13280 5770 13308 17182
rect 13360 13176 13412 13182
rect 13360 13118 13412 13124
rect 13372 12706 13400 13118
rect 13360 12700 13412 12706
rect 13360 12642 13412 12648
rect 13464 9034 13492 17318
rect 13544 14876 13596 14882
rect 13544 14818 13596 14824
rect 13556 14338 13584 14818
rect 13544 14332 13596 14338
rect 13544 14274 13596 14280
rect 13544 12700 13596 12706
rect 13544 12642 13596 12648
rect 13556 12162 13584 12642
rect 13544 12156 13596 12162
rect 13544 12098 13596 12104
rect 13648 9458 13676 22176
rect 13728 19024 13780 19030
rect 13728 18966 13780 18972
rect 13820 19024 13872 19030
rect 13820 18966 13872 18972
rect 13740 18690 13768 18966
rect 13728 18684 13780 18690
rect 13728 18626 13780 18632
rect 13832 18026 13860 18966
rect 14004 18684 14056 18690
rect 14004 18626 14056 18632
rect 13912 18276 13964 18282
rect 13912 18218 13964 18224
rect 13740 18010 13860 18026
rect 13728 18004 13860 18010
rect 13780 17998 13860 18004
rect 13728 17946 13780 17952
rect 13728 16508 13780 16514
rect 13728 16450 13780 16456
rect 13740 16310 13768 16450
rect 13728 16304 13780 16310
rect 13728 16246 13780 16252
rect 13728 13244 13780 13250
rect 13728 13186 13780 13192
rect 13740 12842 13768 13186
rect 13728 12836 13780 12842
rect 13728 12778 13780 12784
rect 13740 12502 13768 12778
rect 13820 12564 13872 12570
rect 13820 12506 13872 12512
rect 13728 12496 13780 12502
rect 13728 12438 13780 12444
rect 13728 11408 13780 11414
rect 13728 11350 13780 11356
rect 13740 11210 13768 11350
rect 13728 11204 13780 11210
rect 13728 11146 13780 11152
rect 13648 9430 13768 9458
rect 13636 9368 13688 9374
rect 13636 9310 13688 9316
rect 13452 9028 13504 9034
rect 13452 8970 13504 8976
rect 13544 8892 13596 8898
rect 13544 8834 13596 8840
rect 13556 8354 13584 8834
rect 13544 8348 13596 8354
rect 13544 8290 13596 8296
rect 13360 8280 13412 8286
rect 13360 8222 13412 8228
rect 13372 7946 13400 8222
rect 13360 7940 13412 7946
rect 13360 7882 13412 7888
rect 13648 7674 13676 9310
rect 13636 7668 13688 7674
rect 13636 7610 13688 7616
rect 13648 7198 13676 7610
rect 13636 7192 13688 7198
rect 13636 7134 13688 7140
rect 13740 6314 13768 9430
rect 13832 7418 13860 12506
rect 13924 7606 13952 18218
rect 14016 18078 14044 18626
rect 14004 18072 14056 18078
rect 14004 18014 14056 18020
rect 14200 18010 14228 22176
rect 14752 20202 14780 22176
rect 14568 20174 14780 20202
rect 14568 18282 14596 20174
rect 14684 20012 14980 20032
rect 14740 20010 14764 20012
rect 14820 20010 14844 20012
rect 14900 20010 14924 20012
rect 14762 19958 14764 20010
rect 14826 19958 14838 20010
rect 14900 19958 14902 20010
rect 14740 19956 14764 19958
rect 14820 19956 14844 19958
rect 14900 19956 14924 19958
rect 14684 19936 14980 19956
rect 14684 18924 14980 18944
rect 14740 18922 14764 18924
rect 14820 18922 14844 18924
rect 14900 18922 14924 18924
rect 14762 18870 14764 18922
rect 14826 18870 14838 18922
rect 14900 18870 14902 18922
rect 14740 18868 14764 18870
rect 14820 18868 14844 18870
rect 14900 18868 14924 18870
rect 14684 18848 14980 18868
rect 14556 18276 14608 18282
rect 14556 18218 14608 18224
rect 15304 18078 15332 22176
rect 15384 19228 15436 19234
rect 15384 19170 15436 19176
rect 15396 18758 15424 19170
rect 15750 19128 15806 19137
rect 15750 19063 15752 19072
rect 15804 19063 15806 19072
rect 15752 19034 15804 19040
rect 15476 19024 15528 19030
rect 15476 18966 15528 18972
rect 15660 19024 15712 19030
rect 15660 18966 15712 18972
rect 15488 18758 15516 18966
rect 15384 18752 15436 18758
rect 15384 18694 15436 18700
rect 15476 18752 15528 18758
rect 15476 18694 15528 18700
rect 15292 18072 15344 18078
rect 15198 18040 15254 18049
rect 14188 18004 14240 18010
rect 14188 17946 14240 17952
rect 15108 18004 15160 18010
rect 15292 18014 15344 18020
rect 15198 17975 15200 17984
rect 15108 17946 15160 17952
rect 15252 17975 15254 17984
rect 15200 17946 15252 17952
rect 14684 17836 14980 17856
rect 14740 17834 14764 17836
rect 14820 17834 14844 17836
rect 14900 17834 14924 17836
rect 14762 17782 14764 17834
rect 14826 17782 14838 17834
rect 14900 17782 14902 17834
rect 14740 17780 14764 17782
rect 14820 17780 14844 17782
rect 14900 17780 14924 17782
rect 14684 17760 14980 17780
rect 14464 17596 14516 17602
rect 14464 17538 14516 17544
rect 14280 17392 14332 17398
rect 14280 17334 14332 17340
rect 14292 12586 14320 17334
rect 14372 16304 14424 16310
rect 14372 16246 14424 16252
rect 14384 15970 14412 16246
rect 14372 15964 14424 15970
rect 14372 15906 14424 15912
rect 14384 14814 14412 15906
rect 14476 15902 14504 17538
rect 14684 16748 14980 16768
rect 14740 16746 14764 16748
rect 14820 16746 14844 16748
rect 14900 16746 14924 16748
rect 14762 16694 14764 16746
rect 14826 16694 14838 16746
rect 14900 16694 14902 16746
rect 14740 16692 14764 16694
rect 14820 16692 14844 16694
rect 14900 16692 14924 16694
rect 14684 16672 14980 16692
rect 14464 15896 14516 15902
rect 14464 15838 14516 15844
rect 14372 14808 14424 14814
rect 14372 14750 14424 14756
rect 14016 12558 14320 12586
rect 14016 12230 14044 12558
rect 14292 12502 14320 12558
rect 14096 12496 14148 12502
rect 14096 12438 14148 12444
rect 14280 12496 14332 12502
rect 14280 12438 14332 12444
rect 14108 12230 14136 12438
rect 14004 12224 14056 12230
rect 14004 12166 14056 12172
rect 14096 12224 14148 12230
rect 14292 12178 14320 12438
rect 14096 12166 14148 12172
rect 14200 12150 14320 12178
rect 14200 11958 14228 12150
rect 14280 12020 14332 12026
rect 14280 11962 14332 11968
rect 14096 11952 14148 11958
rect 14096 11894 14148 11900
rect 14188 11952 14240 11958
rect 14188 11894 14240 11900
rect 14108 11550 14136 11894
rect 14188 11612 14240 11618
rect 14188 11554 14240 11560
rect 14096 11544 14148 11550
rect 14096 11486 14148 11492
rect 14200 10666 14228 11554
rect 14292 11006 14320 11962
rect 14476 11482 14504 15838
rect 14684 15660 14980 15680
rect 14740 15658 14764 15660
rect 14820 15658 14844 15660
rect 14900 15658 14924 15660
rect 14762 15606 14764 15658
rect 14826 15606 14838 15658
rect 14900 15606 14902 15658
rect 14740 15604 14764 15606
rect 14820 15604 14844 15606
rect 14900 15604 14924 15606
rect 14684 15584 14980 15604
rect 14684 14572 14980 14592
rect 14740 14570 14764 14572
rect 14820 14570 14844 14572
rect 14900 14570 14924 14572
rect 14762 14518 14764 14570
rect 14826 14518 14838 14570
rect 14900 14518 14902 14570
rect 14740 14516 14764 14518
rect 14820 14516 14844 14518
rect 14900 14516 14924 14518
rect 14684 14496 14980 14516
rect 14684 13484 14980 13504
rect 14740 13482 14764 13484
rect 14820 13482 14844 13484
rect 14900 13482 14924 13484
rect 14762 13430 14764 13482
rect 14826 13430 14838 13482
rect 14900 13430 14902 13482
rect 14740 13428 14764 13430
rect 14820 13428 14844 13430
rect 14900 13428 14924 13430
rect 14684 13408 14980 13428
rect 14556 12768 14608 12774
rect 14556 12710 14608 12716
rect 14568 12298 14596 12710
rect 15016 12700 15068 12706
rect 15016 12642 15068 12648
rect 14684 12396 14980 12416
rect 14740 12394 14764 12396
rect 14820 12394 14844 12396
rect 14900 12394 14924 12396
rect 14762 12342 14764 12394
rect 14826 12342 14838 12394
rect 14900 12342 14902 12394
rect 14740 12340 14764 12342
rect 14820 12340 14844 12342
rect 14900 12340 14924 12342
rect 14684 12320 14980 12340
rect 15028 12298 15056 12642
rect 14556 12292 14608 12298
rect 14556 12234 14608 12240
rect 15016 12292 15068 12298
rect 15016 12234 15068 12240
rect 14556 11680 14608 11686
rect 14556 11622 14608 11628
rect 14464 11476 14516 11482
rect 14464 11418 14516 11424
rect 14476 11210 14504 11418
rect 14464 11204 14516 11210
rect 14384 11164 14464 11192
rect 14280 11000 14332 11006
rect 14280 10942 14332 10948
rect 14188 10660 14240 10666
rect 14188 10602 14240 10608
rect 14200 9374 14228 10602
rect 14292 10462 14320 10942
rect 14280 10456 14332 10462
rect 14280 10398 14332 10404
rect 14384 9481 14412 11164
rect 14464 11146 14516 11152
rect 14568 11006 14596 11622
rect 14684 11308 14980 11328
rect 14740 11306 14764 11308
rect 14820 11306 14844 11308
rect 14900 11306 14924 11308
rect 14762 11254 14764 11306
rect 14826 11254 14838 11306
rect 14900 11254 14902 11306
rect 14740 11252 14764 11254
rect 14820 11252 14844 11254
rect 14900 11252 14924 11254
rect 14684 11232 14980 11252
rect 14556 11000 14608 11006
rect 14556 10942 14608 10948
rect 14684 10220 14980 10240
rect 14740 10218 14764 10220
rect 14820 10218 14844 10220
rect 14900 10218 14924 10220
rect 14762 10166 14764 10218
rect 14826 10166 14838 10218
rect 14900 10166 14902 10218
rect 14740 10164 14764 10166
rect 14820 10164 14844 10166
rect 14900 10164 14924 10166
rect 14684 10144 14980 10164
rect 15120 9510 15148 17946
rect 15568 16644 15620 16650
rect 15672 16632 15700 18966
rect 15856 18282 15884 22176
rect 16408 18570 16436 22176
rect 16764 19160 16816 19166
rect 16764 19102 16816 19108
rect 16776 18826 16804 19102
rect 16764 18820 16816 18826
rect 16764 18762 16816 18768
rect 16580 18684 16632 18690
rect 16580 18626 16632 18632
rect 16408 18542 16528 18570
rect 16396 18480 16448 18486
rect 16396 18422 16448 18428
rect 15844 18276 15896 18282
rect 15844 18218 15896 18224
rect 16304 18072 16356 18078
rect 16304 18014 16356 18020
rect 15672 16604 15792 16632
rect 15568 16586 15620 16592
rect 15580 16446 15608 16586
rect 15660 16508 15712 16514
rect 15660 16450 15712 16456
rect 15568 16440 15620 16446
rect 15568 16382 15620 16388
rect 15672 15902 15700 16450
rect 15660 15896 15712 15902
rect 15660 15838 15712 15844
rect 15200 15012 15252 15018
rect 15200 14954 15252 14960
rect 15212 14406 15240 14954
rect 15200 14400 15252 14406
rect 15200 14342 15252 14348
rect 15568 13176 15620 13182
rect 15568 13118 15620 13124
rect 15580 12706 15608 13118
rect 15568 12700 15620 12706
rect 15568 12642 15620 12648
rect 15200 12632 15252 12638
rect 15200 12574 15252 12580
rect 15212 11754 15240 12574
rect 15292 12088 15344 12094
rect 15292 12030 15344 12036
rect 15200 11748 15252 11754
rect 15200 11690 15252 11696
rect 15304 10870 15332 12030
rect 15764 11754 15792 16604
rect 15844 15964 15896 15970
rect 15844 15906 15896 15912
rect 15856 15018 15884 15906
rect 15844 15012 15896 15018
rect 15844 14954 15896 14960
rect 15844 12632 15896 12638
rect 15844 12574 15896 12580
rect 15856 12162 15884 12574
rect 15844 12156 15896 12162
rect 15844 12098 15896 12104
rect 15752 11748 15804 11754
rect 15752 11690 15804 11696
rect 15292 10864 15344 10870
rect 15292 10806 15344 10812
rect 15304 9986 15332 10806
rect 16212 10524 16264 10530
rect 16212 10466 16264 10472
rect 16224 10054 16252 10466
rect 16212 10048 16264 10054
rect 16212 9990 16264 9996
rect 15292 9980 15344 9986
rect 15292 9922 15344 9928
rect 15108 9504 15160 9510
rect 14370 9472 14426 9481
rect 15108 9446 15160 9452
rect 14370 9407 14426 9416
rect 14188 9368 14240 9374
rect 14188 9310 14240 9316
rect 15292 9368 15344 9374
rect 15292 9310 15344 9316
rect 14684 9132 14980 9152
rect 14740 9130 14764 9132
rect 14820 9130 14844 9132
rect 14900 9130 14924 9132
rect 14762 9078 14764 9130
rect 14826 9078 14838 9130
rect 14900 9078 14902 9130
rect 14740 9076 14764 9078
rect 14820 9076 14844 9078
rect 14900 9076 14924 9078
rect 14684 9056 14980 9076
rect 15304 8966 15332 9310
rect 15292 8960 15344 8966
rect 15292 8902 15344 8908
rect 15476 8892 15528 8898
rect 15476 8834 15528 8840
rect 14684 8044 14980 8064
rect 14740 8042 14764 8044
rect 14820 8042 14844 8044
rect 14900 8042 14924 8044
rect 14762 7990 14764 8042
rect 14826 7990 14838 8042
rect 14900 7990 14902 8042
rect 14740 7988 14764 7990
rect 14820 7988 14844 7990
rect 14900 7988 14924 7990
rect 14684 7968 14980 7988
rect 15488 7946 15516 8834
rect 15476 7940 15528 7946
rect 15476 7882 15528 7888
rect 16316 7878 16344 18014
rect 16408 16514 16436 18422
rect 16500 17942 16528 18542
rect 16592 18146 16620 18626
rect 16960 18486 16988 22176
rect 17038 18720 17094 18729
rect 17038 18655 17094 18664
rect 16948 18480 17000 18486
rect 16948 18422 17000 18428
rect 16580 18140 16632 18146
rect 16580 18082 16632 18088
rect 16488 17936 16540 17942
rect 16488 17878 16540 17884
rect 17052 17738 17080 18655
rect 17040 17732 17092 17738
rect 17040 17674 17092 17680
rect 17224 17596 17276 17602
rect 17224 17538 17276 17544
rect 16764 17528 16816 17534
rect 16764 17470 16816 17476
rect 17132 17528 17184 17534
rect 17132 17470 17184 17476
rect 16488 16984 16540 16990
rect 16488 16926 16540 16932
rect 16500 16650 16528 16926
rect 16488 16644 16540 16650
rect 16488 16586 16540 16592
rect 16396 16508 16448 16514
rect 16396 16450 16448 16456
rect 16396 14400 16448 14406
rect 16396 14342 16448 14348
rect 16408 12570 16436 14342
rect 16776 13810 16804 17470
rect 17144 16990 17172 17470
rect 17236 17194 17264 17538
rect 17512 17210 17540 22176
rect 17958 21440 18014 21449
rect 17958 21375 18014 21384
rect 17972 19914 18000 21375
rect 17960 19908 18012 19914
rect 17960 19850 18012 19856
rect 17684 19772 17736 19778
rect 17684 19714 17736 19720
rect 17696 19234 17724 19714
rect 18064 19658 18092 22176
rect 18512 19772 18564 19778
rect 18512 19714 18564 19720
rect 17972 19630 18092 19658
rect 17684 19228 17736 19234
rect 17684 19170 17736 19176
rect 17972 18826 18000 19630
rect 18116 19468 18412 19488
rect 18172 19466 18196 19468
rect 18252 19466 18276 19468
rect 18332 19466 18356 19468
rect 18194 19414 18196 19466
rect 18258 19414 18270 19466
rect 18332 19414 18334 19466
rect 18172 19412 18196 19414
rect 18252 19412 18276 19414
rect 18332 19412 18356 19414
rect 18116 19392 18412 19412
rect 17960 18820 18012 18826
rect 17960 18762 18012 18768
rect 18524 18758 18552 19714
rect 18512 18752 18564 18758
rect 18512 18694 18564 18700
rect 17960 18684 18012 18690
rect 17960 18626 18012 18632
rect 17224 17188 17276 17194
rect 17512 17182 17816 17210
rect 17972 17194 18000 18626
rect 18116 18380 18412 18400
rect 18172 18378 18196 18380
rect 18252 18378 18276 18380
rect 18332 18378 18356 18380
rect 18194 18326 18196 18378
rect 18258 18326 18270 18378
rect 18332 18326 18334 18378
rect 18172 18324 18196 18326
rect 18252 18324 18276 18326
rect 18332 18324 18356 18326
rect 18116 18304 18412 18324
rect 18616 17482 18644 22176
rect 18694 21984 18750 21993
rect 18694 21919 18750 21928
rect 18708 19914 18736 21919
rect 18696 19908 18748 19914
rect 18696 19850 18748 19856
rect 18892 19166 18920 22327
rect 19154 22176 19210 22656
rect 19706 22176 19762 22656
rect 20258 22176 20314 22656
rect 20810 22176 20866 22656
rect 21362 22176 21418 22656
rect 21914 22176 21970 22656
rect 22466 22176 22522 22656
rect 18880 19160 18932 19166
rect 18880 19102 18932 19108
rect 18788 19092 18840 19098
rect 18788 19034 18840 19040
rect 18616 17454 18736 17482
rect 18604 17392 18656 17398
rect 18604 17334 18656 17340
rect 18116 17292 18412 17312
rect 18172 17290 18196 17292
rect 18252 17290 18276 17292
rect 18332 17290 18356 17292
rect 18194 17238 18196 17290
rect 18258 17238 18270 17290
rect 18332 17238 18334 17290
rect 18172 17236 18196 17238
rect 18252 17236 18276 17238
rect 18332 17236 18356 17238
rect 18116 17216 18412 17236
rect 17224 17130 17276 17136
rect 17132 16984 17184 16990
rect 17132 16926 17184 16932
rect 17144 16650 17172 16926
rect 17132 16644 17184 16650
rect 17132 16586 17184 16592
rect 16856 14876 16908 14882
rect 16856 14818 16908 14824
rect 16868 14134 16896 14818
rect 16948 14672 17000 14678
rect 16948 14614 17000 14620
rect 17040 14672 17092 14678
rect 17040 14614 17092 14620
rect 16856 14128 16908 14134
rect 16856 14070 16908 14076
rect 16868 13930 16896 14070
rect 16960 13930 16988 14614
rect 16856 13924 16908 13930
rect 16856 13866 16908 13872
rect 16948 13924 17000 13930
rect 16948 13866 17000 13872
rect 17052 13862 17080 14614
rect 17132 14332 17184 14338
rect 17132 14274 17184 14280
rect 17040 13856 17092 13862
rect 16776 13782 16988 13810
rect 17040 13798 17092 13804
rect 17144 13794 17172 14274
rect 17408 14264 17460 14270
rect 17408 14206 17460 14212
rect 16960 13590 16988 13782
rect 17132 13788 17184 13794
rect 17132 13730 17184 13736
rect 17420 13726 17448 14206
rect 17408 13720 17460 13726
rect 17408 13662 17460 13668
rect 16856 13584 16908 13590
rect 16856 13526 16908 13532
rect 16948 13584 17000 13590
rect 16948 13526 17000 13532
rect 16396 12564 16448 12570
rect 16396 12506 16448 12512
rect 16396 11748 16448 11754
rect 16396 11690 16448 11696
rect 16408 10870 16436 11690
rect 16868 11006 16896 13526
rect 17500 12564 17552 12570
rect 17500 12506 17552 12512
rect 16948 12088 17000 12094
rect 16948 12030 17000 12036
rect 16856 11000 16908 11006
rect 16856 10942 16908 10948
rect 16960 10938 16988 12030
rect 17512 11618 17540 12506
rect 17500 11612 17552 11618
rect 17500 11554 17552 11560
rect 17316 11068 17368 11074
rect 17316 11010 17368 11016
rect 17224 11000 17276 11006
rect 17224 10942 17276 10948
rect 16488 10932 16540 10938
rect 16488 10874 16540 10880
rect 16948 10932 17000 10938
rect 16948 10874 17000 10880
rect 16396 10864 16448 10870
rect 16396 10806 16448 10812
rect 16408 9306 16436 10806
rect 16500 10530 16528 10874
rect 16488 10524 16540 10530
rect 16488 10466 16540 10472
rect 16856 10388 16908 10394
rect 16856 10330 16908 10336
rect 16868 9442 16896 10330
rect 16948 10320 17000 10326
rect 16948 10262 17000 10268
rect 16960 9782 16988 10262
rect 16948 9776 17000 9782
rect 16948 9718 17000 9724
rect 16856 9436 16908 9442
rect 16856 9378 16908 9384
rect 16396 9300 16448 9306
rect 16396 9242 16448 9248
rect 16304 7872 16356 7878
rect 16304 7814 16356 7820
rect 14556 7804 14608 7810
rect 14556 7746 14608 7752
rect 14188 7736 14240 7742
rect 14188 7678 14240 7684
rect 14280 7736 14332 7742
rect 14280 7678 14332 7684
rect 13912 7600 13964 7606
rect 13912 7542 13964 7548
rect 13832 7390 13952 7418
rect 13728 6308 13780 6314
rect 13728 6250 13780 6256
rect 13268 5764 13320 5770
rect 13268 5706 13320 5712
rect 4066 5664 4122 5673
rect 4066 5599 4122 5608
rect 4388 5324 4684 5344
rect 4444 5322 4468 5324
rect 4524 5322 4548 5324
rect 4604 5322 4628 5324
rect 4466 5270 4468 5322
rect 4530 5270 4542 5322
rect 4604 5270 4606 5322
rect 4444 5268 4468 5270
rect 4524 5268 4548 5270
rect 4604 5268 4628 5270
rect 4388 5248 4684 5268
rect 11252 5324 11548 5344
rect 11308 5322 11332 5324
rect 11388 5322 11412 5324
rect 11468 5322 11492 5324
rect 11330 5270 11332 5322
rect 11394 5270 11406 5322
rect 11468 5270 11470 5322
rect 11308 5268 11332 5270
rect 11388 5268 11412 5270
rect 11468 5268 11492 5270
rect 11252 5248 11548 5268
rect 7820 4780 8116 4800
rect 7876 4778 7900 4780
rect 7956 4778 7980 4780
rect 8036 4778 8060 4780
rect 7898 4726 7900 4778
rect 7962 4726 7974 4778
rect 8036 4726 8038 4778
rect 7876 4724 7900 4726
rect 7956 4724 7980 4726
rect 8036 4724 8060 4726
rect 7820 4704 8116 4724
rect 4388 4236 4684 4256
rect 4444 4234 4468 4236
rect 4524 4234 4548 4236
rect 4604 4234 4628 4236
rect 4466 4182 4468 4234
rect 4530 4182 4542 4234
rect 4604 4182 4606 4234
rect 4444 4180 4468 4182
rect 4524 4180 4548 4182
rect 4604 4180 4628 4182
rect 4388 4160 4684 4180
rect 11252 4236 11548 4256
rect 11308 4234 11332 4236
rect 11388 4234 11412 4236
rect 11468 4234 11492 4236
rect 11330 4182 11332 4234
rect 11394 4182 11406 4234
rect 11468 4182 11470 4234
rect 11308 4180 11332 4182
rect 11388 4180 11412 4182
rect 11468 4180 11492 4182
rect 11252 4160 11548 4180
rect 7820 3692 8116 3712
rect 7876 3690 7900 3692
rect 7956 3690 7980 3692
rect 8036 3690 8060 3692
rect 7898 3638 7900 3690
rect 7962 3638 7974 3690
rect 8036 3638 8038 3690
rect 7876 3636 7900 3638
rect 7956 3636 7980 3638
rect 8036 3636 8060 3638
rect 7820 3616 8116 3636
rect 4388 3148 4684 3168
rect 4444 3146 4468 3148
rect 4524 3146 4548 3148
rect 4604 3146 4628 3148
rect 4466 3094 4468 3146
rect 4530 3094 4542 3146
rect 4604 3094 4606 3146
rect 4444 3092 4468 3094
rect 4524 3092 4548 3094
rect 4604 3092 4628 3094
rect 4388 3072 4684 3092
rect 11252 3148 11548 3168
rect 11308 3146 11332 3148
rect 11388 3146 11412 3148
rect 11468 3146 11492 3148
rect 11330 3094 11332 3146
rect 11394 3094 11406 3146
rect 11468 3094 11470 3146
rect 11308 3092 11332 3094
rect 11388 3092 11412 3094
rect 11468 3092 11492 3094
rect 11252 3072 11548 3092
rect 7820 2604 8116 2624
rect 7876 2602 7900 2604
rect 7956 2602 7980 2604
rect 8036 2602 8060 2604
rect 7898 2550 7900 2602
rect 7962 2550 7974 2602
rect 8036 2550 8038 2602
rect 7876 2548 7900 2550
rect 7956 2548 7980 2550
rect 8036 2548 8060 2550
rect 7820 2528 8116 2548
rect 4388 2060 4684 2080
rect 4444 2058 4468 2060
rect 4524 2058 4548 2060
rect 4604 2058 4628 2060
rect 4466 2006 4468 2058
rect 4530 2006 4542 2058
rect 4604 2006 4606 2058
rect 4444 2004 4468 2006
rect 4524 2004 4548 2006
rect 4604 2004 4628 2006
rect 4388 1984 4684 2004
rect 11252 2060 11548 2080
rect 11308 2058 11332 2060
rect 11388 2058 11412 2060
rect 11468 2058 11492 2060
rect 11330 2006 11332 2058
rect 11394 2006 11406 2058
rect 11468 2006 11470 2058
rect 11308 2004 11332 2006
rect 11388 2004 11412 2006
rect 11468 2004 11492 2006
rect 11252 1984 11548 2004
rect 13924 1962 13952 7390
rect 14200 6858 14228 7678
rect 14292 7402 14320 7678
rect 14280 7396 14332 7402
rect 14280 7338 14332 7344
rect 14568 7266 14596 7746
rect 14556 7260 14608 7266
rect 14556 7202 14608 7208
rect 14556 7124 14608 7130
rect 14556 7066 14608 7072
rect 14188 6852 14240 6858
rect 14188 6794 14240 6800
rect 14568 6738 14596 7066
rect 14684 6956 14980 6976
rect 14740 6954 14764 6956
rect 14820 6954 14844 6956
rect 14900 6954 14924 6956
rect 14762 6902 14764 6954
rect 14826 6902 14838 6954
rect 14900 6902 14902 6954
rect 14740 6900 14764 6902
rect 14820 6900 14844 6902
rect 14900 6900 14924 6902
rect 14684 6880 14980 6900
rect 14568 6710 14688 6738
rect 14660 6654 14688 6710
rect 14648 6648 14700 6654
rect 14648 6590 14700 6596
rect 14684 5868 14980 5888
rect 14740 5866 14764 5868
rect 14820 5866 14844 5868
rect 14900 5866 14924 5868
rect 14762 5814 14764 5866
rect 14826 5814 14838 5866
rect 14900 5814 14902 5866
rect 14740 5812 14764 5814
rect 14820 5812 14844 5814
rect 14900 5812 14924 5814
rect 14684 5792 14980 5812
rect 14684 4780 14980 4800
rect 14740 4778 14764 4780
rect 14820 4778 14844 4780
rect 14900 4778 14924 4780
rect 14762 4726 14764 4778
rect 14826 4726 14838 4778
rect 14900 4726 14902 4778
rect 14740 4724 14764 4726
rect 14820 4724 14844 4726
rect 14900 4724 14924 4726
rect 14684 4704 14980 4724
rect 16408 4002 16436 9242
rect 16868 8762 16896 9378
rect 16856 8756 16908 8762
rect 16856 8698 16908 8704
rect 16856 7736 16908 7742
rect 16856 7678 16908 7684
rect 16580 7600 16632 7606
rect 16580 7542 16632 7548
rect 16592 7130 16620 7542
rect 16580 7124 16632 7130
rect 16580 7066 16632 7072
rect 16488 6852 16540 6858
rect 16488 6794 16540 6800
rect 16500 5226 16528 6794
rect 16592 6722 16620 7066
rect 16868 6858 16896 7678
rect 16856 6852 16908 6858
rect 16856 6794 16908 6800
rect 16580 6716 16632 6722
rect 16580 6658 16632 6664
rect 16488 5220 16540 5226
rect 16488 5162 16540 5168
rect 16396 3996 16448 4002
rect 16396 3938 16448 3944
rect 14684 3692 14980 3712
rect 14740 3690 14764 3692
rect 14820 3690 14844 3692
rect 14900 3690 14924 3692
rect 14762 3638 14764 3690
rect 14826 3638 14838 3690
rect 14900 3638 14902 3690
rect 14740 3636 14764 3638
rect 14820 3636 14844 3638
rect 14900 3636 14924 3638
rect 14684 3616 14980 3636
rect 14684 2604 14980 2624
rect 14740 2602 14764 2604
rect 14820 2602 14844 2604
rect 14900 2602 14924 2604
rect 14762 2550 14764 2602
rect 14826 2550 14838 2602
rect 14900 2550 14902 2602
rect 14740 2548 14764 2550
rect 14820 2548 14844 2550
rect 14900 2548 14924 2550
rect 14684 2528 14980 2548
rect 13912 1956 13964 1962
rect 13912 1898 13964 1904
rect 16960 1214 16988 9718
rect 16948 1208 17000 1214
rect 16948 1150 17000 1156
rect 17236 97 17264 10942
rect 17328 10666 17356 11010
rect 17512 11006 17540 11554
rect 17500 11000 17552 11006
rect 17500 10942 17552 10948
rect 17316 10660 17368 10666
rect 17316 10602 17368 10608
rect 17512 10122 17540 10942
rect 17500 10116 17552 10122
rect 17500 10058 17552 10064
rect 17788 10054 17816 17182
rect 17960 17188 18012 17194
rect 17960 17130 18012 17136
rect 18616 17058 18644 17334
rect 18604 17052 18656 17058
rect 18604 16994 18656 17000
rect 18052 16848 18104 16854
rect 18052 16790 18104 16796
rect 18064 16650 18092 16790
rect 18052 16644 18104 16650
rect 18052 16586 18104 16592
rect 18116 16204 18412 16224
rect 18172 16202 18196 16204
rect 18252 16202 18276 16204
rect 18332 16202 18356 16204
rect 18194 16150 18196 16202
rect 18258 16150 18270 16202
rect 18332 16150 18334 16202
rect 18172 16148 18196 16150
rect 18252 16148 18276 16150
rect 18332 16148 18356 16150
rect 18116 16128 18412 16148
rect 18116 15116 18412 15136
rect 18172 15114 18196 15116
rect 18252 15114 18276 15116
rect 18332 15114 18356 15116
rect 18194 15062 18196 15114
rect 18258 15062 18270 15114
rect 18332 15062 18334 15114
rect 18172 15060 18196 15062
rect 18252 15060 18276 15062
rect 18332 15060 18356 15062
rect 18116 15040 18412 15060
rect 18512 14400 18564 14406
rect 18512 14342 18564 14348
rect 18116 14028 18412 14048
rect 18172 14026 18196 14028
rect 18252 14026 18276 14028
rect 18332 14026 18356 14028
rect 18194 13974 18196 14026
rect 18258 13974 18270 14026
rect 18332 13974 18334 14026
rect 18172 13972 18196 13974
rect 18252 13972 18276 13974
rect 18332 13972 18356 13974
rect 18116 13952 18412 13972
rect 18524 13794 18552 14342
rect 18708 13930 18736 17454
rect 18800 15222 18828 19034
rect 19062 18720 19118 18729
rect 19062 18655 19118 18664
rect 18880 17664 18932 17670
rect 18880 17606 18932 17612
rect 18892 16514 18920 17606
rect 18880 16508 18932 16514
rect 18880 16450 18932 16456
rect 19076 16106 19104 18655
rect 19168 17890 19196 22176
rect 19246 21032 19302 21041
rect 19246 20967 19302 20976
rect 19260 19030 19288 20967
rect 19720 19930 19748 22176
rect 19720 19902 20024 19930
rect 19340 19772 19392 19778
rect 19340 19714 19392 19720
rect 19708 19772 19760 19778
rect 19708 19714 19760 19720
rect 19248 19024 19300 19030
rect 19248 18966 19300 18972
rect 19352 18078 19380 19714
rect 19524 18684 19576 18690
rect 19524 18626 19576 18632
rect 19536 18214 19564 18626
rect 19720 18622 19748 19714
rect 19800 19704 19852 19710
rect 19800 19646 19852 19652
rect 19890 19672 19946 19681
rect 19812 18690 19840 19646
rect 19890 19607 19946 19616
rect 19800 18684 19852 18690
rect 19800 18626 19852 18632
rect 19708 18616 19760 18622
rect 19708 18558 19760 18564
rect 19720 18282 19840 18298
rect 19904 18282 19932 19607
rect 19708 18276 19840 18282
rect 19760 18270 19840 18276
rect 19708 18218 19760 18224
rect 19524 18208 19576 18214
rect 19524 18150 19576 18156
rect 19708 18140 19760 18146
rect 19708 18082 19760 18088
rect 19340 18072 19392 18078
rect 19340 18014 19392 18020
rect 19616 18072 19668 18078
rect 19616 18014 19668 18020
rect 19524 17936 19576 17942
rect 19168 17862 19472 17890
rect 19524 17878 19576 17884
rect 19248 16984 19300 16990
rect 19246 16952 19248 16961
rect 19340 16984 19392 16990
rect 19300 16952 19302 16961
rect 19340 16926 19392 16932
rect 19246 16887 19302 16896
rect 19064 16100 19116 16106
rect 19064 16042 19116 16048
rect 19352 16038 19380 16926
rect 19340 16032 19392 16038
rect 19340 15974 19392 15980
rect 19156 15896 19208 15902
rect 19156 15838 19208 15844
rect 19168 15494 19196 15838
rect 19156 15488 19208 15494
rect 19156 15430 19208 15436
rect 19340 15420 19392 15426
rect 19340 15362 19392 15368
rect 18788 15216 18840 15222
rect 18788 15158 18840 15164
rect 19352 14950 19380 15362
rect 19340 14944 19392 14950
rect 19340 14886 19392 14892
rect 19154 14232 19210 14241
rect 19154 14167 19210 14176
rect 18696 13924 18748 13930
rect 18696 13866 18748 13872
rect 18512 13788 18564 13794
rect 18512 13730 18564 13736
rect 18788 13720 18840 13726
rect 18788 13662 18840 13668
rect 17868 13584 17920 13590
rect 17868 13526 17920 13532
rect 17880 11074 17908 13526
rect 18800 13318 18828 13662
rect 18788 13312 18840 13318
rect 18788 13254 18840 13260
rect 18696 13244 18748 13250
rect 18696 13186 18748 13192
rect 18116 12940 18412 12960
rect 18172 12938 18196 12940
rect 18252 12938 18276 12940
rect 18332 12938 18356 12940
rect 18194 12886 18196 12938
rect 18258 12886 18270 12938
rect 18332 12886 18334 12938
rect 18172 12884 18196 12886
rect 18252 12884 18276 12886
rect 18332 12884 18356 12886
rect 18116 12864 18412 12884
rect 17960 12496 18012 12502
rect 17960 12438 18012 12444
rect 17972 12298 18000 12438
rect 17960 12292 18012 12298
rect 17960 12234 18012 12240
rect 17960 12156 18012 12162
rect 17960 12098 18012 12104
rect 17972 11754 18000 12098
rect 18116 11852 18412 11872
rect 18172 11850 18196 11852
rect 18252 11850 18276 11852
rect 18332 11850 18356 11852
rect 18194 11798 18196 11850
rect 18258 11798 18270 11850
rect 18332 11798 18334 11850
rect 18172 11796 18196 11798
rect 18252 11796 18276 11798
rect 18332 11796 18356 11798
rect 18116 11776 18412 11796
rect 17960 11748 18012 11754
rect 17960 11690 18012 11696
rect 17868 11068 17920 11074
rect 17868 11010 17920 11016
rect 17776 10048 17828 10054
rect 17776 9990 17828 9996
rect 17880 9034 17908 11010
rect 18116 10764 18412 10784
rect 18172 10762 18196 10764
rect 18252 10762 18276 10764
rect 18332 10762 18356 10764
rect 18194 10710 18196 10762
rect 18258 10710 18270 10762
rect 18332 10710 18334 10762
rect 18172 10708 18196 10710
rect 18252 10708 18276 10710
rect 18332 10708 18356 10710
rect 18116 10688 18412 10708
rect 18708 10666 18736 13186
rect 18880 12836 18932 12842
rect 18880 12778 18932 12784
rect 18788 11408 18840 11414
rect 18788 11350 18840 11356
rect 18800 11210 18828 11350
rect 18788 11204 18840 11210
rect 18788 11146 18840 11152
rect 18696 10660 18748 10666
rect 18696 10602 18748 10608
rect 18052 10388 18104 10394
rect 18052 10330 18104 10336
rect 18064 10122 18092 10330
rect 18052 10116 18104 10122
rect 18052 10058 18104 10064
rect 18512 9980 18564 9986
rect 18512 9922 18564 9928
rect 18116 9676 18412 9696
rect 18172 9674 18196 9676
rect 18252 9674 18276 9676
rect 18332 9674 18356 9676
rect 18194 9622 18196 9674
rect 18258 9622 18270 9674
rect 18332 9622 18334 9674
rect 18172 9620 18196 9622
rect 18252 9620 18276 9622
rect 18332 9620 18356 9622
rect 18116 9600 18412 9620
rect 17960 9232 18012 9238
rect 17960 9174 18012 9180
rect 17868 9028 17920 9034
rect 17868 8970 17920 8976
rect 17592 7736 17644 7742
rect 17592 7678 17644 7684
rect 17604 7402 17632 7678
rect 17592 7396 17644 7402
rect 17592 7338 17644 7344
rect 17880 3633 17908 8970
rect 17972 6858 18000 9174
rect 18524 8966 18552 9922
rect 18696 9436 18748 9442
rect 18696 9378 18748 9384
rect 18512 8960 18564 8966
rect 18512 8902 18564 8908
rect 18116 8588 18412 8608
rect 18172 8586 18196 8588
rect 18252 8586 18276 8588
rect 18332 8586 18356 8588
rect 18194 8534 18196 8586
rect 18258 8534 18270 8586
rect 18332 8534 18334 8586
rect 18172 8532 18196 8534
rect 18252 8532 18276 8534
rect 18332 8532 18356 8534
rect 18116 8512 18412 8532
rect 18524 7946 18552 8902
rect 18052 7940 18104 7946
rect 18052 7882 18104 7888
rect 18512 7940 18564 7946
rect 18512 7882 18564 7888
rect 18064 7742 18092 7882
rect 18052 7736 18104 7742
rect 18052 7678 18104 7684
rect 18116 7500 18412 7520
rect 18172 7498 18196 7500
rect 18252 7498 18276 7500
rect 18332 7498 18356 7500
rect 18194 7446 18196 7498
rect 18258 7446 18270 7498
rect 18332 7446 18334 7498
rect 18172 7444 18196 7446
rect 18252 7444 18276 7446
rect 18332 7444 18356 7446
rect 18116 7424 18412 7444
rect 17960 6852 18012 6858
rect 17960 6794 18012 6800
rect 17972 6518 18000 6794
rect 18512 6784 18564 6790
rect 18512 6726 18564 6732
rect 17960 6512 18012 6518
rect 18524 6489 18552 6726
rect 18604 6580 18656 6586
rect 18604 6522 18656 6528
rect 17960 6454 18012 6460
rect 18510 6480 18566 6489
rect 18116 6412 18412 6432
rect 18510 6415 18566 6424
rect 18172 6410 18196 6412
rect 18252 6410 18276 6412
rect 18332 6410 18356 6412
rect 18194 6358 18196 6410
rect 18258 6358 18270 6410
rect 18332 6358 18334 6410
rect 18172 6356 18196 6358
rect 18252 6356 18276 6358
rect 18332 6356 18356 6358
rect 18116 6336 18412 6356
rect 18616 5537 18644 6522
rect 18602 5528 18658 5537
rect 18602 5463 18658 5472
rect 18116 5324 18412 5344
rect 18172 5322 18196 5324
rect 18252 5322 18276 5324
rect 18332 5322 18356 5324
rect 18194 5270 18196 5322
rect 18258 5270 18270 5322
rect 18332 5270 18334 5322
rect 18172 5268 18196 5270
rect 18252 5268 18276 5270
rect 18332 5268 18356 5270
rect 18116 5248 18412 5268
rect 17960 5220 18012 5226
rect 17960 5162 18012 5168
rect 17972 4585 18000 5162
rect 17958 4576 18014 4585
rect 17958 4511 18014 4520
rect 18116 4236 18412 4256
rect 18172 4234 18196 4236
rect 18252 4234 18276 4236
rect 18332 4234 18356 4236
rect 18194 4182 18196 4234
rect 18258 4182 18270 4234
rect 18332 4182 18334 4234
rect 18172 4180 18196 4182
rect 18252 4180 18276 4182
rect 18332 4180 18356 4182
rect 18116 4160 18412 4180
rect 17866 3624 17922 3633
rect 17866 3559 17922 3568
rect 18116 3148 18412 3168
rect 18172 3146 18196 3148
rect 18252 3146 18276 3148
rect 18332 3146 18356 3148
rect 18194 3094 18196 3146
rect 18258 3094 18270 3146
rect 18332 3094 18334 3146
rect 18172 3092 18196 3094
rect 18252 3092 18276 3094
rect 18332 3092 18356 3094
rect 18116 3072 18412 3092
rect 18116 2060 18412 2080
rect 18172 2058 18196 2060
rect 18252 2058 18276 2060
rect 18332 2058 18356 2060
rect 18194 2006 18196 2058
rect 18258 2006 18270 2058
rect 18332 2006 18334 2058
rect 18172 2004 18196 2006
rect 18252 2004 18276 2006
rect 18332 2004 18356 2006
rect 18116 1984 18412 2004
rect 17960 1956 18012 1962
rect 17960 1898 18012 1904
rect 17972 1457 18000 1898
rect 18708 1865 18736 9378
rect 18786 9336 18842 9345
rect 18786 9271 18842 9280
rect 18800 3225 18828 9271
rect 18786 3216 18842 3225
rect 18786 3151 18842 3160
rect 18694 1856 18750 1865
rect 18694 1791 18750 1800
rect 17958 1448 18014 1457
rect 17958 1383 18014 1392
rect 17960 1208 18012 1214
rect 17960 1150 18012 1156
rect 17972 913 18000 1150
rect 17958 904 18014 913
rect 17958 839 18014 848
rect 18892 505 18920 12778
rect 19064 12632 19116 12638
rect 19064 12574 19116 12580
rect 19076 12298 19104 12574
rect 19064 12292 19116 12298
rect 19064 12234 19116 12240
rect 18972 11952 19024 11958
rect 18972 11894 19024 11900
rect 18984 2273 19012 11894
rect 19168 11754 19196 14167
rect 19248 13244 19300 13250
rect 19248 13186 19300 13192
rect 19260 12337 19288 13186
rect 19246 12328 19302 12337
rect 19246 12263 19302 12272
rect 19156 11748 19208 11754
rect 19156 11690 19208 11696
rect 19444 11210 19472 17862
rect 19536 14898 19564 17878
rect 19628 16582 19656 18014
rect 19616 16576 19668 16582
rect 19616 16518 19668 16524
rect 19536 14870 19656 14898
rect 19524 14808 19576 14814
rect 19524 14750 19576 14756
rect 19536 14406 19564 14750
rect 19524 14400 19576 14406
rect 19524 14342 19576 14348
rect 19432 11204 19484 11210
rect 19432 11146 19484 11152
rect 19248 10864 19300 10870
rect 19248 10806 19300 10812
rect 19260 10546 19288 10806
rect 19168 10530 19288 10546
rect 19156 10524 19288 10530
rect 19208 10518 19288 10524
rect 19156 10466 19208 10472
rect 19156 10320 19208 10326
rect 19156 10262 19208 10268
rect 19062 10016 19118 10025
rect 19062 9951 19118 9960
rect 19076 9374 19104 9951
rect 19168 9578 19196 10262
rect 19260 10122 19288 10518
rect 19248 10116 19300 10122
rect 19248 10058 19300 10064
rect 19156 9572 19208 9578
rect 19156 9514 19208 9520
rect 19432 9436 19484 9442
rect 19432 9378 19484 9384
rect 19064 9368 19116 9374
rect 19064 9310 19116 9316
rect 19444 8898 19472 9378
rect 19432 8892 19484 8898
rect 19432 8834 19484 8840
rect 19444 7946 19472 8834
rect 19628 8762 19656 14870
rect 19720 13930 19748 18082
rect 19812 15986 19840 18270
rect 19892 18276 19944 18282
rect 19892 18218 19944 18224
rect 19892 17936 19944 17942
rect 19892 17878 19944 17884
rect 19904 16938 19932 17878
rect 19996 17040 20024 19902
rect 20076 18820 20128 18826
rect 20076 18762 20128 18768
rect 20088 17194 20116 18762
rect 20272 17942 20300 22176
rect 20626 20624 20682 20633
rect 20626 20559 20682 20568
rect 20640 19914 20668 20559
rect 20718 20080 20774 20089
rect 20718 20015 20774 20024
rect 20628 19908 20680 19914
rect 20628 19850 20680 19856
rect 20732 18826 20760 20015
rect 20720 18820 20772 18826
rect 20720 18762 20772 18768
rect 20350 18312 20406 18321
rect 20350 18247 20406 18256
rect 20260 17936 20312 17942
rect 20260 17878 20312 17884
rect 20364 17738 20392 18247
rect 20824 18162 20852 22176
rect 20994 19264 21050 19273
rect 20994 19199 21050 19208
rect 20548 18134 20852 18162
rect 20444 17936 20496 17942
rect 20444 17878 20496 17884
rect 20352 17732 20404 17738
rect 20352 17674 20404 17680
rect 20168 17596 20220 17602
rect 20168 17538 20220 17544
rect 20076 17188 20128 17194
rect 20076 17130 20128 17136
rect 20180 17058 20208 17538
rect 20352 17188 20404 17194
rect 20352 17130 20404 17136
rect 20168 17052 20220 17058
rect 19996 17012 20116 17040
rect 19904 16910 20024 16938
rect 19812 15958 19932 15986
rect 19800 15896 19852 15902
rect 19800 15838 19852 15844
rect 19812 14882 19840 15838
rect 19800 14876 19852 14882
rect 19800 14818 19852 14824
rect 19708 13924 19760 13930
rect 19708 13866 19760 13872
rect 19708 13720 19760 13726
rect 19708 13662 19760 13668
rect 19720 12881 19748 13662
rect 19706 12872 19762 12881
rect 19706 12807 19762 12816
rect 19904 12774 19932 15958
rect 19892 12768 19944 12774
rect 19892 12710 19944 12716
rect 19996 12298 20024 16910
rect 20088 16836 20116 17012
rect 20168 16994 20220 17000
rect 20088 16808 20300 16836
rect 20168 16644 20220 16650
rect 20168 16586 20220 16592
rect 20180 16417 20208 16586
rect 20166 16408 20222 16417
rect 20166 16343 20222 16352
rect 20076 16032 20128 16038
rect 20074 16000 20076 16009
rect 20128 16000 20130 16009
rect 20074 15935 20130 15944
rect 20074 13280 20130 13289
rect 20074 13215 20130 13224
rect 20168 13244 20220 13250
rect 20088 12842 20116 13215
rect 20168 13186 20220 13192
rect 20076 12836 20128 12842
rect 20076 12778 20128 12784
rect 19984 12292 20036 12298
rect 19984 12234 20036 12240
rect 19892 12156 19944 12162
rect 19892 12098 19944 12104
rect 19904 11521 19932 12098
rect 20180 11929 20208 13186
rect 20272 12298 20300 16808
rect 20260 12292 20312 12298
rect 20260 12234 20312 12240
rect 20166 11920 20222 11929
rect 20166 11855 20222 11864
rect 20260 11544 20312 11550
rect 19890 11512 19946 11521
rect 20260 11486 20312 11492
rect 19890 11447 19946 11456
rect 20272 11142 20300 11486
rect 20260 11136 20312 11142
rect 20260 11078 20312 11084
rect 20364 10666 20392 17130
rect 20456 16961 20484 17878
rect 20442 16952 20498 16961
rect 20442 16887 20498 16896
rect 20444 16848 20496 16854
rect 20444 16790 20496 16796
rect 20456 16514 20484 16790
rect 20444 16508 20496 16514
rect 20444 16450 20496 16456
rect 20442 15592 20498 15601
rect 20442 15527 20498 15536
rect 20456 15018 20484 15527
rect 20444 15012 20496 15018
rect 20444 14954 20496 14960
rect 20442 14640 20498 14649
rect 20442 14575 20498 14584
rect 20456 13930 20484 14575
rect 20444 13924 20496 13930
rect 20444 13866 20496 13872
rect 20548 13386 20576 18134
rect 20628 18072 20680 18078
rect 20628 18014 20680 18020
rect 20536 13380 20588 13386
rect 20536 13322 20588 13328
rect 20640 13114 20668 18014
rect 20812 17936 20864 17942
rect 20812 17878 20864 17884
rect 20902 17904 20958 17913
rect 20718 13688 20774 13697
rect 20718 13623 20774 13632
rect 20732 13386 20760 13623
rect 20720 13380 20772 13386
rect 20720 13322 20772 13328
rect 20628 13108 20680 13114
rect 20628 13050 20680 13056
rect 20628 12768 20680 12774
rect 20628 12710 20680 12716
rect 20444 12156 20496 12162
rect 20444 12098 20496 12104
rect 20456 10977 20484 12098
rect 20536 11068 20588 11074
rect 20536 11010 20588 11016
rect 20442 10968 20498 10977
rect 20442 10903 20498 10912
rect 20352 10660 20404 10666
rect 20352 10602 20404 10608
rect 20548 10569 20576 11010
rect 20534 10560 20590 10569
rect 19708 10524 19760 10530
rect 20534 10495 20590 10504
rect 19708 10466 19760 10472
rect 19720 9986 19748 10466
rect 20260 10456 20312 10462
rect 20260 10398 20312 10404
rect 19708 9980 19760 9986
rect 19708 9922 19760 9928
rect 19720 9034 19748 9922
rect 20272 9617 20300 10398
rect 20536 9980 20588 9986
rect 20536 9922 20588 9928
rect 20258 9608 20314 9617
rect 20258 9543 20314 9552
rect 20548 9209 20576 9922
rect 20534 9200 20590 9209
rect 20534 9135 20590 9144
rect 19708 9028 19760 9034
rect 19708 8970 19760 8976
rect 19984 8892 20036 8898
rect 19984 8834 20036 8840
rect 20536 8892 20588 8898
rect 20536 8834 20588 8840
rect 19616 8756 19668 8762
rect 19616 8698 19668 8704
rect 19996 8257 20024 8834
rect 20548 8665 20576 8834
rect 20534 8656 20590 8665
rect 20534 8591 20590 8600
rect 20640 8490 20668 12710
rect 20628 8484 20680 8490
rect 20628 8426 20680 8432
rect 20260 8280 20312 8286
rect 19982 8248 20038 8257
rect 20260 8222 20312 8228
rect 19982 8183 20038 8192
rect 19432 7940 19484 7946
rect 19432 7882 19484 7888
rect 20272 7849 20300 8222
rect 20258 7840 20314 7849
rect 19984 7804 20036 7810
rect 20258 7775 20314 7784
rect 20536 7804 20588 7810
rect 19984 7746 20036 7752
rect 20536 7746 20588 7752
rect 19996 6897 20024 7746
rect 20548 7305 20576 7746
rect 20534 7296 20590 7305
rect 20534 7231 20590 7240
rect 19982 6888 20038 6897
rect 19982 6823 20038 6832
rect 20536 6716 20588 6722
rect 20536 6658 20588 6664
rect 20548 5945 20576 6658
rect 20720 6512 20772 6518
rect 20720 6454 20772 6460
rect 20732 6314 20760 6454
rect 20720 6308 20772 6314
rect 20720 6250 20772 6256
rect 20534 5936 20590 5945
rect 20534 5871 20590 5880
rect 20536 5628 20588 5634
rect 20536 5570 20588 5576
rect 20548 4993 20576 5570
rect 20534 4984 20590 4993
rect 20534 4919 20590 4928
rect 20824 4682 20852 17878
rect 20902 17839 20958 17848
rect 20916 17738 20944 17839
rect 20904 17732 20956 17738
rect 20904 17674 20956 17680
rect 21008 15562 21036 19199
rect 21180 18480 21232 18486
rect 21180 18422 21232 18428
rect 20996 15556 21048 15562
rect 20996 15498 21048 15504
rect 20902 15048 20958 15057
rect 20902 14983 20958 14992
rect 20916 14474 20944 14983
rect 20904 14468 20956 14474
rect 20904 14410 20956 14416
rect 21192 9034 21220 18422
rect 21376 18078 21404 22176
rect 21928 18146 21956 22176
rect 21916 18140 21968 18146
rect 21916 18082 21968 18088
rect 21364 18072 21416 18078
rect 21364 18014 21416 18020
rect 22480 17942 22508 22176
rect 22468 17936 22520 17942
rect 22468 17878 22520 17884
rect 21730 17360 21786 17369
rect 21730 17295 21732 17304
rect 21784 17295 21786 17304
rect 21732 17266 21784 17272
rect 21180 9028 21232 9034
rect 21180 8970 21232 8976
rect 20812 4676 20864 4682
rect 20812 4618 20864 4624
rect 20536 4540 20588 4546
rect 20536 4482 20588 4488
rect 20548 4177 20576 4482
rect 20534 4168 20590 4177
rect 20534 4103 20590 4112
rect 19064 3996 19116 4002
rect 19064 3938 19116 3944
rect 19076 2817 19104 3938
rect 19062 2808 19118 2817
rect 19062 2743 19118 2752
rect 18970 2264 19026 2273
rect 18970 2199 19026 2208
rect 18878 496 18934 505
rect 18878 431 18934 440
rect 17222 88 17278 97
rect 17222 23 17278 32
<< via2 >>
rect 18878 22336 18934 22392
rect 4066 17032 4122 17088
rect 4388 19466 4444 19468
rect 4468 19466 4524 19468
rect 4548 19466 4604 19468
rect 4628 19466 4684 19468
rect 4388 19414 4414 19466
rect 4414 19414 4444 19466
rect 4468 19414 4478 19466
rect 4478 19414 4524 19466
rect 4548 19414 4594 19466
rect 4594 19414 4604 19466
rect 4628 19414 4658 19466
rect 4658 19414 4684 19466
rect 4388 19412 4444 19414
rect 4468 19412 4524 19414
rect 4548 19412 4604 19414
rect 4628 19412 4684 19414
rect 4388 18378 4444 18380
rect 4468 18378 4524 18380
rect 4548 18378 4604 18380
rect 4628 18378 4684 18380
rect 4388 18326 4414 18378
rect 4414 18326 4444 18378
rect 4468 18326 4478 18378
rect 4478 18326 4524 18378
rect 4548 18326 4594 18378
rect 4594 18326 4604 18378
rect 4628 18326 4658 18378
rect 4658 18326 4684 18378
rect 4388 18324 4444 18326
rect 4468 18324 4524 18326
rect 4548 18324 4604 18326
rect 4628 18324 4684 18326
rect 4388 17290 4444 17292
rect 4468 17290 4524 17292
rect 4548 17290 4604 17292
rect 4628 17290 4684 17292
rect 4388 17238 4414 17290
rect 4414 17238 4444 17290
rect 4468 17238 4478 17290
rect 4478 17238 4524 17290
rect 4548 17238 4594 17290
rect 4594 17238 4604 17290
rect 4628 17238 4658 17290
rect 4658 17238 4684 17290
rect 4388 17236 4444 17238
rect 4468 17236 4524 17238
rect 4548 17236 4604 17238
rect 4628 17236 4684 17238
rect 4388 16202 4444 16204
rect 4468 16202 4524 16204
rect 4548 16202 4604 16204
rect 4628 16202 4684 16204
rect 4388 16150 4414 16202
rect 4414 16150 4444 16202
rect 4468 16150 4478 16202
rect 4478 16150 4524 16202
rect 4548 16150 4594 16202
rect 4594 16150 4604 16202
rect 4628 16150 4658 16202
rect 4658 16150 4684 16202
rect 4388 16148 4444 16150
rect 4468 16148 4524 16150
rect 4548 16148 4604 16150
rect 4628 16148 4684 16150
rect 4388 15114 4444 15116
rect 4468 15114 4524 15116
rect 4548 15114 4604 15116
rect 4628 15114 4684 15116
rect 4388 15062 4414 15114
rect 4414 15062 4444 15114
rect 4468 15062 4478 15114
rect 4478 15062 4524 15114
rect 4548 15062 4594 15114
rect 4594 15062 4604 15114
rect 4628 15062 4658 15114
rect 4658 15062 4684 15114
rect 4388 15060 4444 15062
rect 4468 15060 4524 15062
rect 4548 15060 4604 15062
rect 4628 15060 4684 15062
rect 4388 14026 4444 14028
rect 4468 14026 4524 14028
rect 4548 14026 4604 14028
rect 4628 14026 4684 14028
rect 4388 13974 4414 14026
rect 4414 13974 4444 14026
rect 4468 13974 4478 14026
rect 4478 13974 4524 14026
rect 4548 13974 4594 14026
rect 4594 13974 4604 14026
rect 4628 13974 4658 14026
rect 4658 13974 4684 14026
rect 4388 13972 4444 13974
rect 4468 13972 4524 13974
rect 4548 13972 4604 13974
rect 4628 13972 4684 13974
rect 4388 12938 4444 12940
rect 4468 12938 4524 12940
rect 4548 12938 4604 12940
rect 4628 12938 4684 12940
rect 4388 12886 4414 12938
rect 4414 12886 4444 12938
rect 4468 12886 4478 12938
rect 4478 12886 4524 12938
rect 4548 12886 4594 12938
rect 4594 12886 4604 12938
rect 4628 12886 4658 12938
rect 4658 12886 4684 12938
rect 4388 12884 4444 12886
rect 4468 12884 4524 12886
rect 4548 12884 4604 12886
rect 4628 12884 4684 12886
rect 4388 11850 4444 11852
rect 4468 11850 4524 11852
rect 4548 11850 4604 11852
rect 4628 11850 4684 11852
rect 4388 11798 4414 11850
rect 4414 11798 4444 11850
rect 4468 11798 4478 11850
rect 4478 11798 4524 11850
rect 4548 11798 4594 11850
rect 4594 11798 4604 11850
rect 4628 11798 4658 11850
rect 4658 11798 4684 11850
rect 4388 11796 4444 11798
rect 4468 11796 4524 11798
rect 4548 11796 4604 11798
rect 4628 11796 4684 11798
rect 7820 20010 7876 20012
rect 7900 20010 7956 20012
rect 7980 20010 8036 20012
rect 8060 20010 8116 20012
rect 7820 19958 7846 20010
rect 7846 19958 7876 20010
rect 7900 19958 7910 20010
rect 7910 19958 7956 20010
rect 7980 19958 8026 20010
rect 8026 19958 8036 20010
rect 8060 19958 8090 20010
rect 8090 19958 8116 20010
rect 7820 19956 7876 19958
rect 7900 19956 7956 19958
rect 7980 19956 8036 19958
rect 8060 19956 8116 19958
rect 7820 18922 7876 18924
rect 7900 18922 7956 18924
rect 7980 18922 8036 18924
rect 8060 18922 8116 18924
rect 7820 18870 7846 18922
rect 7846 18870 7876 18922
rect 7900 18870 7910 18922
rect 7910 18870 7956 18922
rect 7980 18870 8026 18922
rect 8026 18870 8036 18922
rect 8060 18870 8090 18922
rect 8090 18870 8116 18922
rect 7820 18868 7876 18870
rect 7900 18868 7956 18870
rect 7980 18868 8036 18870
rect 8060 18868 8116 18870
rect 7820 17834 7876 17836
rect 7900 17834 7956 17836
rect 7980 17834 8036 17836
rect 8060 17834 8116 17836
rect 7820 17782 7846 17834
rect 7846 17782 7876 17834
rect 7900 17782 7910 17834
rect 7910 17782 7956 17834
rect 7980 17782 8026 17834
rect 8026 17782 8036 17834
rect 8060 17782 8090 17834
rect 8090 17782 8116 17834
rect 7820 17780 7876 17782
rect 7900 17780 7956 17782
rect 7980 17780 8036 17782
rect 8060 17780 8116 17782
rect 7820 16746 7876 16748
rect 7900 16746 7956 16748
rect 7980 16746 8036 16748
rect 8060 16746 8116 16748
rect 7820 16694 7846 16746
rect 7846 16694 7876 16746
rect 7900 16694 7910 16746
rect 7910 16694 7956 16746
rect 7980 16694 8026 16746
rect 8026 16694 8036 16746
rect 8060 16694 8090 16746
rect 8090 16694 8116 16746
rect 7820 16692 7876 16694
rect 7900 16692 7956 16694
rect 7980 16692 8036 16694
rect 8060 16692 8116 16694
rect 7820 15658 7876 15660
rect 7900 15658 7956 15660
rect 7980 15658 8036 15660
rect 8060 15658 8116 15660
rect 7820 15606 7846 15658
rect 7846 15606 7876 15658
rect 7900 15606 7910 15658
rect 7910 15606 7956 15658
rect 7980 15606 8026 15658
rect 8026 15606 8036 15658
rect 8060 15606 8090 15658
rect 8090 15606 8116 15658
rect 7820 15604 7876 15606
rect 7900 15604 7956 15606
rect 7980 15604 8036 15606
rect 8060 15604 8116 15606
rect 7820 14570 7876 14572
rect 7900 14570 7956 14572
rect 7980 14570 8036 14572
rect 8060 14570 8116 14572
rect 7820 14518 7846 14570
rect 7846 14518 7876 14570
rect 7900 14518 7910 14570
rect 7910 14518 7956 14570
rect 7980 14518 8026 14570
rect 8026 14518 8036 14570
rect 8060 14518 8090 14570
rect 8090 14518 8116 14570
rect 7820 14516 7876 14518
rect 7900 14516 7956 14518
rect 7980 14516 8036 14518
rect 8060 14516 8116 14518
rect 7820 13482 7876 13484
rect 7900 13482 7956 13484
rect 7980 13482 8036 13484
rect 8060 13482 8116 13484
rect 7820 13430 7846 13482
rect 7846 13430 7876 13482
rect 7900 13430 7910 13482
rect 7910 13430 7956 13482
rect 7980 13430 8026 13482
rect 8026 13430 8036 13482
rect 8060 13430 8090 13482
rect 8090 13430 8116 13482
rect 7820 13428 7876 13430
rect 7900 13428 7956 13430
rect 7980 13428 8036 13430
rect 8060 13428 8116 13430
rect 9034 18120 9090 18176
rect 7820 12394 7876 12396
rect 7900 12394 7956 12396
rect 7980 12394 8036 12396
rect 8060 12394 8116 12396
rect 7820 12342 7846 12394
rect 7846 12342 7876 12394
rect 7900 12342 7910 12394
rect 7910 12342 7956 12394
rect 7980 12342 8026 12394
rect 8026 12342 8036 12394
rect 8060 12342 8090 12394
rect 8090 12342 8116 12394
rect 7820 12340 7876 12342
rect 7900 12340 7956 12342
rect 7980 12340 8036 12342
rect 8060 12340 8116 12342
rect 4388 10762 4444 10764
rect 4468 10762 4524 10764
rect 4548 10762 4604 10764
rect 4628 10762 4684 10764
rect 4388 10710 4414 10762
rect 4414 10710 4444 10762
rect 4468 10710 4478 10762
rect 4478 10710 4524 10762
rect 4548 10710 4594 10762
rect 4594 10710 4604 10762
rect 4628 10710 4658 10762
rect 4658 10710 4684 10762
rect 4388 10708 4444 10710
rect 4468 10708 4524 10710
rect 4548 10708 4604 10710
rect 4628 10708 4684 10710
rect 7820 11306 7876 11308
rect 7900 11306 7956 11308
rect 7980 11306 8036 11308
rect 8060 11306 8116 11308
rect 7820 11254 7846 11306
rect 7846 11254 7876 11306
rect 7900 11254 7910 11306
rect 7910 11254 7956 11306
rect 7980 11254 8026 11306
rect 8026 11254 8036 11306
rect 8060 11254 8090 11306
rect 8090 11254 8116 11306
rect 7820 11252 7876 11254
rect 7900 11252 7956 11254
rect 7980 11252 8036 11254
rect 8060 11252 8116 11254
rect 10230 19072 10286 19128
rect 11252 19466 11308 19468
rect 11332 19466 11388 19468
rect 11412 19466 11468 19468
rect 11492 19466 11548 19468
rect 11252 19414 11278 19466
rect 11278 19414 11308 19466
rect 11332 19414 11342 19466
rect 11342 19414 11388 19466
rect 11412 19414 11458 19466
rect 11458 19414 11468 19466
rect 11492 19414 11522 19466
rect 11522 19414 11548 19466
rect 11252 19412 11308 19414
rect 11332 19412 11388 19414
rect 11412 19412 11468 19414
rect 11492 19412 11548 19414
rect 10782 18664 10838 18720
rect 10414 18120 10470 18176
rect 9770 16896 9826 16952
rect 7820 10218 7876 10220
rect 7900 10218 7956 10220
rect 7980 10218 8036 10220
rect 8060 10218 8116 10220
rect 7820 10166 7846 10218
rect 7846 10166 7876 10218
rect 7900 10166 7910 10218
rect 7910 10166 7956 10218
rect 7980 10166 8026 10218
rect 8026 10166 8036 10218
rect 8060 10166 8090 10218
rect 8090 10166 8116 10218
rect 7820 10164 7876 10166
rect 7900 10164 7956 10166
rect 7980 10164 8036 10166
rect 8060 10164 8116 10166
rect 4388 9674 4444 9676
rect 4468 9674 4524 9676
rect 4548 9674 4604 9676
rect 4628 9674 4684 9676
rect 4388 9622 4414 9674
rect 4414 9622 4444 9674
rect 4468 9622 4478 9674
rect 4478 9622 4524 9674
rect 4548 9622 4594 9674
rect 4594 9622 4604 9674
rect 4628 9622 4658 9674
rect 4658 9622 4684 9674
rect 4388 9620 4444 9622
rect 4468 9620 4524 9622
rect 4548 9620 4604 9622
rect 4628 9620 4684 9622
rect 4388 8586 4444 8588
rect 4468 8586 4524 8588
rect 4548 8586 4604 8588
rect 4628 8586 4684 8588
rect 4388 8534 4414 8586
rect 4414 8534 4444 8586
rect 4468 8534 4478 8586
rect 4478 8534 4524 8586
rect 4548 8534 4594 8586
rect 4594 8534 4604 8586
rect 4628 8534 4658 8586
rect 4658 8534 4684 8586
rect 4388 8532 4444 8534
rect 4468 8532 4524 8534
rect 4548 8532 4604 8534
rect 4628 8532 4684 8534
rect 7820 9130 7876 9132
rect 7900 9130 7956 9132
rect 7980 9130 8036 9132
rect 8060 9130 8116 9132
rect 7820 9078 7846 9130
rect 7846 9078 7876 9130
rect 7900 9078 7910 9130
rect 7910 9078 7956 9130
rect 7980 9078 8026 9130
rect 8026 9078 8036 9130
rect 8060 9078 8090 9130
rect 8090 9078 8116 9130
rect 7820 9076 7876 9078
rect 7900 9076 7956 9078
rect 7980 9076 8036 9078
rect 8060 9076 8116 9078
rect 7820 8042 7876 8044
rect 7900 8042 7956 8044
rect 7980 8042 8036 8044
rect 8060 8042 8116 8044
rect 7820 7990 7846 8042
rect 7846 7990 7876 8042
rect 7900 7990 7910 8042
rect 7910 7990 7956 8042
rect 7980 7990 8026 8042
rect 8026 7990 8036 8042
rect 8060 7990 8090 8042
rect 8090 7990 8116 8042
rect 7820 7988 7876 7990
rect 7900 7988 7956 7990
rect 7980 7988 8036 7990
rect 8060 7988 8116 7990
rect 4388 7498 4444 7500
rect 4468 7498 4524 7500
rect 4548 7498 4604 7500
rect 4628 7498 4684 7500
rect 4388 7446 4414 7498
rect 4414 7446 4444 7498
rect 4468 7446 4478 7498
rect 4478 7446 4524 7498
rect 4548 7446 4594 7498
rect 4594 7446 4604 7498
rect 4628 7446 4658 7498
rect 4658 7446 4684 7498
rect 4388 7444 4444 7446
rect 4468 7444 4524 7446
rect 4548 7444 4604 7446
rect 4628 7444 4684 7446
rect 7820 6954 7876 6956
rect 7900 6954 7956 6956
rect 7980 6954 8036 6956
rect 8060 6954 8116 6956
rect 7820 6902 7846 6954
rect 7846 6902 7876 6954
rect 7900 6902 7910 6954
rect 7910 6902 7956 6954
rect 7980 6902 8026 6954
rect 8026 6902 8036 6954
rect 8060 6902 8090 6954
rect 8090 6902 8116 6954
rect 7820 6900 7876 6902
rect 7900 6900 7956 6902
rect 7980 6900 8036 6902
rect 8060 6900 8116 6902
rect 10598 18004 10654 18040
rect 10598 17984 10600 18004
rect 10600 17984 10652 18004
rect 10652 17984 10654 18004
rect 11252 18378 11308 18380
rect 11332 18378 11388 18380
rect 11412 18378 11468 18380
rect 11492 18378 11548 18380
rect 11252 18326 11278 18378
rect 11278 18326 11308 18378
rect 11332 18326 11342 18378
rect 11342 18326 11388 18378
rect 11412 18326 11458 18378
rect 11458 18326 11468 18378
rect 11492 18326 11522 18378
rect 11522 18326 11548 18378
rect 11252 18324 11308 18326
rect 11332 18324 11388 18326
rect 11412 18324 11468 18326
rect 11492 18324 11548 18326
rect 11252 17290 11308 17292
rect 11332 17290 11388 17292
rect 11412 17290 11468 17292
rect 11492 17290 11548 17292
rect 11252 17238 11278 17290
rect 11278 17238 11308 17290
rect 11332 17238 11342 17290
rect 11342 17238 11388 17290
rect 11412 17238 11458 17290
rect 11458 17238 11468 17290
rect 11492 17238 11522 17290
rect 11522 17238 11548 17290
rect 11252 17236 11308 17238
rect 11332 17236 11388 17238
rect 11412 17236 11468 17238
rect 11492 17236 11548 17238
rect 11252 16202 11308 16204
rect 11332 16202 11388 16204
rect 11412 16202 11468 16204
rect 11492 16202 11548 16204
rect 11252 16150 11278 16202
rect 11278 16150 11308 16202
rect 11332 16150 11342 16202
rect 11342 16150 11388 16202
rect 11412 16150 11458 16202
rect 11458 16150 11468 16202
rect 11492 16150 11522 16202
rect 11522 16150 11548 16202
rect 11252 16148 11308 16150
rect 11332 16148 11388 16150
rect 11412 16148 11468 16150
rect 11492 16148 11548 16150
rect 11252 15114 11308 15116
rect 11332 15114 11388 15116
rect 11412 15114 11468 15116
rect 11492 15114 11548 15116
rect 11252 15062 11278 15114
rect 11278 15062 11308 15114
rect 11332 15062 11342 15114
rect 11342 15062 11388 15114
rect 11412 15062 11458 15114
rect 11458 15062 11468 15114
rect 11492 15062 11522 15114
rect 11522 15062 11548 15114
rect 11252 15060 11308 15062
rect 11332 15060 11388 15062
rect 11412 15060 11468 15062
rect 11492 15060 11548 15062
rect 11252 14026 11308 14028
rect 11332 14026 11388 14028
rect 11412 14026 11468 14028
rect 11492 14026 11548 14028
rect 11252 13974 11278 14026
rect 11278 13974 11308 14026
rect 11332 13974 11342 14026
rect 11342 13974 11388 14026
rect 11412 13974 11458 14026
rect 11458 13974 11468 14026
rect 11492 13974 11522 14026
rect 11522 13974 11548 14026
rect 11252 13972 11308 13974
rect 11332 13972 11388 13974
rect 11412 13972 11468 13974
rect 11492 13972 11548 13974
rect 11252 12938 11308 12940
rect 11332 12938 11388 12940
rect 11412 12938 11468 12940
rect 11492 12938 11548 12940
rect 11252 12886 11278 12938
rect 11278 12886 11308 12938
rect 11332 12886 11342 12938
rect 11342 12886 11388 12938
rect 11412 12886 11458 12938
rect 11458 12886 11468 12938
rect 11492 12886 11522 12938
rect 11522 12886 11548 12938
rect 11252 12884 11308 12886
rect 11332 12884 11388 12886
rect 11412 12884 11468 12886
rect 11492 12884 11548 12886
rect 11252 11850 11308 11852
rect 11332 11850 11388 11852
rect 11412 11850 11468 11852
rect 11492 11850 11548 11852
rect 11252 11798 11278 11850
rect 11278 11798 11308 11850
rect 11332 11798 11342 11850
rect 11342 11798 11388 11850
rect 11412 11798 11458 11850
rect 11458 11798 11468 11850
rect 11492 11798 11522 11850
rect 11522 11798 11548 11850
rect 11252 11796 11308 11798
rect 11332 11796 11388 11798
rect 11412 11796 11468 11798
rect 11492 11796 11548 11798
rect 11252 10762 11308 10764
rect 11332 10762 11388 10764
rect 11412 10762 11468 10764
rect 11492 10762 11548 10764
rect 11252 10710 11278 10762
rect 11278 10710 11308 10762
rect 11332 10710 11342 10762
rect 11342 10710 11388 10762
rect 11412 10710 11458 10762
rect 11458 10710 11468 10762
rect 11492 10710 11522 10762
rect 11522 10710 11548 10762
rect 11252 10708 11308 10710
rect 11332 10708 11388 10710
rect 11412 10708 11468 10710
rect 11492 10708 11548 10710
rect 11252 9674 11308 9676
rect 11332 9674 11388 9676
rect 11412 9674 11468 9676
rect 11492 9674 11548 9676
rect 11252 9622 11278 9674
rect 11278 9622 11308 9674
rect 11332 9622 11342 9674
rect 11342 9622 11388 9674
rect 11412 9622 11458 9674
rect 11458 9622 11468 9674
rect 11492 9622 11522 9674
rect 11522 9622 11548 9674
rect 11252 9620 11308 9622
rect 11332 9620 11388 9622
rect 11412 9620 11468 9622
rect 11492 9620 11548 9622
rect 11252 8586 11308 8588
rect 11332 8586 11388 8588
rect 11412 8586 11468 8588
rect 11492 8586 11548 8588
rect 11252 8534 11278 8586
rect 11278 8534 11308 8586
rect 11332 8534 11342 8586
rect 11342 8534 11388 8586
rect 11412 8534 11458 8586
rect 11458 8534 11468 8586
rect 11492 8534 11522 8586
rect 11522 8534 11548 8586
rect 11252 8532 11308 8534
rect 11332 8532 11388 8534
rect 11412 8532 11468 8534
rect 11492 8532 11548 8534
rect 11252 7498 11308 7500
rect 11332 7498 11388 7500
rect 11412 7498 11468 7500
rect 11492 7498 11548 7500
rect 11252 7446 11278 7498
rect 11278 7446 11308 7498
rect 11332 7446 11342 7498
rect 11342 7446 11388 7498
rect 11412 7446 11458 7498
rect 11458 7446 11468 7498
rect 11492 7446 11522 7498
rect 11522 7446 11548 7498
rect 11252 7444 11308 7446
rect 11332 7444 11388 7446
rect 11412 7444 11468 7446
rect 11492 7444 11548 7446
rect 4388 6410 4444 6412
rect 4468 6410 4524 6412
rect 4548 6410 4604 6412
rect 4628 6410 4684 6412
rect 4388 6358 4414 6410
rect 4414 6358 4444 6410
rect 4468 6358 4478 6410
rect 4478 6358 4524 6410
rect 4548 6358 4594 6410
rect 4594 6358 4604 6410
rect 4628 6358 4658 6410
rect 4658 6358 4684 6410
rect 4388 6356 4444 6358
rect 4468 6356 4524 6358
rect 4548 6356 4604 6358
rect 4628 6356 4684 6358
rect 11252 6410 11308 6412
rect 11332 6410 11388 6412
rect 11412 6410 11468 6412
rect 11492 6410 11548 6412
rect 11252 6358 11278 6410
rect 11278 6358 11308 6410
rect 11332 6358 11342 6410
rect 11342 6358 11388 6410
rect 11412 6358 11458 6410
rect 11458 6358 11468 6410
rect 11492 6358 11522 6410
rect 11522 6358 11548 6410
rect 11252 6356 11308 6358
rect 11332 6356 11388 6358
rect 11412 6356 11468 6358
rect 11492 6356 11548 6358
rect 7820 5866 7876 5868
rect 7900 5866 7956 5868
rect 7980 5866 8036 5868
rect 8060 5866 8116 5868
rect 7820 5814 7846 5866
rect 7846 5814 7876 5866
rect 7900 5814 7910 5866
rect 7910 5814 7956 5866
rect 7980 5814 8026 5866
rect 8026 5814 8036 5866
rect 8060 5814 8090 5866
rect 8090 5814 8116 5866
rect 7820 5812 7876 5814
rect 7900 5812 7956 5814
rect 7980 5812 8036 5814
rect 8060 5812 8116 5814
rect 14684 20010 14740 20012
rect 14764 20010 14820 20012
rect 14844 20010 14900 20012
rect 14924 20010 14980 20012
rect 14684 19958 14710 20010
rect 14710 19958 14740 20010
rect 14764 19958 14774 20010
rect 14774 19958 14820 20010
rect 14844 19958 14890 20010
rect 14890 19958 14900 20010
rect 14924 19958 14954 20010
rect 14954 19958 14980 20010
rect 14684 19956 14740 19958
rect 14764 19956 14820 19958
rect 14844 19956 14900 19958
rect 14924 19956 14980 19958
rect 14684 18922 14740 18924
rect 14764 18922 14820 18924
rect 14844 18922 14900 18924
rect 14924 18922 14980 18924
rect 14684 18870 14710 18922
rect 14710 18870 14740 18922
rect 14764 18870 14774 18922
rect 14774 18870 14820 18922
rect 14844 18870 14890 18922
rect 14890 18870 14900 18922
rect 14924 18870 14954 18922
rect 14954 18870 14980 18922
rect 14684 18868 14740 18870
rect 14764 18868 14820 18870
rect 14844 18868 14900 18870
rect 14924 18868 14980 18870
rect 15750 19092 15806 19128
rect 15750 19072 15752 19092
rect 15752 19072 15804 19092
rect 15804 19072 15806 19092
rect 15198 18004 15254 18040
rect 15198 17984 15200 18004
rect 15200 17984 15252 18004
rect 15252 17984 15254 18004
rect 14684 17834 14740 17836
rect 14764 17834 14820 17836
rect 14844 17834 14900 17836
rect 14924 17834 14980 17836
rect 14684 17782 14710 17834
rect 14710 17782 14740 17834
rect 14764 17782 14774 17834
rect 14774 17782 14820 17834
rect 14844 17782 14890 17834
rect 14890 17782 14900 17834
rect 14924 17782 14954 17834
rect 14954 17782 14980 17834
rect 14684 17780 14740 17782
rect 14764 17780 14820 17782
rect 14844 17780 14900 17782
rect 14924 17780 14980 17782
rect 14684 16746 14740 16748
rect 14764 16746 14820 16748
rect 14844 16746 14900 16748
rect 14924 16746 14980 16748
rect 14684 16694 14710 16746
rect 14710 16694 14740 16746
rect 14764 16694 14774 16746
rect 14774 16694 14820 16746
rect 14844 16694 14890 16746
rect 14890 16694 14900 16746
rect 14924 16694 14954 16746
rect 14954 16694 14980 16746
rect 14684 16692 14740 16694
rect 14764 16692 14820 16694
rect 14844 16692 14900 16694
rect 14924 16692 14980 16694
rect 14684 15658 14740 15660
rect 14764 15658 14820 15660
rect 14844 15658 14900 15660
rect 14924 15658 14980 15660
rect 14684 15606 14710 15658
rect 14710 15606 14740 15658
rect 14764 15606 14774 15658
rect 14774 15606 14820 15658
rect 14844 15606 14890 15658
rect 14890 15606 14900 15658
rect 14924 15606 14954 15658
rect 14954 15606 14980 15658
rect 14684 15604 14740 15606
rect 14764 15604 14820 15606
rect 14844 15604 14900 15606
rect 14924 15604 14980 15606
rect 14684 14570 14740 14572
rect 14764 14570 14820 14572
rect 14844 14570 14900 14572
rect 14924 14570 14980 14572
rect 14684 14518 14710 14570
rect 14710 14518 14740 14570
rect 14764 14518 14774 14570
rect 14774 14518 14820 14570
rect 14844 14518 14890 14570
rect 14890 14518 14900 14570
rect 14924 14518 14954 14570
rect 14954 14518 14980 14570
rect 14684 14516 14740 14518
rect 14764 14516 14820 14518
rect 14844 14516 14900 14518
rect 14924 14516 14980 14518
rect 14684 13482 14740 13484
rect 14764 13482 14820 13484
rect 14844 13482 14900 13484
rect 14924 13482 14980 13484
rect 14684 13430 14710 13482
rect 14710 13430 14740 13482
rect 14764 13430 14774 13482
rect 14774 13430 14820 13482
rect 14844 13430 14890 13482
rect 14890 13430 14900 13482
rect 14924 13430 14954 13482
rect 14954 13430 14980 13482
rect 14684 13428 14740 13430
rect 14764 13428 14820 13430
rect 14844 13428 14900 13430
rect 14924 13428 14980 13430
rect 14684 12394 14740 12396
rect 14764 12394 14820 12396
rect 14844 12394 14900 12396
rect 14924 12394 14980 12396
rect 14684 12342 14710 12394
rect 14710 12342 14740 12394
rect 14764 12342 14774 12394
rect 14774 12342 14820 12394
rect 14844 12342 14890 12394
rect 14890 12342 14900 12394
rect 14924 12342 14954 12394
rect 14954 12342 14980 12394
rect 14684 12340 14740 12342
rect 14764 12340 14820 12342
rect 14844 12340 14900 12342
rect 14924 12340 14980 12342
rect 14684 11306 14740 11308
rect 14764 11306 14820 11308
rect 14844 11306 14900 11308
rect 14924 11306 14980 11308
rect 14684 11254 14710 11306
rect 14710 11254 14740 11306
rect 14764 11254 14774 11306
rect 14774 11254 14820 11306
rect 14844 11254 14890 11306
rect 14890 11254 14900 11306
rect 14924 11254 14954 11306
rect 14954 11254 14980 11306
rect 14684 11252 14740 11254
rect 14764 11252 14820 11254
rect 14844 11252 14900 11254
rect 14924 11252 14980 11254
rect 14684 10218 14740 10220
rect 14764 10218 14820 10220
rect 14844 10218 14900 10220
rect 14924 10218 14980 10220
rect 14684 10166 14710 10218
rect 14710 10166 14740 10218
rect 14764 10166 14774 10218
rect 14774 10166 14820 10218
rect 14844 10166 14890 10218
rect 14890 10166 14900 10218
rect 14924 10166 14954 10218
rect 14954 10166 14980 10218
rect 14684 10164 14740 10166
rect 14764 10164 14820 10166
rect 14844 10164 14900 10166
rect 14924 10164 14980 10166
rect 14370 9416 14426 9472
rect 14684 9130 14740 9132
rect 14764 9130 14820 9132
rect 14844 9130 14900 9132
rect 14924 9130 14980 9132
rect 14684 9078 14710 9130
rect 14710 9078 14740 9130
rect 14764 9078 14774 9130
rect 14774 9078 14820 9130
rect 14844 9078 14890 9130
rect 14890 9078 14900 9130
rect 14924 9078 14954 9130
rect 14954 9078 14980 9130
rect 14684 9076 14740 9078
rect 14764 9076 14820 9078
rect 14844 9076 14900 9078
rect 14924 9076 14980 9078
rect 14684 8042 14740 8044
rect 14764 8042 14820 8044
rect 14844 8042 14900 8044
rect 14924 8042 14980 8044
rect 14684 7990 14710 8042
rect 14710 7990 14740 8042
rect 14764 7990 14774 8042
rect 14774 7990 14820 8042
rect 14844 7990 14890 8042
rect 14890 7990 14900 8042
rect 14924 7990 14954 8042
rect 14954 7990 14980 8042
rect 14684 7988 14740 7990
rect 14764 7988 14820 7990
rect 14844 7988 14900 7990
rect 14924 7988 14980 7990
rect 17038 18664 17094 18720
rect 17958 21384 18014 21440
rect 18116 19466 18172 19468
rect 18196 19466 18252 19468
rect 18276 19466 18332 19468
rect 18356 19466 18412 19468
rect 18116 19414 18142 19466
rect 18142 19414 18172 19466
rect 18196 19414 18206 19466
rect 18206 19414 18252 19466
rect 18276 19414 18322 19466
rect 18322 19414 18332 19466
rect 18356 19414 18386 19466
rect 18386 19414 18412 19466
rect 18116 19412 18172 19414
rect 18196 19412 18252 19414
rect 18276 19412 18332 19414
rect 18356 19412 18412 19414
rect 18116 18378 18172 18380
rect 18196 18378 18252 18380
rect 18276 18378 18332 18380
rect 18356 18378 18412 18380
rect 18116 18326 18142 18378
rect 18142 18326 18172 18378
rect 18196 18326 18206 18378
rect 18206 18326 18252 18378
rect 18276 18326 18322 18378
rect 18322 18326 18332 18378
rect 18356 18326 18386 18378
rect 18386 18326 18412 18378
rect 18116 18324 18172 18326
rect 18196 18324 18252 18326
rect 18276 18324 18332 18326
rect 18356 18324 18412 18326
rect 18694 21928 18750 21984
rect 18116 17290 18172 17292
rect 18196 17290 18252 17292
rect 18276 17290 18332 17292
rect 18356 17290 18412 17292
rect 18116 17238 18142 17290
rect 18142 17238 18172 17290
rect 18196 17238 18206 17290
rect 18206 17238 18252 17290
rect 18276 17238 18322 17290
rect 18322 17238 18332 17290
rect 18356 17238 18386 17290
rect 18386 17238 18412 17290
rect 18116 17236 18172 17238
rect 18196 17236 18252 17238
rect 18276 17236 18332 17238
rect 18356 17236 18412 17238
rect 4066 5608 4122 5664
rect 4388 5322 4444 5324
rect 4468 5322 4524 5324
rect 4548 5322 4604 5324
rect 4628 5322 4684 5324
rect 4388 5270 4414 5322
rect 4414 5270 4444 5322
rect 4468 5270 4478 5322
rect 4478 5270 4524 5322
rect 4548 5270 4594 5322
rect 4594 5270 4604 5322
rect 4628 5270 4658 5322
rect 4658 5270 4684 5322
rect 4388 5268 4444 5270
rect 4468 5268 4524 5270
rect 4548 5268 4604 5270
rect 4628 5268 4684 5270
rect 11252 5322 11308 5324
rect 11332 5322 11388 5324
rect 11412 5322 11468 5324
rect 11492 5322 11548 5324
rect 11252 5270 11278 5322
rect 11278 5270 11308 5322
rect 11332 5270 11342 5322
rect 11342 5270 11388 5322
rect 11412 5270 11458 5322
rect 11458 5270 11468 5322
rect 11492 5270 11522 5322
rect 11522 5270 11548 5322
rect 11252 5268 11308 5270
rect 11332 5268 11388 5270
rect 11412 5268 11468 5270
rect 11492 5268 11548 5270
rect 7820 4778 7876 4780
rect 7900 4778 7956 4780
rect 7980 4778 8036 4780
rect 8060 4778 8116 4780
rect 7820 4726 7846 4778
rect 7846 4726 7876 4778
rect 7900 4726 7910 4778
rect 7910 4726 7956 4778
rect 7980 4726 8026 4778
rect 8026 4726 8036 4778
rect 8060 4726 8090 4778
rect 8090 4726 8116 4778
rect 7820 4724 7876 4726
rect 7900 4724 7956 4726
rect 7980 4724 8036 4726
rect 8060 4724 8116 4726
rect 4388 4234 4444 4236
rect 4468 4234 4524 4236
rect 4548 4234 4604 4236
rect 4628 4234 4684 4236
rect 4388 4182 4414 4234
rect 4414 4182 4444 4234
rect 4468 4182 4478 4234
rect 4478 4182 4524 4234
rect 4548 4182 4594 4234
rect 4594 4182 4604 4234
rect 4628 4182 4658 4234
rect 4658 4182 4684 4234
rect 4388 4180 4444 4182
rect 4468 4180 4524 4182
rect 4548 4180 4604 4182
rect 4628 4180 4684 4182
rect 11252 4234 11308 4236
rect 11332 4234 11388 4236
rect 11412 4234 11468 4236
rect 11492 4234 11548 4236
rect 11252 4182 11278 4234
rect 11278 4182 11308 4234
rect 11332 4182 11342 4234
rect 11342 4182 11388 4234
rect 11412 4182 11458 4234
rect 11458 4182 11468 4234
rect 11492 4182 11522 4234
rect 11522 4182 11548 4234
rect 11252 4180 11308 4182
rect 11332 4180 11388 4182
rect 11412 4180 11468 4182
rect 11492 4180 11548 4182
rect 7820 3690 7876 3692
rect 7900 3690 7956 3692
rect 7980 3690 8036 3692
rect 8060 3690 8116 3692
rect 7820 3638 7846 3690
rect 7846 3638 7876 3690
rect 7900 3638 7910 3690
rect 7910 3638 7956 3690
rect 7980 3638 8026 3690
rect 8026 3638 8036 3690
rect 8060 3638 8090 3690
rect 8090 3638 8116 3690
rect 7820 3636 7876 3638
rect 7900 3636 7956 3638
rect 7980 3636 8036 3638
rect 8060 3636 8116 3638
rect 4388 3146 4444 3148
rect 4468 3146 4524 3148
rect 4548 3146 4604 3148
rect 4628 3146 4684 3148
rect 4388 3094 4414 3146
rect 4414 3094 4444 3146
rect 4468 3094 4478 3146
rect 4478 3094 4524 3146
rect 4548 3094 4594 3146
rect 4594 3094 4604 3146
rect 4628 3094 4658 3146
rect 4658 3094 4684 3146
rect 4388 3092 4444 3094
rect 4468 3092 4524 3094
rect 4548 3092 4604 3094
rect 4628 3092 4684 3094
rect 11252 3146 11308 3148
rect 11332 3146 11388 3148
rect 11412 3146 11468 3148
rect 11492 3146 11548 3148
rect 11252 3094 11278 3146
rect 11278 3094 11308 3146
rect 11332 3094 11342 3146
rect 11342 3094 11388 3146
rect 11412 3094 11458 3146
rect 11458 3094 11468 3146
rect 11492 3094 11522 3146
rect 11522 3094 11548 3146
rect 11252 3092 11308 3094
rect 11332 3092 11388 3094
rect 11412 3092 11468 3094
rect 11492 3092 11548 3094
rect 7820 2602 7876 2604
rect 7900 2602 7956 2604
rect 7980 2602 8036 2604
rect 8060 2602 8116 2604
rect 7820 2550 7846 2602
rect 7846 2550 7876 2602
rect 7900 2550 7910 2602
rect 7910 2550 7956 2602
rect 7980 2550 8026 2602
rect 8026 2550 8036 2602
rect 8060 2550 8090 2602
rect 8090 2550 8116 2602
rect 7820 2548 7876 2550
rect 7900 2548 7956 2550
rect 7980 2548 8036 2550
rect 8060 2548 8116 2550
rect 4388 2058 4444 2060
rect 4468 2058 4524 2060
rect 4548 2058 4604 2060
rect 4628 2058 4684 2060
rect 4388 2006 4414 2058
rect 4414 2006 4444 2058
rect 4468 2006 4478 2058
rect 4478 2006 4524 2058
rect 4548 2006 4594 2058
rect 4594 2006 4604 2058
rect 4628 2006 4658 2058
rect 4658 2006 4684 2058
rect 4388 2004 4444 2006
rect 4468 2004 4524 2006
rect 4548 2004 4604 2006
rect 4628 2004 4684 2006
rect 11252 2058 11308 2060
rect 11332 2058 11388 2060
rect 11412 2058 11468 2060
rect 11492 2058 11548 2060
rect 11252 2006 11278 2058
rect 11278 2006 11308 2058
rect 11332 2006 11342 2058
rect 11342 2006 11388 2058
rect 11412 2006 11458 2058
rect 11458 2006 11468 2058
rect 11492 2006 11522 2058
rect 11522 2006 11548 2058
rect 11252 2004 11308 2006
rect 11332 2004 11388 2006
rect 11412 2004 11468 2006
rect 11492 2004 11548 2006
rect 14684 6954 14740 6956
rect 14764 6954 14820 6956
rect 14844 6954 14900 6956
rect 14924 6954 14980 6956
rect 14684 6902 14710 6954
rect 14710 6902 14740 6954
rect 14764 6902 14774 6954
rect 14774 6902 14820 6954
rect 14844 6902 14890 6954
rect 14890 6902 14900 6954
rect 14924 6902 14954 6954
rect 14954 6902 14980 6954
rect 14684 6900 14740 6902
rect 14764 6900 14820 6902
rect 14844 6900 14900 6902
rect 14924 6900 14980 6902
rect 14684 5866 14740 5868
rect 14764 5866 14820 5868
rect 14844 5866 14900 5868
rect 14924 5866 14980 5868
rect 14684 5814 14710 5866
rect 14710 5814 14740 5866
rect 14764 5814 14774 5866
rect 14774 5814 14820 5866
rect 14844 5814 14890 5866
rect 14890 5814 14900 5866
rect 14924 5814 14954 5866
rect 14954 5814 14980 5866
rect 14684 5812 14740 5814
rect 14764 5812 14820 5814
rect 14844 5812 14900 5814
rect 14924 5812 14980 5814
rect 14684 4778 14740 4780
rect 14764 4778 14820 4780
rect 14844 4778 14900 4780
rect 14924 4778 14980 4780
rect 14684 4726 14710 4778
rect 14710 4726 14740 4778
rect 14764 4726 14774 4778
rect 14774 4726 14820 4778
rect 14844 4726 14890 4778
rect 14890 4726 14900 4778
rect 14924 4726 14954 4778
rect 14954 4726 14980 4778
rect 14684 4724 14740 4726
rect 14764 4724 14820 4726
rect 14844 4724 14900 4726
rect 14924 4724 14980 4726
rect 14684 3690 14740 3692
rect 14764 3690 14820 3692
rect 14844 3690 14900 3692
rect 14924 3690 14980 3692
rect 14684 3638 14710 3690
rect 14710 3638 14740 3690
rect 14764 3638 14774 3690
rect 14774 3638 14820 3690
rect 14844 3638 14890 3690
rect 14890 3638 14900 3690
rect 14924 3638 14954 3690
rect 14954 3638 14980 3690
rect 14684 3636 14740 3638
rect 14764 3636 14820 3638
rect 14844 3636 14900 3638
rect 14924 3636 14980 3638
rect 14684 2602 14740 2604
rect 14764 2602 14820 2604
rect 14844 2602 14900 2604
rect 14924 2602 14980 2604
rect 14684 2550 14710 2602
rect 14710 2550 14740 2602
rect 14764 2550 14774 2602
rect 14774 2550 14820 2602
rect 14844 2550 14890 2602
rect 14890 2550 14900 2602
rect 14924 2550 14954 2602
rect 14954 2550 14980 2602
rect 14684 2548 14740 2550
rect 14764 2548 14820 2550
rect 14844 2548 14900 2550
rect 14924 2548 14980 2550
rect 18116 16202 18172 16204
rect 18196 16202 18252 16204
rect 18276 16202 18332 16204
rect 18356 16202 18412 16204
rect 18116 16150 18142 16202
rect 18142 16150 18172 16202
rect 18196 16150 18206 16202
rect 18206 16150 18252 16202
rect 18276 16150 18322 16202
rect 18322 16150 18332 16202
rect 18356 16150 18386 16202
rect 18386 16150 18412 16202
rect 18116 16148 18172 16150
rect 18196 16148 18252 16150
rect 18276 16148 18332 16150
rect 18356 16148 18412 16150
rect 18116 15114 18172 15116
rect 18196 15114 18252 15116
rect 18276 15114 18332 15116
rect 18356 15114 18412 15116
rect 18116 15062 18142 15114
rect 18142 15062 18172 15114
rect 18196 15062 18206 15114
rect 18206 15062 18252 15114
rect 18276 15062 18322 15114
rect 18322 15062 18332 15114
rect 18356 15062 18386 15114
rect 18386 15062 18412 15114
rect 18116 15060 18172 15062
rect 18196 15060 18252 15062
rect 18276 15060 18332 15062
rect 18356 15060 18412 15062
rect 18116 14026 18172 14028
rect 18196 14026 18252 14028
rect 18276 14026 18332 14028
rect 18356 14026 18412 14028
rect 18116 13974 18142 14026
rect 18142 13974 18172 14026
rect 18196 13974 18206 14026
rect 18206 13974 18252 14026
rect 18276 13974 18322 14026
rect 18322 13974 18332 14026
rect 18356 13974 18386 14026
rect 18386 13974 18412 14026
rect 18116 13972 18172 13974
rect 18196 13972 18252 13974
rect 18276 13972 18332 13974
rect 18356 13972 18412 13974
rect 19062 18664 19118 18720
rect 19246 20976 19302 21032
rect 19890 19616 19946 19672
rect 19246 16932 19248 16952
rect 19248 16932 19300 16952
rect 19300 16932 19302 16952
rect 19246 16896 19302 16932
rect 19154 14176 19210 14232
rect 18116 12938 18172 12940
rect 18196 12938 18252 12940
rect 18276 12938 18332 12940
rect 18356 12938 18412 12940
rect 18116 12886 18142 12938
rect 18142 12886 18172 12938
rect 18196 12886 18206 12938
rect 18206 12886 18252 12938
rect 18276 12886 18322 12938
rect 18322 12886 18332 12938
rect 18356 12886 18386 12938
rect 18386 12886 18412 12938
rect 18116 12884 18172 12886
rect 18196 12884 18252 12886
rect 18276 12884 18332 12886
rect 18356 12884 18412 12886
rect 18116 11850 18172 11852
rect 18196 11850 18252 11852
rect 18276 11850 18332 11852
rect 18356 11850 18412 11852
rect 18116 11798 18142 11850
rect 18142 11798 18172 11850
rect 18196 11798 18206 11850
rect 18206 11798 18252 11850
rect 18276 11798 18322 11850
rect 18322 11798 18332 11850
rect 18356 11798 18386 11850
rect 18386 11798 18412 11850
rect 18116 11796 18172 11798
rect 18196 11796 18252 11798
rect 18276 11796 18332 11798
rect 18356 11796 18412 11798
rect 18116 10762 18172 10764
rect 18196 10762 18252 10764
rect 18276 10762 18332 10764
rect 18356 10762 18412 10764
rect 18116 10710 18142 10762
rect 18142 10710 18172 10762
rect 18196 10710 18206 10762
rect 18206 10710 18252 10762
rect 18276 10710 18322 10762
rect 18322 10710 18332 10762
rect 18356 10710 18386 10762
rect 18386 10710 18412 10762
rect 18116 10708 18172 10710
rect 18196 10708 18252 10710
rect 18276 10708 18332 10710
rect 18356 10708 18412 10710
rect 18116 9674 18172 9676
rect 18196 9674 18252 9676
rect 18276 9674 18332 9676
rect 18356 9674 18412 9676
rect 18116 9622 18142 9674
rect 18142 9622 18172 9674
rect 18196 9622 18206 9674
rect 18206 9622 18252 9674
rect 18276 9622 18322 9674
rect 18322 9622 18332 9674
rect 18356 9622 18386 9674
rect 18386 9622 18412 9674
rect 18116 9620 18172 9622
rect 18196 9620 18252 9622
rect 18276 9620 18332 9622
rect 18356 9620 18412 9622
rect 18116 8586 18172 8588
rect 18196 8586 18252 8588
rect 18276 8586 18332 8588
rect 18356 8586 18412 8588
rect 18116 8534 18142 8586
rect 18142 8534 18172 8586
rect 18196 8534 18206 8586
rect 18206 8534 18252 8586
rect 18276 8534 18322 8586
rect 18322 8534 18332 8586
rect 18356 8534 18386 8586
rect 18386 8534 18412 8586
rect 18116 8532 18172 8534
rect 18196 8532 18252 8534
rect 18276 8532 18332 8534
rect 18356 8532 18412 8534
rect 18116 7498 18172 7500
rect 18196 7498 18252 7500
rect 18276 7498 18332 7500
rect 18356 7498 18412 7500
rect 18116 7446 18142 7498
rect 18142 7446 18172 7498
rect 18196 7446 18206 7498
rect 18206 7446 18252 7498
rect 18276 7446 18322 7498
rect 18322 7446 18332 7498
rect 18356 7446 18386 7498
rect 18386 7446 18412 7498
rect 18116 7444 18172 7446
rect 18196 7444 18252 7446
rect 18276 7444 18332 7446
rect 18356 7444 18412 7446
rect 18510 6424 18566 6480
rect 18116 6410 18172 6412
rect 18196 6410 18252 6412
rect 18276 6410 18332 6412
rect 18356 6410 18412 6412
rect 18116 6358 18142 6410
rect 18142 6358 18172 6410
rect 18196 6358 18206 6410
rect 18206 6358 18252 6410
rect 18276 6358 18322 6410
rect 18322 6358 18332 6410
rect 18356 6358 18386 6410
rect 18386 6358 18412 6410
rect 18116 6356 18172 6358
rect 18196 6356 18252 6358
rect 18276 6356 18332 6358
rect 18356 6356 18412 6358
rect 18602 5472 18658 5528
rect 18116 5322 18172 5324
rect 18196 5322 18252 5324
rect 18276 5322 18332 5324
rect 18356 5322 18412 5324
rect 18116 5270 18142 5322
rect 18142 5270 18172 5322
rect 18196 5270 18206 5322
rect 18206 5270 18252 5322
rect 18276 5270 18322 5322
rect 18322 5270 18332 5322
rect 18356 5270 18386 5322
rect 18386 5270 18412 5322
rect 18116 5268 18172 5270
rect 18196 5268 18252 5270
rect 18276 5268 18332 5270
rect 18356 5268 18412 5270
rect 17958 4520 18014 4576
rect 18116 4234 18172 4236
rect 18196 4234 18252 4236
rect 18276 4234 18332 4236
rect 18356 4234 18412 4236
rect 18116 4182 18142 4234
rect 18142 4182 18172 4234
rect 18196 4182 18206 4234
rect 18206 4182 18252 4234
rect 18276 4182 18322 4234
rect 18322 4182 18332 4234
rect 18356 4182 18386 4234
rect 18386 4182 18412 4234
rect 18116 4180 18172 4182
rect 18196 4180 18252 4182
rect 18276 4180 18332 4182
rect 18356 4180 18412 4182
rect 17866 3568 17922 3624
rect 18116 3146 18172 3148
rect 18196 3146 18252 3148
rect 18276 3146 18332 3148
rect 18356 3146 18412 3148
rect 18116 3094 18142 3146
rect 18142 3094 18172 3146
rect 18196 3094 18206 3146
rect 18206 3094 18252 3146
rect 18276 3094 18322 3146
rect 18322 3094 18332 3146
rect 18356 3094 18386 3146
rect 18386 3094 18412 3146
rect 18116 3092 18172 3094
rect 18196 3092 18252 3094
rect 18276 3092 18332 3094
rect 18356 3092 18412 3094
rect 18116 2058 18172 2060
rect 18196 2058 18252 2060
rect 18276 2058 18332 2060
rect 18356 2058 18412 2060
rect 18116 2006 18142 2058
rect 18142 2006 18172 2058
rect 18196 2006 18206 2058
rect 18206 2006 18252 2058
rect 18276 2006 18322 2058
rect 18322 2006 18332 2058
rect 18356 2006 18386 2058
rect 18386 2006 18412 2058
rect 18116 2004 18172 2006
rect 18196 2004 18252 2006
rect 18276 2004 18332 2006
rect 18356 2004 18412 2006
rect 18786 9280 18842 9336
rect 18786 3160 18842 3216
rect 18694 1800 18750 1856
rect 17958 1392 18014 1448
rect 17958 848 18014 904
rect 19246 12272 19302 12328
rect 19062 9960 19118 10016
rect 20626 20568 20682 20624
rect 20718 20024 20774 20080
rect 20350 18256 20406 18312
rect 20994 19208 21050 19264
rect 19706 12816 19762 12872
rect 20166 16352 20222 16408
rect 20074 15980 20076 16000
rect 20076 15980 20128 16000
rect 20128 15980 20130 16000
rect 20074 15944 20130 15980
rect 20074 13224 20130 13280
rect 20166 11864 20222 11920
rect 19890 11456 19946 11512
rect 20442 16896 20498 16952
rect 20442 15536 20498 15592
rect 20442 14584 20498 14640
rect 20718 13632 20774 13688
rect 20442 10912 20498 10968
rect 20534 10504 20590 10560
rect 20258 9552 20314 9608
rect 20534 9144 20590 9200
rect 20534 8600 20590 8656
rect 19982 8192 20038 8248
rect 20258 7784 20314 7840
rect 20534 7240 20590 7296
rect 19982 6832 20038 6888
rect 20534 5880 20590 5936
rect 20534 4928 20590 4984
rect 20902 17848 20958 17904
rect 20902 14992 20958 15048
rect 21730 17324 21786 17360
rect 21730 17304 21732 17324
rect 21732 17304 21784 17324
rect 21784 17304 21786 17324
rect 20534 4112 20590 4168
rect 19062 2752 19118 2808
rect 18970 2208 19026 2264
rect 18878 440 18934 496
rect 17222 32 17278 88
<< metal3 >>
rect 18873 22394 18939 22397
rect 22320 22394 22800 22424
rect 18873 22392 22800 22394
rect 18873 22336 18878 22392
rect 18934 22336 22800 22392
rect 18873 22334 22800 22336
rect 18873 22331 18939 22334
rect 22320 22304 22800 22334
rect 18689 21986 18755 21989
rect 22320 21986 22800 22016
rect 18689 21984 22800 21986
rect 18689 21928 18694 21984
rect 18750 21928 22800 21984
rect 18689 21926 22800 21928
rect 18689 21923 18755 21926
rect 22320 21896 22800 21926
rect 17953 21442 18019 21445
rect 22320 21442 22800 21472
rect 17953 21440 22800 21442
rect 17953 21384 17958 21440
rect 18014 21384 22800 21440
rect 17953 21382 22800 21384
rect 17953 21379 18019 21382
rect 22320 21352 22800 21382
rect 19241 21034 19307 21037
rect 22320 21034 22800 21064
rect 19241 21032 22800 21034
rect 19241 20976 19246 21032
rect 19302 20976 22800 21032
rect 19241 20974 22800 20976
rect 19241 20971 19307 20974
rect 22320 20944 22800 20974
rect 20621 20626 20687 20629
rect 22320 20626 22800 20656
rect 20621 20624 22800 20626
rect 20621 20568 20626 20624
rect 20682 20568 22800 20624
rect 20621 20566 22800 20568
rect 20621 20563 20687 20566
rect 22320 20536 22800 20566
rect 20713 20082 20779 20085
rect 22320 20082 22800 20112
rect 20713 20080 22800 20082
rect 20713 20024 20718 20080
rect 20774 20024 22800 20080
rect 20713 20022 22800 20024
rect 20713 20019 20779 20022
rect 7808 20016 8128 20017
rect 7808 19952 7816 20016
rect 7880 19952 7896 20016
rect 7960 19952 7976 20016
rect 8040 19952 8056 20016
rect 8120 19952 8128 20016
rect 7808 19951 8128 19952
rect 14672 20016 14992 20017
rect 14672 19952 14680 20016
rect 14744 19952 14760 20016
rect 14824 19952 14840 20016
rect 14904 19952 14920 20016
rect 14984 19952 14992 20016
rect 22320 19992 22800 20022
rect 14672 19951 14992 19952
rect 19885 19674 19951 19677
rect 22320 19674 22800 19704
rect 19885 19672 22800 19674
rect 19885 19616 19890 19672
rect 19946 19616 22800 19672
rect 19885 19614 22800 19616
rect 19885 19611 19951 19614
rect 22320 19584 22800 19614
rect 4376 19472 4696 19473
rect 4376 19408 4384 19472
rect 4448 19408 4464 19472
rect 4528 19408 4544 19472
rect 4608 19408 4624 19472
rect 4688 19408 4696 19472
rect 4376 19407 4696 19408
rect 11240 19472 11560 19473
rect 11240 19408 11248 19472
rect 11312 19408 11328 19472
rect 11392 19408 11408 19472
rect 11472 19408 11488 19472
rect 11552 19408 11560 19472
rect 11240 19407 11560 19408
rect 18104 19472 18424 19473
rect 18104 19408 18112 19472
rect 18176 19408 18192 19472
rect 18256 19408 18272 19472
rect 18336 19408 18352 19472
rect 18416 19408 18424 19472
rect 18104 19407 18424 19408
rect 20989 19266 21055 19269
rect 22320 19266 22800 19296
rect 20989 19264 22800 19266
rect 20989 19208 20994 19264
rect 21050 19208 22800 19264
rect 20989 19206 22800 19208
rect 20989 19203 21055 19206
rect 22320 19176 22800 19206
rect 10225 19130 10291 19133
rect 15745 19130 15811 19133
rect 10225 19128 15811 19130
rect 10225 19072 10230 19128
rect 10286 19072 15750 19128
rect 15806 19072 15811 19128
rect 10225 19070 15811 19072
rect 10225 19067 10291 19070
rect 15745 19067 15811 19070
rect 7808 18928 8128 18929
rect 7808 18864 7816 18928
rect 7880 18864 7896 18928
rect 7960 18864 7976 18928
rect 8040 18864 8056 18928
rect 8120 18864 8128 18928
rect 7808 18863 8128 18864
rect 14672 18928 14992 18929
rect 14672 18864 14680 18928
rect 14744 18864 14760 18928
rect 14824 18864 14840 18928
rect 14904 18864 14920 18928
rect 14984 18864 14992 18928
rect 14672 18863 14992 18864
rect 10777 18722 10843 18725
rect 17033 18722 17099 18725
rect 10777 18720 17099 18722
rect 10777 18664 10782 18720
rect 10838 18664 17038 18720
rect 17094 18664 17099 18720
rect 10777 18662 17099 18664
rect 10777 18659 10843 18662
rect 17033 18659 17099 18662
rect 19057 18722 19123 18725
rect 22320 18722 22800 18752
rect 19057 18720 22800 18722
rect 19057 18664 19062 18720
rect 19118 18664 22800 18720
rect 19057 18662 22800 18664
rect 19057 18659 19123 18662
rect 22320 18632 22800 18662
rect 4376 18384 4696 18385
rect 4376 18320 4384 18384
rect 4448 18320 4464 18384
rect 4528 18320 4544 18384
rect 4608 18320 4624 18384
rect 4688 18320 4696 18384
rect 4376 18319 4696 18320
rect 11240 18384 11560 18385
rect 11240 18320 11248 18384
rect 11312 18320 11328 18384
rect 11392 18320 11408 18384
rect 11472 18320 11488 18384
rect 11552 18320 11560 18384
rect 11240 18319 11560 18320
rect 18104 18384 18424 18385
rect 18104 18320 18112 18384
rect 18176 18320 18192 18384
rect 18256 18320 18272 18384
rect 18336 18320 18352 18384
rect 18416 18320 18424 18384
rect 18104 18319 18424 18320
rect 20345 18314 20411 18317
rect 22320 18314 22800 18344
rect 20345 18312 22800 18314
rect 20345 18256 20350 18312
rect 20406 18256 22800 18312
rect 20345 18254 22800 18256
rect 20345 18251 20411 18254
rect 22320 18224 22800 18254
rect 9029 18178 9095 18181
rect 10409 18178 10475 18181
rect 9029 18176 10475 18178
rect 9029 18120 9034 18176
rect 9090 18120 10414 18176
rect 10470 18120 10475 18176
rect 9029 18118 10475 18120
rect 9029 18115 9095 18118
rect 10409 18115 10475 18118
rect 10593 18042 10659 18045
rect 15193 18042 15259 18045
rect 10593 18040 15259 18042
rect 10593 17984 10598 18040
rect 10654 17984 15198 18040
rect 15254 17984 15259 18040
rect 10593 17982 15259 17984
rect 10593 17979 10659 17982
rect 15193 17979 15259 17982
rect 20897 17906 20963 17909
rect 22320 17906 22800 17936
rect 20897 17904 22800 17906
rect 20897 17848 20902 17904
rect 20958 17848 22800 17904
rect 20897 17846 22800 17848
rect 20897 17843 20963 17846
rect 7808 17840 8128 17841
rect 7808 17776 7816 17840
rect 7880 17776 7896 17840
rect 7960 17776 7976 17840
rect 8040 17776 8056 17840
rect 8120 17776 8128 17840
rect 7808 17775 8128 17776
rect 14672 17840 14992 17841
rect 14672 17776 14680 17840
rect 14744 17776 14760 17840
rect 14824 17776 14840 17840
rect 14904 17776 14920 17840
rect 14984 17776 14992 17840
rect 22320 17816 22800 17846
rect 14672 17775 14992 17776
rect 21725 17362 21791 17365
rect 22320 17362 22800 17392
rect 21725 17360 22800 17362
rect 21725 17304 21730 17360
rect 21786 17304 22800 17360
rect 21725 17302 22800 17304
rect 21725 17299 21791 17302
rect 4376 17296 4696 17297
rect 4376 17232 4384 17296
rect 4448 17232 4464 17296
rect 4528 17232 4544 17296
rect 4608 17232 4624 17296
rect 4688 17232 4696 17296
rect 4376 17231 4696 17232
rect 11240 17296 11560 17297
rect 11240 17232 11248 17296
rect 11312 17232 11328 17296
rect 11392 17232 11408 17296
rect 11472 17232 11488 17296
rect 11552 17232 11560 17296
rect 11240 17231 11560 17232
rect 18104 17296 18424 17297
rect 18104 17232 18112 17296
rect 18176 17232 18192 17296
rect 18256 17232 18272 17296
rect 18336 17232 18352 17296
rect 18416 17232 18424 17296
rect 22320 17272 22800 17302
rect 18104 17231 18424 17232
rect 0 17090 480 17120
rect 4061 17090 4127 17093
rect 0 17088 4127 17090
rect 0 17032 4066 17088
rect 4122 17032 4127 17088
rect 0 17030 4127 17032
rect 0 17000 480 17030
rect 4061 17027 4127 17030
rect 9765 16954 9831 16957
rect 19241 16954 19307 16957
rect 9765 16952 19307 16954
rect 9765 16896 9770 16952
rect 9826 16896 19246 16952
rect 19302 16896 19307 16952
rect 9765 16894 19307 16896
rect 9765 16891 9831 16894
rect 19241 16891 19307 16894
rect 20437 16954 20503 16957
rect 22320 16954 22800 16984
rect 20437 16952 22800 16954
rect 20437 16896 20442 16952
rect 20498 16896 22800 16952
rect 20437 16894 22800 16896
rect 20437 16891 20503 16894
rect 22320 16864 22800 16894
rect 7808 16752 8128 16753
rect 7808 16688 7816 16752
rect 7880 16688 7896 16752
rect 7960 16688 7976 16752
rect 8040 16688 8056 16752
rect 8120 16688 8128 16752
rect 7808 16687 8128 16688
rect 14672 16752 14992 16753
rect 14672 16688 14680 16752
rect 14744 16688 14760 16752
rect 14824 16688 14840 16752
rect 14904 16688 14920 16752
rect 14984 16688 14992 16752
rect 14672 16687 14992 16688
rect 20161 16410 20227 16413
rect 22320 16410 22800 16440
rect 20161 16408 22800 16410
rect 20161 16352 20166 16408
rect 20222 16352 22800 16408
rect 20161 16350 22800 16352
rect 20161 16347 20227 16350
rect 22320 16320 22800 16350
rect 4376 16208 4696 16209
rect 4376 16144 4384 16208
rect 4448 16144 4464 16208
rect 4528 16144 4544 16208
rect 4608 16144 4624 16208
rect 4688 16144 4696 16208
rect 4376 16143 4696 16144
rect 11240 16208 11560 16209
rect 11240 16144 11248 16208
rect 11312 16144 11328 16208
rect 11392 16144 11408 16208
rect 11472 16144 11488 16208
rect 11552 16144 11560 16208
rect 11240 16143 11560 16144
rect 18104 16208 18424 16209
rect 18104 16144 18112 16208
rect 18176 16144 18192 16208
rect 18256 16144 18272 16208
rect 18336 16144 18352 16208
rect 18416 16144 18424 16208
rect 18104 16143 18424 16144
rect 20069 16002 20135 16005
rect 22320 16002 22800 16032
rect 20069 16000 22800 16002
rect 20069 15944 20074 16000
rect 20130 15944 22800 16000
rect 20069 15942 22800 15944
rect 20069 15939 20135 15942
rect 22320 15912 22800 15942
rect 7808 15664 8128 15665
rect 7808 15600 7816 15664
rect 7880 15600 7896 15664
rect 7960 15600 7976 15664
rect 8040 15600 8056 15664
rect 8120 15600 8128 15664
rect 7808 15599 8128 15600
rect 14672 15664 14992 15665
rect 14672 15600 14680 15664
rect 14744 15600 14760 15664
rect 14824 15600 14840 15664
rect 14904 15600 14920 15664
rect 14984 15600 14992 15664
rect 14672 15599 14992 15600
rect 20437 15594 20503 15597
rect 22320 15594 22800 15624
rect 20437 15592 22800 15594
rect 20437 15536 20442 15592
rect 20498 15536 22800 15592
rect 20437 15534 22800 15536
rect 20437 15531 20503 15534
rect 22320 15504 22800 15534
rect 4376 15120 4696 15121
rect 4376 15056 4384 15120
rect 4448 15056 4464 15120
rect 4528 15056 4544 15120
rect 4608 15056 4624 15120
rect 4688 15056 4696 15120
rect 4376 15055 4696 15056
rect 11240 15120 11560 15121
rect 11240 15056 11248 15120
rect 11312 15056 11328 15120
rect 11392 15056 11408 15120
rect 11472 15056 11488 15120
rect 11552 15056 11560 15120
rect 11240 15055 11560 15056
rect 18104 15120 18424 15121
rect 18104 15056 18112 15120
rect 18176 15056 18192 15120
rect 18256 15056 18272 15120
rect 18336 15056 18352 15120
rect 18416 15056 18424 15120
rect 18104 15055 18424 15056
rect 20897 15050 20963 15053
rect 22320 15050 22800 15080
rect 20897 15048 22800 15050
rect 20897 14992 20902 15048
rect 20958 14992 22800 15048
rect 20897 14990 22800 14992
rect 20897 14987 20963 14990
rect 22320 14960 22800 14990
rect 20437 14642 20503 14645
rect 22320 14642 22800 14672
rect 20437 14640 22800 14642
rect 20437 14584 20442 14640
rect 20498 14584 22800 14640
rect 20437 14582 22800 14584
rect 20437 14579 20503 14582
rect 7808 14576 8128 14577
rect 7808 14512 7816 14576
rect 7880 14512 7896 14576
rect 7960 14512 7976 14576
rect 8040 14512 8056 14576
rect 8120 14512 8128 14576
rect 7808 14511 8128 14512
rect 14672 14576 14992 14577
rect 14672 14512 14680 14576
rect 14744 14512 14760 14576
rect 14824 14512 14840 14576
rect 14904 14512 14920 14576
rect 14984 14512 14992 14576
rect 22320 14552 22800 14582
rect 14672 14511 14992 14512
rect 19149 14234 19215 14237
rect 22320 14234 22800 14264
rect 19149 14232 22800 14234
rect 19149 14176 19154 14232
rect 19210 14176 22800 14232
rect 19149 14174 22800 14176
rect 19149 14171 19215 14174
rect 22320 14144 22800 14174
rect 4376 14032 4696 14033
rect 4376 13968 4384 14032
rect 4448 13968 4464 14032
rect 4528 13968 4544 14032
rect 4608 13968 4624 14032
rect 4688 13968 4696 14032
rect 4376 13967 4696 13968
rect 11240 14032 11560 14033
rect 11240 13968 11248 14032
rect 11312 13968 11328 14032
rect 11392 13968 11408 14032
rect 11472 13968 11488 14032
rect 11552 13968 11560 14032
rect 11240 13967 11560 13968
rect 18104 14032 18424 14033
rect 18104 13968 18112 14032
rect 18176 13968 18192 14032
rect 18256 13968 18272 14032
rect 18336 13968 18352 14032
rect 18416 13968 18424 14032
rect 18104 13967 18424 13968
rect 20713 13690 20779 13693
rect 22320 13690 22800 13720
rect 20713 13688 22800 13690
rect 20713 13632 20718 13688
rect 20774 13632 22800 13688
rect 20713 13630 22800 13632
rect 20713 13627 20779 13630
rect 22320 13600 22800 13630
rect 7808 13488 8128 13489
rect 7808 13424 7816 13488
rect 7880 13424 7896 13488
rect 7960 13424 7976 13488
rect 8040 13424 8056 13488
rect 8120 13424 8128 13488
rect 7808 13423 8128 13424
rect 14672 13488 14992 13489
rect 14672 13424 14680 13488
rect 14744 13424 14760 13488
rect 14824 13424 14840 13488
rect 14904 13424 14920 13488
rect 14984 13424 14992 13488
rect 14672 13423 14992 13424
rect 20069 13282 20135 13285
rect 22320 13282 22800 13312
rect 20069 13280 22800 13282
rect 20069 13224 20074 13280
rect 20130 13224 22800 13280
rect 20069 13222 22800 13224
rect 20069 13219 20135 13222
rect 22320 13192 22800 13222
rect 4376 12944 4696 12945
rect 4376 12880 4384 12944
rect 4448 12880 4464 12944
rect 4528 12880 4544 12944
rect 4608 12880 4624 12944
rect 4688 12880 4696 12944
rect 4376 12879 4696 12880
rect 11240 12944 11560 12945
rect 11240 12880 11248 12944
rect 11312 12880 11328 12944
rect 11392 12880 11408 12944
rect 11472 12880 11488 12944
rect 11552 12880 11560 12944
rect 11240 12879 11560 12880
rect 18104 12944 18424 12945
rect 18104 12880 18112 12944
rect 18176 12880 18192 12944
rect 18256 12880 18272 12944
rect 18336 12880 18352 12944
rect 18416 12880 18424 12944
rect 18104 12879 18424 12880
rect 19701 12874 19767 12877
rect 22320 12874 22800 12904
rect 19701 12872 22800 12874
rect 19701 12816 19706 12872
rect 19762 12816 22800 12872
rect 19701 12814 22800 12816
rect 19701 12811 19767 12814
rect 22320 12784 22800 12814
rect 7808 12400 8128 12401
rect 7808 12336 7816 12400
rect 7880 12336 7896 12400
rect 7960 12336 7976 12400
rect 8040 12336 8056 12400
rect 8120 12336 8128 12400
rect 7808 12335 8128 12336
rect 14672 12400 14992 12401
rect 14672 12336 14680 12400
rect 14744 12336 14760 12400
rect 14824 12336 14840 12400
rect 14904 12336 14920 12400
rect 14984 12336 14992 12400
rect 14672 12335 14992 12336
rect 19241 12330 19307 12333
rect 22320 12330 22800 12360
rect 19241 12328 22800 12330
rect 19241 12272 19246 12328
rect 19302 12272 22800 12328
rect 19241 12270 22800 12272
rect 19241 12267 19307 12270
rect 22320 12240 22800 12270
rect 20161 11922 20227 11925
rect 22320 11922 22800 11952
rect 20161 11920 22800 11922
rect 20161 11864 20166 11920
rect 20222 11864 22800 11920
rect 20161 11862 22800 11864
rect 20161 11859 20227 11862
rect 4376 11856 4696 11857
rect 4376 11792 4384 11856
rect 4448 11792 4464 11856
rect 4528 11792 4544 11856
rect 4608 11792 4624 11856
rect 4688 11792 4696 11856
rect 4376 11791 4696 11792
rect 11240 11856 11560 11857
rect 11240 11792 11248 11856
rect 11312 11792 11328 11856
rect 11392 11792 11408 11856
rect 11472 11792 11488 11856
rect 11552 11792 11560 11856
rect 11240 11791 11560 11792
rect 18104 11856 18424 11857
rect 18104 11792 18112 11856
rect 18176 11792 18192 11856
rect 18256 11792 18272 11856
rect 18336 11792 18352 11856
rect 18416 11792 18424 11856
rect 22320 11832 22800 11862
rect 18104 11791 18424 11792
rect 19885 11514 19951 11517
rect 22320 11514 22800 11544
rect 19885 11512 22800 11514
rect 19885 11456 19890 11512
rect 19946 11456 22800 11512
rect 19885 11454 22800 11456
rect 19885 11451 19951 11454
rect 22320 11424 22800 11454
rect 7808 11312 8128 11313
rect 7808 11248 7816 11312
rect 7880 11248 7896 11312
rect 7960 11248 7976 11312
rect 8040 11248 8056 11312
rect 8120 11248 8128 11312
rect 7808 11247 8128 11248
rect 14672 11312 14992 11313
rect 14672 11248 14680 11312
rect 14744 11248 14760 11312
rect 14824 11248 14840 11312
rect 14904 11248 14920 11312
rect 14984 11248 14992 11312
rect 14672 11247 14992 11248
rect 20437 10970 20503 10973
rect 22320 10970 22800 11000
rect 20437 10968 22800 10970
rect 20437 10912 20442 10968
rect 20498 10912 22800 10968
rect 20437 10910 22800 10912
rect 20437 10907 20503 10910
rect 22320 10880 22800 10910
rect 4376 10768 4696 10769
rect 4376 10704 4384 10768
rect 4448 10704 4464 10768
rect 4528 10704 4544 10768
rect 4608 10704 4624 10768
rect 4688 10704 4696 10768
rect 4376 10703 4696 10704
rect 11240 10768 11560 10769
rect 11240 10704 11248 10768
rect 11312 10704 11328 10768
rect 11392 10704 11408 10768
rect 11472 10704 11488 10768
rect 11552 10704 11560 10768
rect 11240 10703 11560 10704
rect 18104 10768 18424 10769
rect 18104 10704 18112 10768
rect 18176 10704 18192 10768
rect 18256 10704 18272 10768
rect 18336 10704 18352 10768
rect 18416 10704 18424 10768
rect 18104 10703 18424 10704
rect 20529 10562 20595 10565
rect 22320 10562 22800 10592
rect 20529 10560 22800 10562
rect 20529 10504 20534 10560
rect 20590 10504 22800 10560
rect 20529 10502 22800 10504
rect 20529 10499 20595 10502
rect 22320 10472 22800 10502
rect 7808 10224 8128 10225
rect 7808 10160 7816 10224
rect 7880 10160 7896 10224
rect 7960 10160 7976 10224
rect 8040 10160 8056 10224
rect 8120 10160 8128 10224
rect 7808 10159 8128 10160
rect 14672 10224 14992 10225
rect 14672 10160 14680 10224
rect 14744 10160 14760 10224
rect 14824 10160 14840 10224
rect 14904 10160 14920 10224
rect 14984 10160 14992 10224
rect 14672 10159 14992 10160
rect 19057 10018 19123 10021
rect 22320 10018 22800 10048
rect 19057 10016 22800 10018
rect 19057 9960 19062 10016
rect 19118 9960 22800 10016
rect 19057 9958 22800 9960
rect 19057 9955 19123 9958
rect 22320 9928 22800 9958
rect 4376 9680 4696 9681
rect 4376 9616 4384 9680
rect 4448 9616 4464 9680
rect 4528 9616 4544 9680
rect 4608 9616 4624 9680
rect 4688 9616 4696 9680
rect 4376 9615 4696 9616
rect 11240 9680 11560 9681
rect 11240 9616 11248 9680
rect 11312 9616 11328 9680
rect 11392 9616 11408 9680
rect 11472 9616 11488 9680
rect 11552 9616 11560 9680
rect 11240 9615 11560 9616
rect 18104 9680 18424 9681
rect 18104 9616 18112 9680
rect 18176 9616 18192 9680
rect 18256 9616 18272 9680
rect 18336 9616 18352 9680
rect 18416 9616 18424 9680
rect 18104 9615 18424 9616
rect 20253 9610 20319 9613
rect 22320 9610 22800 9640
rect 20253 9608 22800 9610
rect 20253 9552 20258 9608
rect 20314 9552 22800 9608
rect 20253 9550 22800 9552
rect 20253 9547 20319 9550
rect 22320 9520 22800 9550
rect 14365 9474 14431 9477
rect 14230 9472 14431 9474
rect 14230 9416 14370 9472
rect 14426 9416 14431 9472
rect 14230 9414 14431 9416
rect 14230 9338 14290 9414
rect 14365 9411 14431 9414
rect 18781 9338 18847 9341
rect 14230 9336 18847 9338
rect 14230 9280 18786 9336
rect 18842 9280 18847 9336
rect 14230 9278 18847 9280
rect 18781 9275 18847 9278
rect 20529 9202 20595 9205
rect 22320 9202 22800 9232
rect 20529 9200 22800 9202
rect 20529 9144 20534 9200
rect 20590 9144 22800 9200
rect 20529 9142 22800 9144
rect 20529 9139 20595 9142
rect 7808 9136 8128 9137
rect 7808 9072 7816 9136
rect 7880 9072 7896 9136
rect 7960 9072 7976 9136
rect 8040 9072 8056 9136
rect 8120 9072 8128 9136
rect 7808 9071 8128 9072
rect 14672 9136 14992 9137
rect 14672 9072 14680 9136
rect 14744 9072 14760 9136
rect 14824 9072 14840 9136
rect 14904 9072 14920 9136
rect 14984 9072 14992 9136
rect 22320 9112 22800 9142
rect 14672 9071 14992 9072
rect 20529 8658 20595 8661
rect 22320 8658 22800 8688
rect 20529 8656 22800 8658
rect 20529 8600 20534 8656
rect 20590 8600 22800 8656
rect 20529 8598 22800 8600
rect 20529 8595 20595 8598
rect 4376 8592 4696 8593
rect 4376 8528 4384 8592
rect 4448 8528 4464 8592
rect 4528 8528 4544 8592
rect 4608 8528 4624 8592
rect 4688 8528 4696 8592
rect 4376 8527 4696 8528
rect 11240 8592 11560 8593
rect 11240 8528 11248 8592
rect 11312 8528 11328 8592
rect 11392 8528 11408 8592
rect 11472 8528 11488 8592
rect 11552 8528 11560 8592
rect 11240 8527 11560 8528
rect 18104 8592 18424 8593
rect 18104 8528 18112 8592
rect 18176 8528 18192 8592
rect 18256 8528 18272 8592
rect 18336 8528 18352 8592
rect 18416 8528 18424 8592
rect 22320 8568 22800 8598
rect 18104 8527 18424 8528
rect 19977 8250 20043 8253
rect 22320 8250 22800 8280
rect 19977 8248 22800 8250
rect 19977 8192 19982 8248
rect 20038 8192 22800 8248
rect 19977 8190 22800 8192
rect 19977 8187 20043 8190
rect 22320 8160 22800 8190
rect 7808 8048 8128 8049
rect 7808 7984 7816 8048
rect 7880 7984 7896 8048
rect 7960 7984 7976 8048
rect 8040 7984 8056 8048
rect 8120 7984 8128 8048
rect 7808 7983 8128 7984
rect 14672 8048 14992 8049
rect 14672 7984 14680 8048
rect 14744 7984 14760 8048
rect 14824 7984 14840 8048
rect 14904 7984 14920 8048
rect 14984 7984 14992 8048
rect 14672 7983 14992 7984
rect 20253 7842 20319 7845
rect 22320 7842 22800 7872
rect 20253 7840 22800 7842
rect 20253 7784 20258 7840
rect 20314 7784 22800 7840
rect 20253 7782 22800 7784
rect 20253 7779 20319 7782
rect 22320 7752 22800 7782
rect 4376 7504 4696 7505
rect 4376 7440 4384 7504
rect 4448 7440 4464 7504
rect 4528 7440 4544 7504
rect 4608 7440 4624 7504
rect 4688 7440 4696 7504
rect 4376 7439 4696 7440
rect 11240 7504 11560 7505
rect 11240 7440 11248 7504
rect 11312 7440 11328 7504
rect 11392 7440 11408 7504
rect 11472 7440 11488 7504
rect 11552 7440 11560 7504
rect 11240 7439 11560 7440
rect 18104 7504 18424 7505
rect 18104 7440 18112 7504
rect 18176 7440 18192 7504
rect 18256 7440 18272 7504
rect 18336 7440 18352 7504
rect 18416 7440 18424 7504
rect 18104 7439 18424 7440
rect 20529 7298 20595 7301
rect 22320 7298 22800 7328
rect 20529 7296 22800 7298
rect 20529 7240 20534 7296
rect 20590 7240 22800 7296
rect 20529 7238 22800 7240
rect 20529 7235 20595 7238
rect 22320 7208 22800 7238
rect 7808 6960 8128 6961
rect 7808 6896 7816 6960
rect 7880 6896 7896 6960
rect 7960 6896 7976 6960
rect 8040 6896 8056 6960
rect 8120 6896 8128 6960
rect 7808 6895 8128 6896
rect 14672 6960 14992 6961
rect 14672 6896 14680 6960
rect 14744 6896 14760 6960
rect 14824 6896 14840 6960
rect 14904 6896 14920 6960
rect 14984 6896 14992 6960
rect 14672 6895 14992 6896
rect 19977 6890 20043 6893
rect 22320 6890 22800 6920
rect 19977 6888 22800 6890
rect 19977 6832 19982 6888
rect 20038 6832 22800 6888
rect 19977 6830 22800 6832
rect 19977 6827 20043 6830
rect 22320 6800 22800 6830
rect 18505 6482 18571 6485
rect 22320 6482 22800 6512
rect 18505 6480 22800 6482
rect 18505 6424 18510 6480
rect 18566 6424 22800 6480
rect 18505 6422 22800 6424
rect 18505 6419 18571 6422
rect 4376 6416 4696 6417
rect 4376 6352 4384 6416
rect 4448 6352 4464 6416
rect 4528 6352 4544 6416
rect 4608 6352 4624 6416
rect 4688 6352 4696 6416
rect 4376 6351 4696 6352
rect 11240 6416 11560 6417
rect 11240 6352 11248 6416
rect 11312 6352 11328 6416
rect 11392 6352 11408 6416
rect 11472 6352 11488 6416
rect 11552 6352 11560 6416
rect 11240 6351 11560 6352
rect 18104 6416 18424 6417
rect 18104 6352 18112 6416
rect 18176 6352 18192 6416
rect 18256 6352 18272 6416
rect 18336 6352 18352 6416
rect 18416 6352 18424 6416
rect 22320 6392 22800 6422
rect 18104 6351 18424 6352
rect 20529 5938 20595 5941
rect 22320 5938 22800 5968
rect 20529 5936 22800 5938
rect 20529 5880 20534 5936
rect 20590 5880 22800 5936
rect 20529 5878 22800 5880
rect 20529 5875 20595 5878
rect 7808 5872 8128 5873
rect 7808 5808 7816 5872
rect 7880 5808 7896 5872
rect 7960 5808 7976 5872
rect 8040 5808 8056 5872
rect 8120 5808 8128 5872
rect 7808 5807 8128 5808
rect 14672 5872 14992 5873
rect 14672 5808 14680 5872
rect 14744 5808 14760 5872
rect 14824 5808 14840 5872
rect 14904 5808 14920 5872
rect 14984 5808 14992 5872
rect 22320 5848 22800 5878
rect 14672 5807 14992 5808
rect 0 5666 480 5696
rect 4061 5666 4127 5669
rect 0 5664 4127 5666
rect 0 5608 4066 5664
rect 4122 5608 4127 5664
rect 0 5606 4127 5608
rect 0 5576 480 5606
rect 4061 5603 4127 5606
rect 18597 5530 18663 5533
rect 22320 5530 22800 5560
rect 18597 5528 22800 5530
rect 18597 5472 18602 5528
rect 18658 5472 22800 5528
rect 18597 5470 22800 5472
rect 18597 5467 18663 5470
rect 22320 5440 22800 5470
rect 4376 5328 4696 5329
rect 4376 5264 4384 5328
rect 4448 5264 4464 5328
rect 4528 5264 4544 5328
rect 4608 5264 4624 5328
rect 4688 5264 4696 5328
rect 4376 5263 4696 5264
rect 11240 5328 11560 5329
rect 11240 5264 11248 5328
rect 11312 5264 11328 5328
rect 11392 5264 11408 5328
rect 11472 5264 11488 5328
rect 11552 5264 11560 5328
rect 11240 5263 11560 5264
rect 18104 5328 18424 5329
rect 18104 5264 18112 5328
rect 18176 5264 18192 5328
rect 18256 5264 18272 5328
rect 18336 5264 18352 5328
rect 18416 5264 18424 5328
rect 18104 5263 18424 5264
rect 20529 4986 20595 4989
rect 22320 4986 22800 5016
rect 20529 4984 22800 4986
rect 20529 4928 20534 4984
rect 20590 4928 22800 4984
rect 20529 4926 22800 4928
rect 20529 4923 20595 4926
rect 22320 4896 22800 4926
rect 7808 4784 8128 4785
rect 7808 4720 7816 4784
rect 7880 4720 7896 4784
rect 7960 4720 7976 4784
rect 8040 4720 8056 4784
rect 8120 4720 8128 4784
rect 7808 4719 8128 4720
rect 14672 4784 14992 4785
rect 14672 4720 14680 4784
rect 14744 4720 14760 4784
rect 14824 4720 14840 4784
rect 14904 4720 14920 4784
rect 14984 4720 14992 4784
rect 14672 4719 14992 4720
rect 17953 4578 18019 4581
rect 22320 4578 22800 4608
rect 17953 4576 22800 4578
rect 17953 4520 17958 4576
rect 18014 4520 22800 4576
rect 17953 4518 22800 4520
rect 17953 4515 18019 4518
rect 22320 4488 22800 4518
rect 4376 4240 4696 4241
rect 4376 4176 4384 4240
rect 4448 4176 4464 4240
rect 4528 4176 4544 4240
rect 4608 4176 4624 4240
rect 4688 4176 4696 4240
rect 4376 4175 4696 4176
rect 11240 4240 11560 4241
rect 11240 4176 11248 4240
rect 11312 4176 11328 4240
rect 11392 4176 11408 4240
rect 11472 4176 11488 4240
rect 11552 4176 11560 4240
rect 11240 4175 11560 4176
rect 18104 4240 18424 4241
rect 18104 4176 18112 4240
rect 18176 4176 18192 4240
rect 18256 4176 18272 4240
rect 18336 4176 18352 4240
rect 18416 4176 18424 4240
rect 18104 4175 18424 4176
rect 20529 4170 20595 4173
rect 22320 4170 22800 4200
rect 20529 4168 22800 4170
rect 20529 4112 20534 4168
rect 20590 4112 22800 4168
rect 20529 4110 22800 4112
rect 20529 4107 20595 4110
rect 22320 4080 22800 4110
rect 7808 3696 8128 3697
rect 7808 3632 7816 3696
rect 7880 3632 7896 3696
rect 7960 3632 7976 3696
rect 8040 3632 8056 3696
rect 8120 3632 8128 3696
rect 7808 3631 8128 3632
rect 14672 3696 14992 3697
rect 14672 3632 14680 3696
rect 14744 3632 14760 3696
rect 14824 3632 14840 3696
rect 14904 3632 14920 3696
rect 14984 3632 14992 3696
rect 14672 3631 14992 3632
rect 17861 3626 17927 3629
rect 22320 3626 22800 3656
rect 17861 3624 22800 3626
rect 17861 3568 17866 3624
rect 17922 3568 22800 3624
rect 17861 3566 22800 3568
rect 17861 3563 17927 3566
rect 22320 3536 22800 3566
rect 18781 3218 18847 3221
rect 22320 3218 22800 3248
rect 18781 3216 22800 3218
rect 18781 3160 18786 3216
rect 18842 3160 22800 3216
rect 18781 3158 22800 3160
rect 18781 3155 18847 3158
rect 4376 3152 4696 3153
rect 4376 3088 4384 3152
rect 4448 3088 4464 3152
rect 4528 3088 4544 3152
rect 4608 3088 4624 3152
rect 4688 3088 4696 3152
rect 4376 3087 4696 3088
rect 11240 3152 11560 3153
rect 11240 3088 11248 3152
rect 11312 3088 11328 3152
rect 11392 3088 11408 3152
rect 11472 3088 11488 3152
rect 11552 3088 11560 3152
rect 11240 3087 11560 3088
rect 18104 3152 18424 3153
rect 18104 3088 18112 3152
rect 18176 3088 18192 3152
rect 18256 3088 18272 3152
rect 18336 3088 18352 3152
rect 18416 3088 18424 3152
rect 22320 3128 22800 3158
rect 18104 3087 18424 3088
rect 19057 2810 19123 2813
rect 22320 2810 22800 2840
rect 19057 2808 22800 2810
rect 19057 2752 19062 2808
rect 19118 2752 22800 2808
rect 19057 2750 22800 2752
rect 19057 2747 19123 2750
rect 22320 2720 22800 2750
rect 7808 2608 8128 2609
rect 7808 2544 7816 2608
rect 7880 2544 7896 2608
rect 7960 2544 7976 2608
rect 8040 2544 8056 2608
rect 8120 2544 8128 2608
rect 7808 2543 8128 2544
rect 14672 2608 14992 2609
rect 14672 2544 14680 2608
rect 14744 2544 14760 2608
rect 14824 2544 14840 2608
rect 14904 2544 14920 2608
rect 14984 2544 14992 2608
rect 14672 2543 14992 2544
rect 18965 2266 19031 2269
rect 22320 2266 22800 2296
rect 18965 2264 22800 2266
rect 18965 2208 18970 2264
rect 19026 2208 22800 2264
rect 18965 2206 22800 2208
rect 18965 2203 19031 2206
rect 22320 2176 22800 2206
rect 4376 2064 4696 2065
rect 4376 2000 4384 2064
rect 4448 2000 4464 2064
rect 4528 2000 4544 2064
rect 4608 2000 4624 2064
rect 4688 2000 4696 2064
rect 4376 1999 4696 2000
rect 11240 2064 11560 2065
rect 11240 2000 11248 2064
rect 11312 2000 11328 2064
rect 11392 2000 11408 2064
rect 11472 2000 11488 2064
rect 11552 2000 11560 2064
rect 11240 1999 11560 2000
rect 18104 2064 18424 2065
rect 18104 2000 18112 2064
rect 18176 2000 18192 2064
rect 18256 2000 18272 2064
rect 18336 2000 18352 2064
rect 18416 2000 18424 2064
rect 18104 1999 18424 2000
rect 18689 1858 18755 1861
rect 22320 1858 22800 1888
rect 18689 1856 22800 1858
rect 18689 1800 18694 1856
rect 18750 1800 22800 1856
rect 18689 1798 22800 1800
rect 18689 1795 18755 1798
rect 22320 1768 22800 1798
rect 17953 1450 18019 1453
rect 22320 1450 22800 1480
rect 17953 1448 22800 1450
rect 17953 1392 17958 1448
rect 18014 1392 22800 1448
rect 17953 1390 22800 1392
rect 17953 1387 18019 1390
rect 22320 1360 22800 1390
rect 17953 906 18019 909
rect 22320 906 22800 936
rect 17953 904 22800 906
rect 17953 848 17958 904
rect 18014 848 22800 904
rect 17953 846 22800 848
rect 17953 843 18019 846
rect 22320 816 22800 846
rect 18873 498 18939 501
rect 22320 498 22800 528
rect 18873 496 22800 498
rect 18873 440 18878 496
rect 18934 440 22800 496
rect 18873 438 22800 440
rect 18873 435 18939 438
rect 22320 408 22800 438
rect 17217 90 17283 93
rect 22320 90 22800 120
rect 17217 88 22800 90
rect 17217 32 17222 88
rect 17278 32 22800 88
rect 17217 30 22800 32
rect 17217 27 17283 30
rect 22320 0 22800 30
<< via3 >>
rect 7816 20012 7880 20016
rect 7816 19956 7820 20012
rect 7820 19956 7876 20012
rect 7876 19956 7880 20012
rect 7816 19952 7880 19956
rect 7896 20012 7960 20016
rect 7896 19956 7900 20012
rect 7900 19956 7956 20012
rect 7956 19956 7960 20012
rect 7896 19952 7960 19956
rect 7976 20012 8040 20016
rect 7976 19956 7980 20012
rect 7980 19956 8036 20012
rect 8036 19956 8040 20012
rect 7976 19952 8040 19956
rect 8056 20012 8120 20016
rect 8056 19956 8060 20012
rect 8060 19956 8116 20012
rect 8116 19956 8120 20012
rect 8056 19952 8120 19956
rect 14680 20012 14744 20016
rect 14680 19956 14684 20012
rect 14684 19956 14740 20012
rect 14740 19956 14744 20012
rect 14680 19952 14744 19956
rect 14760 20012 14824 20016
rect 14760 19956 14764 20012
rect 14764 19956 14820 20012
rect 14820 19956 14824 20012
rect 14760 19952 14824 19956
rect 14840 20012 14904 20016
rect 14840 19956 14844 20012
rect 14844 19956 14900 20012
rect 14900 19956 14904 20012
rect 14840 19952 14904 19956
rect 14920 20012 14984 20016
rect 14920 19956 14924 20012
rect 14924 19956 14980 20012
rect 14980 19956 14984 20012
rect 14920 19952 14984 19956
rect 4384 19468 4448 19472
rect 4384 19412 4388 19468
rect 4388 19412 4444 19468
rect 4444 19412 4448 19468
rect 4384 19408 4448 19412
rect 4464 19468 4528 19472
rect 4464 19412 4468 19468
rect 4468 19412 4524 19468
rect 4524 19412 4528 19468
rect 4464 19408 4528 19412
rect 4544 19468 4608 19472
rect 4544 19412 4548 19468
rect 4548 19412 4604 19468
rect 4604 19412 4608 19468
rect 4544 19408 4608 19412
rect 4624 19468 4688 19472
rect 4624 19412 4628 19468
rect 4628 19412 4684 19468
rect 4684 19412 4688 19468
rect 4624 19408 4688 19412
rect 11248 19468 11312 19472
rect 11248 19412 11252 19468
rect 11252 19412 11308 19468
rect 11308 19412 11312 19468
rect 11248 19408 11312 19412
rect 11328 19468 11392 19472
rect 11328 19412 11332 19468
rect 11332 19412 11388 19468
rect 11388 19412 11392 19468
rect 11328 19408 11392 19412
rect 11408 19468 11472 19472
rect 11408 19412 11412 19468
rect 11412 19412 11468 19468
rect 11468 19412 11472 19468
rect 11408 19408 11472 19412
rect 11488 19468 11552 19472
rect 11488 19412 11492 19468
rect 11492 19412 11548 19468
rect 11548 19412 11552 19468
rect 11488 19408 11552 19412
rect 18112 19468 18176 19472
rect 18112 19412 18116 19468
rect 18116 19412 18172 19468
rect 18172 19412 18176 19468
rect 18112 19408 18176 19412
rect 18192 19468 18256 19472
rect 18192 19412 18196 19468
rect 18196 19412 18252 19468
rect 18252 19412 18256 19468
rect 18192 19408 18256 19412
rect 18272 19468 18336 19472
rect 18272 19412 18276 19468
rect 18276 19412 18332 19468
rect 18332 19412 18336 19468
rect 18272 19408 18336 19412
rect 18352 19468 18416 19472
rect 18352 19412 18356 19468
rect 18356 19412 18412 19468
rect 18412 19412 18416 19468
rect 18352 19408 18416 19412
rect 7816 18924 7880 18928
rect 7816 18868 7820 18924
rect 7820 18868 7876 18924
rect 7876 18868 7880 18924
rect 7816 18864 7880 18868
rect 7896 18924 7960 18928
rect 7896 18868 7900 18924
rect 7900 18868 7956 18924
rect 7956 18868 7960 18924
rect 7896 18864 7960 18868
rect 7976 18924 8040 18928
rect 7976 18868 7980 18924
rect 7980 18868 8036 18924
rect 8036 18868 8040 18924
rect 7976 18864 8040 18868
rect 8056 18924 8120 18928
rect 8056 18868 8060 18924
rect 8060 18868 8116 18924
rect 8116 18868 8120 18924
rect 8056 18864 8120 18868
rect 14680 18924 14744 18928
rect 14680 18868 14684 18924
rect 14684 18868 14740 18924
rect 14740 18868 14744 18924
rect 14680 18864 14744 18868
rect 14760 18924 14824 18928
rect 14760 18868 14764 18924
rect 14764 18868 14820 18924
rect 14820 18868 14824 18924
rect 14760 18864 14824 18868
rect 14840 18924 14904 18928
rect 14840 18868 14844 18924
rect 14844 18868 14900 18924
rect 14900 18868 14904 18924
rect 14840 18864 14904 18868
rect 14920 18924 14984 18928
rect 14920 18868 14924 18924
rect 14924 18868 14980 18924
rect 14980 18868 14984 18924
rect 14920 18864 14984 18868
rect 4384 18380 4448 18384
rect 4384 18324 4388 18380
rect 4388 18324 4444 18380
rect 4444 18324 4448 18380
rect 4384 18320 4448 18324
rect 4464 18380 4528 18384
rect 4464 18324 4468 18380
rect 4468 18324 4524 18380
rect 4524 18324 4528 18380
rect 4464 18320 4528 18324
rect 4544 18380 4608 18384
rect 4544 18324 4548 18380
rect 4548 18324 4604 18380
rect 4604 18324 4608 18380
rect 4544 18320 4608 18324
rect 4624 18380 4688 18384
rect 4624 18324 4628 18380
rect 4628 18324 4684 18380
rect 4684 18324 4688 18380
rect 4624 18320 4688 18324
rect 11248 18380 11312 18384
rect 11248 18324 11252 18380
rect 11252 18324 11308 18380
rect 11308 18324 11312 18380
rect 11248 18320 11312 18324
rect 11328 18380 11392 18384
rect 11328 18324 11332 18380
rect 11332 18324 11388 18380
rect 11388 18324 11392 18380
rect 11328 18320 11392 18324
rect 11408 18380 11472 18384
rect 11408 18324 11412 18380
rect 11412 18324 11468 18380
rect 11468 18324 11472 18380
rect 11408 18320 11472 18324
rect 11488 18380 11552 18384
rect 11488 18324 11492 18380
rect 11492 18324 11548 18380
rect 11548 18324 11552 18380
rect 11488 18320 11552 18324
rect 18112 18380 18176 18384
rect 18112 18324 18116 18380
rect 18116 18324 18172 18380
rect 18172 18324 18176 18380
rect 18112 18320 18176 18324
rect 18192 18380 18256 18384
rect 18192 18324 18196 18380
rect 18196 18324 18252 18380
rect 18252 18324 18256 18380
rect 18192 18320 18256 18324
rect 18272 18380 18336 18384
rect 18272 18324 18276 18380
rect 18276 18324 18332 18380
rect 18332 18324 18336 18380
rect 18272 18320 18336 18324
rect 18352 18380 18416 18384
rect 18352 18324 18356 18380
rect 18356 18324 18412 18380
rect 18412 18324 18416 18380
rect 18352 18320 18416 18324
rect 7816 17836 7880 17840
rect 7816 17780 7820 17836
rect 7820 17780 7876 17836
rect 7876 17780 7880 17836
rect 7816 17776 7880 17780
rect 7896 17836 7960 17840
rect 7896 17780 7900 17836
rect 7900 17780 7956 17836
rect 7956 17780 7960 17836
rect 7896 17776 7960 17780
rect 7976 17836 8040 17840
rect 7976 17780 7980 17836
rect 7980 17780 8036 17836
rect 8036 17780 8040 17836
rect 7976 17776 8040 17780
rect 8056 17836 8120 17840
rect 8056 17780 8060 17836
rect 8060 17780 8116 17836
rect 8116 17780 8120 17836
rect 8056 17776 8120 17780
rect 14680 17836 14744 17840
rect 14680 17780 14684 17836
rect 14684 17780 14740 17836
rect 14740 17780 14744 17836
rect 14680 17776 14744 17780
rect 14760 17836 14824 17840
rect 14760 17780 14764 17836
rect 14764 17780 14820 17836
rect 14820 17780 14824 17836
rect 14760 17776 14824 17780
rect 14840 17836 14904 17840
rect 14840 17780 14844 17836
rect 14844 17780 14900 17836
rect 14900 17780 14904 17836
rect 14840 17776 14904 17780
rect 14920 17836 14984 17840
rect 14920 17780 14924 17836
rect 14924 17780 14980 17836
rect 14980 17780 14984 17836
rect 14920 17776 14984 17780
rect 4384 17292 4448 17296
rect 4384 17236 4388 17292
rect 4388 17236 4444 17292
rect 4444 17236 4448 17292
rect 4384 17232 4448 17236
rect 4464 17292 4528 17296
rect 4464 17236 4468 17292
rect 4468 17236 4524 17292
rect 4524 17236 4528 17292
rect 4464 17232 4528 17236
rect 4544 17292 4608 17296
rect 4544 17236 4548 17292
rect 4548 17236 4604 17292
rect 4604 17236 4608 17292
rect 4544 17232 4608 17236
rect 4624 17292 4688 17296
rect 4624 17236 4628 17292
rect 4628 17236 4684 17292
rect 4684 17236 4688 17292
rect 4624 17232 4688 17236
rect 11248 17292 11312 17296
rect 11248 17236 11252 17292
rect 11252 17236 11308 17292
rect 11308 17236 11312 17292
rect 11248 17232 11312 17236
rect 11328 17292 11392 17296
rect 11328 17236 11332 17292
rect 11332 17236 11388 17292
rect 11388 17236 11392 17292
rect 11328 17232 11392 17236
rect 11408 17292 11472 17296
rect 11408 17236 11412 17292
rect 11412 17236 11468 17292
rect 11468 17236 11472 17292
rect 11408 17232 11472 17236
rect 11488 17292 11552 17296
rect 11488 17236 11492 17292
rect 11492 17236 11548 17292
rect 11548 17236 11552 17292
rect 11488 17232 11552 17236
rect 18112 17292 18176 17296
rect 18112 17236 18116 17292
rect 18116 17236 18172 17292
rect 18172 17236 18176 17292
rect 18112 17232 18176 17236
rect 18192 17292 18256 17296
rect 18192 17236 18196 17292
rect 18196 17236 18252 17292
rect 18252 17236 18256 17292
rect 18192 17232 18256 17236
rect 18272 17292 18336 17296
rect 18272 17236 18276 17292
rect 18276 17236 18332 17292
rect 18332 17236 18336 17292
rect 18272 17232 18336 17236
rect 18352 17292 18416 17296
rect 18352 17236 18356 17292
rect 18356 17236 18412 17292
rect 18412 17236 18416 17292
rect 18352 17232 18416 17236
rect 7816 16748 7880 16752
rect 7816 16692 7820 16748
rect 7820 16692 7876 16748
rect 7876 16692 7880 16748
rect 7816 16688 7880 16692
rect 7896 16748 7960 16752
rect 7896 16692 7900 16748
rect 7900 16692 7956 16748
rect 7956 16692 7960 16748
rect 7896 16688 7960 16692
rect 7976 16748 8040 16752
rect 7976 16692 7980 16748
rect 7980 16692 8036 16748
rect 8036 16692 8040 16748
rect 7976 16688 8040 16692
rect 8056 16748 8120 16752
rect 8056 16692 8060 16748
rect 8060 16692 8116 16748
rect 8116 16692 8120 16748
rect 8056 16688 8120 16692
rect 14680 16748 14744 16752
rect 14680 16692 14684 16748
rect 14684 16692 14740 16748
rect 14740 16692 14744 16748
rect 14680 16688 14744 16692
rect 14760 16748 14824 16752
rect 14760 16692 14764 16748
rect 14764 16692 14820 16748
rect 14820 16692 14824 16748
rect 14760 16688 14824 16692
rect 14840 16748 14904 16752
rect 14840 16692 14844 16748
rect 14844 16692 14900 16748
rect 14900 16692 14904 16748
rect 14840 16688 14904 16692
rect 14920 16748 14984 16752
rect 14920 16692 14924 16748
rect 14924 16692 14980 16748
rect 14980 16692 14984 16748
rect 14920 16688 14984 16692
rect 4384 16204 4448 16208
rect 4384 16148 4388 16204
rect 4388 16148 4444 16204
rect 4444 16148 4448 16204
rect 4384 16144 4448 16148
rect 4464 16204 4528 16208
rect 4464 16148 4468 16204
rect 4468 16148 4524 16204
rect 4524 16148 4528 16204
rect 4464 16144 4528 16148
rect 4544 16204 4608 16208
rect 4544 16148 4548 16204
rect 4548 16148 4604 16204
rect 4604 16148 4608 16204
rect 4544 16144 4608 16148
rect 4624 16204 4688 16208
rect 4624 16148 4628 16204
rect 4628 16148 4684 16204
rect 4684 16148 4688 16204
rect 4624 16144 4688 16148
rect 11248 16204 11312 16208
rect 11248 16148 11252 16204
rect 11252 16148 11308 16204
rect 11308 16148 11312 16204
rect 11248 16144 11312 16148
rect 11328 16204 11392 16208
rect 11328 16148 11332 16204
rect 11332 16148 11388 16204
rect 11388 16148 11392 16204
rect 11328 16144 11392 16148
rect 11408 16204 11472 16208
rect 11408 16148 11412 16204
rect 11412 16148 11468 16204
rect 11468 16148 11472 16204
rect 11408 16144 11472 16148
rect 11488 16204 11552 16208
rect 11488 16148 11492 16204
rect 11492 16148 11548 16204
rect 11548 16148 11552 16204
rect 11488 16144 11552 16148
rect 18112 16204 18176 16208
rect 18112 16148 18116 16204
rect 18116 16148 18172 16204
rect 18172 16148 18176 16204
rect 18112 16144 18176 16148
rect 18192 16204 18256 16208
rect 18192 16148 18196 16204
rect 18196 16148 18252 16204
rect 18252 16148 18256 16204
rect 18192 16144 18256 16148
rect 18272 16204 18336 16208
rect 18272 16148 18276 16204
rect 18276 16148 18332 16204
rect 18332 16148 18336 16204
rect 18272 16144 18336 16148
rect 18352 16204 18416 16208
rect 18352 16148 18356 16204
rect 18356 16148 18412 16204
rect 18412 16148 18416 16204
rect 18352 16144 18416 16148
rect 7816 15660 7880 15664
rect 7816 15604 7820 15660
rect 7820 15604 7876 15660
rect 7876 15604 7880 15660
rect 7816 15600 7880 15604
rect 7896 15660 7960 15664
rect 7896 15604 7900 15660
rect 7900 15604 7956 15660
rect 7956 15604 7960 15660
rect 7896 15600 7960 15604
rect 7976 15660 8040 15664
rect 7976 15604 7980 15660
rect 7980 15604 8036 15660
rect 8036 15604 8040 15660
rect 7976 15600 8040 15604
rect 8056 15660 8120 15664
rect 8056 15604 8060 15660
rect 8060 15604 8116 15660
rect 8116 15604 8120 15660
rect 8056 15600 8120 15604
rect 14680 15660 14744 15664
rect 14680 15604 14684 15660
rect 14684 15604 14740 15660
rect 14740 15604 14744 15660
rect 14680 15600 14744 15604
rect 14760 15660 14824 15664
rect 14760 15604 14764 15660
rect 14764 15604 14820 15660
rect 14820 15604 14824 15660
rect 14760 15600 14824 15604
rect 14840 15660 14904 15664
rect 14840 15604 14844 15660
rect 14844 15604 14900 15660
rect 14900 15604 14904 15660
rect 14840 15600 14904 15604
rect 14920 15660 14984 15664
rect 14920 15604 14924 15660
rect 14924 15604 14980 15660
rect 14980 15604 14984 15660
rect 14920 15600 14984 15604
rect 4384 15116 4448 15120
rect 4384 15060 4388 15116
rect 4388 15060 4444 15116
rect 4444 15060 4448 15116
rect 4384 15056 4448 15060
rect 4464 15116 4528 15120
rect 4464 15060 4468 15116
rect 4468 15060 4524 15116
rect 4524 15060 4528 15116
rect 4464 15056 4528 15060
rect 4544 15116 4608 15120
rect 4544 15060 4548 15116
rect 4548 15060 4604 15116
rect 4604 15060 4608 15116
rect 4544 15056 4608 15060
rect 4624 15116 4688 15120
rect 4624 15060 4628 15116
rect 4628 15060 4684 15116
rect 4684 15060 4688 15116
rect 4624 15056 4688 15060
rect 11248 15116 11312 15120
rect 11248 15060 11252 15116
rect 11252 15060 11308 15116
rect 11308 15060 11312 15116
rect 11248 15056 11312 15060
rect 11328 15116 11392 15120
rect 11328 15060 11332 15116
rect 11332 15060 11388 15116
rect 11388 15060 11392 15116
rect 11328 15056 11392 15060
rect 11408 15116 11472 15120
rect 11408 15060 11412 15116
rect 11412 15060 11468 15116
rect 11468 15060 11472 15116
rect 11408 15056 11472 15060
rect 11488 15116 11552 15120
rect 11488 15060 11492 15116
rect 11492 15060 11548 15116
rect 11548 15060 11552 15116
rect 11488 15056 11552 15060
rect 18112 15116 18176 15120
rect 18112 15060 18116 15116
rect 18116 15060 18172 15116
rect 18172 15060 18176 15116
rect 18112 15056 18176 15060
rect 18192 15116 18256 15120
rect 18192 15060 18196 15116
rect 18196 15060 18252 15116
rect 18252 15060 18256 15116
rect 18192 15056 18256 15060
rect 18272 15116 18336 15120
rect 18272 15060 18276 15116
rect 18276 15060 18332 15116
rect 18332 15060 18336 15116
rect 18272 15056 18336 15060
rect 18352 15116 18416 15120
rect 18352 15060 18356 15116
rect 18356 15060 18412 15116
rect 18412 15060 18416 15116
rect 18352 15056 18416 15060
rect 7816 14572 7880 14576
rect 7816 14516 7820 14572
rect 7820 14516 7876 14572
rect 7876 14516 7880 14572
rect 7816 14512 7880 14516
rect 7896 14572 7960 14576
rect 7896 14516 7900 14572
rect 7900 14516 7956 14572
rect 7956 14516 7960 14572
rect 7896 14512 7960 14516
rect 7976 14572 8040 14576
rect 7976 14516 7980 14572
rect 7980 14516 8036 14572
rect 8036 14516 8040 14572
rect 7976 14512 8040 14516
rect 8056 14572 8120 14576
rect 8056 14516 8060 14572
rect 8060 14516 8116 14572
rect 8116 14516 8120 14572
rect 8056 14512 8120 14516
rect 14680 14572 14744 14576
rect 14680 14516 14684 14572
rect 14684 14516 14740 14572
rect 14740 14516 14744 14572
rect 14680 14512 14744 14516
rect 14760 14572 14824 14576
rect 14760 14516 14764 14572
rect 14764 14516 14820 14572
rect 14820 14516 14824 14572
rect 14760 14512 14824 14516
rect 14840 14572 14904 14576
rect 14840 14516 14844 14572
rect 14844 14516 14900 14572
rect 14900 14516 14904 14572
rect 14840 14512 14904 14516
rect 14920 14572 14984 14576
rect 14920 14516 14924 14572
rect 14924 14516 14980 14572
rect 14980 14516 14984 14572
rect 14920 14512 14984 14516
rect 4384 14028 4448 14032
rect 4384 13972 4388 14028
rect 4388 13972 4444 14028
rect 4444 13972 4448 14028
rect 4384 13968 4448 13972
rect 4464 14028 4528 14032
rect 4464 13972 4468 14028
rect 4468 13972 4524 14028
rect 4524 13972 4528 14028
rect 4464 13968 4528 13972
rect 4544 14028 4608 14032
rect 4544 13972 4548 14028
rect 4548 13972 4604 14028
rect 4604 13972 4608 14028
rect 4544 13968 4608 13972
rect 4624 14028 4688 14032
rect 4624 13972 4628 14028
rect 4628 13972 4684 14028
rect 4684 13972 4688 14028
rect 4624 13968 4688 13972
rect 11248 14028 11312 14032
rect 11248 13972 11252 14028
rect 11252 13972 11308 14028
rect 11308 13972 11312 14028
rect 11248 13968 11312 13972
rect 11328 14028 11392 14032
rect 11328 13972 11332 14028
rect 11332 13972 11388 14028
rect 11388 13972 11392 14028
rect 11328 13968 11392 13972
rect 11408 14028 11472 14032
rect 11408 13972 11412 14028
rect 11412 13972 11468 14028
rect 11468 13972 11472 14028
rect 11408 13968 11472 13972
rect 11488 14028 11552 14032
rect 11488 13972 11492 14028
rect 11492 13972 11548 14028
rect 11548 13972 11552 14028
rect 11488 13968 11552 13972
rect 18112 14028 18176 14032
rect 18112 13972 18116 14028
rect 18116 13972 18172 14028
rect 18172 13972 18176 14028
rect 18112 13968 18176 13972
rect 18192 14028 18256 14032
rect 18192 13972 18196 14028
rect 18196 13972 18252 14028
rect 18252 13972 18256 14028
rect 18192 13968 18256 13972
rect 18272 14028 18336 14032
rect 18272 13972 18276 14028
rect 18276 13972 18332 14028
rect 18332 13972 18336 14028
rect 18272 13968 18336 13972
rect 18352 14028 18416 14032
rect 18352 13972 18356 14028
rect 18356 13972 18412 14028
rect 18412 13972 18416 14028
rect 18352 13968 18416 13972
rect 7816 13484 7880 13488
rect 7816 13428 7820 13484
rect 7820 13428 7876 13484
rect 7876 13428 7880 13484
rect 7816 13424 7880 13428
rect 7896 13484 7960 13488
rect 7896 13428 7900 13484
rect 7900 13428 7956 13484
rect 7956 13428 7960 13484
rect 7896 13424 7960 13428
rect 7976 13484 8040 13488
rect 7976 13428 7980 13484
rect 7980 13428 8036 13484
rect 8036 13428 8040 13484
rect 7976 13424 8040 13428
rect 8056 13484 8120 13488
rect 8056 13428 8060 13484
rect 8060 13428 8116 13484
rect 8116 13428 8120 13484
rect 8056 13424 8120 13428
rect 14680 13484 14744 13488
rect 14680 13428 14684 13484
rect 14684 13428 14740 13484
rect 14740 13428 14744 13484
rect 14680 13424 14744 13428
rect 14760 13484 14824 13488
rect 14760 13428 14764 13484
rect 14764 13428 14820 13484
rect 14820 13428 14824 13484
rect 14760 13424 14824 13428
rect 14840 13484 14904 13488
rect 14840 13428 14844 13484
rect 14844 13428 14900 13484
rect 14900 13428 14904 13484
rect 14840 13424 14904 13428
rect 14920 13484 14984 13488
rect 14920 13428 14924 13484
rect 14924 13428 14980 13484
rect 14980 13428 14984 13484
rect 14920 13424 14984 13428
rect 4384 12940 4448 12944
rect 4384 12884 4388 12940
rect 4388 12884 4444 12940
rect 4444 12884 4448 12940
rect 4384 12880 4448 12884
rect 4464 12940 4528 12944
rect 4464 12884 4468 12940
rect 4468 12884 4524 12940
rect 4524 12884 4528 12940
rect 4464 12880 4528 12884
rect 4544 12940 4608 12944
rect 4544 12884 4548 12940
rect 4548 12884 4604 12940
rect 4604 12884 4608 12940
rect 4544 12880 4608 12884
rect 4624 12940 4688 12944
rect 4624 12884 4628 12940
rect 4628 12884 4684 12940
rect 4684 12884 4688 12940
rect 4624 12880 4688 12884
rect 11248 12940 11312 12944
rect 11248 12884 11252 12940
rect 11252 12884 11308 12940
rect 11308 12884 11312 12940
rect 11248 12880 11312 12884
rect 11328 12940 11392 12944
rect 11328 12884 11332 12940
rect 11332 12884 11388 12940
rect 11388 12884 11392 12940
rect 11328 12880 11392 12884
rect 11408 12940 11472 12944
rect 11408 12884 11412 12940
rect 11412 12884 11468 12940
rect 11468 12884 11472 12940
rect 11408 12880 11472 12884
rect 11488 12940 11552 12944
rect 11488 12884 11492 12940
rect 11492 12884 11548 12940
rect 11548 12884 11552 12940
rect 11488 12880 11552 12884
rect 18112 12940 18176 12944
rect 18112 12884 18116 12940
rect 18116 12884 18172 12940
rect 18172 12884 18176 12940
rect 18112 12880 18176 12884
rect 18192 12940 18256 12944
rect 18192 12884 18196 12940
rect 18196 12884 18252 12940
rect 18252 12884 18256 12940
rect 18192 12880 18256 12884
rect 18272 12940 18336 12944
rect 18272 12884 18276 12940
rect 18276 12884 18332 12940
rect 18332 12884 18336 12940
rect 18272 12880 18336 12884
rect 18352 12940 18416 12944
rect 18352 12884 18356 12940
rect 18356 12884 18412 12940
rect 18412 12884 18416 12940
rect 18352 12880 18416 12884
rect 7816 12396 7880 12400
rect 7816 12340 7820 12396
rect 7820 12340 7876 12396
rect 7876 12340 7880 12396
rect 7816 12336 7880 12340
rect 7896 12396 7960 12400
rect 7896 12340 7900 12396
rect 7900 12340 7956 12396
rect 7956 12340 7960 12396
rect 7896 12336 7960 12340
rect 7976 12396 8040 12400
rect 7976 12340 7980 12396
rect 7980 12340 8036 12396
rect 8036 12340 8040 12396
rect 7976 12336 8040 12340
rect 8056 12396 8120 12400
rect 8056 12340 8060 12396
rect 8060 12340 8116 12396
rect 8116 12340 8120 12396
rect 8056 12336 8120 12340
rect 14680 12396 14744 12400
rect 14680 12340 14684 12396
rect 14684 12340 14740 12396
rect 14740 12340 14744 12396
rect 14680 12336 14744 12340
rect 14760 12396 14824 12400
rect 14760 12340 14764 12396
rect 14764 12340 14820 12396
rect 14820 12340 14824 12396
rect 14760 12336 14824 12340
rect 14840 12396 14904 12400
rect 14840 12340 14844 12396
rect 14844 12340 14900 12396
rect 14900 12340 14904 12396
rect 14840 12336 14904 12340
rect 14920 12396 14984 12400
rect 14920 12340 14924 12396
rect 14924 12340 14980 12396
rect 14980 12340 14984 12396
rect 14920 12336 14984 12340
rect 4384 11852 4448 11856
rect 4384 11796 4388 11852
rect 4388 11796 4444 11852
rect 4444 11796 4448 11852
rect 4384 11792 4448 11796
rect 4464 11852 4528 11856
rect 4464 11796 4468 11852
rect 4468 11796 4524 11852
rect 4524 11796 4528 11852
rect 4464 11792 4528 11796
rect 4544 11852 4608 11856
rect 4544 11796 4548 11852
rect 4548 11796 4604 11852
rect 4604 11796 4608 11852
rect 4544 11792 4608 11796
rect 4624 11852 4688 11856
rect 4624 11796 4628 11852
rect 4628 11796 4684 11852
rect 4684 11796 4688 11852
rect 4624 11792 4688 11796
rect 11248 11852 11312 11856
rect 11248 11796 11252 11852
rect 11252 11796 11308 11852
rect 11308 11796 11312 11852
rect 11248 11792 11312 11796
rect 11328 11852 11392 11856
rect 11328 11796 11332 11852
rect 11332 11796 11388 11852
rect 11388 11796 11392 11852
rect 11328 11792 11392 11796
rect 11408 11852 11472 11856
rect 11408 11796 11412 11852
rect 11412 11796 11468 11852
rect 11468 11796 11472 11852
rect 11408 11792 11472 11796
rect 11488 11852 11552 11856
rect 11488 11796 11492 11852
rect 11492 11796 11548 11852
rect 11548 11796 11552 11852
rect 11488 11792 11552 11796
rect 18112 11852 18176 11856
rect 18112 11796 18116 11852
rect 18116 11796 18172 11852
rect 18172 11796 18176 11852
rect 18112 11792 18176 11796
rect 18192 11852 18256 11856
rect 18192 11796 18196 11852
rect 18196 11796 18252 11852
rect 18252 11796 18256 11852
rect 18192 11792 18256 11796
rect 18272 11852 18336 11856
rect 18272 11796 18276 11852
rect 18276 11796 18332 11852
rect 18332 11796 18336 11852
rect 18272 11792 18336 11796
rect 18352 11852 18416 11856
rect 18352 11796 18356 11852
rect 18356 11796 18412 11852
rect 18412 11796 18416 11852
rect 18352 11792 18416 11796
rect 7816 11308 7880 11312
rect 7816 11252 7820 11308
rect 7820 11252 7876 11308
rect 7876 11252 7880 11308
rect 7816 11248 7880 11252
rect 7896 11308 7960 11312
rect 7896 11252 7900 11308
rect 7900 11252 7956 11308
rect 7956 11252 7960 11308
rect 7896 11248 7960 11252
rect 7976 11308 8040 11312
rect 7976 11252 7980 11308
rect 7980 11252 8036 11308
rect 8036 11252 8040 11308
rect 7976 11248 8040 11252
rect 8056 11308 8120 11312
rect 8056 11252 8060 11308
rect 8060 11252 8116 11308
rect 8116 11252 8120 11308
rect 8056 11248 8120 11252
rect 14680 11308 14744 11312
rect 14680 11252 14684 11308
rect 14684 11252 14740 11308
rect 14740 11252 14744 11308
rect 14680 11248 14744 11252
rect 14760 11308 14824 11312
rect 14760 11252 14764 11308
rect 14764 11252 14820 11308
rect 14820 11252 14824 11308
rect 14760 11248 14824 11252
rect 14840 11308 14904 11312
rect 14840 11252 14844 11308
rect 14844 11252 14900 11308
rect 14900 11252 14904 11308
rect 14840 11248 14904 11252
rect 14920 11308 14984 11312
rect 14920 11252 14924 11308
rect 14924 11252 14980 11308
rect 14980 11252 14984 11308
rect 14920 11248 14984 11252
rect 4384 10764 4448 10768
rect 4384 10708 4388 10764
rect 4388 10708 4444 10764
rect 4444 10708 4448 10764
rect 4384 10704 4448 10708
rect 4464 10764 4528 10768
rect 4464 10708 4468 10764
rect 4468 10708 4524 10764
rect 4524 10708 4528 10764
rect 4464 10704 4528 10708
rect 4544 10764 4608 10768
rect 4544 10708 4548 10764
rect 4548 10708 4604 10764
rect 4604 10708 4608 10764
rect 4544 10704 4608 10708
rect 4624 10764 4688 10768
rect 4624 10708 4628 10764
rect 4628 10708 4684 10764
rect 4684 10708 4688 10764
rect 4624 10704 4688 10708
rect 11248 10764 11312 10768
rect 11248 10708 11252 10764
rect 11252 10708 11308 10764
rect 11308 10708 11312 10764
rect 11248 10704 11312 10708
rect 11328 10764 11392 10768
rect 11328 10708 11332 10764
rect 11332 10708 11388 10764
rect 11388 10708 11392 10764
rect 11328 10704 11392 10708
rect 11408 10764 11472 10768
rect 11408 10708 11412 10764
rect 11412 10708 11468 10764
rect 11468 10708 11472 10764
rect 11408 10704 11472 10708
rect 11488 10764 11552 10768
rect 11488 10708 11492 10764
rect 11492 10708 11548 10764
rect 11548 10708 11552 10764
rect 11488 10704 11552 10708
rect 18112 10764 18176 10768
rect 18112 10708 18116 10764
rect 18116 10708 18172 10764
rect 18172 10708 18176 10764
rect 18112 10704 18176 10708
rect 18192 10764 18256 10768
rect 18192 10708 18196 10764
rect 18196 10708 18252 10764
rect 18252 10708 18256 10764
rect 18192 10704 18256 10708
rect 18272 10764 18336 10768
rect 18272 10708 18276 10764
rect 18276 10708 18332 10764
rect 18332 10708 18336 10764
rect 18272 10704 18336 10708
rect 18352 10764 18416 10768
rect 18352 10708 18356 10764
rect 18356 10708 18412 10764
rect 18412 10708 18416 10764
rect 18352 10704 18416 10708
rect 7816 10220 7880 10224
rect 7816 10164 7820 10220
rect 7820 10164 7876 10220
rect 7876 10164 7880 10220
rect 7816 10160 7880 10164
rect 7896 10220 7960 10224
rect 7896 10164 7900 10220
rect 7900 10164 7956 10220
rect 7956 10164 7960 10220
rect 7896 10160 7960 10164
rect 7976 10220 8040 10224
rect 7976 10164 7980 10220
rect 7980 10164 8036 10220
rect 8036 10164 8040 10220
rect 7976 10160 8040 10164
rect 8056 10220 8120 10224
rect 8056 10164 8060 10220
rect 8060 10164 8116 10220
rect 8116 10164 8120 10220
rect 8056 10160 8120 10164
rect 14680 10220 14744 10224
rect 14680 10164 14684 10220
rect 14684 10164 14740 10220
rect 14740 10164 14744 10220
rect 14680 10160 14744 10164
rect 14760 10220 14824 10224
rect 14760 10164 14764 10220
rect 14764 10164 14820 10220
rect 14820 10164 14824 10220
rect 14760 10160 14824 10164
rect 14840 10220 14904 10224
rect 14840 10164 14844 10220
rect 14844 10164 14900 10220
rect 14900 10164 14904 10220
rect 14840 10160 14904 10164
rect 14920 10220 14984 10224
rect 14920 10164 14924 10220
rect 14924 10164 14980 10220
rect 14980 10164 14984 10220
rect 14920 10160 14984 10164
rect 4384 9676 4448 9680
rect 4384 9620 4388 9676
rect 4388 9620 4444 9676
rect 4444 9620 4448 9676
rect 4384 9616 4448 9620
rect 4464 9676 4528 9680
rect 4464 9620 4468 9676
rect 4468 9620 4524 9676
rect 4524 9620 4528 9676
rect 4464 9616 4528 9620
rect 4544 9676 4608 9680
rect 4544 9620 4548 9676
rect 4548 9620 4604 9676
rect 4604 9620 4608 9676
rect 4544 9616 4608 9620
rect 4624 9676 4688 9680
rect 4624 9620 4628 9676
rect 4628 9620 4684 9676
rect 4684 9620 4688 9676
rect 4624 9616 4688 9620
rect 11248 9676 11312 9680
rect 11248 9620 11252 9676
rect 11252 9620 11308 9676
rect 11308 9620 11312 9676
rect 11248 9616 11312 9620
rect 11328 9676 11392 9680
rect 11328 9620 11332 9676
rect 11332 9620 11388 9676
rect 11388 9620 11392 9676
rect 11328 9616 11392 9620
rect 11408 9676 11472 9680
rect 11408 9620 11412 9676
rect 11412 9620 11468 9676
rect 11468 9620 11472 9676
rect 11408 9616 11472 9620
rect 11488 9676 11552 9680
rect 11488 9620 11492 9676
rect 11492 9620 11548 9676
rect 11548 9620 11552 9676
rect 11488 9616 11552 9620
rect 18112 9676 18176 9680
rect 18112 9620 18116 9676
rect 18116 9620 18172 9676
rect 18172 9620 18176 9676
rect 18112 9616 18176 9620
rect 18192 9676 18256 9680
rect 18192 9620 18196 9676
rect 18196 9620 18252 9676
rect 18252 9620 18256 9676
rect 18192 9616 18256 9620
rect 18272 9676 18336 9680
rect 18272 9620 18276 9676
rect 18276 9620 18332 9676
rect 18332 9620 18336 9676
rect 18272 9616 18336 9620
rect 18352 9676 18416 9680
rect 18352 9620 18356 9676
rect 18356 9620 18412 9676
rect 18412 9620 18416 9676
rect 18352 9616 18416 9620
rect 7816 9132 7880 9136
rect 7816 9076 7820 9132
rect 7820 9076 7876 9132
rect 7876 9076 7880 9132
rect 7816 9072 7880 9076
rect 7896 9132 7960 9136
rect 7896 9076 7900 9132
rect 7900 9076 7956 9132
rect 7956 9076 7960 9132
rect 7896 9072 7960 9076
rect 7976 9132 8040 9136
rect 7976 9076 7980 9132
rect 7980 9076 8036 9132
rect 8036 9076 8040 9132
rect 7976 9072 8040 9076
rect 8056 9132 8120 9136
rect 8056 9076 8060 9132
rect 8060 9076 8116 9132
rect 8116 9076 8120 9132
rect 8056 9072 8120 9076
rect 14680 9132 14744 9136
rect 14680 9076 14684 9132
rect 14684 9076 14740 9132
rect 14740 9076 14744 9132
rect 14680 9072 14744 9076
rect 14760 9132 14824 9136
rect 14760 9076 14764 9132
rect 14764 9076 14820 9132
rect 14820 9076 14824 9132
rect 14760 9072 14824 9076
rect 14840 9132 14904 9136
rect 14840 9076 14844 9132
rect 14844 9076 14900 9132
rect 14900 9076 14904 9132
rect 14840 9072 14904 9076
rect 14920 9132 14984 9136
rect 14920 9076 14924 9132
rect 14924 9076 14980 9132
rect 14980 9076 14984 9132
rect 14920 9072 14984 9076
rect 4384 8588 4448 8592
rect 4384 8532 4388 8588
rect 4388 8532 4444 8588
rect 4444 8532 4448 8588
rect 4384 8528 4448 8532
rect 4464 8588 4528 8592
rect 4464 8532 4468 8588
rect 4468 8532 4524 8588
rect 4524 8532 4528 8588
rect 4464 8528 4528 8532
rect 4544 8588 4608 8592
rect 4544 8532 4548 8588
rect 4548 8532 4604 8588
rect 4604 8532 4608 8588
rect 4544 8528 4608 8532
rect 4624 8588 4688 8592
rect 4624 8532 4628 8588
rect 4628 8532 4684 8588
rect 4684 8532 4688 8588
rect 4624 8528 4688 8532
rect 11248 8588 11312 8592
rect 11248 8532 11252 8588
rect 11252 8532 11308 8588
rect 11308 8532 11312 8588
rect 11248 8528 11312 8532
rect 11328 8588 11392 8592
rect 11328 8532 11332 8588
rect 11332 8532 11388 8588
rect 11388 8532 11392 8588
rect 11328 8528 11392 8532
rect 11408 8588 11472 8592
rect 11408 8532 11412 8588
rect 11412 8532 11468 8588
rect 11468 8532 11472 8588
rect 11408 8528 11472 8532
rect 11488 8588 11552 8592
rect 11488 8532 11492 8588
rect 11492 8532 11548 8588
rect 11548 8532 11552 8588
rect 11488 8528 11552 8532
rect 18112 8588 18176 8592
rect 18112 8532 18116 8588
rect 18116 8532 18172 8588
rect 18172 8532 18176 8588
rect 18112 8528 18176 8532
rect 18192 8588 18256 8592
rect 18192 8532 18196 8588
rect 18196 8532 18252 8588
rect 18252 8532 18256 8588
rect 18192 8528 18256 8532
rect 18272 8588 18336 8592
rect 18272 8532 18276 8588
rect 18276 8532 18332 8588
rect 18332 8532 18336 8588
rect 18272 8528 18336 8532
rect 18352 8588 18416 8592
rect 18352 8532 18356 8588
rect 18356 8532 18412 8588
rect 18412 8532 18416 8588
rect 18352 8528 18416 8532
rect 7816 8044 7880 8048
rect 7816 7988 7820 8044
rect 7820 7988 7876 8044
rect 7876 7988 7880 8044
rect 7816 7984 7880 7988
rect 7896 8044 7960 8048
rect 7896 7988 7900 8044
rect 7900 7988 7956 8044
rect 7956 7988 7960 8044
rect 7896 7984 7960 7988
rect 7976 8044 8040 8048
rect 7976 7988 7980 8044
rect 7980 7988 8036 8044
rect 8036 7988 8040 8044
rect 7976 7984 8040 7988
rect 8056 8044 8120 8048
rect 8056 7988 8060 8044
rect 8060 7988 8116 8044
rect 8116 7988 8120 8044
rect 8056 7984 8120 7988
rect 14680 8044 14744 8048
rect 14680 7988 14684 8044
rect 14684 7988 14740 8044
rect 14740 7988 14744 8044
rect 14680 7984 14744 7988
rect 14760 8044 14824 8048
rect 14760 7988 14764 8044
rect 14764 7988 14820 8044
rect 14820 7988 14824 8044
rect 14760 7984 14824 7988
rect 14840 8044 14904 8048
rect 14840 7988 14844 8044
rect 14844 7988 14900 8044
rect 14900 7988 14904 8044
rect 14840 7984 14904 7988
rect 14920 8044 14984 8048
rect 14920 7988 14924 8044
rect 14924 7988 14980 8044
rect 14980 7988 14984 8044
rect 14920 7984 14984 7988
rect 4384 7500 4448 7504
rect 4384 7444 4388 7500
rect 4388 7444 4444 7500
rect 4444 7444 4448 7500
rect 4384 7440 4448 7444
rect 4464 7500 4528 7504
rect 4464 7444 4468 7500
rect 4468 7444 4524 7500
rect 4524 7444 4528 7500
rect 4464 7440 4528 7444
rect 4544 7500 4608 7504
rect 4544 7444 4548 7500
rect 4548 7444 4604 7500
rect 4604 7444 4608 7500
rect 4544 7440 4608 7444
rect 4624 7500 4688 7504
rect 4624 7444 4628 7500
rect 4628 7444 4684 7500
rect 4684 7444 4688 7500
rect 4624 7440 4688 7444
rect 11248 7500 11312 7504
rect 11248 7444 11252 7500
rect 11252 7444 11308 7500
rect 11308 7444 11312 7500
rect 11248 7440 11312 7444
rect 11328 7500 11392 7504
rect 11328 7444 11332 7500
rect 11332 7444 11388 7500
rect 11388 7444 11392 7500
rect 11328 7440 11392 7444
rect 11408 7500 11472 7504
rect 11408 7444 11412 7500
rect 11412 7444 11468 7500
rect 11468 7444 11472 7500
rect 11408 7440 11472 7444
rect 11488 7500 11552 7504
rect 11488 7444 11492 7500
rect 11492 7444 11548 7500
rect 11548 7444 11552 7500
rect 11488 7440 11552 7444
rect 18112 7500 18176 7504
rect 18112 7444 18116 7500
rect 18116 7444 18172 7500
rect 18172 7444 18176 7500
rect 18112 7440 18176 7444
rect 18192 7500 18256 7504
rect 18192 7444 18196 7500
rect 18196 7444 18252 7500
rect 18252 7444 18256 7500
rect 18192 7440 18256 7444
rect 18272 7500 18336 7504
rect 18272 7444 18276 7500
rect 18276 7444 18332 7500
rect 18332 7444 18336 7500
rect 18272 7440 18336 7444
rect 18352 7500 18416 7504
rect 18352 7444 18356 7500
rect 18356 7444 18412 7500
rect 18412 7444 18416 7500
rect 18352 7440 18416 7444
rect 7816 6956 7880 6960
rect 7816 6900 7820 6956
rect 7820 6900 7876 6956
rect 7876 6900 7880 6956
rect 7816 6896 7880 6900
rect 7896 6956 7960 6960
rect 7896 6900 7900 6956
rect 7900 6900 7956 6956
rect 7956 6900 7960 6956
rect 7896 6896 7960 6900
rect 7976 6956 8040 6960
rect 7976 6900 7980 6956
rect 7980 6900 8036 6956
rect 8036 6900 8040 6956
rect 7976 6896 8040 6900
rect 8056 6956 8120 6960
rect 8056 6900 8060 6956
rect 8060 6900 8116 6956
rect 8116 6900 8120 6956
rect 8056 6896 8120 6900
rect 14680 6956 14744 6960
rect 14680 6900 14684 6956
rect 14684 6900 14740 6956
rect 14740 6900 14744 6956
rect 14680 6896 14744 6900
rect 14760 6956 14824 6960
rect 14760 6900 14764 6956
rect 14764 6900 14820 6956
rect 14820 6900 14824 6956
rect 14760 6896 14824 6900
rect 14840 6956 14904 6960
rect 14840 6900 14844 6956
rect 14844 6900 14900 6956
rect 14900 6900 14904 6956
rect 14840 6896 14904 6900
rect 14920 6956 14984 6960
rect 14920 6900 14924 6956
rect 14924 6900 14980 6956
rect 14980 6900 14984 6956
rect 14920 6896 14984 6900
rect 4384 6412 4448 6416
rect 4384 6356 4388 6412
rect 4388 6356 4444 6412
rect 4444 6356 4448 6412
rect 4384 6352 4448 6356
rect 4464 6412 4528 6416
rect 4464 6356 4468 6412
rect 4468 6356 4524 6412
rect 4524 6356 4528 6412
rect 4464 6352 4528 6356
rect 4544 6412 4608 6416
rect 4544 6356 4548 6412
rect 4548 6356 4604 6412
rect 4604 6356 4608 6412
rect 4544 6352 4608 6356
rect 4624 6412 4688 6416
rect 4624 6356 4628 6412
rect 4628 6356 4684 6412
rect 4684 6356 4688 6412
rect 4624 6352 4688 6356
rect 11248 6412 11312 6416
rect 11248 6356 11252 6412
rect 11252 6356 11308 6412
rect 11308 6356 11312 6412
rect 11248 6352 11312 6356
rect 11328 6412 11392 6416
rect 11328 6356 11332 6412
rect 11332 6356 11388 6412
rect 11388 6356 11392 6412
rect 11328 6352 11392 6356
rect 11408 6412 11472 6416
rect 11408 6356 11412 6412
rect 11412 6356 11468 6412
rect 11468 6356 11472 6412
rect 11408 6352 11472 6356
rect 11488 6412 11552 6416
rect 11488 6356 11492 6412
rect 11492 6356 11548 6412
rect 11548 6356 11552 6412
rect 11488 6352 11552 6356
rect 18112 6412 18176 6416
rect 18112 6356 18116 6412
rect 18116 6356 18172 6412
rect 18172 6356 18176 6412
rect 18112 6352 18176 6356
rect 18192 6412 18256 6416
rect 18192 6356 18196 6412
rect 18196 6356 18252 6412
rect 18252 6356 18256 6412
rect 18192 6352 18256 6356
rect 18272 6412 18336 6416
rect 18272 6356 18276 6412
rect 18276 6356 18332 6412
rect 18332 6356 18336 6412
rect 18272 6352 18336 6356
rect 18352 6412 18416 6416
rect 18352 6356 18356 6412
rect 18356 6356 18412 6412
rect 18412 6356 18416 6412
rect 18352 6352 18416 6356
rect 7816 5868 7880 5872
rect 7816 5812 7820 5868
rect 7820 5812 7876 5868
rect 7876 5812 7880 5868
rect 7816 5808 7880 5812
rect 7896 5868 7960 5872
rect 7896 5812 7900 5868
rect 7900 5812 7956 5868
rect 7956 5812 7960 5868
rect 7896 5808 7960 5812
rect 7976 5868 8040 5872
rect 7976 5812 7980 5868
rect 7980 5812 8036 5868
rect 8036 5812 8040 5868
rect 7976 5808 8040 5812
rect 8056 5868 8120 5872
rect 8056 5812 8060 5868
rect 8060 5812 8116 5868
rect 8116 5812 8120 5868
rect 8056 5808 8120 5812
rect 14680 5868 14744 5872
rect 14680 5812 14684 5868
rect 14684 5812 14740 5868
rect 14740 5812 14744 5868
rect 14680 5808 14744 5812
rect 14760 5868 14824 5872
rect 14760 5812 14764 5868
rect 14764 5812 14820 5868
rect 14820 5812 14824 5868
rect 14760 5808 14824 5812
rect 14840 5868 14904 5872
rect 14840 5812 14844 5868
rect 14844 5812 14900 5868
rect 14900 5812 14904 5868
rect 14840 5808 14904 5812
rect 14920 5868 14984 5872
rect 14920 5812 14924 5868
rect 14924 5812 14980 5868
rect 14980 5812 14984 5868
rect 14920 5808 14984 5812
rect 4384 5324 4448 5328
rect 4384 5268 4388 5324
rect 4388 5268 4444 5324
rect 4444 5268 4448 5324
rect 4384 5264 4448 5268
rect 4464 5324 4528 5328
rect 4464 5268 4468 5324
rect 4468 5268 4524 5324
rect 4524 5268 4528 5324
rect 4464 5264 4528 5268
rect 4544 5324 4608 5328
rect 4544 5268 4548 5324
rect 4548 5268 4604 5324
rect 4604 5268 4608 5324
rect 4544 5264 4608 5268
rect 4624 5324 4688 5328
rect 4624 5268 4628 5324
rect 4628 5268 4684 5324
rect 4684 5268 4688 5324
rect 4624 5264 4688 5268
rect 11248 5324 11312 5328
rect 11248 5268 11252 5324
rect 11252 5268 11308 5324
rect 11308 5268 11312 5324
rect 11248 5264 11312 5268
rect 11328 5324 11392 5328
rect 11328 5268 11332 5324
rect 11332 5268 11388 5324
rect 11388 5268 11392 5324
rect 11328 5264 11392 5268
rect 11408 5324 11472 5328
rect 11408 5268 11412 5324
rect 11412 5268 11468 5324
rect 11468 5268 11472 5324
rect 11408 5264 11472 5268
rect 11488 5324 11552 5328
rect 11488 5268 11492 5324
rect 11492 5268 11548 5324
rect 11548 5268 11552 5324
rect 11488 5264 11552 5268
rect 18112 5324 18176 5328
rect 18112 5268 18116 5324
rect 18116 5268 18172 5324
rect 18172 5268 18176 5324
rect 18112 5264 18176 5268
rect 18192 5324 18256 5328
rect 18192 5268 18196 5324
rect 18196 5268 18252 5324
rect 18252 5268 18256 5324
rect 18192 5264 18256 5268
rect 18272 5324 18336 5328
rect 18272 5268 18276 5324
rect 18276 5268 18332 5324
rect 18332 5268 18336 5324
rect 18272 5264 18336 5268
rect 18352 5324 18416 5328
rect 18352 5268 18356 5324
rect 18356 5268 18412 5324
rect 18412 5268 18416 5324
rect 18352 5264 18416 5268
rect 7816 4780 7880 4784
rect 7816 4724 7820 4780
rect 7820 4724 7876 4780
rect 7876 4724 7880 4780
rect 7816 4720 7880 4724
rect 7896 4780 7960 4784
rect 7896 4724 7900 4780
rect 7900 4724 7956 4780
rect 7956 4724 7960 4780
rect 7896 4720 7960 4724
rect 7976 4780 8040 4784
rect 7976 4724 7980 4780
rect 7980 4724 8036 4780
rect 8036 4724 8040 4780
rect 7976 4720 8040 4724
rect 8056 4780 8120 4784
rect 8056 4724 8060 4780
rect 8060 4724 8116 4780
rect 8116 4724 8120 4780
rect 8056 4720 8120 4724
rect 14680 4780 14744 4784
rect 14680 4724 14684 4780
rect 14684 4724 14740 4780
rect 14740 4724 14744 4780
rect 14680 4720 14744 4724
rect 14760 4780 14824 4784
rect 14760 4724 14764 4780
rect 14764 4724 14820 4780
rect 14820 4724 14824 4780
rect 14760 4720 14824 4724
rect 14840 4780 14904 4784
rect 14840 4724 14844 4780
rect 14844 4724 14900 4780
rect 14900 4724 14904 4780
rect 14840 4720 14904 4724
rect 14920 4780 14984 4784
rect 14920 4724 14924 4780
rect 14924 4724 14980 4780
rect 14980 4724 14984 4780
rect 14920 4720 14984 4724
rect 4384 4236 4448 4240
rect 4384 4180 4388 4236
rect 4388 4180 4444 4236
rect 4444 4180 4448 4236
rect 4384 4176 4448 4180
rect 4464 4236 4528 4240
rect 4464 4180 4468 4236
rect 4468 4180 4524 4236
rect 4524 4180 4528 4236
rect 4464 4176 4528 4180
rect 4544 4236 4608 4240
rect 4544 4180 4548 4236
rect 4548 4180 4604 4236
rect 4604 4180 4608 4236
rect 4544 4176 4608 4180
rect 4624 4236 4688 4240
rect 4624 4180 4628 4236
rect 4628 4180 4684 4236
rect 4684 4180 4688 4236
rect 4624 4176 4688 4180
rect 11248 4236 11312 4240
rect 11248 4180 11252 4236
rect 11252 4180 11308 4236
rect 11308 4180 11312 4236
rect 11248 4176 11312 4180
rect 11328 4236 11392 4240
rect 11328 4180 11332 4236
rect 11332 4180 11388 4236
rect 11388 4180 11392 4236
rect 11328 4176 11392 4180
rect 11408 4236 11472 4240
rect 11408 4180 11412 4236
rect 11412 4180 11468 4236
rect 11468 4180 11472 4236
rect 11408 4176 11472 4180
rect 11488 4236 11552 4240
rect 11488 4180 11492 4236
rect 11492 4180 11548 4236
rect 11548 4180 11552 4236
rect 11488 4176 11552 4180
rect 18112 4236 18176 4240
rect 18112 4180 18116 4236
rect 18116 4180 18172 4236
rect 18172 4180 18176 4236
rect 18112 4176 18176 4180
rect 18192 4236 18256 4240
rect 18192 4180 18196 4236
rect 18196 4180 18252 4236
rect 18252 4180 18256 4236
rect 18192 4176 18256 4180
rect 18272 4236 18336 4240
rect 18272 4180 18276 4236
rect 18276 4180 18332 4236
rect 18332 4180 18336 4236
rect 18272 4176 18336 4180
rect 18352 4236 18416 4240
rect 18352 4180 18356 4236
rect 18356 4180 18412 4236
rect 18412 4180 18416 4236
rect 18352 4176 18416 4180
rect 7816 3692 7880 3696
rect 7816 3636 7820 3692
rect 7820 3636 7876 3692
rect 7876 3636 7880 3692
rect 7816 3632 7880 3636
rect 7896 3692 7960 3696
rect 7896 3636 7900 3692
rect 7900 3636 7956 3692
rect 7956 3636 7960 3692
rect 7896 3632 7960 3636
rect 7976 3692 8040 3696
rect 7976 3636 7980 3692
rect 7980 3636 8036 3692
rect 8036 3636 8040 3692
rect 7976 3632 8040 3636
rect 8056 3692 8120 3696
rect 8056 3636 8060 3692
rect 8060 3636 8116 3692
rect 8116 3636 8120 3692
rect 8056 3632 8120 3636
rect 14680 3692 14744 3696
rect 14680 3636 14684 3692
rect 14684 3636 14740 3692
rect 14740 3636 14744 3692
rect 14680 3632 14744 3636
rect 14760 3692 14824 3696
rect 14760 3636 14764 3692
rect 14764 3636 14820 3692
rect 14820 3636 14824 3692
rect 14760 3632 14824 3636
rect 14840 3692 14904 3696
rect 14840 3636 14844 3692
rect 14844 3636 14900 3692
rect 14900 3636 14904 3692
rect 14840 3632 14904 3636
rect 14920 3692 14984 3696
rect 14920 3636 14924 3692
rect 14924 3636 14980 3692
rect 14980 3636 14984 3692
rect 14920 3632 14984 3636
rect 4384 3148 4448 3152
rect 4384 3092 4388 3148
rect 4388 3092 4444 3148
rect 4444 3092 4448 3148
rect 4384 3088 4448 3092
rect 4464 3148 4528 3152
rect 4464 3092 4468 3148
rect 4468 3092 4524 3148
rect 4524 3092 4528 3148
rect 4464 3088 4528 3092
rect 4544 3148 4608 3152
rect 4544 3092 4548 3148
rect 4548 3092 4604 3148
rect 4604 3092 4608 3148
rect 4544 3088 4608 3092
rect 4624 3148 4688 3152
rect 4624 3092 4628 3148
rect 4628 3092 4684 3148
rect 4684 3092 4688 3148
rect 4624 3088 4688 3092
rect 11248 3148 11312 3152
rect 11248 3092 11252 3148
rect 11252 3092 11308 3148
rect 11308 3092 11312 3148
rect 11248 3088 11312 3092
rect 11328 3148 11392 3152
rect 11328 3092 11332 3148
rect 11332 3092 11388 3148
rect 11388 3092 11392 3148
rect 11328 3088 11392 3092
rect 11408 3148 11472 3152
rect 11408 3092 11412 3148
rect 11412 3092 11468 3148
rect 11468 3092 11472 3148
rect 11408 3088 11472 3092
rect 11488 3148 11552 3152
rect 11488 3092 11492 3148
rect 11492 3092 11548 3148
rect 11548 3092 11552 3148
rect 11488 3088 11552 3092
rect 18112 3148 18176 3152
rect 18112 3092 18116 3148
rect 18116 3092 18172 3148
rect 18172 3092 18176 3148
rect 18112 3088 18176 3092
rect 18192 3148 18256 3152
rect 18192 3092 18196 3148
rect 18196 3092 18252 3148
rect 18252 3092 18256 3148
rect 18192 3088 18256 3092
rect 18272 3148 18336 3152
rect 18272 3092 18276 3148
rect 18276 3092 18332 3148
rect 18332 3092 18336 3148
rect 18272 3088 18336 3092
rect 18352 3148 18416 3152
rect 18352 3092 18356 3148
rect 18356 3092 18412 3148
rect 18412 3092 18416 3148
rect 18352 3088 18416 3092
rect 7816 2604 7880 2608
rect 7816 2548 7820 2604
rect 7820 2548 7876 2604
rect 7876 2548 7880 2604
rect 7816 2544 7880 2548
rect 7896 2604 7960 2608
rect 7896 2548 7900 2604
rect 7900 2548 7956 2604
rect 7956 2548 7960 2604
rect 7896 2544 7960 2548
rect 7976 2604 8040 2608
rect 7976 2548 7980 2604
rect 7980 2548 8036 2604
rect 8036 2548 8040 2604
rect 7976 2544 8040 2548
rect 8056 2604 8120 2608
rect 8056 2548 8060 2604
rect 8060 2548 8116 2604
rect 8116 2548 8120 2604
rect 8056 2544 8120 2548
rect 14680 2604 14744 2608
rect 14680 2548 14684 2604
rect 14684 2548 14740 2604
rect 14740 2548 14744 2604
rect 14680 2544 14744 2548
rect 14760 2604 14824 2608
rect 14760 2548 14764 2604
rect 14764 2548 14820 2604
rect 14820 2548 14824 2604
rect 14760 2544 14824 2548
rect 14840 2604 14904 2608
rect 14840 2548 14844 2604
rect 14844 2548 14900 2604
rect 14900 2548 14904 2604
rect 14840 2544 14904 2548
rect 14920 2604 14984 2608
rect 14920 2548 14924 2604
rect 14924 2548 14980 2604
rect 14980 2548 14984 2604
rect 14920 2544 14984 2548
rect 4384 2060 4448 2064
rect 4384 2004 4388 2060
rect 4388 2004 4444 2060
rect 4444 2004 4448 2060
rect 4384 2000 4448 2004
rect 4464 2060 4528 2064
rect 4464 2004 4468 2060
rect 4468 2004 4524 2060
rect 4524 2004 4528 2060
rect 4464 2000 4528 2004
rect 4544 2060 4608 2064
rect 4544 2004 4548 2060
rect 4548 2004 4604 2060
rect 4604 2004 4608 2060
rect 4544 2000 4608 2004
rect 4624 2060 4688 2064
rect 4624 2004 4628 2060
rect 4628 2004 4684 2060
rect 4684 2004 4688 2060
rect 4624 2000 4688 2004
rect 11248 2060 11312 2064
rect 11248 2004 11252 2060
rect 11252 2004 11308 2060
rect 11308 2004 11312 2060
rect 11248 2000 11312 2004
rect 11328 2060 11392 2064
rect 11328 2004 11332 2060
rect 11332 2004 11388 2060
rect 11388 2004 11392 2060
rect 11328 2000 11392 2004
rect 11408 2060 11472 2064
rect 11408 2004 11412 2060
rect 11412 2004 11468 2060
rect 11468 2004 11472 2060
rect 11408 2000 11472 2004
rect 11488 2060 11552 2064
rect 11488 2004 11492 2060
rect 11492 2004 11548 2060
rect 11548 2004 11552 2060
rect 11488 2000 11552 2004
rect 18112 2060 18176 2064
rect 18112 2004 18116 2060
rect 18116 2004 18172 2060
rect 18172 2004 18176 2060
rect 18112 2000 18176 2004
rect 18192 2060 18256 2064
rect 18192 2004 18196 2060
rect 18196 2004 18252 2060
rect 18252 2004 18256 2060
rect 18192 2000 18256 2004
rect 18272 2060 18336 2064
rect 18272 2004 18276 2060
rect 18276 2004 18332 2060
rect 18332 2004 18336 2060
rect 18272 2000 18336 2004
rect 18352 2060 18416 2064
rect 18352 2004 18356 2060
rect 18356 2004 18412 2060
rect 18412 2004 18416 2060
rect 18352 2000 18416 2004
<< metal4 >>
rect 4376 19472 4696 20032
rect 4376 19408 4384 19472
rect 4448 19408 4464 19472
rect 4528 19408 4544 19472
rect 4608 19408 4624 19472
rect 4688 19408 4696 19472
rect 4376 18384 4696 19408
rect 4376 18320 4384 18384
rect 4448 18320 4464 18384
rect 4528 18320 4544 18384
rect 4608 18320 4624 18384
rect 4688 18320 4696 18384
rect 4376 17296 4696 18320
rect 4376 17232 4384 17296
rect 4448 17232 4464 17296
rect 4528 17232 4544 17296
rect 4608 17232 4624 17296
rect 4688 17232 4696 17296
rect 4376 16208 4696 17232
rect 4376 16144 4384 16208
rect 4448 16144 4464 16208
rect 4528 16144 4544 16208
rect 4608 16144 4624 16208
rect 4688 16144 4696 16208
rect 4376 15120 4696 16144
rect 4376 15056 4384 15120
rect 4448 15056 4464 15120
rect 4528 15056 4544 15120
rect 4608 15056 4624 15120
rect 4688 15056 4696 15120
rect 4376 14032 4696 15056
rect 4376 13968 4384 14032
rect 4448 13968 4464 14032
rect 4528 13968 4544 14032
rect 4608 13968 4624 14032
rect 4688 13968 4696 14032
rect 4376 12944 4696 13968
rect 4376 12880 4384 12944
rect 4448 12880 4464 12944
rect 4528 12880 4544 12944
rect 4608 12880 4624 12944
rect 4688 12880 4696 12944
rect 4376 11856 4696 12880
rect 4376 11792 4384 11856
rect 4448 11792 4464 11856
rect 4528 11792 4544 11856
rect 4608 11792 4624 11856
rect 4688 11792 4696 11856
rect 4376 10768 4696 11792
rect 4376 10704 4384 10768
rect 4448 10704 4464 10768
rect 4528 10704 4544 10768
rect 4608 10704 4624 10768
rect 4688 10704 4696 10768
rect 4376 9680 4696 10704
rect 4376 9616 4384 9680
rect 4448 9616 4464 9680
rect 4528 9616 4544 9680
rect 4608 9616 4624 9680
rect 4688 9616 4696 9680
rect 4376 8592 4696 9616
rect 4376 8528 4384 8592
rect 4448 8528 4464 8592
rect 4528 8528 4544 8592
rect 4608 8528 4624 8592
rect 4688 8528 4696 8592
rect 4376 7504 4696 8528
rect 4376 7440 4384 7504
rect 4448 7440 4464 7504
rect 4528 7440 4544 7504
rect 4608 7440 4624 7504
rect 4688 7440 4696 7504
rect 4376 6416 4696 7440
rect 4376 6352 4384 6416
rect 4448 6352 4464 6416
rect 4528 6352 4544 6416
rect 4608 6352 4624 6416
rect 4688 6352 4696 6416
rect 4376 5328 4696 6352
rect 4376 5264 4384 5328
rect 4448 5264 4464 5328
rect 4528 5264 4544 5328
rect 4608 5264 4624 5328
rect 4688 5264 4696 5328
rect 4376 4240 4696 5264
rect 4376 4176 4384 4240
rect 4448 4176 4464 4240
rect 4528 4176 4544 4240
rect 4608 4176 4624 4240
rect 4688 4176 4696 4240
rect 4376 3152 4696 4176
rect 4376 3088 4384 3152
rect 4448 3088 4464 3152
rect 4528 3088 4544 3152
rect 4608 3088 4624 3152
rect 4688 3088 4696 3152
rect 4376 2064 4696 3088
rect 4376 2000 4384 2064
rect 4448 2000 4464 2064
rect 4528 2000 4544 2064
rect 4608 2000 4624 2064
rect 4688 2000 4696 2064
rect 4376 1984 4696 2000
rect 7808 20016 8128 20032
rect 7808 19952 7816 20016
rect 7880 19952 7896 20016
rect 7960 19952 7976 20016
rect 8040 19952 8056 20016
rect 8120 19952 8128 20016
rect 7808 18928 8128 19952
rect 7808 18864 7816 18928
rect 7880 18864 7896 18928
rect 7960 18864 7976 18928
rect 8040 18864 8056 18928
rect 8120 18864 8128 18928
rect 7808 17840 8128 18864
rect 7808 17776 7816 17840
rect 7880 17776 7896 17840
rect 7960 17776 7976 17840
rect 8040 17776 8056 17840
rect 8120 17776 8128 17840
rect 7808 16752 8128 17776
rect 7808 16688 7816 16752
rect 7880 16688 7896 16752
rect 7960 16688 7976 16752
rect 8040 16688 8056 16752
rect 8120 16688 8128 16752
rect 7808 15664 8128 16688
rect 7808 15600 7816 15664
rect 7880 15600 7896 15664
rect 7960 15600 7976 15664
rect 8040 15600 8056 15664
rect 8120 15600 8128 15664
rect 7808 14576 8128 15600
rect 7808 14512 7816 14576
rect 7880 14512 7896 14576
rect 7960 14512 7976 14576
rect 8040 14512 8056 14576
rect 8120 14512 8128 14576
rect 7808 13488 8128 14512
rect 7808 13424 7816 13488
rect 7880 13424 7896 13488
rect 7960 13424 7976 13488
rect 8040 13424 8056 13488
rect 8120 13424 8128 13488
rect 7808 12400 8128 13424
rect 7808 12336 7816 12400
rect 7880 12336 7896 12400
rect 7960 12336 7976 12400
rect 8040 12336 8056 12400
rect 8120 12336 8128 12400
rect 7808 11312 8128 12336
rect 7808 11248 7816 11312
rect 7880 11248 7896 11312
rect 7960 11248 7976 11312
rect 8040 11248 8056 11312
rect 8120 11248 8128 11312
rect 7808 10224 8128 11248
rect 7808 10160 7816 10224
rect 7880 10160 7896 10224
rect 7960 10160 7976 10224
rect 8040 10160 8056 10224
rect 8120 10160 8128 10224
rect 7808 9136 8128 10160
rect 7808 9072 7816 9136
rect 7880 9072 7896 9136
rect 7960 9072 7976 9136
rect 8040 9072 8056 9136
rect 8120 9072 8128 9136
rect 7808 8048 8128 9072
rect 7808 7984 7816 8048
rect 7880 7984 7896 8048
rect 7960 7984 7976 8048
rect 8040 7984 8056 8048
rect 8120 7984 8128 8048
rect 7808 6960 8128 7984
rect 7808 6896 7816 6960
rect 7880 6896 7896 6960
rect 7960 6896 7976 6960
rect 8040 6896 8056 6960
rect 8120 6896 8128 6960
rect 7808 5872 8128 6896
rect 7808 5808 7816 5872
rect 7880 5808 7896 5872
rect 7960 5808 7976 5872
rect 8040 5808 8056 5872
rect 8120 5808 8128 5872
rect 7808 4784 8128 5808
rect 7808 4720 7816 4784
rect 7880 4720 7896 4784
rect 7960 4720 7976 4784
rect 8040 4720 8056 4784
rect 8120 4720 8128 4784
rect 7808 3696 8128 4720
rect 7808 3632 7816 3696
rect 7880 3632 7896 3696
rect 7960 3632 7976 3696
rect 8040 3632 8056 3696
rect 8120 3632 8128 3696
rect 7808 2608 8128 3632
rect 7808 2544 7816 2608
rect 7880 2544 7896 2608
rect 7960 2544 7976 2608
rect 8040 2544 8056 2608
rect 8120 2544 8128 2608
rect 7808 1984 8128 2544
rect 11240 19472 11560 20032
rect 11240 19408 11248 19472
rect 11312 19408 11328 19472
rect 11392 19408 11408 19472
rect 11472 19408 11488 19472
rect 11552 19408 11560 19472
rect 11240 18384 11560 19408
rect 11240 18320 11248 18384
rect 11312 18320 11328 18384
rect 11392 18320 11408 18384
rect 11472 18320 11488 18384
rect 11552 18320 11560 18384
rect 11240 17296 11560 18320
rect 11240 17232 11248 17296
rect 11312 17232 11328 17296
rect 11392 17232 11408 17296
rect 11472 17232 11488 17296
rect 11552 17232 11560 17296
rect 11240 16208 11560 17232
rect 11240 16144 11248 16208
rect 11312 16144 11328 16208
rect 11392 16144 11408 16208
rect 11472 16144 11488 16208
rect 11552 16144 11560 16208
rect 11240 15120 11560 16144
rect 11240 15056 11248 15120
rect 11312 15056 11328 15120
rect 11392 15056 11408 15120
rect 11472 15056 11488 15120
rect 11552 15056 11560 15120
rect 11240 14032 11560 15056
rect 11240 13968 11248 14032
rect 11312 13968 11328 14032
rect 11392 13968 11408 14032
rect 11472 13968 11488 14032
rect 11552 13968 11560 14032
rect 11240 12944 11560 13968
rect 11240 12880 11248 12944
rect 11312 12880 11328 12944
rect 11392 12880 11408 12944
rect 11472 12880 11488 12944
rect 11552 12880 11560 12944
rect 11240 11856 11560 12880
rect 11240 11792 11248 11856
rect 11312 11792 11328 11856
rect 11392 11792 11408 11856
rect 11472 11792 11488 11856
rect 11552 11792 11560 11856
rect 11240 10768 11560 11792
rect 11240 10704 11248 10768
rect 11312 10704 11328 10768
rect 11392 10704 11408 10768
rect 11472 10704 11488 10768
rect 11552 10704 11560 10768
rect 11240 9680 11560 10704
rect 11240 9616 11248 9680
rect 11312 9616 11328 9680
rect 11392 9616 11408 9680
rect 11472 9616 11488 9680
rect 11552 9616 11560 9680
rect 11240 8592 11560 9616
rect 11240 8528 11248 8592
rect 11312 8528 11328 8592
rect 11392 8528 11408 8592
rect 11472 8528 11488 8592
rect 11552 8528 11560 8592
rect 11240 7504 11560 8528
rect 11240 7440 11248 7504
rect 11312 7440 11328 7504
rect 11392 7440 11408 7504
rect 11472 7440 11488 7504
rect 11552 7440 11560 7504
rect 11240 6416 11560 7440
rect 11240 6352 11248 6416
rect 11312 6352 11328 6416
rect 11392 6352 11408 6416
rect 11472 6352 11488 6416
rect 11552 6352 11560 6416
rect 11240 5328 11560 6352
rect 11240 5264 11248 5328
rect 11312 5264 11328 5328
rect 11392 5264 11408 5328
rect 11472 5264 11488 5328
rect 11552 5264 11560 5328
rect 11240 4240 11560 5264
rect 11240 4176 11248 4240
rect 11312 4176 11328 4240
rect 11392 4176 11408 4240
rect 11472 4176 11488 4240
rect 11552 4176 11560 4240
rect 11240 3152 11560 4176
rect 11240 3088 11248 3152
rect 11312 3088 11328 3152
rect 11392 3088 11408 3152
rect 11472 3088 11488 3152
rect 11552 3088 11560 3152
rect 11240 2064 11560 3088
rect 11240 2000 11248 2064
rect 11312 2000 11328 2064
rect 11392 2000 11408 2064
rect 11472 2000 11488 2064
rect 11552 2000 11560 2064
rect 11240 1984 11560 2000
rect 14672 20016 14992 20032
rect 14672 19952 14680 20016
rect 14744 19952 14760 20016
rect 14824 19952 14840 20016
rect 14904 19952 14920 20016
rect 14984 19952 14992 20016
rect 14672 18928 14992 19952
rect 14672 18864 14680 18928
rect 14744 18864 14760 18928
rect 14824 18864 14840 18928
rect 14904 18864 14920 18928
rect 14984 18864 14992 18928
rect 14672 17840 14992 18864
rect 14672 17776 14680 17840
rect 14744 17776 14760 17840
rect 14824 17776 14840 17840
rect 14904 17776 14920 17840
rect 14984 17776 14992 17840
rect 14672 16752 14992 17776
rect 14672 16688 14680 16752
rect 14744 16688 14760 16752
rect 14824 16688 14840 16752
rect 14904 16688 14920 16752
rect 14984 16688 14992 16752
rect 14672 15664 14992 16688
rect 14672 15600 14680 15664
rect 14744 15600 14760 15664
rect 14824 15600 14840 15664
rect 14904 15600 14920 15664
rect 14984 15600 14992 15664
rect 14672 14576 14992 15600
rect 14672 14512 14680 14576
rect 14744 14512 14760 14576
rect 14824 14512 14840 14576
rect 14904 14512 14920 14576
rect 14984 14512 14992 14576
rect 14672 13488 14992 14512
rect 14672 13424 14680 13488
rect 14744 13424 14760 13488
rect 14824 13424 14840 13488
rect 14904 13424 14920 13488
rect 14984 13424 14992 13488
rect 14672 12400 14992 13424
rect 14672 12336 14680 12400
rect 14744 12336 14760 12400
rect 14824 12336 14840 12400
rect 14904 12336 14920 12400
rect 14984 12336 14992 12400
rect 14672 11312 14992 12336
rect 14672 11248 14680 11312
rect 14744 11248 14760 11312
rect 14824 11248 14840 11312
rect 14904 11248 14920 11312
rect 14984 11248 14992 11312
rect 14672 10224 14992 11248
rect 14672 10160 14680 10224
rect 14744 10160 14760 10224
rect 14824 10160 14840 10224
rect 14904 10160 14920 10224
rect 14984 10160 14992 10224
rect 14672 9136 14992 10160
rect 14672 9072 14680 9136
rect 14744 9072 14760 9136
rect 14824 9072 14840 9136
rect 14904 9072 14920 9136
rect 14984 9072 14992 9136
rect 14672 8048 14992 9072
rect 14672 7984 14680 8048
rect 14744 7984 14760 8048
rect 14824 7984 14840 8048
rect 14904 7984 14920 8048
rect 14984 7984 14992 8048
rect 14672 6960 14992 7984
rect 14672 6896 14680 6960
rect 14744 6896 14760 6960
rect 14824 6896 14840 6960
rect 14904 6896 14920 6960
rect 14984 6896 14992 6960
rect 14672 5872 14992 6896
rect 14672 5808 14680 5872
rect 14744 5808 14760 5872
rect 14824 5808 14840 5872
rect 14904 5808 14920 5872
rect 14984 5808 14992 5872
rect 14672 4784 14992 5808
rect 14672 4720 14680 4784
rect 14744 4720 14760 4784
rect 14824 4720 14840 4784
rect 14904 4720 14920 4784
rect 14984 4720 14992 4784
rect 14672 3696 14992 4720
rect 14672 3632 14680 3696
rect 14744 3632 14760 3696
rect 14824 3632 14840 3696
rect 14904 3632 14920 3696
rect 14984 3632 14992 3696
rect 14672 2608 14992 3632
rect 14672 2544 14680 2608
rect 14744 2544 14760 2608
rect 14824 2544 14840 2608
rect 14904 2544 14920 2608
rect 14984 2544 14992 2608
rect 14672 1984 14992 2544
rect 18104 19472 18424 20032
rect 18104 19408 18112 19472
rect 18176 19408 18192 19472
rect 18256 19408 18272 19472
rect 18336 19408 18352 19472
rect 18416 19408 18424 19472
rect 18104 18384 18424 19408
rect 18104 18320 18112 18384
rect 18176 18320 18192 18384
rect 18256 18320 18272 18384
rect 18336 18320 18352 18384
rect 18416 18320 18424 18384
rect 18104 17296 18424 18320
rect 18104 17232 18112 17296
rect 18176 17232 18192 17296
rect 18256 17232 18272 17296
rect 18336 17232 18352 17296
rect 18416 17232 18424 17296
rect 18104 16208 18424 17232
rect 18104 16144 18112 16208
rect 18176 16144 18192 16208
rect 18256 16144 18272 16208
rect 18336 16144 18352 16208
rect 18416 16144 18424 16208
rect 18104 15120 18424 16144
rect 18104 15056 18112 15120
rect 18176 15056 18192 15120
rect 18256 15056 18272 15120
rect 18336 15056 18352 15120
rect 18416 15056 18424 15120
rect 18104 14032 18424 15056
rect 18104 13968 18112 14032
rect 18176 13968 18192 14032
rect 18256 13968 18272 14032
rect 18336 13968 18352 14032
rect 18416 13968 18424 14032
rect 18104 12944 18424 13968
rect 18104 12880 18112 12944
rect 18176 12880 18192 12944
rect 18256 12880 18272 12944
rect 18336 12880 18352 12944
rect 18416 12880 18424 12944
rect 18104 11856 18424 12880
rect 18104 11792 18112 11856
rect 18176 11792 18192 11856
rect 18256 11792 18272 11856
rect 18336 11792 18352 11856
rect 18416 11792 18424 11856
rect 18104 10768 18424 11792
rect 18104 10704 18112 10768
rect 18176 10704 18192 10768
rect 18256 10704 18272 10768
rect 18336 10704 18352 10768
rect 18416 10704 18424 10768
rect 18104 9680 18424 10704
rect 18104 9616 18112 9680
rect 18176 9616 18192 9680
rect 18256 9616 18272 9680
rect 18336 9616 18352 9680
rect 18416 9616 18424 9680
rect 18104 8592 18424 9616
rect 18104 8528 18112 8592
rect 18176 8528 18192 8592
rect 18256 8528 18272 8592
rect 18336 8528 18352 8592
rect 18416 8528 18424 8592
rect 18104 7504 18424 8528
rect 18104 7440 18112 7504
rect 18176 7440 18192 7504
rect 18256 7440 18272 7504
rect 18336 7440 18352 7504
rect 18416 7440 18424 7504
rect 18104 6416 18424 7440
rect 18104 6352 18112 6416
rect 18176 6352 18192 6416
rect 18256 6352 18272 6416
rect 18336 6352 18352 6416
rect 18416 6352 18424 6416
rect 18104 5328 18424 6352
rect 18104 5264 18112 5328
rect 18176 5264 18192 5328
rect 18256 5264 18272 5328
rect 18336 5264 18352 5328
rect 18416 5264 18424 5328
rect 18104 4240 18424 5264
rect 18104 4176 18112 4240
rect 18176 4176 18192 4240
rect 18256 4176 18272 4240
rect 18336 4176 18352 4240
rect 18416 4176 18424 4240
rect 18104 3152 18424 4176
rect 18104 3088 18112 3152
rect 18176 3088 18192 3152
rect 18256 3088 18272 3152
rect 18336 3088 18352 3152
rect 18416 3088 18424 3152
rect 18104 2064 18424 3088
rect 18104 2000 18112 2064
rect 18176 2000 18192 2064
rect 18256 2000 18272 2064
rect 18336 2000 18352 2064
rect 18416 2000 18424 2064
rect 18104 1984 18424 2000
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1104 0 -1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606256979
transform 1 0 1104 0 1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 1380 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1606256979
transform 1 0 2484 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1606256979
transform 1 0 1380 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1606256979
transform 1 0 2484 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3956 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606256979
transform 1 0 3956 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 3588 0 -1 2576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1606256979
transform 1 0 4048 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_27
timestamp 1606256979
transform 1 0 3588 0 1 2576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_32
timestamp 1606256979
transform 1 0 4048 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606256979
transform 1 0 6808 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1606256979
transform 1 0 5152 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 6256 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_44
timestamp 1606256979
transform 1 0 5152 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_56
timestamp 1606256979
transform 1 0 6256 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1606256979
transform 1 0 6900 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1606256979
transform 1 0 8004 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_68
timestamp 1606256979
transform 1 0 7360 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_80
timestamp 1606256979
transform 1 0 8464 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606256979
transform 1 0 9660 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606256979
transform 1 0 9568 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1606256979
transform 1 0 9108 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1606256979
transform 1 0 9752 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1606256979
transform 1 0 9660 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606256979
transform 1 0 12512 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1606256979
transform 1 0 10856 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1606256979
transform 1 0 11960 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1606256979
transform 1 0 12604 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_105
timestamp 1606256979
transform 1 0 10764 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_117
timestamp 1606256979
transform 1 0 11868 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1606256979
transform 1 0 13708 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_129
timestamp 1606256979
transform 1 0 12972 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_141
timestamp 1606256979
transform 1 0 14076 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606256979
transform 1 0 15364 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606256979
transform 1 0 15180 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1606256979
transform 1 0 14812 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1606256979
transform 1 0 15456 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_154
timestamp 1606256979
transform 1 0 15272 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_166
timestamp 1606256979
transform 1 0 16376 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606256979
transform 1 0 18216 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1606256979
transform 1 0 16560 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1606256979
transform 1 0 17664 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1606256979
transform 1 0 18308 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_178
timestamp 1606256979
transform 1 0 17480 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1606256979
transform 1 0 19412 0 -1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_190
timestamp 1606256979
transform 1 0 18584 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_202
timestamp 1606256979
transform 1 0 19688 0 1 2576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606256979
transform -1 0 21620 0 -1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606256979
transform -1 0 21620 0 1 2576
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606256979
transform 1 0 21068 0 -1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606256979
transform 1 0 20792 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1606256979
transform 1 0 20516 0 -1 2576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 21160 0 -1 2576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1606256979
transform 1 0 20884 0 1 2576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_219 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 21252 0 1 2576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606256979
transform 1 0 1104 0 -1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1606256979
transform 1 0 1380 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1606256979
transform 1 0 2484 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_27
timestamp 1606256979
transform 1 0 3588 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_39
timestamp 1606256979
transform 1 0 4692 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606256979
transform 1 0 6716 0 -1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 5796 0 -1 3664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_59
timestamp 1606256979
transform 1 0 6532 0 -1 3664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_62
timestamp 1606256979
transform 1 0 6808 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_74
timestamp 1606256979
transform 1 0 7912 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_86
timestamp 1606256979
transform 1 0 9016 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_98
timestamp 1606256979
transform 1 0 10120 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606256979
transform 1 0 12328 0 -1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_110
timestamp 1606256979
transform 1 0 11224 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_123
timestamp 1606256979
transform 1 0 12420 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_135
timestamp 1606256979
transform 1 0 13524 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_147
timestamp 1606256979
transform 1 0 14628 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_159
timestamp 1606256979
transform 1 0 15732 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606256979
transform 1 0 17940 0 -1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_171
timestamp 1606256979
transform 1 0 16836 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_184
timestamp 1606256979
transform 1 0 18032 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_196
timestamp 1606256979
transform 1 0 19136 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_208
timestamp 1606256979
transform 1 0 20240 0 -1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606256979
transform -1 0 21620 0 -1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606256979
transform 1 0 1104 0 1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1606256979
transform 1 0 1380 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1606256979
transform 1 0 2484 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606256979
transform 1 0 3956 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1606256979
transform 1 0 3588 0 1 3664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_32
timestamp 1606256979
transform 1 0 4048 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_44
timestamp 1606256979
transform 1 0 5152 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_56
timestamp 1606256979
transform 1 0 6256 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_68
timestamp 1606256979
transform 1 0 7360 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_80
timestamp 1606256979
transform 1 0 8464 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606256979
transform 1 0 9568 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1606256979
transform 1 0 9660 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_105
timestamp 1606256979
transform 1 0 10764 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_117
timestamp 1606256979
transform 1 0 11868 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_129
timestamp 1606256979
transform 1 0 12972 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_141
timestamp 1606256979
transform 1 0 14076 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606256979
transform 1 0 15180 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_154
timestamp 1606256979
transform 1 0 15272 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_166
timestamp 1606256979
transform 1 0 16376 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_178
timestamp 1606256979
transform 1 0 17480 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_190
timestamp 1606256979
transform 1 0 18584 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_202
timestamp 1606256979
transform 1 0 19688 0 1 3664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606256979
transform -1 0 21620 0 1 3664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606256979
transform 1 0 20792 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_215
timestamp 1606256979
transform 1 0 20884 0 1 3664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_219
timestamp 1606256979
transform 1 0 21252 0 1 3664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606256979
transform 1 0 1104 0 -1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1606256979
transform 1 0 1380 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1606256979
transform 1 0 2484 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_27
timestamp 1606256979
transform 1 0 3588 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_39
timestamp 1606256979
transform 1 0 4692 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606256979
transform 1 0 6716 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_51
timestamp 1606256979
transform 1 0 5796 0 -1 4752
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_59
timestamp 1606256979
transform 1 0 6532 0 -1 4752
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_62
timestamp 1606256979
transform 1 0 6808 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_74
timestamp 1606256979
transform 1 0 7912 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_86
timestamp 1606256979
transform 1 0 9016 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_98
timestamp 1606256979
transform 1 0 10120 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606256979
transform 1 0 12328 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_110
timestamp 1606256979
transform 1 0 11224 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_123
timestamp 1606256979
transform 1 0 12420 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_135
timestamp 1606256979
transform 1 0 13524 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_147
timestamp 1606256979
transform 1 0 14628 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_159
timestamp 1606256979
transform 1 0 15732 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606256979
transform 1 0 17940 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_171
timestamp 1606256979
transform 1 0 16836 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_184
timestamp 1606256979
transform 1 0 18032 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_196
timestamp 1606256979
transform 1 0 19136 0 -1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_208
timestamp 1606256979
transform 1 0 20240 0 -1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _68_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 20516 0 -1 4752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606256979
transform -1 0 21620 0 -1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1606256979
transform 1 0 20884 0 -1 4752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1606256979
transform 1 0 21252 0 -1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606256979
transform 1 0 1104 0 1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1606256979
transform 1 0 1380 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1606256979
transform 1 0 2484 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606256979
transform 1 0 3956 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_27
timestamp 1606256979
transform 1 0 3588 0 1 4752
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_32
timestamp 1606256979
transform 1 0 4048 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_44
timestamp 1606256979
transform 1 0 5152 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_56
timestamp 1606256979
transform 1 0 6256 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_68
timestamp 1606256979
transform 1 0 7360 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_80
timestamp 1606256979
transform 1 0 8464 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606256979
transform 1 0 9568 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1606256979
transform 1 0 9660 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_105
timestamp 1606256979
transform 1 0 10764 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_117
timestamp 1606256979
transform 1 0 11868 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_129
timestamp 1606256979
transform 1 0 12972 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_141
timestamp 1606256979
transform 1 0 14076 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606256979
transform 1 0 15180 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_154
timestamp 1606256979
transform 1 0 15272 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_166
timestamp 1606256979
transform 1 0 16376 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_178
timestamp 1606256979
transform 1 0 17480 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_190
timestamp 1606256979
transform 1 0 18584 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_202
timestamp 1606256979
transform 1 0 19688 0 1 4752
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606256979
transform -1 0 21620 0 1 4752
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606256979
transform 1 0 20792 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_215
timestamp 1606256979
transform 1 0 20884 0 1 4752
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_219
timestamp 1606256979
transform 1 0 21252 0 1 4752
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606256979
transform 1 0 1104 0 -1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606256979
transform 1 0 1104 0 1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1606256979
transform 1 0 1380 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1606256979
transform 1 0 2484 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1606256979
transform 1 0 1380 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1606256979
transform 1 0 2484 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606256979
transform 1 0 3956 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_27
timestamp 1606256979
transform 1 0 3588 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_39
timestamp 1606256979
transform 1 0 4692 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_27
timestamp 1606256979
transform 1 0 3588 0 1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_32
timestamp 1606256979
transform 1 0 4048 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606256979
transform 1 0 6716 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_51
timestamp 1606256979
transform 1 0 5796 0 -1 5840
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_59
timestamp 1606256979
transform 1 0 6532 0 -1 5840
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_62
timestamp 1606256979
transform 1 0 6808 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_44
timestamp 1606256979
transform 1 0 5152 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_56
timestamp 1606256979
transform 1 0 6256 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_74
timestamp 1606256979
transform 1 0 7912 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_68
timestamp 1606256979
transform 1 0 7360 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_80
timestamp 1606256979
transform 1 0 8464 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606256979
transform 1 0 9568 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_86
timestamp 1606256979
transform 1 0 9016 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_98
timestamp 1606256979
transform 1 0 10120 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1606256979
transform 1 0 9660 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606256979
transform 1 0 12328 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_110
timestamp 1606256979
transform 1 0 11224 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_123
timestamp 1606256979
transform 1 0 12420 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_105
timestamp 1606256979
transform 1 0 10764 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_117
timestamp 1606256979
transform 1 0 11868 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_135
timestamp 1606256979
transform 1 0 13524 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_129
timestamp 1606256979
transform 1 0 12972 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_141
timestamp 1606256979
transform 1 0 14076 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606256979
transform 1 0 15180 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_147
timestamp 1606256979
transform 1 0 14628 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_159
timestamp 1606256979
transform 1 0 15732 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_154
timestamp 1606256979
transform 1 0 15272 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_166
timestamp 1606256979
transform 1 0 16376 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606256979
transform 1 0 17940 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_171
timestamp 1606256979
transform 1 0 16836 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_184
timestamp 1606256979
transform 1 0 18032 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_178
timestamp 1606256979
transform 1 0 17480 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_196
timestamp 1606256979
transform 1 0 19136 0 -1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_208
timestamp 1606256979
transform 1 0 20240 0 -1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_190
timestamp 1606256979
transform 1 0 18584 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_202
timestamp 1606256979
transform 1 0 19688 0 1 5840
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _86_
timestamp 1606256979
transform 1 0 20516 0 -1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606256979
transform -1 0 21620 0 -1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606256979
transform -1 0 21620 0 1 5840
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606256979
transform 1 0 20792 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1606256979
transform 1 0 20884 0 -1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1606256979
transform 1 0 21252 0 -1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_215
timestamp 1606256979
transform 1 0 20884 0 1 5840
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_219
timestamp 1606256979
transform 1 0 21252 0 1 5840
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606256979
transform 1 0 1104 0 -1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1606256979
transform 1 0 1380 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1606256979
transform 1 0 2484 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_27
timestamp 1606256979
transform 1 0 3588 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_39
timestamp 1606256979
transform 1 0 4692 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606256979
transform 1 0 6716 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_51
timestamp 1606256979
transform 1 0 5796 0 -1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_59
timestamp 1606256979
transform 1 0 6532 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_62
timestamp 1606256979
transform 1 0 6808 0 -1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 7268 0 -1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_66
timestamp 1606256979
transform 1 0 7176 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_83
timestamp 1606256979
transform 1 0 8740 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 10580 0 -1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_95
timestamp 1606256979
transform 1 0 9844 0 -1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606256979
transform 1 0 12328 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_112
timestamp 1606256979
transform 1 0 11408 0 -1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_120
timestamp 1606256979
transform 1 0 12144 0 -1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1606256979
transform 1 0 12420 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1606256979
transform 1 0 14076 0 -1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_8_135
timestamp 1606256979
transform 1 0 13524 0 -1 6928
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_150
timestamp 1606256979
transform 1 0 14904 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_162
timestamp 1606256979
transform 1 0 16008 0 -1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1606256979
transform 1 0 16836 0 -1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606256979
transform 1 0 17940 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_170
timestamp 1606256979
transform 1 0 16744 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_180
timestamp 1606256979
transform 1 0 17664 0 -1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_184
timestamp 1606256979
transform 1 0 18032 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_196
timestamp 1606256979
transform 1 0 19136 0 -1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_208
timestamp 1606256979
transform 1 0 20240 0 -1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _84_
timestamp 1606256979
transform 1 0 20516 0 -1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606256979
transform -1 0 21620 0 -1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1606256979
transform 1 0 20884 0 -1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1606256979
transform 1 0 21252 0 -1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606256979
transform 1 0 1104 0 1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1606256979
transform 1 0 1380 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1606256979
transform 1 0 2484 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606256979
transform 1 0 3956 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1606256979
transform 1 0 3588 0 1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_32
timestamp 1606256979
transform 1 0 4048 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_44
timestamp 1606256979
transform 1 0 5152 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_56
timestamp 1606256979
transform 1 0 6256 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_68
timestamp 1606256979
transform 1 0 7360 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_80
timestamp 1606256979
transform 1 0 8464 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _31_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 9752 0 1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10212 0 1 6928
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606256979
transform 1 0 9568 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_93
timestamp 1606256979
transform 1 0 9660 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_97
timestamp 1606256979
transform 1 0 10028 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 11224 0 1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_108
timestamp 1606256979
transform 1 0 11040 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12880 0 1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_126
timestamp 1606256979
transform 1 0 12696 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_144
timestamp 1606256979
transform 1 0 14352 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1606256979
transform 1 0 14536 0 1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 16192 0 1 6928
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606256979
transform 1 0 15180 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_149
timestamp 1606256979
transform 1 0 14812 0 1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_154
timestamp 1606256979
transform 1 0 15272 0 1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_162
timestamp 1606256979
transform 1 0 16008 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_180
timestamp 1606256979
transform 1 0 17664 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_192
timestamp 1606256979
transform 1 0 18768 0 1 6928
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_204
timestamp 1606256979
transform 1 0 19872 0 1 6928
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606256979
transform -1 0 21620 0 1 6928
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606256979
transform 1 0 20792 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_212
timestamp 1606256979
transform 1 0 20608 0 1 6928
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_215
timestamp 1606256979
transform 1 0 20884 0 1 6928
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_219
timestamp 1606256979
transform 1 0 21252 0 1 6928
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606256979
transform 1 0 1104 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1606256979
transform 1 0 1380 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1606256979
transform 1 0 2484 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_27
timestamp 1606256979
transform 1 0 3588 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_39
timestamp 1606256979
transform 1 0 4692 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606256979
transform 1 0 6716 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_51
timestamp 1606256979
transform 1 0 5796 0 -1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_59
timestamp 1606256979
transform 1 0 6532 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_62
timestamp 1606256979
transform 1 0 6808 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_74
timestamp 1606256979
transform 1 0 7912 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9200 0 -1 8016
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_86
timestamp 1606256979
transform 1 0 9016 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_104
timestamp 1606256979
transform 1 0 10672 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 10856 0 -1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606256979
transform 1 0 12328 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_112
timestamp 1606256979
transform 1 0 11408 0 -1 8016
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_120
timestamp 1606256979
transform 1 0 12144 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_123
timestamp 1606256979
transform 1 0 12420 0 -1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1606256979
transform 1 0 13708 0 -1 8016
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_135
timestamp 1606256979
transform 1 0 13524 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 14720 0 -1 8016
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16376 0 -1 8016
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_146
timestamp 1606256979
transform 1 0 14536 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_164
timestamp 1606256979
transform 1 0 16192 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1606256979
transform 1 0 17388 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 18032 0 -1 8016
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606256979
transform 1 0 17940 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_175
timestamp 1606256979
transform 1 0 17204 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_180
timestamp 1606256979
transform 1 0 17664 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _82_
timestamp 1606256979
transform 1 0 19964 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_200
timestamp 1606256979
transform 1 0 19504 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_204
timestamp 1606256979
transform 1 0 19872 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _81_
timestamp 1606256979
transform 1 0 20516 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606256979
transform -1 0 21620 0 -1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_209
timestamp 1606256979
transform 1 0 20332 0 -1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_215
timestamp 1606256979
transform 1 0 20884 0 -1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_219
timestamp 1606256979
transform 1 0 21252 0 -1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606256979
transform 1 0 1104 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1606256979
transform 1 0 1380 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1606256979
transform 1 0 2484 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606256979
transform 1 0 3956 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1606256979
transform 1 0 3588 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_32
timestamp 1606256979
transform 1 0 4048 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_44
timestamp 1606256979
transform 1 0 5152 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_56
timestamp 1606256979
transform 1 0 6256 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_68
timestamp 1606256979
transform 1 0 7360 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_80
timestamp 1606256979
transform 1 0 8464 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606256979
transform 1 0 9568 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1606256979
transform 1 0 9660 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _87_
timestamp 1606256979
transform 1 0 11224 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_105
timestamp 1606256979
transform 1 0 10764 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_109
timestamp 1606256979
transform 1 0 11132 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_114
timestamp 1606256979
transform 1 0 11592 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 13340 0 1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_126
timestamp 1606256979
transform 1 0 12696 0 1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_132
timestamp 1606256979
transform 1 0 13248 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_139
timestamp 1606256979
transform 1 0 13892 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606256979
transform 1 0 15180 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_151
timestamp 1606256979
transform 1 0 14996 0 1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_154
timestamp 1606256979
transform 1 0 15272 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_166
timestamp 1606256979
transform 1 0 16376 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_178
timestamp 1606256979
transform 1 0 17480 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1606256979
transform 1 0 20240 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_190
timestamp 1606256979
transform 1 0 18584 0 1 8016
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_202
timestamp 1606256979
transform 1 0 19688 0 1 8016
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606256979
transform -1 0 21620 0 1 8016
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606256979
transform 1 0 20792 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_212
timestamp 1606256979
transform 1 0 20608 0 1 8016
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_215
timestamp 1606256979
transform 1 0 20884 0 1 8016
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_219
timestamp 1606256979
transform 1 0 21252 0 1 8016
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606256979
transform 1 0 1104 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1606256979
transform 1 0 1380 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1606256979
transform 1 0 2484 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_27
timestamp 1606256979
transform 1 0 3588 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_39
timestamp 1606256979
transform 1 0 4692 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606256979
transform 1 0 6716 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_51
timestamp 1606256979
transform 1 0 5796 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_59
timestamp 1606256979
transform 1 0 6532 0 -1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_62
timestamp 1606256979
transform 1 0 6808 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_74
timestamp 1606256979
transform 1 0 7912 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_86
timestamp 1606256979
transform 1 0 9016 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_98
timestamp 1606256979
transform 1 0 10120 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1606256979
transform 1 0 11040 0 -1 9104
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606256979
transform 1 0 12328 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_106
timestamp 1606256979
transform 1 0 10856 0 -1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_117
timestamp 1606256979
transform 1 0 11868 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_121
timestamp 1606256979
transform 1 0 12236 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_123
timestamp 1606256979
transform 1 0 12420 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _85_
timestamp 1606256979
transform 1 0 13248 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_131
timestamp 1606256979
transform 1 0 13156 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_136
timestamp 1606256979
transform 1 0 13616 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 15456 0 -1 9104
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_12_148
timestamp 1606256979
transform 1 0 14720 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_162
timestamp 1606256979
transform 1 0 16008 0 -1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 18308 0 -1 9104
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606256979
transform 1 0 17940 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_174
timestamp 1606256979
transform 1 0 17112 0 -1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_182
timestamp 1606256979
transform 1 0 17848 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_184
timestamp 1606256979
transform 1 0 18032 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1606256979
transform 1 0 19964 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_203
timestamp 1606256979
transform 1 0 19780 0 -1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1606256979
transform 1 0 20516 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606256979
transform -1 0 21620 0 -1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_209
timestamp 1606256979
transform 1 0 20332 0 -1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1606256979
transform 1 0 20884 0 -1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1606256979
transform 1 0 21252 0 -1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606256979
transform 1 0 1104 0 1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606256979
transform 1 0 1104 0 -1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1606256979
transform 1 0 1380 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1606256979
transform 1 0 2484 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1606256979
transform 1 0 1380 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1606256979
transform 1 0 2484 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606256979
transform 1 0 3956 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_27
timestamp 1606256979
transform 1 0 3588 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_32
timestamp 1606256979
transform 1 0 4048 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_27
timestamp 1606256979
transform 1 0 3588 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_39
timestamp 1606256979
transform 1 0 4692 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606256979
transform 1 0 6716 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_44
timestamp 1606256979
transform 1 0 5152 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_56
timestamp 1606256979
transform 1 0 6256 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_51
timestamp 1606256979
transform 1 0 5796 0 -1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_59
timestamp 1606256979
transform 1 0 6532 0 -1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_62
timestamp 1606256979
transform 1 0 6808 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 7912 0 1 9104
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 8096 0 -1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_13_68
timestamp 1606256979
transform 1 0 7360 0 1 9104
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_74
timestamp 1606256979
transform 1 0 7912 0 -1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10580 0 -1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606256979
transform 1 0 9568 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_90
timestamp 1606256979
transform 1 0 9384 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1606256979
transform 1 0 9660 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_92
timestamp 1606256979
transform 1 0 9568 0 -1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_100
timestamp 1606256979
transform 1 0 10304 0 -1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1606256979
transform 1 0 11776 0 1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1606256979
transform 1 0 12328 0 1 9104
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1606256979
transform 1 0 10764 0 1 9104
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606256979
transform 1 0 12328 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_114
timestamp 1606256979
transform 1 0 11592 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_119
timestamp 1606256979
transform 1 0 12052 0 1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_112
timestamp 1606256979
transform 1 0 11408 0 -1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_120
timestamp 1606256979
transform 1 0 12144 0 -1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_123
timestamp 1606256979
transform 1 0 12420 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13524 0 1 9104
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_13_131
timestamp 1606256979
transform 1 0 13156 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_135
timestamp 1606256979
transform 1 0 13524 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _83_
timestamp 1606256979
transform 1 0 15272 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15916 0 -1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606256979
transform 1 0 15180 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_151
timestamp 1606256979
transform 1 0 14996 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_158
timestamp 1606256979
transform 1 0 15640 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_147
timestamp 1606256979
transform 1 0 14628 0 -1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_159
timestamp 1606256979
transform 1 0 15732 0 -1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1606256979
transform 1 0 18032 0 -1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606256979
transform 1 0 17940 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_170
timestamp 1606256979
transform 1 0 16744 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_182
timestamp 1606256979
transform 1 0 17848 0 1 9104
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_177
timestamp 1606256979
transform 1 0 17388 0 -1 10192
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_187
timestamp 1606256979
transform 1 0 18308 0 -1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 18492 0 -1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1606256979
transform 1 0 18676 0 1 9104
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_190
timestamp 1606256979
transform 1 0 18584 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_200
timestamp 1606256979
transform 1 0 19504 0 1 9104
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_205
timestamp 1606256979
transform 1 0 19964 0 -1 10192
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1606256979
transform 1 0 20516 0 -1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606256979
transform -1 0 21620 0 1 9104
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606256979
transform -1 0 21620 0 -1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606256979
transform 1 0 20792 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_212
timestamp 1606256979
transform 1 0 20608 0 1 9104
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_215
timestamp 1606256979
transform 1 0 20884 0 1 9104
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_219
timestamp 1606256979
transform 1 0 21252 0 1 9104
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1606256979
transform 1 0 20884 0 -1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1606256979
transform 1 0 21252 0 -1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606256979
transform 1 0 1104 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1606256979
transform 1 0 1380 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1606256979
transform 1 0 2484 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606256979
transform 1 0 3956 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1606256979
transform 1 0 3588 0 1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_32
timestamp 1606256979
transform 1 0 4048 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_44
timestamp 1606256979
transform 1 0 5152 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_56
timestamp 1606256979
transform 1 0 6256 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7176 0 1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_64
timestamp 1606256979
transform 1 0 6992 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_82
timestamp 1606256979
transform 1 0 8648 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1606256979
transform 1 0 10212 0 1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606256979
transform 1 0 9568 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_90
timestamp 1606256979
transform 1 0 9384 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_93
timestamp 1606256979
transform 1 0 9660 0 1 10192
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11224 0 1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_108
timestamp 1606256979
transform 1 0 11040 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_119
timestamp 1606256979
transform 1 0 12052 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 12788 0 1 10192
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_15_143
timestamp 1606256979
transform 1 0 14260 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606256979
transform 1 0 15180 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_151
timestamp 1606256979
transform 1 0 14996 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_154
timestamp 1606256979
transform 1 0 15272 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_166
timestamp 1606256979
transform 1 0 16376 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1606256979
transform 1 0 16468 0 1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_15_176
timestamp 1606256979
transform 1 0 17296 0 1 10192
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1606256979
transform 1 0 20240 0 1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1606256979
transform 1 0 18676 0 1 10192
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_15_188
timestamp 1606256979
transform 1 0 18400 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_200
timestamp 1606256979
transform 1 0 19504 0 1 10192
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606256979
transform -1 0 21620 0 1 10192
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606256979
transform 1 0 20792 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_212
timestamp 1606256979
transform 1 0 20608 0 1 10192
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_215
timestamp 1606256979
transform 1 0 20884 0 1 10192
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_219
timestamp 1606256979
transform 1 0 21252 0 1 10192
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606256979
transform 1 0 1104 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1606256979
transform 1 0 1380 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1606256979
transform 1 0 2484 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_27
timestamp 1606256979
transform 1 0 3588 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_39
timestamp 1606256979
transform 1 0 4692 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606256979
transform 1 0 6716 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_51
timestamp 1606256979
transform 1 0 5796 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_59
timestamp 1606256979
transform 1 0 6532 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_62
timestamp 1606256979
transform 1 0 6808 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1606256979
transform 1 0 8188 0 -1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_16_74
timestamp 1606256979
transform 1 0 7912 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_86
timestamp 1606256979
transform 1 0 9016 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_98
timestamp 1606256979
transform 1 0 10120 0 -1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_104
timestamp 1606256979
transform 1 0 10672 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 10764 0 -1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606256979
transform 1 0 12328 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_111
timestamp 1606256979
transform 1 0 11316 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_119
timestamp 1606256979
transform 1 0 12052 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_123
timestamp 1606256979
transform 1 0 12420 0 -1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1606256979
transform 1 0 13708 0 -1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_135
timestamp 1606256979
transform 1 0 13524 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1606256979
transform 1 0 14720 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15916 0 -1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_146
timestamp 1606256979
transform 1 0 14536 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_151
timestamp 1606256979
transform 1 0 14996 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_159
timestamp 1606256979
transform 1 0 15732 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16928 0 -1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606256979
transform 1 0 17940 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1606256979
transform 1 0 16744 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_181
timestamp 1606256979
transform 1 0 17756 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_184
timestamp 1606256979
transform 1 0 18032 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1606256979
transform 1 0 18768 0 -1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_201
timestamp 1606256979
transform 1 0 19596 0 -1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1606256979
transform 1 0 20516 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606256979
transform -1 0 21620 0 -1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_209
timestamp 1606256979
transform 1 0 20332 0 -1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1606256979
transform 1 0 20884 0 -1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1606256979
transform 1 0 21252 0 -1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606256979
transform 1 0 1104 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1606256979
transform 1 0 1380 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1606256979
transform 1 0 2484 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606256979
transform 1 0 3956 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_27
timestamp 1606256979
transform 1 0 3588 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_32
timestamp 1606256979
transform 1 0 4048 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1606256979
transform 1 0 6808 0 1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_17_44
timestamp 1606256979
transform 1 0 5152 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_56
timestamp 1606256979
transform 1 0 6256 0 1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1606256979
transform 1 0 7912 0 1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_17_71
timestamp 1606256979
transform 1 0 7636 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_83
timestamp 1606256979
transform 1 0 8740 0 1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1606256979
transform 1 0 10304 0 1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606256979
transform 1 0 9568 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_91
timestamp 1606256979
transform 1 0 9476 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_93
timestamp 1606256979
transform 1 0 9660 0 1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_99
timestamp 1606256979
transform 1 0 10212 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1606256979
transform 1 0 11316 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_109
timestamp 1606256979
transform 1 0 11132 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_114
timestamp 1606256979
transform 1 0 11592 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1606256979
transform 1 0 13616 0 1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_right_track_0.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 13340 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_126
timestamp 1606256979
transform 1 0 12696 0 1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_132
timestamp 1606256979
transform 1 0 13248 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_145
timestamp 1606256979
transform 1 0 14444 0 1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606256979
transform 1 0 15180 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_154
timestamp 1606256979
transform 1 0 15272 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_166
timestamp 1606256979
transform 1 0 16376 0 1 11280
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1606256979
transform 1 0 18032 0 1 11280
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_17_178
timestamp 1606256979
transform 1 0 17480 0 1 11280
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1606256979
transform 1 0 19044 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1606256979
transform 1 0 20240 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_193
timestamp 1606256979
transform 1 0 18860 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_198
timestamp 1606256979
transform 1 0 19320 0 1 11280
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_206
timestamp 1606256979
transform 1 0 20056 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606256979
transform -1 0 21620 0 1 11280
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606256979
transform 1 0 20792 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_212
timestamp 1606256979
transform 1 0 20608 0 1 11280
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_215
timestamp 1606256979
transform 1 0 20884 0 1 11280
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_219
timestamp 1606256979
transform 1 0 21252 0 1 11280
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606256979
transform 1 0 1104 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1606256979
transform 1 0 1380 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1606256979
transform 1 0 2484 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_27
timestamp 1606256979
transform 1 0 3588 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_39
timestamp 1606256979
transform 1 0 4692 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606256979
transform 1 0 6716 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_51
timestamp 1606256979
transform 1 0 5796 0 -1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_59
timestamp 1606256979
transform 1 0 6532 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_62
timestamp 1606256979
transform 1 0 6808 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6992 0 -1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 8648 0 -1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_18_80
timestamp 1606256979
transform 1 0 8464 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1606256979
transform 1 0 10304 0 -1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_98
timestamp 1606256979
transform 1 0 10120 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12420 0 -1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606256979
transform 1 0 12328 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1606256979
transform 1 0 11132 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_121
timestamp 1606256979
transform 1 0 12236 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1606256979
transform 1 0 14076 0 -1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_139
timestamp 1606256979
transform 1 0 13892 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15272 0 -1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_150
timestamp 1606256979
transform 1 0 14904 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1606256979
transform 1 0 18032 0 -1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606256979
transform 1 0 17940 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_170
timestamp 1606256979
transform 1 0 16744 0 -1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_182
timestamp 1606256979
transform 1 0 17848 0 -1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1606256979
transform 1 0 19872 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_193
timestamp 1606256979
transform 1 0 18860 0 -1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_201
timestamp 1606256979
transform 1 0 19596 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_208
timestamp 1606256979
transform 1 0 20240 0 -1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1606256979
transform 1 0 20424 0 -1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606256979
transform -1 0 21620 0 -1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_214
timestamp 1606256979
transform 1 0 20792 0 -1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606256979
transform 1 0 1104 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606256979
transform 1 0 1104 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1606256979
transform 1 0 1380 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1606256979
transform 1 0 2484 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1606256979
transform 1 0 1380 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1606256979
transform 1 0 2484 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 3864 0 -1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606256979
transform 1 0 3956 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_27
timestamp 1606256979
transform 1 0 3588 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_32
timestamp 1606256979
transform 1 0 4048 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_27
timestamp 1606256979
transform 1 0 3588 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1606256979
transform 1 0 5612 0 -1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606256979
transform 1 0 6716 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_44
timestamp 1606256979
transform 1 0 5152 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_56
timestamp 1606256979
transform 1 0 6256 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_46
timestamp 1606256979
transform 1 0 5336 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_58
timestamp 1606256979
transform 1 0 6440 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_62
timestamp 1606256979
transform 1 0 6808 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_right_track_0.prog_clk
timestamp 1606256979
transform 1 0 7636 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_68
timestamp 1606256979
transform 1 0 7360 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1606256979
transform 1 0 7912 0 1 12368
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_74
timestamp 1606256979
transform 1 0 7912 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 9844 0 1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606256979
transform 1 0 9568 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_right_track_0.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 10028 0 -1 13456
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_19_86
timestamp 1606256979
transform 1 0 9016 0 1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_93
timestamp 1606256979
transform 1 0 9660 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_86
timestamp 1606256979
transform 1 0 9016 0 -1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_94
timestamp 1606256979
transform 1 0 9752 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 11316 0 1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606256979
transform 1 0 12328 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_right_track_0.prog_clk
timestamp 1606256979
transform 1 0 12420 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_117
timestamp 1606256979
transform 1 0 11868 0 1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_117
timestamp 1606256979
transform 1 0 11868 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_121
timestamp 1606256979
transform 1 0 12236 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_123
timestamp 1606256979
transform 1 0 12420 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12880 0 1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1606256979
transform 1 0 14076 0 1 12368
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_126
timestamp 1606256979
transform 1 0 12696 0 1 12368
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_137
timestamp 1606256979
transform 1 0 13708 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_135
timestamp 1606256979
transform 1 0 13524 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 15272 0 1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606256979
transform 1 0 15180 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_150
timestamp 1606256979
transform 1 0 14904 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_160
timestamp 1606256979
transform 1 0 15824 0 1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_147
timestamp 1606256979
transform 1 0 14628 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_159
timestamp 1606256979
transform 1 0 15732 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606256979
transform 1 0 16560 0 1 12368
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 18308 0 -1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606256979
transform 1 0 17940 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_184
timestamp 1606256979
transform 1 0 18032 0 1 12368
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_171
timestamp 1606256979
transform 1 0 16836 0 -1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_184
timestamp 1606256979
transform 1 0 18032 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1606256979
transform 1 0 19872 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1606256979
transform 1 0 19412 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1606256979
transform 1 0 19964 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19044 0 1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_192
timestamp 1606256979
transform 1 0 18768 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_201
timestamp 1606256979
transform 1 0 19596 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_208
timestamp 1606256979
transform 1 0 20240 0 1 12368
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_193
timestamp 1606256979
transform 1 0 18860 0 -1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_203
timestamp 1606256979
transform 1 0 19780 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1606256979
transform 1 0 20516 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606256979
transform -1 0 21620 0 1 12368
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606256979
transform -1 0 21620 0 -1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606256979
transform 1 0 20792 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_215
timestamp 1606256979
transform 1 0 20884 0 1 12368
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_219
timestamp 1606256979
transform 1 0 21252 0 1 12368
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_209
timestamp 1606256979
transform 1 0 20332 0 -1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1606256979
transform 1 0 20884 0 -1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1606256979
transform 1 0 21252 0 -1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606256979
transform 1 0 1104 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1606256979
transform 1 0 1380 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1606256979
transform 1 0 2484 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4784 0 1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606256979
transform 1 0 3956 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_27
timestamp 1606256979
transform 1 0 3588 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_32
timestamp 1606256979
transform 1 0 4048 0 1 13456
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1606256979
transform 1 0 6440 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_56
timestamp 1606256979
transform 1 0 6256 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_61
timestamp 1606256979
transform 1 0 6716 0 1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7268 0 1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_83
timestamp 1606256979
transform 1 0 8740 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606256979
transform 1 0 9568 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_right_track_0.prog_clk
timestamp 1606256979
transform 1 0 8924 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_88
timestamp 1606256979
transform 1 0 9200 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1606256979
transform 1 0 9660 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 10948 0 1 13456
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1606256979
transform 1 0 12604 0 1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_105
timestamp 1606256979
transform 1 0 10764 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1606256979
transform 1 0 12420 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1606256979
transform 1 0 13616 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_134
timestamp 1606256979
transform 1 0 13432 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_139
timestamp 1606256979
transform 1 0 13892 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606256979
transform 1 0 15180 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_151
timestamp 1606256979
transform 1 0 14996 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_154
timestamp 1606256979
transform 1 0 15272 0 1 13456
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_166
timestamp 1606256979
transform 1 0 16376 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1606256979
transform 1 0 16468 0 1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1606256979
transform 1 0 17480 0 1 13456
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_176
timestamp 1606256979
transform 1 0 17296 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_187
timestamp 1606256979
transform 1 0 18308 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1606256979
transform 1 0 20240 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1606256979
transform 1 0 19688 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1606256979
transform 1 0 18768 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_191
timestamp 1606256979
transform 1 0 18676 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_196
timestamp 1606256979
transform 1 0 19136 0 1 13456
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_206
timestamp 1606256979
transform 1 0 20056 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606256979
transform -1 0 21620 0 1 13456
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606256979
transform 1 0 20792 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_212
timestamp 1606256979
transform 1 0 20608 0 1 13456
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_215
timestamp 1606256979
transform 1 0 20884 0 1 13456
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_219
timestamp 1606256979
transform 1 0 21252 0 1 13456
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2208 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606256979
transform 1 0 1104 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1606256979
transform 1 0 1380 0 -1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_11
timestamp 1606256979
transform 1 0 2116 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_28
timestamp 1606256979
transform 1 0 3680 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_40
timestamp 1606256979
transform 1 0 4784 0 -1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1606256979
transform 1 0 5704 0 -1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606256979
transform 1 0 6716 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_48
timestamp 1606256979
transform 1 0 5520 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_59
timestamp 1606256979
transform 1 0 6532 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_62
timestamp 1606256979
transform 1 0 6808 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8280 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_22_74
timestamp 1606256979
transform 1 0 7912 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_94
timestamp 1606256979
transform 1 0 9752 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12420 0 -1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606256979
transform 1 0 12328 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_106
timestamp 1606256979
transform 1 0 10856 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_118
timestamp 1606256979
transform 1 0 11960 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13892 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_22_132
timestamp 1606256979
transform 1 0 13248 0 -1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_138
timestamp 1606256979
transform 1 0 13800 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15548 0 -1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_155
timestamp 1606256979
transform 1 0 15364 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1606256979
transform 1 0 17388 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606256979
transform 1 0 17940 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_173
timestamp 1606256979
transform 1 0 17020 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_180
timestamp 1606256979
transform 1 0 17664 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_184
timestamp 1606256979
transform 1 0 18032 0 -1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19228 0 -1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19964 0 -1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_196
timestamp 1606256979
transform 1 0 19136 0 -1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_203
timestamp 1606256979
transform 1 0 19780 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1606256979
transform 1 0 20700 0 -1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606256979
transform -1 0 21620 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_211
timestamp 1606256979
transform 1 0 20516 0 -1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_217
timestamp 1606256979
transform 1 0 21068 0 -1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 1564 0 1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606256979
transform 1 0 1104 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1606256979
transform 1 0 1380 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1606256979
transform 1 0 3404 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4048 0 1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606256979
transform 1 0 3956 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_21
timestamp 1606256979
transform 1 0 3036 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_28
timestamp 1606256979
transform 1 0 3680 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_41
timestamp 1606256979
transform 1 0 4876 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_53
timestamp 1606256979
transform 1 0 5980 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1606256979
transform 1 0 7912 0 1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_65
timestamp 1606256979
transform 1 0 7084 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_73
timestamp 1606256979
transform 1 0 7820 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_83
timestamp 1606256979
transform 1 0 8740 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1606256979
transform 1 0 10672 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9660 0 1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606256979
transform 1 0 9568 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_91
timestamp 1606256979
transform 1 0 9476 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_102
timestamp 1606256979
transform 1 0 10488 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11960 0 1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_23_107
timestamp 1606256979
transform 1 0 10948 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_115
timestamp 1606256979
transform 1 0 11684 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 13524 0 1 14544
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_right_track_0.prog_clk
timestamp 1606256979
transform 1 0 13156 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_127
timestamp 1606256979
transform 1 0 12788 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_134
timestamp 1606256979
transform 1 0 13432 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606256979
transform 1 0 15180 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_151
timestamp 1606256979
transform 1 0 14996 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_154
timestamp 1606256979
transform 1 0 15272 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1606256979
transform 1 0 16376 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16560 0 1 14544
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_23_177
timestamp 1606256979
transform 1 0 17388 0 1 14544
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1606256979
transform 1 0 20240 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 18768 0 1 14544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_23_189
timestamp 1606256979
transform 1 0 18492 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_198
timestamp 1606256979
transform 1 0 19320 0 1 14544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_206
timestamp 1606256979
transform 1 0 20056 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606256979
transform -1 0 21620 0 1 14544
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606256979
transform 1 0 20792 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_212
timestamp 1606256979
transform 1 0 20608 0 1 14544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1606256979
transform 1 0 20884 0 1 14544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_219
timestamp 1606256979
transform 1 0 21252 0 1 14544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606256979
transform 1 0 1104 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1606256979
transform 1 0 1380 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_15
timestamp 1606256979
transform 1 0 2484 0 -1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4876 0 -1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1606256979
transform 1 0 3036 0 -1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_24_30
timestamp 1606256979
transform 1 0 3864 0 -1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_38
timestamp 1606256979
transform 1 0 4600 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606256979
transform 1 0 6716 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_57
timestamp 1606256979
transform 1 0 6348 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_62
timestamp 1606256979
transform 1 0 6808 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_right_track_0.prog_clk
timestamp 1606256979
transform 1 0 7176 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_69
timestamp 1606256979
transform 1 0 7452 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_81
timestamp 1606256979
transform 1 0 8556 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1606256979
transform 1 0 9660 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606256979
transform 1 0 12328 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1606256979
transform 1 0 10764 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_117
timestamp 1606256979
transform 1 0 11868 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_121
timestamp 1606256979
transform 1 0 12236 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1606256979
transform 1 0 12420 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_135
timestamp 1606256979
transform 1 0 13524 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_147
timestamp 1606256979
transform 1 0 14628 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_159
timestamp 1606256979
transform 1 0 15732 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606256979
transform 1 0 17940 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_171
timestamp 1606256979
transform 1 0 16836 0 -1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_184
timestamp 1606256979
transform 1 0 18032 0 -1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 18860 0 -1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19596 0 -1 15632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_192
timestamp 1606256979
transform 1 0 18768 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_199
timestamp 1606256979
transform 1 0 19412 0 -1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_207
timestamp 1606256979
transform 1 0 20148 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1606256979
transform 1 0 20516 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606256979
transform -1 0 21620 0 -1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1606256979
transform 1 0 20884 0 -1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1606256979
transform 1 0 21252 0 -1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 1748 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606256979
transform 1 0 1104 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1606256979
transform 1 0 1380 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606256979
transform 1 0 3956 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_23
timestamp 1606256979
transform 1 0 3220 0 1 15632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_32
timestamp 1606256979
transform 1 0 4048 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 5612 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_44
timestamp 1606256979
transform 1 0 5152 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_48
timestamp 1606256979
transform 1 0 5520 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1606256979
transform 1 0 7268 0 1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_65
timestamp 1606256979
transform 1 0 7084 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_76
timestamp 1606256979
transform 1 0 8096 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _40_
timestamp 1606256979
transform 1 0 10120 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606256979
transform 1 0 9568 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_88
timestamp 1606256979
transform 1 0 9200 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_93
timestamp 1606256979
transform 1 0 9660 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_97
timestamp 1606256979
transform 1 0 10028 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_101
timestamp 1606256979
transform 1 0 10396 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 11500 0 1 15632
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1606256979
transform 1 0 14076 0 1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_25_129
timestamp 1606256979
transform 1 0 12972 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1606256979
transform 1 0 15272 0 1 15632
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606256979
transform 1 0 15180 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_150
timestamp 1606256979
transform 1 0 14904 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_163
timestamp 1606256979
transform 1 0 16100 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_175
timestamp 1606256979
transform 1 0 17204 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_187
timestamp 1606256979
transform 1 0 18308 0 1 15632
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1606256979
transform 1 0 20240 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1606256979
transform 1 0 19688 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_25_199
timestamp 1606256979
transform 1 0 19412 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_206
timestamp 1606256979
transform 1 0 20056 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606256979
transform -1 0 21620 0 1 15632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606256979
transform 1 0 20792 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_212
timestamp 1606256979
transform 1 0 20608 0 1 15632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1606256979
transform 1 0 20884 0 1 15632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_219
timestamp 1606256979
transform 1 0 21252 0 1 15632
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1606256979
transform 1 0 2944 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606256979
transform 1 0 1104 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606256979
transform 1 0 1104 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1606256979
transform 1 0 1380 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1606256979
transform 1 0 2484 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1606256979
transform 1 0 1380 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_15
timestamp 1606256979
transform 1 0 2484 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_19
timestamp 1606256979
transform 1 0 2852 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4048 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 3864 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606256979
transform 1 0 3956 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_27
timestamp 1606256979
transform 1 0 3588 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_36
timestamp 1606256979
transform 1 0 4416 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_29
timestamp 1606256979
transform 1 0 3772 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_41
timestamp 1606256979
transform 1 0 4876 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 6532 0 1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606256979
transform 1 0 6716 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_48
timestamp 1606256979
transform 1 0 5520 0 -1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_60
timestamp 1606256979
transform 1 0 6624 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_62
timestamp 1606256979
transform 1 0 6808 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_53
timestamp 1606256979
transform 1 0 5980 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1606256979
transform 1 0 7912 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 8648 0 -1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1606256979
transform 1 0 8556 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1606256979
transform 1 0 6900 0 -1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_72
timestamp 1606256979
transform 1 0 7728 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_77
timestamp 1606256979
transform 1 0 8188 0 -1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_81
timestamp 1606256979
transform 1 0 8556 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_75
timestamp 1606256979
transform 1 0 8004 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10304 0 -1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1606256979
transform 1 0 9752 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606256979
transform 1 0 9568 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_98
timestamp 1606256979
transform 1 0 10120 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_90
timestamp 1606256979
transform 1 0 9384 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_93
timestamp 1606256979
transform 1 0 9660 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_103
timestamp 1606256979
transform 1 0 10580 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1606256979
transform 1 0 12512 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1606256979
transform 1 0 11776 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606256979
transform 1 0 12328 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_116
timestamp 1606256979
transform 1 0 11776 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_123
timestamp 1606256979
transform 1 0 12420 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_115
timestamp 1606256979
transform 1 0 11684 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_125
timestamp 1606256979
transform 1 0 12604 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 12972 0 -1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1606256979
transform 1 0 12788 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_26_127
timestamp 1606256979
transform 1 0 12788 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_145
timestamp 1606256979
transform 1 0 14444 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_136
timestamp 1606256979
transform 1 0 13616 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1606256979
transform 1 0 14996 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 15548 0 -1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606256979
transform 1 0 15180 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_154
timestamp 1606256979
transform 1 0 15272 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_148
timestamp 1606256979
transform 1 0 14720 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_152
timestamp 1606256979
transform 1 0 15088 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_154
timestamp 1606256979
transform 1 0 15272 0 1 16720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_166
timestamp 1606256979
transform 1 0 16376 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1606256979
transform 1 0 18032 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 16468 0 1 16720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1606256979
transform 1 0 18124 0 1 16720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606256979
transform 1 0 17940 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_173
timestamp 1606256979
transform 1 0 17020 0 -1 16720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_181
timestamp 1606256979
transform 1 0 17756 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_187
timestamp 1606256979
transform 1 0 18308 0 -1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_183
timestamp 1606256979
transform 1 0 17940 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1606256979
transform 1 0 19964 0 -1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19228 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19964 0 1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 18768 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_191
timestamp 1606256979
transform 1 0 18676 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_198
timestamp 1606256979
transform 1 0 19320 0 -1 16720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_204
timestamp 1606256979
transform 1 0 19872 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_194
timestamp 1606256979
transform 1 0 18952 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_203
timestamp 1606256979
transform 1 0 19780 0 1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_211
timestamp 1606256979
transform 1 0 20516 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_209
timestamp 1606256979
transform 1 0 20332 0 -1 16720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1606256979
transform 1 0 20516 0 -1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_215
timestamp 1606256979
transform 1 0 20884 0 1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1606256979
transform 1 0 20884 0 -1 16720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606256979
transform 1 0 20792 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_219
timestamp 1606256979
transform 1 0 21252 0 1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1606256979
transform 1 0 21252 0 -1 16720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606256979
transform -1 0 21620 0 1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606256979
transform -1 0 21620 0 -1 16720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 1564 0 -1 17808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606256979
transform 1 0 1104 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1606256979
transform 1 0 1380 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1606256979
transform 1 0 3312 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 4876 0 -1 17808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_28_21
timestamp 1606256979
transform 1 0 3036 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_27
timestamp 1606256979
transform 1 0 3588 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_39
timestamp 1606256979
transform 1 0 4692 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606256979
transform 1 0 6716 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_57
timestamp 1606256979
transform 1 0 6348 0 -1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_62
timestamp 1606256979
transform 1 0 6808 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_74
timestamp 1606256979
transform 1 0 7912 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_86
timestamp 1606256979
transform 1 0 9016 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_98
timestamp 1606256979
transform 1 0 10120 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606256979
transform 1 0 12328 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_110
timestamp 1606256979
transform 1 0 11224 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_123
timestamp 1606256979
transform 1 0 12420 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_135
timestamp 1606256979
transform 1 0 13524 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_147
timestamp 1606256979
transform 1 0 14628 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_159
timestamp 1606256979
transform 1 0 15732 0 -1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1606256979
transform 1 0 16560 0 -1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606256979
transform 1 0 17940 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_167
timestamp 1606256979
transform 1 0 16468 0 -1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_177
timestamp 1606256979
transform 1 0 17388 0 -1 17808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_184
timestamp 1606256979
transform 1 0 18032 0 -1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1606256979
transform 1 0 20148 0 -1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19320 0 -1 17808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_196
timestamp 1606256979
transform 1 0 19136 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_204
timestamp 1606256979
transform 1 0 19872 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1606256979
transform 1 0 20700 0 -1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606256979
transform -1 0 21620 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_211
timestamp 1606256979
transform 1 0 20516 0 -1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_217
timestamp 1606256979
transform 1 0 21068 0 -1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606256979
transform 1 0 1104 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1606256979
transform 1 0 1380 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1606256979
transform 1 0 2484 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606256979
transform 1 0 3956 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_27
timestamp 1606256979
transform 1 0 3588 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_32
timestamp 1606256979
transform 1 0 4048 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 5152 0 1 17808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_50
timestamp 1606256979
transform 1 0 5704 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_62
timestamp 1606256979
transform 1 0 6808 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1606256979
transform 1 0 7636 0 1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_29_70
timestamp 1606256979
transform 1 0 7544 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_80
timestamp 1606256979
transform 1 0 8464 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1606256979
transform 1 0 10396 0 1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606256979
transform 1 0 9568 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_93
timestamp 1606256979
transform 1 0 9660 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_110
timestamp 1606256979
transform 1 0 11224 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_122
timestamp 1606256979
transform 1 0 12328 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1606256979
transform 1 0 13340 0 1 17808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_29_130
timestamp 1606256979
transform 1 0 13064 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_142
timestamp 1606256979
transform 1 0 14168 0 1 17808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606256979
transform 1 0 15180 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_150
timestamp 1606256979
transform 1 0 14904 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_154
timestamp 1606256979
transform 1 0 15272 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1606256979
transform 1 0 16376 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1606256979
transform 1 0 16560 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1606256979
transform 1 0 16836 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_183
timestamp 1606256979
transform 1 0 17940 0 1 17808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1606256979
transform 1 0 19596 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1606256979
transform 1 0 20240 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_195
timestamp 1606256979
transform 1 0 19044 0 1 17808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_29_205
timestamp 1606256979
transform 1 0 19964 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606256979
transform -1 0 21620 0 1 17808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606256979
transform 1 0 20792 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_212
timestamp 1606256979
transform 1 0 20608 0 1 17808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_215
timestamp 1606256979
transform 1 0 20884 0 1 17808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_219
timestamp 1606256979
transform 1 0 21252 0 1 17808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 2392 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606256979
transform 1 0 1104 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1606256979
transform 1 0 1380 0 -1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_11
timestamp 1606256979
transform 1 0 2116 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1606256979
transform 1 0 4692 0 -1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_30_30
timestamp 1606256979
transform 1 0 3864 0 -1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_38
timestamp 1606256979
transform 1 0 4600 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1606256979
transform 1 0 5704 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606256979
transform 1 0 6716 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_48
timestamp 1606256979
transform 1 0 5520 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_53
timestamp 1606256979
transform 1 0 5980 0 -1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_62
timestamp 1606256979
transform 1 0 6808 0 -1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1606256979
transform 1 0 8372 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1606256979
transform 1 0 7360 0 -1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_77
timestamp 1606256979
transform 1 0 8188 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_82
timestamp 1606256979
transform 1 0 8648 0 -1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1606256979
transform 1 0 10212 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 10672 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1606256979
transform 1 0 9200 0 -1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_97
timestamp 1606256979
transform 1 0 10028 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_102
timestamp 1606256979
transform 1 0 10488 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1606256979
transform 1 0 12420 0 -1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606256979
transform 1 0 12328 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_120
timestamp 1606256979
transform 1 0 12144 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 13432 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_132
timestamp 1606256979
transform 1 0 13248 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 15088 0 -1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_150
timestamp 1606256979
transform 1 0 14904 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1606256979
transform 1 0 16744 0 -1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 18032 0 -1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606256979
transform 1 0 17940 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_168
timestamp 1606256979
transform 1 0 16560 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_179
timestamp 1606256979
transform 1 0 17572 0 -1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19504 0 -1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_190
timestamp 1606256979
transform 1 0 18584 0 -1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_198
timestamp 1606256979
transform 1 0 19320 0 -1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_206
timestamp 1606256979
transform 1 0 20056 0 -1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1606256979
transform 1 0 20516 0 -1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606256979
transform -1 0 21620 0 -1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_210
timestamp 1606256979
transform 1 0 20424 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1606256979
transform 1 0 20884 0 -1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1606256979
transform 1 0 21252 0 -1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606256979
transform 1 0 1104 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1606256979
transform 1 0 1380 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1606256979
transform 1 0 2484 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 4048 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606256979
transform 1 0 3956 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_27
timestamp 1606256979
transform 1 0 3588 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 6072 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_31_48
timestamp 1606256979
transform 1 0 5520 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606256979
transform 1 0 7728 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_70
timestamp 1606256979
transform 1 0 7544 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 9660 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606256979
transform 1 0 9568 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_88
timestamp 1606256979
transform 1 0 9200 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606256979
transform 1 0 12328 0 1 18896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_31_109
timestamp 1606256979
transform 1 0 11132 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_121
timestamp 1606256979
transform 1 0 12236 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1606256979
transform 1 0 13984 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_138
timestamp 1606256979
transform 1 0 13800 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_143
timestamp 1606256979
transform 1 0 14260 0 1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1606256979
transform 1 0 15272 0 1 18896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606256979
transform 1 0 15180 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_151
timestamp 1606256979
transform 1 0 14996 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_163
timestamp 1606256979
transform 1 0 16100 0 1 18896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 16836 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606256979
transform 1 0 17940 0 1 18896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_177
timestamp 1606256979
transform 1 0 17388 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1606256979
transform 1 0 20240 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19504 0 1 18896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_195
timestamp 1606256979
transform 1 0 19044 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_199
timestamp 1606256979
transform 1 0 19412 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_206
timestamp 1606256979
transform 1 0 20056 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606256979
transform -1 0 21620 0 1 18896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606256979
transform 1 0 20792 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_212
timestamp 1606256979
transform 1 0 20608 0 1 18896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1606256979
transform 1 0 20884 0 1 18896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_219
timestamp 1606256979
transform 1 0 21252 0 1 18896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606256979
transform 1 0 1104 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1606256979
transform 1 0 1380 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1606256979
transform 1 0 2484 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1606256979
transform 1 0 4600 0 -1 19984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606256979
transform 1 0 3956 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1606256979
transform 1 0 3588 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_32
timestamp 1606256979
transform 1 0 4048 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606256979
transform 1 0 6808 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_47
timestamp 1606256979
transform 1 0 5428 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_59
timestamp 1606256979
transform 1 0 6532 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1606256979
transform 1 0 6900 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_75
timestamp 1606256979
transform 1 0 8004 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606256979
transform 1 0 9660 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_87
timestamp 1606256979
transform 1 0 9108 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1606256979
transform 1 0 9752 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606256979
transform 1 0 12512 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_106
timestamp 1606256979
transform 1 0 10856 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_118
timestamp 1606256979
transform 1 0 11960 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_125
timestamp 1606256979
transform 1 0 12604 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_137
timestamp 1606256979
transform 1 0 13708 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606256979
transform 1 0 15364 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_149
timestamp 1606256979
transform 1 0 14812 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1606256979
transform 1 0 15456 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1606256979
transform 1 0 17664 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606256979
transform 1 0 18216 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1606256979
transform 1 0 16560 0 -1 19984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_184
timestamp 1606256979
transform 1 0 18032 0 -1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_187
timestamp 1606256979
transform 1 0 18308 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1606256979
transform 1 0 18400 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1606256979
transform 1 0 19504 0 -1 19984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_192
timestamp 1606256979
transform 1 0 18768 0 -1 19984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_206
timestamp 1606256979
transform 1 0 20056 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1606256979
transform 1 0 20516 0 -1 19984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606256979
transform -1 0 21620 0 -1 19984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1606256979
transform 1 0 21068 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_210
timestamp 1606256979
transform 1 0 20424 0 -1 19984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1606256979
transform 1 0 20884 0 -1 19984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1606256979
transform 1 0 21160 0 -1 19984
box -38 -48 222 592
<< labels >>
rlabel metal3 s 0 5576 480 5696 6 ccff_head
port 0 nsew default input
rlabel metal3 s 0 17000 480 17120 6 ccff_tail
port 1 nsew default tristate
rlabel metal3 s 22320 4080 22800 4200 6 chanx_right_in[0]
port 2 nsew default input
rlabel metal3 s 22320 8568 22800 8688 6 chanx_right_in[10]
port 3 nsew default input
rlabel metal3 s 22320 9112 22800 9232 6 chanx_right_in[11]
port 4 nsew default input
rlabel metal3 s 22320 9520 22800 9640 6 chanx_right_in[12]
port 5 nsew default input
rlabel metal3 s 22320 9928 22800 10048 6 chanx_right_in[13]
port 6 nsew default input
rlabel metal3 s 22320 10472 22800 10592 6 chanx_right_in[14]
port 7 nsew default input
rlabel metal3 s 22320 10880 22800 11000 6 chanx_right_in[15]
port 8 nsew default input
rlabel metal3 s 22320 11424 22800 11544 6 chanx_right_in[16]
port 9 nsew default input
rlabel metal3 s 22320 11832 22800 11952 6 chanx_right_in[17]
port 10 nsew default input
rlabel metal3 s 22320 12240 22800 12360 6 chanx_right_in[18]
port 11 nsew default input
rlabel metal3 s 22320 12784 22800 12904 6 chanx_right_in[19]
port 12 nsew default input
rlabel metal3 s 22320 4488 22800 4608 6 chanx_right_in[1]
port 13 nsew default input
rlabel metal3 s 22320 4896 22800 5016 6 chanx_right_in[2]
port 14 nsew default input
rlabel metal3 s 22320 5440 22800 5560 6 chanx_right_in[3]
port 15 nsew default input
rlabel metal3 s 22320 5848 22800 5968 6 chanx_right_in[4]
port 16 nsew default input
rlabel metal3 s 22320 6392 22800 6512 6 chanx_right_in[5]
port 17 nsew default input
rlabel metal3 s 22320 6800 22800 6920 6 chanx_right_in[6]
port 18 nsew default input
rlabel metal3 s 22320 7208 22800 7328 6 chanx_right_in[7]
port 19 nsew default input
rlabel metal3 s 22320 7752 22800 7872 6 chanx_right_in[8]
port 20 nsew default input
rlabel metal3 s 22320 8160 22800 8280 6 chanx_right_in[9]
port 21 nsew default input
rlabel metal3 s 22320 13192 22800 13312 6 chanx_right_out[0]
port 22 nsew default tristate
rlabel metal3 s 22320 17816 22800 17936 6 chanx_right_out[10]
port 23 nsew default tristate
rlabel metal3 s 22320 18224 22800 18344 6 chanx_right_out[11]
port 24 nsew default tristate
rlabel metal3 s 22320 18632 22800 18752 6 chanx_right_out[12]
port 25 nsew default tristate
rlabel metal3 s 22320 19176 22800 19296 6 chanx_right_out[13]
port 26 nsew default tristate
rlabel metal3 s 22320 19584 22800 19704 6 chanx_right_out[14]
port 27 nsew default tristate
rlabel metal3 s 22320 19992 22800 20112 6 chanx_right_out[15]
port 28 nsew default tristate
rlabel metal3 s 22320 20536 22800 20656 6 chanx_right_out[16]
port 29 nsew default tristate
rlabel metal3 s 22320 20944 22800 21064 6 chanx_right_out[17]
port 30 nsew default tristate
rlabel metal3 s 22320 21352 22800 21472 6 chanx_right_out[18]
port 31 nsew default tristate
rlabel metal3 s 22320 21896 22800 22016 6 chanx_right_out[19]
port 32 nsew default tristate
rlabel metal3 s 22320 13600 22800 13720 6 chanx_right_out[1]
port 33 nsew default tristate
rlabel metal3 s 22320 14144 22800 14264 6 chanx_right_out[2]
port 34 nsew default tristate
rlabel metal3 s 22320 14552 22800 14672 6 chanx_right_out[3]
port 35 nsew default tristate
rlabel metal3 s 22320 14960 22800 15080 6 chanx_right_out[4]
port 36 nsew default tristate
rlabel metal3 s 22320 15504 22800 15624 6 chanx_right_out[5]
port 37 nsew default tristate
rlabel metal3 s 22320 15912 22800 16032 6 chanx_right_out[6]
port 38 nsew default tristate
rlabel metal3 s 22320 16320 22800 16440 6 chanx_right_out[7]
port 39 nsew default tristate
rlabel metal3 s 22320 16864 22800 16984 6 chanx_right_out[8]
port 40 nsew default tristate
rlabel metal3 s 22320 17272 22800 17392 6 chanx_right_out[9]
port 41 nsew default tristate
rlabel metal2 s 846 22176 902 22656 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 6366 22176 6422 22656 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 6918 22176 6974 22656 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 7470 22176 7526 22656 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 8022 22176 8078 22656 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 8574 22176 8630 22656 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 9126 22176 9182 22656 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 9678 22176 9734 22656 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 10230 22176 10286 22656 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 10782 22176 10838 22656 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 11334 22176 11390 22656 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 1398 22176 1454 22656 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 1950 22176 2006 22656 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 2502 22176 2558 22656 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 3054 22176 3110 22656 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 3606 22176 3662 22656 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 4158 22176 4214 22656 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 4710 22176 4766 22656 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 5262 22176 5318 22656 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 5814 22176 5870 22656 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 11978 22176 12034 22656 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 17498 22176 17554 22656 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 18050 22176 18106 22656 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 18602 22176 18658 22656 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 19154 22176 19210 22656 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 19706 22176 19762 22656 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 20258 22176 20314 22656 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 20810 22176 20866 22656 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 21362 22176 21418 22656 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 21914 22176 21970 22656 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 22466 22176 22522 22656 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 12530 22176 12586 22656 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 13082 22176 13138 22656 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 13634 22176 13690 22656 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 14186 22176 14242 22656 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 14738 22176 14794 22656 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 15290 22176 15346 22656 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 15842 22176 15898 22656 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 16394 22176 16450 22656 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 16946 22176 17002 22656 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 22320 22304 22800 22424 6 prog_clk_0_E_in
port 82 nsew default input
rlabel metal3 s 22320 2176 22800 2296 6 right_bottom_grid_pin_11_
port 83 nsew default input
rlabel metal3 s 22320 2720 22800 2840 6 right_bottom_grid_pin_13_
port 84 nsew default input
rlabel metal3 s 22320 3128 22800 3248 6 right_bottom_grid_pin_15_
port 85 nsew default input
rlabel metal3 s 22320 3536 22800 3656 6 right_bottom_grid_pin_17_
port 86 nsew default input
rlabel metal3 s 22320 0 22800 120 6 right_bottom_grid_pin_1_
port 87 nsew default input
rlabel metal3 s 22320 408 22800 528 6 right_bottom_grid_pin_3_
port 88 nsew default input
rlabel metal3 s 22320 816 22800 936 6 right_bottom_grid_pin_5_
port 89 nsew default input
rlabel metal3 s 22320 1360 22800 1480 6 right_bottom_grid_pin_7_
port 90 nsew default input
rlabel metal3 s 22320 1768 22800 1888 6 right_bottom_grid_pin_9_
port 91 nsew default input
rlabel metal2 s 294 22176 350 22656 6 top_left_grid_pin_1_
port 92 nsew default input
rlabel metal4 s 4376 1984 4696 20032 6 VPWR
port 93 nsew default input
rlabel metal4 s 7808 1984 8128 20032 6 VGND
port 94 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22656
<< end >>
