VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_8__0_
  CLASS BLOCK ;
  FOREIGN sb_8__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 114.000 BY 114.000 ;
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 111.600 57.160 114.000 57.760 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 2.400 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 2.400 21.720 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 2.400 45.520 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 2.400 47.560 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 2.400 50.280 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 2.400 52.320 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 2.400 54.360 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 2.400 57.080 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 2.400 59.120 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 2.400 61.840 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 2.400 63.880 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 2.400 66.600 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 2.400 24.440 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 2.400 26.480 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 2.400 29.200 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 2.400 31.240 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.400 33.960 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 2.400 36.000 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 2.400 38.040 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 2.400 40.760 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 2.400 42.800 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 2.400 68.640 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 2.400 91.760 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 2.400 94.480 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 2.400 96.520 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 2.400 99.240 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 2.400 101.280 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 2.400 103.320 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 2.400 106.040 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 2.400 108.080 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 2.400 110.800 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 2.400 112.840 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 2.400 70.680 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 2.400 73.400 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 2.400 75.440 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 2.400 78.160 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 2.400 80.200 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 2.400 82.920 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 2.400 84.960 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 2.400 87.000 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 2.400 89.720 ;
    END
  END chanx_left_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.410 111.600 19.690 114.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.870 111.600 43.150 114.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.170 111.600 45.450 114.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.470 111.600 47.750 114.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.770 111.600 50.050 114.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.070 111.600 52.350 114.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.370 111.600 54.650 114.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.670 111.600 56.950 114.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 111.600 59.250 114.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.270 111.600 61.550 114.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.570 111.600 63.850 114.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.710 111.600 21.990 114.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 111.600 24.290 114.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.310 111.600 26.590 114.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 111.600 28.890 114.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.910 111.600 31.190 114.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.210 111.600 33.490 114.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.510 111.600 35.790 114.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.810 111.600 38.090 114.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.570 111.600 40.850 114.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.870 111.600 66.150 114.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.330 111.600 89.610 114.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.630 111.600 91.910 114.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.930 111.600 94.210 114.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 96.230 111.600 96.510 114.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.530 111.600 98.810 114.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.830 111.600 101.110 114.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.130 111.600 103.410 114.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.430 111.600 105.710 114.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.730 111.600 108.010 114.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.030 111.600 110.310 114.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.170 111.600 68.450 114.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.470 111.600 70.750 114.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.770 111.600 73.050 114.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.070 111.600 75.350 114.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.830 111.600 78.110 114.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.130 111.600 80.410 114.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.430 111.600 82.710 114.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 84.730 111.600 85.010 114.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.030 111.600 87.310 114.000 ;
    END
  END chany_top_out[9]
  PIN left_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 2.400 12.880 ;
    END
  END left_bottom_grid_pin_11_
  PIN left_bottom_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 2.400 14.920 ;
    END
  END left_bottom_grid_pin_13_
  PIN left_bottom_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 2.400 17.640 ;
    END
  END left_bottom_grid_pin_15_
  PIN left_bottom_grid_pin_17_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 2.400 19.680 ;
    END
  END left_bottom_grid_pin_17_
  PIN left_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 2.400 1.320 ;
    END
  END left_bottom_grid_pin_1_
  PIN left_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 2.400 3.360 ;
    END
  END left_bottom_grid_pin_3_
  PIN left_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 2.400 5.400 ;
    END
  END left_bottom_grid_pin_5_
  PIN left_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 2.400 8.120 ;
    END
  END left_bottom_grid_pin_7_
  PIN left_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 2.400 10.160 ;
    END
  END left_bottom_grid_pin_9_
  PIN prog_clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 2.400 ;
    END
  END prog_clk
  PIN top_left_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.010 111.600 1.290 114.000 ;
    END
  END top_left_grid_pin_42_
  PIN top_left_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.310 111.600 3.590 114.000 ;
    END
  END top_left_grid_pin_43_
  PIN top_left_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.610 111.600 5.890 114.000 ;
    END
  END top_left_grid_pin_44_
  PIN top_left_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.910 111.600 8.190 114.000 ;
    END
  END top_left_grid_pin_45_
  PIN top_left_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 111.600 10.490 114.000 ;
    END
  END top_left_grid_pin_46_
  PIN top_left_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.510 111.600 12.790 114.000 ;
    END
  END top_left_grid_pin_47_
  PIN top_left_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.810 111.600 15.090 114.000 ;
    END
  END top_left_grid_pin_48_
  PIN top_left_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 111.600 17.390 114.000 ;
    END
  END top_left_grid_pin_49_
  PIN top_right_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.330 111.600 112.610 114.000 ;
    END
  END top_right_grid_pin_1_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.880 10.640 23.480 100.880 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.040 10.640 40.640 100.880 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 108.100 100.725 ;
      LAYER met1 ;
        RECT 0.990 2.760 112.630 100.880 ;
      LAYER met2 ;
        RECT 1.570 111.320 3.030 112.725 ;
        RECT 3.870 111.320 5.330 112.725 ;
        RECT 6.170 111.320 7.630 112.725 ;
        RECT 8.470 111.320 9.930 112.725 ;
        RECT 10.770 111.320 12.230 112.725 ;
        RECT 13.070 111.320 14.530 112.725 ;
        RECT 15.370 111.320 16.830 112.725 ;
        RECT 17.670 111.320 19.130 112.725 ;
        RECT 19.970 111.320 21.430 112.725 ;
        RECT 22.270 111.320 23.730 112.725 ;
        RECT 24.570 111.320 26.030 112.725 ;
        RECT 26.870 111.320 28.330 112.725 ;
        RECT 29.170 111.320 30.630 112.725 ;
        RECT 31.470 111.320 32.930 112.725 ;
        RECT 33.770 111.320 35.230 112.725 ;
        RECT 36.070 111.320 37.530 112.725 ;
        RECT 38.370 111.320 40.290 112.725 ;
        RECT 41.130 111.320 42.590 112.725 ;
        RECT 43.430 111.320 44.890 112.725 ;
        RECT 45.730 111.320 47.190 112.725 ;
        RECT 48.030 111.320 49.490 112.725 ;
        RECT 50.330 111.320 51.790 112.725 ;
        RECT 52.630 111.320 54.090 112.725 ;
        RECT 54.930 111.320 56.390 112.725 ;
        RECT 57.230 111.320 58.690 112.725 ;
        RECT 59.530 111.320 60.990 112.725 ;
        RECT 61.830 111.320 63.290 112.725 ;
        RECT 64.130 111.320 65.590 112.725 ;
        RECT 66.430 111.320 67.890 112.725 ;
        RECT 68.730 111.320 70.190 112.725 ;
        RECT 71.030 111.320 72.490 112.725 ;
        RECT 73.330 111.320 74.790 112.725 ;
        RECT 75.630 111.320 77.550 112.725 ;
        RECT 78.390 111.320 79.850 112.725 ;
        RECT 80.690 111.320 82.150 112.725 ;
        RECT 82.990 111.320 84.450 112.725 ;
        RECT 85.290 111.320 86.750 112.725 ;
        RECT 87.590 111.320 89.050 112.725 ;
        RECT 89.890 111.320 91.350 112.725 ;
        RECT 92.190 111.320 93.650 112.725 ;
        RECT 94.490 111.320 95.950 112.725 ;
        RECT 96.790 111.320 98.250 112.725 ;
        RECT 99.090 111.320 100.550 112.725 ;
        RECT 101.390 111.320 102.850 112.725 ;
        RECT 103.690 111.320 105.150 112.725 ;
        RECT 105.990 111.320 107.450 112.725 ;
        RECT 108.290 111.320 109.750 112.725 ;
        RECT 110.590 111.320 112.050 112.725 ;
        RECT 1.020 2.680 112.600 111.320 ;
        RECT 1.020 0.835 28.330 2.680 ;
        RECT 29.170 0.835 85.370 2.680 ;
        RECT 86.210 0.835 112.600 2.680 ;
      LAYER met3 ;
        RECT 2.800 111.840 111.600 112.705 ;
        RECT 2.400 111.200 111.600 111.840 ;
        RECT 2.800 109.800 111.600 111.200 ;
        RECT 2.400 108.480 111.600 109.800 ;
        RECT 2.800 107.080 111.600 108.480 ;
        RECT 2.400 106.440 111.600 107.080 ;
        RECT 2.800 105.040 111.600 106.440 ;
        RECT 2.400 103.720 111.600 105.040 ;
        RECT 2.800 102.320 111.600 103.720 ;
        RECT 2.400 101.680 111.600 102.320 ;
        RECT 2.800 100.280 111.600 101.680 ;
        RECT 2.400 99.640 111.600 100.280 ;
        RECT 2.800 98.240 111.600 99.640 ;
        RECT 2.400 96.920 111.600 98.240 ;
        RECT 2.800 95.520 111.600 96.920 ;
        RECT 2.400 94.880 111.600 95.520 ;
        RECT 2.800 93.480 111.600 94.880 ;
        RECT 2.400 92.160 111.600 93.480 ;
        RECT 2.800 90.760 111.600 92.160 ;
        RECT 2.400 90.120 111.600 90.760 ;
        RECT 2.800 88.720 111.600 90.120 ;
        RECT 2.400 87.400 111.600 88.720 ;
        RECT 2.800 86.000 111.600 87.400 ;
        RECT 2.400 85.360 111.600 86.000 ;
        RECT 2.800 83.960 111.600 85.360 ;
        RECT 2.400 83.320 111.600 83.960 ;
        RECT 2.800 81.920 111.600 83.320 ;
        RECT 2.400 80.600 111.600 81.920 ;
        RECT 2.800 79.200 111.600 80.600 ;
        RECT 2.400 78.560 111.600 79.200 ;
        RECT 2.800 77.160 111.600 78.560 ;
        RECT 2.400 75.840 111.600 77.160 ;
        RECT 2.800 74.440 111.600 75.840 ;
        RECT 2.400 73.800 111.600 74.440 ;
        RECT 2.800 72.400 111.600 73.800 ;
        RECT 2.400 71.080 111.600 72.400 ;
        RECT 2.800 69.680 111.600 71.080 ;
        RECT 2.400 69.040 111.600 69.680 ;
        RECT 2.800 67.640 111.600 69.040 ;
        RECT 2.400 67.000 111.600 67.640 ;
        RECT 2.800 65.600 111.600 67.000 ;
        RECT 2.400 64.280 111.600 65.600 ;
        RECT 2.800 62.880 111.600 64.280 ;
        RECT 2.400 62.240 111.600 62.880 ;
        RECT 2.800 60.840 111.600 62.240 ;
        RECT 2.400 59.520 111.600 60.840 ;
        RECT 2.800 58.160 111.600 59.520 ;
        RECT 2.800 58.120 111.200 58.160 ;
        RECT 2.400 57.480 111.200 58.120 ;
        RECT 2.800 56.760 111.200 57.480 ;
        RECT 2.800 56.080 111.600 56.760 ;
        RECT 2.400 54.760 111.600 56.080 ;
        RECT 2.800 53.360 111.600 54.760 ;
        RECT 2.400 52.720 111.600 53.360 ;
        RECT 2.800 51.320 111.600 52.720 ;
        RECT 2.400 50.680 111.600 51.320 ;
        RECT 2.800 49.280 111.600 50.680 ;
        RECT 2.400 47.960 111.600 49.280 ;
        RECT 2.800 46.560 111.600 47.960 ;
        RECT 2.400 45.920 111.600 46.560 ;
        RECT 2.800 44.520 111.600 45.920 ;
        RECT 2.400 43.200 111.600 44.520 ;
        RECT 2.800 41.800 111.600 43.200 ;
        RECT 2.400 41.160 111.600 41.800 ;
        RECT 2.800 39.760 111.600 41.160 ;
        RECT 2.400 38.440 111.600 39.760 ;
        RECT 2.800 37.040 111.600 38.440 ;
        RECT 2.400 36.400 111.600 37.040 ;
        RECT 2.800 35.000 111.600 36.400 ;
        RECT 2.400 34.360 111.600 35.000 ;
        RECT 2.800 32.960 111.600 34.360 ;
        RECT 2.400 31.640 111.600 32.960 ;
        RECT 2.800 30.240 111.600 31.640 ;
        RECT 2.400 29.600 111.600 30.240 ;
        RECT 2.800 28.200 111.600 29.600 ;
        RECT 2.400 26.880 111.600 28.200 ;
        RECT 2.800 25.480 111.600 26.880 ;
        RECT 2.400 24.840 111.600 25.480 ;
        RECT 2.800 23.440 111.600 24.840 ;
        RECT 2.400 22.120 111.600 23.440 ;
        RECT 2.800 20.720 111.600 22.120 ;
        RECT 2.400 20.080 111.600 20.720 ;
        RECT 2.800 18.680 111.600 20.080 ;
        RECT 2.400 18.040 111.600 18.680 ;
        RECT 2.800 16.640 111.600 18.040 ;
        RECT 2.400 15.320 111.600 16.640 ;
        RECT 2.800 13.920 111.600 15.320 ;
        RECT 2.400 13.280 111.600 13.920 ;
        RECT 2.800 11.880 111.600 13.280 ;
        RECT 2.400 10.560 111.600 11.880 ;
        RECT 2.800 9.160 111.600 10.560 ;
        RECT 2.400 8.520 111.600 9.160 ;
        RECT 2.800 7.120 111.600 8.520 ;
        RECT 2.400 5.800 111.600 7.120 ;
        RECT 2.800 4.400 111.600 5.800 ;
        RECT 2.400 3.760 111.600 4.400 ;
        RECT 2.800 2.360 111.600 3.760 ;
        RECT 2.400 1.720 111.600 2.360 ;
        RECT 2.800 0.855 111.600 1.720 ;
      LAYER met4 ;
        RECT 56.200 10.640 92.120 100.880 ;
  END
END sb_8__0_
END LIBRARY

