magic
tech EFS8A
magscale 1 2
timestamp 1604337537
<< locali >>
rect 1777 3927 1811 4097
rect 10057 3995 10091 4233
rect 19993 3451 20027 3689
rect 3249 2499 3283 2601
<< viali >>
rect 1409 14365 1443 14399
rect 2237 14297 2271 14331
rect 1961 14229 1995 14263
rect 2053 14025 2087 14059
rect 2789 13889 2823 13923
rect 1409 13821 1443 13855
rect 2329 13821 2363 13855
rect 3065 13753 3099 13787
rect 1593 13685 1627 13719
rect 7849 13481 7883 13515
rect 1409 13345 1443 13379
rect 2513 13345 2547 13379
rect 3157 13277 3191 13311
rect 2053 13209 2087 13243
rect 3801 13209 3835 13243
rect 1593 13141 1627 13175
rect 2329 13141 2363 13175
rect 2697 13141 2731 13175
rect 3433 13141 3467 13175
rect 4353 13141 4387 13175
rect 2605 12937 2639 12971
rect 3709 12937 3743 12971
rect 1685 12869 1719 12903
rect 3985 12869 4019 12903
rect 7941 12869 7975 12903
rect 2145 12801 2179 12835
rect 2237 12801 2271 12835
rect 3433 12801 3467 12835
rect 4445 12801 4479 12835
rect 7389 12733 7423 12767
rect 8493 12733 8527 12767
rect 2145 12665 2179 12699
rect 4445 12665 4479 12699
rect 4537 12665 4571 12699
rect 8217 12665 8251 12699
rect 3065 12597 3099 12631
rect 4905 12597 4939 12631
rect 6837 12597 6871 12631
rect 7757 12597 7791 12631
rect 8401 12597 8435 12631
rect 9413 12597 9447 12631
rect 2053 12393 2087 12427
rect 2513 12393 2547 12427
rect 3249 12393 3283 12427
rect 5273 12325 5307 12359
rect 5457 12325 5491 12359
rect 5917 12325 5951 12359
rect 10048 12325 10082 12359
rect 1869 12257 1903 12291
rect 6725 12257 6759 12291
rect 2145 12189 2179 12223
rect 4353 12189 4387 12223
rect 5549 12189 5583 12223
rect 6469 12189 6503 12223
rect 9781 12189 9815 12223
rect 1593 12121 1627 12155
rect 2973 12053 3007 12087
rect 3709 12053 3743 12087
rect 4629 12053 4663 12087
rect 4997 12053 5031 12087
rect 7849 12053 7883 12087
rect 11161 12053 11195 12087
rect 1501 11849 1535 11883
rect 5549 11849 5583 11883
rect 8953 11849 8987 11883
rect 1961 11713 1995 11747
rect 5733 11713 5767 11747
rect 3249 11645 3283 11679
rect 3505 11645 3539 11679
rect 7573 11645 7607 11679
rect 2053 11577 2087 11611
rect 7389 11577 7423 11611
rect 7818 11577 7852 11611
rect 1961 11509 1995 11543
rect 2421 11509 2455 11543
rect 3065 11509 3099 11543
rect 4629 11509 4663 11543
rect 5273 11509 5307 11543
rect 6561 11509 6595 11543
rect 7021 11509 7055 11543
rect 9781 11509 9815 11543
rect 10057 11509 10091 11543
rect 10517 11509 10551 11543
rect 11161 11509 11195 11543
rect 12449 11509 12483 11543
rect 2881 11305 2915 11339
rect 4261 11305 4295 11339
rect 4997 11305 5031 11339
rect 6745 11305 6779 11339
rect 8585 11305 8619 11339
rect 9413 11305 9447 11339
rect 1768 11237 1802 11271
rect 5610 11237 5644 11271
rect 11152 11237 11186 11271
rect 4077 11169 4111 11203
rect 8401 11169 8435 11203
rect 9689 11169 9723 11203
rect 16221 11169 16255 11203
rect 1501 11101 1535 11135
rect 5365 11101 5399 11135
rect 8677 11101 8711 11135
rect 9045 11101 9079 11135
rect 10885 11101 10919 11135
rect 13369 11101 13403 11135
rect 16497 11101 16531 11135
rect 3893 11033 3927 11067
rect 8125 11033 8159 11067
rect 10149 11033 10183 11067
rect 3525 10965 3559 10999
rect 7573 10965 7607 10999
rect 12265 10965 12299 10999
rect 12909 10965 12943 10999
rect 5641 10761 5675 10795
rect 6653 10761 6687 10795
rect 8125 10761 8159 10795
rect 10057 10761 10091 10795
rect 6929 10693 6963 10727
rect 12541 10693 12575 10727
rect 16221 10693 16255 10727
rect 7297 10625 7331 10659
rect 1777 10557 1811 10591
rect 4261 10557 4295 10591
rect 8677 10557 8711 10591
rect 8944 10557 8978 10591
rect 11897 10557 11931 10591
rect 13093 10557 13127 10591
rect 16681 10557 16715 10591
rect 17417 10557 17451 10591
rect 2044 10489 2078 10523
rect 3801 10489 3835 10523
rect 4528 10489 4562 10523
rect 7481 10489 7515 10523
rect 10885 10489 10919 10523
rect 11253 10489 11287 10523
rect 12173 10489 12207 10523
rect 12817 10489 12851 10523
rect 16957 10489 16991 10523
rect 1685 10421 1719 10455
rect 3157 10421 3191 10455
rect 4169 10421 4203 10455
rect 6285 10421 6319 10455
rect 7389 10421 7423 10455
rect 8493 10421 8527 10455
rect 13001 10421 13035 10455
rect 2789 10217 2823 10251
rect 3065 10217 3099 10251
rect 3801 10217 3835 10251
rect 5457 10217 5491 10251
rect 7021 10217 7055 10251
rect 8033 10217 8067 10251
rect 8585 10217 8619 10251
rect 8953 10217 8987 10251
rect 9505 10217 9539 10251
rect 10977 10217 11011 10251
rect 2237 10149 2271 10183
rect 4905 10149 4939 10183
rect 6285 10149 6319 10183
rect 6469 10149 6503 10183
rect 10149 10149 10183 10183
rect 10333 10149 10367 10183
rect 10425 10149 10459 10183
rect 12072 10149 12106 10183
rect 4721 10081 4755 10115
rect 5825 10081 5859 10115
rect 6561 10081 6595 10115
rect 7389 10081 7423 10115
rect 8125 10081 8159 10115
rect 2145 10013 2179 10047
rect 2329 10013 2363 10047
rect 4997 10013 5031 10047
rect 8033 10013 8067 10047
rect 11805 10013 11839 10047
rect 15301 10013 15335 10047
rect 1777 9945 1811 9979
rect 4445 9945 4479 9979
rect 7573 9945 7607 9979
rect 9873 9945 9907 9979
rect 3525 9877 3559 9911
rect 6009 9877 6043 9911
rect 11253 9877 11287 9911
rect 13185 9877 13219 9911
rect 13737 9877 13771 9911
rect 5457 9673 5491 9707
rect 6285 9673 6319 9707
rect 7849 9673 7883 9707
rect 12173 9673 12207 9707
rect 2605 9605 2639 9639
rect 3893 9605 3927 9639
rect 4445 9605 4479 9639
rect 8125 9605 8159 9639
rect 10885 9605 10919 9639
rect 4997 9537 5031 9571
rect 5917 9537 5951 9571
rect 8309 9537 8343 9571
rect 10241 9537 10275 9571
rect 1409 9469 1443 9503
rect 2881 9469 2915 9503
rect 4721 9469 4755 9503
rect 6837 9469 6871 9503
rect 7481 9469 7515 9503
rect 8565 9469 8599 9503
rect 11897 9469 11931 9503
rect 12725 9469 12759 9503
rect 12992 9469 13026 9503
rect 18061 9469 18095 9503
rect 18797 9469 18831 9503
rect 3157 9401 3191 9435
rect 4905 9401 4939 9435
rect 10701 9401 10735 9435
rect 11161 9401 11195 9435
rect 11437 9401 11471 9435
rect 18337 9401 18371 9435
rect 1593 9333 1627 9367
rect 1961 9333 1995 9367
rect 2421 9333 2455 9367
rect 3065 9333 3099 9367
rect 4169 9333 4203 9367
rect 7021 9333 7055 9367
rect 9689 9333 9723 9367
rect 11345 9333 11379 9367
rect 14105 9333 14139 9367
rect 15209 9333 15243 9367
rect 2881 9129 2915 9163
rect 5089 9129 5123 9163
rect 5549 9129 5583 9163
rect 8493 9129 8527 9163
rect 9045 9129 9079 9163
rect 9413 9129 9447 9163
rect 11427 9129 11461 9163
rect 13461 9129 13495 9163
rect 14289 9129 14323 9163
rect 15853 9129 15887 9163
rect 4629 9061 4663 9095
rect 7358 9061 7392 9095
rect 10057 9061 10091 9095
rect 10241 9061 10275 9095
rect 11713 9061 11747 9095
rect 11897 9061 11931 9095
rect 13277 9061 13311 9095
rect 15669 9061 15703 9095
rect 1768 8993 1802 9027
rect 3893 8993 3927 9027
rect 4721 8993 4755 9027
rect 5641 8993 5675 9027
rect 10333 8993 10367 9027
rect 12449 8993 12483 9027
rect 13553 8993 13587 9027
rect 13921 8993 13955 9027
rect 18337 8993 18371 9027
rect 1501 8925 1535 8959
rect 4537 8925 4571 8959
rect 7113 8925 7147 8959
rect 11989 8925 12023 8959
rect 15945 8925 15979 8959
rect 16865 8925 16899 8959
rect 4169 8857 4203 8891
rect 10885 8857 10919 8891
rect 12817 8857 12851 8891
rect 3525 8789 3559 8823
rect 5825 8789 5859 8823
rect 6561 8789 6595 8823
rect 6837 8789 6871 8823
rect 9781 8789 9815 8823
rect 11253 8789 11287 8823
rect 13001 8789 13035 8823
rect 15393 8789 15427 8823
rect 18521 8789 18555 8823
rect 1777 8585 1811 8619
rect 8217 8585 8251 8619
rect 8769 8585 8803 8619
rect 9137 8585 9171 8619
rect 11713 8585 11747 8619
rect 12633 8585 12667 8619
rect 15669 8585 15703 8619
rect 16037 8585 16071 8619
rect 16681 8585 16715 8619
rect 18337 8585 18371 8619
rect 5549 8517 5583 8551
rect 12265 8517 12299 8551
rect 2237 8449 2271 8483
rect 2697 8449 2731 8483
rect 3065 8381 3099 8415
rect 3249 8381 3283 8415
rect 5733 8381 5767 8415
rect 6837 8381 6871 8415
rect 9321 8381 9355 8415
rect 12449 8381 12483 8415
rect 13737 8381 13771 8415
rect 2237 8313 2271 8347
rect 2329 8313 2363 8347
rect 3516 8313 3550 8347
rect 5273 8313 5307 8347
rect 6193 8313 6227 8347
rect 7104 8313 7138 8347
rect 9566 8313 9600 8347
rect 11437 8313 11471 8347
rect 13093 8313 13127 8347
rect 14004 8313 14038 8347
rect 16221 8313 16255 8347
rect 4629 8245 4663 8279
rect 6561 8245 6595 8279
rect 10701 8245 10735 8279
rect 13553 8245 13587 8279
rect 15117 8245 15151 8279
rect 1409 8041 1443 8075
rect 1869 8041 1903 8075
rect 2329 8041 2363 8075
rect 8309 8041 8343 8075
rect 11437 8041 11471 8075
rect 13829 8041 13863 8075
rect 16681 8041 16715 8075
rect 2973 7973 3007 8007
rect 4629 7973 4663 8007
rect 10057 7973 10091 8007
rect 10241 7973 10275 8007
rect 10333 7973 10367 8007
rect 15546 7973 15580 8007
rect 3065 7905 3099 7939
rect 5089 7905 5123 7939
rect 5917 7905 5951 7939
rect 6184 7905 6218 7939
rect 8401 7905 8435 7939
rect 11796 7905 11830 7939
rect 15301 7905 15335 7939
rect 18337 7905 18371 7939
rect 20913 7905 20947 7939
rect 2973 7837 3007 7871
rect 4537 7837 4571 7871
rect 4721 7837 4755 7871
rect 11529 7837 11563 7871
rect 14013 7837 14047 7871
rect 18613 7837 18647 7871
rect 21189 7837 21223 7871
rect 2513 7769 2547 7803
rect 3525 7769 3559 7803
rect 8585 7769 8619 7803
rect 9781 7769 9815 7803
rect 3801 7701 3835 7735
rect 4169 7701 4203 7735
rect 5825 7701 5859 7735
rect 7297 7701 7331 7735
rect 7941 7701 7975 7735
rect 9045 7701 9079 7735
rect 9321 7701 9355 7735
rect 10793 7701 10827 7735
rect 12909 7701 12943 7735
rect 14473 7701 14507 7735
rect 18153 7701 18187 7735
rect 2329 7497 2363 7531
rect 3801 7497 3835 7531
rect 4445 7497 4479 7531
rect 4813 7497 4847 7531
rect 6653 7497 6687 7531
rect 7205 7497 7239 7531
rect 10149 7497 10183 7531
rect 12633 7497 12667 7531
rect 13829 7497 13863 7531
rect 20913 7497 20947 7531
rect 5273 7429 5307 7463
rect 7757 7429 7791 7463
rect 9137 7429 9171 7463
rect 10793 7429 10827 7463
rect 2421 7361 2455 7395
rect 5733 7361 5767 7395
rect 7573 7361 7607 7395
rect 8125 7361 8159 7395
rect 10517 7361 10551 7395
rect 11345 7361 11379 7395
rect 13277 7361 13311 7395
rect 14381 7361 14415 7395
rect 17877 7361 17911 7395
rect 18061 7361 18095 7395
rect 2677 7293 2711 7327
rect 8677 7293 8711 7327
rect 9229 7293 9263 7327
rect 9781 7293 9815 7327
rect 11069 7293 11103 7327
rect 12449 7293 12483 7327
rect 14933 7293 14967 7327
rect 15393 7293 15427 7327
rect 15485 7293 15519 7327
rect 18317 7293 18351 7327
rect 21373 7293 21407 7327
rect 22109 7293 22143 7327
rect 5825 7225 5859 7259
rect 8309 7225 8343 7259
rect 11253 7225 11287 7259
rect 14105 7225 14139 7259
rect 15752 7225 15786 7259
rect 21649 7225 21683 7259
rect 1409 7157 1443 7191
rect 1961 7157 1995 7191
rect 5733 7157 5767 7191
rect 6285 7157 6319 7191
rect 8217 7157 8251 7191
rect 9413 7157 9447 7191
rect 11713 7157 11747 7191
rect 12173 7157 12207 7191
rect 13553 7157 13587 7191
rect 14289 7157 14323 7191
rect 16865 7157 16899 7191
rect 19441 7157 19475 7191
rect 2329 6953 2363 6987
rect 3525 6953 3559 6987
rect 3893 6953 3927 6987
rect 6653 6953 6687 6987
rect 7757 6953 7791 6987
rect 8217 6953 8251 6987
rect 9321 6953 9355 6987
rect 10241 6953 10275 6987
rect 13553 6953 13587 6987
rect 13921 6953 13955 6987
rect 15025 6953 15059 6987
rect 15945 6953 15979 6987
rect 18337 6953 18371 6987
rect 2973 6885 3007 6919
rect 4629 6885 4663 6919
rect 4721 6885 4755 6919
rect 6193 6885 6227 6919
rect 6285 6885 6319 6919
rect 11498 6885 11532 6919
rect 16672 6885 16706 6919
rect 4445 6817 4479 6851
rect 5273 6817 5307 6851
rect 8953 6817 8987 6851
rect 10057 6817 10091 6851
rect 10701 6817 10735 6851
rect 13185 6817 13219 6851
rect 13737 6817 13771 6851
rect 15301 6817 15335 6851
rect 16313 6817 16347 6851
rect 19441 6817 19475 6851
rect 1409 6749 1443 6783
rect 2973 6749 3007 6783
rect 3065 6749 3099 6783
rect 6101 6749 6135 6783
rect 7757 6749 7791 6783
rect 7849 6749 7883 6783
rect 10333 6749 10367 6783
rect 11069 6749 11103 6783
rect 11253 6749 11287 6783
rect 16405 6749 16439 6783
rect 4169 6681 4203 6715
rect 5733 6681 5767 6715
rect 8585 6681 8619 6715
rect 15485 6681 15519 6715
rect 17785 6681 17819 6715
rect 1961 6613 1995 6647
rect 2513 6613 2547 6647
rect 7113 6613 7147 6647
rect 7297 6613 7331 6647
rect 9781 6613 9815 6647
rect 12633 6613 12667 6647
rect 14289 6613 14323 6647
rect 14657 6613 14691 6647
rect 19625 6613 19659 6647
rect 2697 6409 2731 6443
rect 4261 6409 4295 6443
rect 5181 6409 5215 6443
rect 6009 6409 6043 6443
rect 9321 6409 9355 6443
rect 11805 6409 11839 6443
rect 12725 6409 12759 6443
rect 15209 6409 15243 6443
rect 16681 6409 16715 6443
rect 17785 6409 17819 6443
rect 19441 6409 19475 6443
rect 14197 6341 14231 6375
rect 15761 6341 15795 6375
rect 17417 6341 17451 6375
rect 18153 6341 18187 6375
rect 25513 6341 25547 6375
rect 2881 6273 2915 6307
rect 9505 6273 9539 6307
rect 12265 6273 12299 6307
rect 16129 6273 16163 6307
rect 16313 6273 16347 6307
rect 17049 6273 17083 6307
rect 18705 6273 18739 6307
rect 24041 6273 24075 6307
rect 1593 6205 1627 6239
rect 5365 6205 5399 6239
rect 7021 6205 7055 6239
rect 7288 6205 7322 6239
rect 9772 6205 9806 6239
rect 11529 6205 11563 6239
rect 12817 6205 12851 6239
rect 13073 6205 13107 6239
rect 19625 6205 19659 6239
rect 20361 6205 20395 6239
rect 24133 6205 24167 6239
rect 24400 6205 24434 6239
rect 1869 6137 1903 6171
rect 3148 6137 3182 6171
rect 18429 6137 18463 6171
rect 18613 6137 18647 6171
rect 19901 6137 19935 6171
rect 2421 6069 2455 6103
rect 4813 6069 4847 6103
rect 5549 6069 5583 6103
rect 6561 6069 6595 6103
rect 8401 6069 8435 6103
rect 8953 6069 8987 6103
rect 10885 6069 10919 6103
rect 14749 6069 14783 6103
rect 15485 6069 15519 6103
rect 16221 6069 16255 6103
rect 1961 5865 1995 5899
rect 2421 5865 2455 5899
rect 3893 5865 3927 5899
rect 8953 5865 8987 5899
rect 9873 5865 9907 5899
rect 10241 5865 10275 5899
rect 17233 5865 17267 5899
rect 18153 5865 18187 5899
rect 24133 5865 24167 5899
rect 1777 5797 1811 5831
rect 2789 5797 2823 5831
rect 2973 5797 3007 5831
rect 7573 5797 7607 5831
rect 7757 5797 7791 5831
rect 10692 5797 10726 5831
rect 13461 5797 13495 5831
rect 13553 5797 13587 5831
rect 14289 5797 14323 5831
rect 15546 5797 15580 5831
rect 4977 5729 5011 5763
rect 7849 5729 7883 5763
rect 10432 5729 10466 5763
rect 13277 5729 13311 5763
rect 18521 5729 18555 5763
rect 20913 5729 20947 5763
rect 2053 5661 2087 5695
rect 4721 5661 4755 5695
rect 7113 5661 7147 5695
rect 15301 5661 15335 5695
rect 17601 5661 17635 5695
rect 18797 5661 18831 5695
rect 19809 5661 19843 5695
rect 1501 5593 1535 5627
rect 3525 5593 3559 5627
rect 7297 5593 7331 5627
rect 13921 5593 13955 5627
rect 4261 5525 4295 5559
rect 6101 5525 6135 5559
rect 6745 5525 6779 5559
rect 8309 5525 8343 5559
rect 8585 5525 8619 5559
rect 9413 5525 9447 5559
rect 11805 5525 11839 5559
rect 12449 5525 12483 5559
rect 13001 5525 13035 5559
rect 15025 5525 15059 5559
rect 16681 5525 16715 5559
rect 21097 5525 21131 5559
rect 1685 5321 1719 5355
rect 3249 5321 3283 5355
rect 3985 5321 4019 5355
rect 4629 5321 4663 5355
rect 6285 5321 6319 5355
rect 10609 5321 10643 5355
rect 11069 5321 11103 5355
rect 11713 5321 11747 5355
rect 13829 5321 13863 5355
rect 14381 5321 14415 5355
rect 14841 5321 14875 5355
rect 16865 5321 16899 5355
rect 18981 5321 19015 5355
rect 21189 5321 21223 5355
rect 4997 5253 5031 5287
rect 5273 5253 5307 5287
rect 9689 5253 9723 5287
rect 5641 5185 5675 5219
rect 5825 5185 5859 5219
rect 7113 5185 7147 5219
rect 14933 5185 14967 5219
rect 1869 5117 1903 5151
rect 9505 5117 9539 5151
rect 10241 5117 10275 5151
rect 11161 5117 11195 5151
rect 12449 5117 12483 5151
rect 12705 5117 12739 5151
rect 15200 5117 15234 5151
rect 17601 5117 17635 5151
rect 18061 5117 18095 5151
rect 18613 5117 18647 5151
rect 19165 5117 19199 5151
rect 19717 5117 19751 5151
rect 20269 5117 20303 5151
rect 20821 5117 20855 5151
rect 21373 5117 21407 5151
rect 21925 5117 21959 5151
rect 22477 5117 22511 5151
rect 23029 5117 23063 5151
rect 2114 5049 2148 5083
rect 4261 5049 4295 5083
rect 5733 5049 5767 5083
rect 7358 5049 7392 5083
rect 9965 5049 9999 5083
rect 10149 5049 10183 5083
rect 6561 4981 6595 5015
rect 8493 4981 8527 5015
rect 9045 4981 9079 5015
rect 11345 4981 11379 5015
rect 12173 4981 12207 5015
rect 16313 4981 16347 5015
rect 17233 4981 17267 5015
rect 18245 4981 18279 5015
rect 19349 4981 19383 5015
rect 20453 4981 20487 5015
rect 21557 4981 21591 5015
rect 22661 4981 22695 5015
rect 1409 4777 1443 4811
rect 3801 4777 3835 4811
rect 5457 4777 5491 4811
rect 6745 4777 6779 4811
rect 7389 4777 7423 4811
rect 7849 4777 7883 4811
rect 8585 4777 8619 4811
rect 10885 4777 10919 4811
rect 11805 4777 11839 4811
rect 12541 4777 12575 4811
rect 14381 4777 14415 4811
rect 15117 4777 15151 4811
rect 15761 4777 15795 4811
rect 17877 4777 17911 4811
rect 2973 4709 3007 4743
rect 3525 4709 3559 4743
rect 4344 4709 4378 4743
rect 7205 4709 7239 4743
rect 7481 4709 7515 4743
rect 10241 4709 10275 4743
rect 11621 4709 11655 4743
rect 11897 4709 11931 4743
rect 13461 4709 13495 4743
rect 13553 4709 13587 4743
rect 18245 4709 18279 4743
rect 18981 4709 19015 4743
rect 4077 4641 4111 4675
rect 8401 4641 8435 4675
rect 10057 4641 10091 4675
rect 15945 4641 15979 4675
rect 16212 4641 16246 4675
rect 20913 4641 20947 4675
rect 22477 4641 22511 4675
rect 22753 4641 22787 4675
rect 23765 4641 23799 4675
rect 2881 4573 2915 4607
rect 3065 4573 3099 4607
rect 10333 4573 10367 4607
rect 13369 4573 13403 4607
rect 14657 4573 14691 4607
rect 18889 4573 18923 4607
rect 19073 4573 19107 4607
rect 13001 4505 13035 4539
rect 2145 4437 2179 4471
rect 2513 4437 2547 4471
rect 6009 4437 6043 4471
rect 6929 4437 6963 4471
rect 8309 4437 8343 4471
rect 9321 4437 9355 4471
rect 9781 4437 9815 4471
rect 11345 4437 11379 4471
rect 13921 4437 13955 4471
rect 17325 4437 17359 4471
rect 18521 4437 18555 4471
rect 21097 4437 21131 4471
rect 23949 4437 23983 4471
rect 7113 4233 7147 4267
rect 7757 4233 7791 4267
rect 9321 4233 9355 4267
rect 10057 4233 10091 4267
rect 10701 4233 10735 4267
rect 11805 4233 11839 4267
rect 12541 4233 12575 4267
rect 13461 4233 13495 4267
rect 16773 4233 16807 4267
rect 18889 4233 18923 4267
rect 19165 4233 19199 4267
rect 22845 4233 22879 4267
rect 24593 4233 24627 4267
rect 3065 4165 3099 4199
rect 1777 4097 1811 4131
rect 2697 4097 2731 4131
rect 4261 4097 4295 4131
rect 6193 4097 6227 4131
rect 6561 4097 6595 4131
rect 7481 4097 7515 4131
rect 8309 4097 8343 4131
rect 9873 4097 9907 4131
rect 5089 4029 5123 4063
rect 5549 4029 5583 4063
rect 10885 4165 10919 4199
rect 15853 4165 15887 4199
rect 11437 4097 11471 4131
rect 12173 4097 12207 4131
rect 12909 4097 12943 4131
rect 13093 4097 13127 4131
rect 13921 4097 13955 4131
rect 14657 4097 14691 4131
rect 17785 4097 17819 4131
rect 18337 4097 18371 4131
rect 14381 4029 14415 4063
rect 16129 4029 16163 4063
rect 17141 4029 17175 4063
rect 18061 4029 18095 4063
rect 19349 4029 19383 4063
rect 19901 4029 19935 4063
rect 20453 4029 20487 4063
rect 21741 4029 21775 4063
rect 22477 4029 22511 4063
rect 23673 4029 23707 4063
rect 24225 4029 24259 4063
rect 24777 4029 24811 4063
rect 25329 4029 25363 4063
rect 2421 3961 2455 3995
rect 2605 3961 2639 3995
rect 3525 3961 3559 3995
rect 3985 3961 4019 3995
rect 4169 3961 4203 3995
rect 5825 3961 5859 3995
rect 8033 3961 8067 3995
rect 8217 3961 8251 3995
rect 8769 3961 8803 3995
rect 9597 3961 9631 3995
rect 10057 3961 10091 3995
rect 10333 3961 10367 3995
rect 11161 3961 11195 3995
rect 11345 3961 11379 3995
rect 13001 3961 13035 3995
rect 14565 3961 14599 3995
rect 15301 3961 15335 3995
rect 16405 3961 16439 3995
rect 22017 3961 22051 3995
rect 1777 3893 1811 3927
rect 1869 3893 1903 3927
rect 2135 3893 2169 3927
rect 3699 3893 3733 3927
rect 4721 3893 4755 3927
rect 5263 3893 5297 3927
rect 5733 3893 5767 3927
rect 9137 3893 9171 3927
rect 9781 3893 9815 3927
rect 14095 3893 14129 3927
rect 15577 3893 15611 3927
rect 16313 3893 16347 3927
rect 19533 3893 19567 3927
rect 20269 3893 20303 3927
rect 20637 3893 20671 3927
rect 21005 3893 21039 3927
rect 23857 3893 23891 3927
rect 24961 3893 24995 3927
rect 2053 3689 2087 3723
rect 3433 3689 3467 3723
rect 3801 3689 3835 3723
rect 7113 3689 7147 3723
rect 8033 3689 8067 3723
rect 9229 3689 9263 3723
rect 10425 3689 10459 3723
rect 10885 3689 10919 3723
rect 12541 3689 12575 3723
rect 13277 3689 13311 3723
rect 14013 3689 14047 3723
rect 14473 3689 14507 3723
rect 16129 3689 16163 3723
rect 16405 3689 16439 3723
rect 19073 3689 19107 3723
rect 19809 3689 19843 3723
rect 19993 3689 20027 3723
rect 2973 3621 3007 3655
rect 4445 3621 4479 3655
rect 4629 3621 4663 3655
rect 5549 3621 5583 3655
rect 8493 3621 8527 3655
rect 9965 3621 9999 3655
rect 11529 3621 11563 3655
rect 11713 3621 11747 3655
rect 14749 3621 14783 3655
rect 17040 3621 17074 3655
rect 18705 3621 18739 3655
rect 3065 3553 3099 3587
rect 6000 3553 6034 3587
rect 8217 3553 8251 3587
rect 9689 3553 9723 3587
rect 13093 3553 13127 3587
rect 15301 3553 15335 3587
rect 16773 3553 16807 3587
rect 19257 3553 19291 3587
rect 1409 3485 1443 3519
rect 2973 3485 3007 3519
rect 4721 3485 4755 3519
rect 5733 3485 5767 3519
rect 11805 3485 11839 3519
rect 13369 3485 13403 3519
rect 15577 3485 15611 3519
rect 23029 3621 23063 3655
rect 20913 3553 20947 3587
rect 22753 3553 22787 3587
rect 24041 3553 24075 3587
rect 25145 3553 25179 3587
rect 2513 3417 2547 3451
rect 11253 3417 11287 3451
rect 19441 3417 19475 3451
rect 19993 3417 20027 3451
rect 4169 3349 4203 3383
rect 5089 3349 5123 3383
rect 7665 3349 7699 3383
rect 12817 3349 12851 3383
rect 18153 3349 18187 3383
rect 20177 3349 20211 3383
rect 21097 3349 21131 3383
rect 24225 3349 24259 3383
rect 25329 3349 25363 3383
rect 2789 3145 2823 3179
rect 5641 3145 5675 3179
rect 9137 3145 9171 3179
rect 10977 3145 11011 3179
rect 11621 3145 11655 3179
rect 11897 3145 11931 3179
rect 13829 3145 13863 3179
rect 14381 3145 14415 3179
rect 15945 3145 15979 3179
rect 16497 3145 16531 3179
rect 17417 3145 17451 3179
rect 17785 3145 17819 3179
rect 19993 3145 20027 3179
rect 21649 3145 21683 3179
rect 22753 3145 22787 3179
rect 23489 3145 23523 3179
rect 25513 3145 25547 3179
rect 3709 3077 3743 3111
rect 1685 3009 1719 3043
rect 3157 3009 3191 3043
rect 3341 3009 3375 3043
rect 15393 3009 15427 3043
rect 16313 3009 16347 3043
rect 16957 3009 16991 3043
rect 18061 3009 18095 3043
rect 1409 2941 1443 2975
rect 4261 2941 4295 2975
rect 6193 2941 6227 2975
rect 6561 2941 6595 2975
rect 7113 2941 7147 2975
rect 7380 2941 7414 2975
rect 9505 2941 9539 2975
rect 9597 2941 9631 2975
rect 12449 2941 12483 2975
rect 12716 2941 12750 2975
rect 14841 2941 14875 2975
rect 15117 2941 15151 2975
rect 17049 2941 17083 2975
rect 20545 2941 20579 2975
rect 21281 2941 21315 2975
rect 21833 2941 21867 2975
rect 22385 2941 22419 2975
rect 23673 2941 23707 2975
rect 24409 2941 24443 2975
rect 24869 2941 24903 2975
rect 24961 2941 24995 2975
rect 2237 2873 2271 2907
rect 4528 2873 4562 2907
rect 9842 2873 9876 2907
rect 16957 2873 16991 2907
rect 18306 2873 18340 2907
rect 20361 2873 20395 2907
rect 20821 2873 20855 2907
rect 23949 2873 23983 2907
rect 2605 2805 2639 2839
rect 3249 2805 3283 2839
rect 4169 2805 4203 2839
rect 8493 2805 8527 2839
rect 19441 2805 19475 2839
rect 22017 2805 22051 2839
rect 25145 2805 25179 2839
rect 2237 2601 2271 2635
rect 3249 2601 3283 2635
rect 3525 2601 3559 2635
rect 5457 2601 5491 2635
rect 6285 2601 6319 2635
rect 6745 2601 6779 2635
rect 8585 2601 8619 2635
rect 11161 2601 11195 2635
rect 12449 2601 12483 2635
rect 14013 2601 14047 2635
rect 16497 2601 16531 2635
rect 18061 2601 18095 2635
rect 19809 2601 19843 2635
rect 21373 2601 21407 2635
rect 1409 2533 1443 2567
rect 2789 2533 2823 2567
rect 2973 2533 3007 2567
rect 4344 2533 4378 2567
rect 7450 2533 7484 2567
rect 9229 2533 9263 2567
rect 10048 2533 10082 2567
rect 12081 2533 12115 2567
rect 12878 2533 12912 2567
rect 14565 2533 14599 2567
rect 17049 2533 17083 2567
rect 18613 2533 18647 2567
rect 24317 2533 24351 2567
rect 3065 2465 3099 2499
rect 3249 2465 3283 2499
rect 7205 2465 7239 2499
rect 9505 2465 9539 2499
rect 9781 2465 9815 2499
rect 12633 2465 12667 2499
rect 15485 2465 15519 2499
rect 16773 2465 16807 2499
rect 17509 2465 17543 2499
rect 18337 2465 18371 2499
rect 19073 2465 19107 2499
rect 19625 2465 19659 2499
rect 20177 2465 20211 2499
rect 21189 2465 21223 2499
rect 21741 2465 21775 2499
rect 22293 2465 22327 2499
rect 22845 2465 22879 2499
rect 24041 2465 24075 2499
rect 24869 2465 24903 2499
rect 25329 2465 25363 2499
rect 25881 2465 25915 2499
rect 1961 2397 1995 2431
rect 3893 2397 3927 2431
rect 4077 2397 4111 2431
rect 15761 2397 15795 2431
rect 20545 2397 20579 2431
rect 2513 2329 2547 2363
rect 25513 2329 25547 2363
rect 14933 2261 14967 2295
rect 19441 2261 19475 2295
rect 22477 2261 22511 2295
<< metal1 >>
rect 2958 26256 2964 26308
rect 3016 26296 3022 26308
rect 15746 26296 15752 26308
rect 3016 26268 15752 26296
rect 3016 26256 3022 26268
rect 15746 26256 15752 26268
rect 15804 26256 15810 26308
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 3418 24896 3424 24948
rect 3476 24936 3482 24948
rect 13262 24936 13268 24948
rect 3476 24908 13268 24936
rect 3476 24896 3482 24908
rect 13262 24896 13268 24908
rect 13320 24896 13326 24948
rect 3510 24828 3516 24880
rect 3568 24868 3574 24880
rect 13998 24868 14004 24880
rect 3568 24840 14004 24868
rect 3568 24828 3574 24840
rect 13998 24828 14004 24840
rect 14056 24828 14062 24880
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1397 14399 1455 14405
rect 1397 14365 1409 14399
rect 1443 14396 1455 14399
rect 2406 14396 2412 14408
rect 1443 14368 2412 14396
rect 1443 14365 1455 14368
rect 1397 14359 1455 14365
rect 2406 14356 2412 14368
rect 2464 14356 2470 14408
rect 2225 14331 2283 14337
rect 2225 14328 2237 14331
rect 1412 14300 2237 14328
rect 1412 14272 1440 14300
rect 2225 14297 2237 14300
rect 2271 14297 2283 14331
rect 2225 14291 2283 14297
rect 1394 14220 1400 14272
rect 1452 14220 1458 14272
rect 1946 14260 1952 14272
rect 1907 14232 1952 14260
rect 1946 14220 1952 14232
rect 2004 14220 2010 14272
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 2038 14056 2044 14068
rect 1999 14028 2044 14056
rect 2038 14016 2044 14028
rect 2096 14016 2102 14068
rect 2777 13923 2835 13929
rect 2777 13889 2789 13923
rect 2823 13920 2835 13923
rect 2866 13920 2872 13932
rect 2823 13892 2872 13920
rect 2823 13889 2835 13892
rect 2777 13883 2835 13889
rect 2866 13880 2872 13892
rect 2924 13880 2930 13932
rect 1397 13855 1455 13861
rect 1397 13821 1409 13855
rect 1443 13852 1455 13855
rect 2038 13852 2044 13864
rect 1443 13824 2044 13852
rect 1443 13821 1455 13824
rect 1397 13815 1455 13821
rect 2038 13812 2044 13824
rect 2096 13812 2102 13864
rect 2222 13812 2228 13864
rect 2280 13852 2286 13864
rect 2317 13855 2375 13861
rect 2317 13852 2329 13855
rect 2280 13824 2329 13852
rect 2280 13812 2286 13824
rect 2317 13821 2329 13824
rect 2363 13821 2375 13855
rect 2317 13815 2375 13821
rect 2130 13744 2136 13796
rect 2188 13784 2194 13796
rect 3053 13787 3111 13793
rect 3053 13784 3065 13787
rect 2188 13756 3065 13784
rect 2188 13744 2194 13756
rect 3053 13753 3065 13756
rect 3099 13753 3111 13787
rect 3053 13747 3111 13753
rect 1578 13716 1584 13728
rect 1539 13688 1584 13716
rect 1578 13676 1584 13688
rect 1636 13676 1642 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 7834 13512 7840 13524
rect 7795 13484 7840 13512
rect 7834 13472 7840 13484
rect 7892 13472 7898 13524
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 2501 13379 2559 13385
rect 1443 13348 2084 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 2056 13249 2084 13348
rect 2501 13345 2513 13379
rect 2547 13376 2559 13379
rect 2590 13376 2596 13388
rect 2547 13348 2596 13376
rect 2547 13345 2559 13348
rect 2501 13339 2559 13345
rect 2590 13336 2596 13348
rect 2648 13376 2654 13388
rect 4982 13376 4988 13388
rect 2648 13348 4988 13376
rect 2648 13336 2654 13348
rect 4982 13336 4988 13348
rect 5040 13336 5046 13388
rect 3145 13311 3203 13317
rect 3145 13277 3157 13311
rect 3191 13308 3203 13311
rect 4154 13308 4160 13320
rect 3191 13280 4160 13308
rect 3191 13277 3203 13280
rect 3145 13271 3203 13277
rect 4154 13268 4160 13280
rect 4212 13268 4218 13320
rect 2041 13243 2099 13249
rect 2041 13209 2053 13243
rect 2087 13240 2099 13243
rect 2498 13240 2504 13252
rect 2087 13212 2504 13240
rect 2087 13209 2099 13212
rect 2041 13203 2099 13209
rect 2498 13200 2504 13212
rect 2556 13200 2562 13252
rect 2958 13200 2964 13252
rect 3016 13240 3022 13252
rect 3789 13243 3847 13249
rect 3789 13240 3801 13243
rect 3016 13212 3801 13240
rect 3016 13200 3022 13212
rect 3789 13209 3801 13212
rect 3835 13209 3847 13243
rect 3789 13203 3847 13209
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13172 1639 13175
rect 1854 13172 1860 13184
rect 1627 13144 1860 13172
rect 1627 13141 1639 13144
rect 1581 13135 1639 13141
rect 1854 13132 1860 13144
rect 1912 13132 1918 13184
rect 2314 13172 2320 13184
rect 2275 13144 2320 13172
rect 2314 13132 2320 13144
rect 2372 13132 2378 13184
rect 2682 13172 2688 13184
rect 2643 13144 2688 13172
rect 2682 13132 2688 13144
rect 2740 13132 2746 13184
rect 3418 13172 3424 13184
rect 3379 13144 3424 13172
rect 3418 13132 3424 13144
rect 3476 13132 3482 13184
rect 4341 13175 4399 13181
rect 4341 13141 4353 13175
rect 4387 13172 4399 13175
rect 4798 13172 4804 13184
rect 4387 13144 4804 13172
rect 4387 13141 4399 13144
rect 4341 13135 4399 13141
rect 4798 13132 4804 13144
rect 4856 13132 4862 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 2590 12968 2596 12980
rect 2551 12940 2596 12968
rect 2590 12928 2596 12940
rect 2648 12928 2654 12980
rect 3694 12968 3700 12980
rect 3655 12940 3700 12968
rect 3694 12928 3700 12940
rect 3752 12928 3758 12980
rect 6086 12968 6092 12980
rect 3896 12940 6092 12968
rect 1673 12903 1731 12909
rect 1673 12869 1685 12903
rect 1719 12900 1731 12903
rect 3896 12900 3924 12940
rect 6086 12928 6092 12940
rect 6144 12928 6150 12980
rect 1719 12872 3924 12900
rect 3973 12903 4031 12909
rect 1719 12869 1731 12872
rect 1673 12863 1731 12869
rect 3973 12869 3985 12903
rect 4019 12900 4031 12903
rect 4706 12900 4712 12912
rect 4019 12872 4712 12900
rect 4019 12869 4031 12872
rect 3973 12863 4031 12869
rect 4706 12860 4712 12872
rect 4764 12860 4770 12912
rect 7929 12903 7987 12909
rect 7929 12869 7941 12903
rect 7975 12900 7987 12903
rect 8294 12900 8300 12912
rect 7975 12872 8300 12900
rect 7975 12869 7987 12872
rect 7929 12863 7987 12869
rect 8294 12860 8300 12872
rect 8352 12860 8358 12912
rect 2130 12832 2136 12844
rect 2091 12804 2136 12832
rect 2130 12792 2136 12804
rect 2188 12792 2194 12844
rect 2225 12835 2283 12841
rect 2225 12801 2237 12835
rect 2271 12832 2283 12835
rect 2314 12832 2320 12844
rect 2271 12804 2320 12832
rect 2271 12801 2283 12804
rect 2225 12795 2283 12801
rect 2314 12792 2320 12804
rect 2372 12832 2378 12844
rect 2774 12832 2780 12844
rect 2372 12804 2780 12832
rect 2372 12792 2378 12804
rect 2774 12792 2780 12804
rect 2832 12792 2838 12844
rect 3421 12835 3479 12841
rect 3421 12801 3433 12835
rect 3467 12832 3479 12835
rect 4433 12835 4491 12841
rect 4433 12832 4445 12835
rect 3467 12804 4445 12832
rect 3467 12801 3479 12804
rect 3421 12795 3479 12801
rect 4433 12801 4445 12804
rect 4479 12832 4491 12835
rect 5442 12832 5448 12844
rect 4479 12804 5448 12832
rect 4479 12801 4491 12804
rect 4433 12795 4491 12801
rect 5442 12792 5448 12804
rect 5500 12792 5506 12844
rect 7377 12767 7435 12773
rect 7377 12733 7389 12767
rect 7423 12764 7435 12767
rect 8481 12767 8539 12773
rect 8481 12764 8493 12767
rect 7423 12736 8493 12764
rect 7423 12733 7435 12736
rect 7377 12727 7435 12733
rect 8481 12733 8493 12736
rect 8527 12764 8539 12767
rect 8938 12764 8944 12776
rect 8527 12736 8944 12764
rect 8527 12733 8539 12736
rect 8481 12727 8539 12733
rect 8938 12724 8944 12736
rect 8996 12724 9002 12776
rect 2038 12656 2044 12708
rect 2096 12696 2102 12708
rect 2133 12699 2191 12705
rect 2133 12696 2145 12699
rect 2096 12668 2145 12696
rect 2096 12656 2102 12668
rect 2133 12665 2145 12668
rect 2179 12696 2191 12699
rect 3418 12696 3424 12708
rect 2179 12668 3424 12696
rect 2179 12665 2191 12668
rect 2133 12659 2191 12665
rect 3418 12656 3424 12668
rect 3476 12656 3482 12708
rect 3694 12656 3700 12708
rect 3752 12696 3758 12708
rect 4433 12699 4491 12705
rect 4433 12696 4445 12699
rect 3752 12668 4445 12696
rect 3752 12656 3758 12668
rect 4433 12665 4445 12668
rect 4479 12665 4491 12699
rect 4433 12659 4491 12665
rect 4525 12699 4583 12705
rect 4525 12665 4537 12699
rect 4571 12696 4583 12699
rect 4614 12696 4620 12708
rect 4571 12668 4620 12696
rect 4571 12665 4583 12668
rect 4525 12659 4583 12665
rect 4614 12656 4620 12668
rect 4672 12656 4678 12708
rect 7834 12656 7840 12708
rect 7892 12696 7898 12708
rect 8205 12699 8263 12705
rect 8205 12696 8217 12699
rect 7892 12668 8217 12696
rect 7892 12656 7898 12668
rect 8205 12665 8217 12668
rect 8251 12665 8263 12699
rect 8205 12659 8263 12665
rect 3050 12628 3056 12640
rect 3011 12600 3056 12628
rect 3050 12588 3056 12600
rect 3108 12588 3114 12640
rect 4890 12628 4896 12640
rect 4851 12600 4896 12628
rect 4890 12588 4896 12600
rect 4948 12588 4954 12640
rect 6638 12588 6644 12640
rect 6696 12628 6702 12640
rect 6825 12631 6883 12637
rect 6825 12628 6837 12631
rect 6696 12600 6837 12628
rect 6696 12588 6702 12600
rect 6825 12597 6837 12600
rect 6871 12597 6883 12631
rect 6825 12591 6883 12597
rect 7745 12631 7803 12637
rect 7745 12597 7757 12631
rect 7791 12628 7803 12631
rect 8389 12631 8447 12637
rect 8389 12628 8401 12631
rect 7791 12600 8401 12628
rect 7791 12597 7803 12600
rect 7745 12591 7803 12597
rect 8389 12597 8401 12600
rect 8435 12628 8447 12631
rect 9122 12628 9128 12640
rect 8435 12600 9128 12628
rect 8435 12597 8447 12600
rect 8389 12591 8447 12597
rect 9122 12588 9128 12600
rect 9180 12588 9186 12640
rect 9401 12631 9459 12637
rect 9401 12597 9413 12631
rect 9447 12628 9459 12631
rect 9582 12628 9588 12640
rect 9447 12600 9588 12628
rect 9447 12597 9459 12600
rect 9401 12591 9459 12597
rect 9582 12588 9588 12600
rect 9640 12588 9646 12640
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1946 12384 1952 12436
rect 2004 12424 2010 12436
rect 2041 12427 2099 12433
rect 2041 12424 2053 12427
rect 2004 12396 2053 12424
rect 2004 12384 2010 12396
rect 2041 12393 2053 12396
rect 2087 12393 2099 12427
rect 2041 12387 2099 12393
rect 2406 12384 2412 12436
rect 2464 12424 2470 12436
rect 2501 12427 2559 12433
rect 2501 12424 2513 12427
rect 2464 12396 2513 12424
rect 2464 12384 2470 12396
rect 2501 12393 2513 12396
rect 2547 12393 2559 12427
rect 2501 12387 2559 12393
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 3237 12427 3295 12433
rect 3237 12424 3249 12427
rect 2832 12396 3249 12424
rect 2832 12384 2838 12396
rect 3237 12393 3249 12396
rect 3283 12424 3295 12427
rect 3326 12424 3332 12436
rect 3283 12396 3332 12424
rect 3283 12393 3295 12396
rect 3237 12387 3295 12393
rect 3326 12384 3332 12396
rect 3384 12384 3390 12436
rect 3142 12316 3148 12368
rect 3200 12356 3206 12368
rect 3602 12356 3608 12368
rect 3200 12328 3608 12356
rect 3200 12316 3206 12328
rect 3602 12316 3608 12328
rect 3660 12316 3666 12368
rect 3878 12316 3884 12368
rect 3936 12356 3942 12368
rect 5258 12356 5264 12368
rect 3936 12328 5264 12356
rect 3936 12316 3942 12328
rect 5258 12316 5264 12328
rect 5316 12316 5322 12368
rect 5350 12316 5356 12368
rect 5408 12356 5414 12368
rect 5445 12359 5503 12365
rect 5445 12356 5457 12359
rect 5408 12328 5457 12356
rect 5408 12316 5414 12328
rect 5445 12325 5457 12328
rect 5491 12325 5503 12359
rect 5902 12356 5908 12368
rect 5863 12328 5908 12356
rect 5445 12319 5503 12325
rect 5902 12316 5908 12328
rect 5960 12316 5966 12368
rect 10036 12359 10094 12365
rect 10036 12325 10048 12359
rect 10082 12356 10094 12359
rect 10134 12356 10140 12368
rect 10082 12328 10140 12356
rect 10082 12325 10094 12328
rect 10036 12319 10094 12325
rect 10134 12316 10140 12328
rect 10192 12316 10198 12368
rect 1394 12248 1400 12300
rect 1452 12288 1458 12300
rect 1857 12291 1915 12297
rect 1857 12288 1869 12291
rect 1452 12260 1869 12288
rect 1452 12248 1458 12260
rect 1857 12257 1869 12260
rect 1903 12288 1915 12291
rect 2314 12288 2320 12300
rect 1903 12260 2320 12288
rect 1903 12257 1915 12260
rect 1857 12251 1915 12257
rect 2314 12248 2320 12260
rect 2372 12248 2378 12300
rect 6713 12291 6771 12297
rect 6713 12288 6725 12291
rect 5552 12260 6725 12288
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12189 2191 12223
rect 2133 12183 2191 12189
rect 4341 12223 4399 12229
rect 4341 12189 4353 12223
rect 4387 12220 4399 12223
rect 4614 12220 4620 12232
rect 4387 12192 4620 12220
rect 4387 12189 4399 12192
rect 4341 12183 4399 12189
rect 1581 12155 1639 12161
rect 1581 12121 1593 12155
rect 1627 12152 1639 12155
rect 2038 12152 2044 12164
rect 1627 12124 2044 12152
rect 1627 12121 1639 12124
rect 1581 12115 1639 12121
rect 2038 12112 2044 12124
rect 2096 12112 2102 12164
rect 2148 12084 2176 12183
rect 4614 12180 4620 12192
rect 4672 12180 4678 12232
rect 5442 12180 5448 12232
rect 5500 12220 5506 12232
rect 5552 12229 5580 12260
rect 6713 12257 6725 12260
rect 6759 12257 6771 12291
rect 6713 12251 6771 12257
rect 5537 12223 5595 12229
rect 5537 12220 5549 12223
rect 5500 12192 5549 12220
rect 5500 12180 5506 12192
rect 5537 12189 5549 12192
rect 5583 12189 5595 12223
rect 6454 12220 6460 12232
rect 6415 12192 6460 12220
rect 5537 12183 5595 12189
rect 6454 12180 6460 12192
rect 6512 12180 6518 12232
rect 9766 12220 9772 12232
rect 9727 12192 9772 12220
rect 9766 12180 9772 12192
rect 9824 12180 9830 12232
rect 2961 12087 3019 12093
rect 2961 12084 2973 12087
rect 2148 12056 2973 12084
rect 2961 12053 2973 12056
rect 3007 12084 3019 12087
rect 3142 12084 3148 12096
rect 3007 12056 3148 12084
rect 3007 12053 3019 12056
rect 2961 12047 3019 12053
rect 3142 12044 3148 12056
rect 3200 12044 3206 12096
rect 3697 12087 3755 12093
rect 3697 12053 3709 12087
rect 3743 12084 3755 12087
rect 4062 12084 4068 12096
rect 3743 12056 4068 12084
rect 3743 12053 3755 12056
rect 3697 12047 3755 12053
rect 4062 12044 4068 12056
rect 4120 12044 4126 12096
rect 4246 12044 4252 12096
rect 4304 12084 4310 12096
rect 4617 12087 4675 12093
rect 4617 12084 4629 12087
rect 4304 12056 4629 12084
rect 4304 12044 4310 12056
rect 4617 12053 4629 12056
rect 4663 12053 4675 12087
rect 4982 12084 4988 12096
rect 4943 12056 4988 12084
rect 4617 12047 4675 12053
rect 4982 12044 4988 12056
rect 5040 12044 5046 12096
rect 7466 12044 7472 12096
rect 7524 12084 7530 12096
rect 7837 12087 7895 12093
rect 7837 12084 7849 12087
rect 7524 12056 7849 12084
rect 7524 12044 7530 12056
rect 7837 12053 7849 12056
rect 7883 12053 7895 12087
rect 11146 12084 11152 12096
rect 11107 12056 11152 12084
rect 7837 12047 7895 12053
rect 11146 12044 11152 12056
rect 11204 12044 11210 12096
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1489 11883 1547 11889
rect 1489 11849 1501 11883
rect 1535 11880 1547 11883
rect 2130 11880 2136 11892
rect 1535 11852 2136 11880
rect 1535 11849 1547 11852
rect 1489 11843 1547 11849
rect 2130 11840 2136 11852
rect 2188 11840 2194 11892
rect 5258 11840 5264 11892
rect 5316 11880 5322 11892
rect 5537 11883 5595 11889
rect 5537 11880 5549 11883
rect 5316 11852 5549 11880
rect 5316 11840 5322 11852
rect 5537 11849 5549 11852
rect 5583 11849 5595 11883
rect 8938 11880 8944 11892
rect 8899 11852 8944 11880
rect 5537 11843 5595 11849
rect 8938 11840 8944 11852
rect 8996 11840 9002 11892
rect 11238 11840 11244 11892
rect 11296 11880 11302 11892
rect 16390 11880 16396 11892
rect 11296 11852 16396 11880
rect 11296 11840 11302 11852
rect 16390 11840 16396 11852
rect 16448 11840 16454 11892
rect 1949 11747 2007 11753
rect 1949 11713 1961 11747
rect 1995 11744 2007 11747
rect 2406 11744 2412 11756
rect 1995 11716 2412 11744
rect 1995 11713 2007 11716
rect 1949 11707 2007 11713
rect 2406 11704 2412 11716
rect 2464 11704 2470 11756
rect 5534 11704 5540 11756
rect 5592 11744 5598 11756
rect 5721 11747 5779 11753
rect 5721 11744 5733 11747
rect 5592 11716 5733 11744
rect 5592 11704 5598 11716
rect 5721 11713 5733 11716
rect 5767 11713 5779 11747
rect 5721 11707 5779 11713
rect 3237 11679 3295 11685
rect 3237 11645 3249 11679
rect 3283 11645 3295 11679
rect 3237 11639 3295 11645
rect 2038 11608 2044 11620
rect 1951 11580 2044 11608
rect 2038 11568 2044 11580
rect 2096 11608 2102 11620
rect 3142 11608 3148 11620
rect 2096 11580 3148 11608
rect 2096 11568 2102 11580
rect 3142 11568 3148 11580
rect 3200 11568 3206 11620
rect 1486 11500 1492 11552
rect 1544 11540 1550 11552
rect 1949 11543 2007 11549
rect 1949 11540 1961 11543
rect 1544 11512 1961 11540
rect 1544 11500 1550 11512
rect 1949 11509 1961 11512
rect 1995 11540 2007 11543
rect 2409 11543 2467 11549
rect 2409 11540 2421 11543
rect 1995 11512 2421 11540
rect 1995 11509 2007 11512
rect 1949 11503 2007 11509
rect 2409 11509 2421 11512
rect 2455 11509 2467 11543
rect 2409 11503 2467 11509
rect 2774 11500 2780 11552
rect 2832 11540 2838 11552
rect 3053 11543 3111 11549
rect 3053 11540 3065 11543
rect 2832 11512 3065 11540
rect 2832 11500 2838 11512
rect 3053 11509 3065 11512
rect 3099 11540 3111 11543
rect 3252 11540 3280 11639
rect 3326 11636 3332 11688
rect 3384 11676 3390 11688
rect 3493 11679 3551 11685
rect 3493 11676 3505 11679
rect 3384 11648 3505 11676
rect 3384 11636 3390 11648
rect 3493 11645 3505 11648
rect 3539 11645 3551 11679
rect 7561 11679 7619 11685
rect 7561 11676 7573 11679
rect 3493 11639 3551 11645
rect 7392 11648 7573 11676
rect 7392 11617 7420 11648
rect 7561 11645 7573 11648
rect 7607 11645 7619 11679
rect 7561 11639 7619 11645
rect 7377 11611 7435 11617
rect 7377 11608 7389 11611
rect 6748 11580 7389 11608
rect 6748 11552 6776 11580
rect 7377 11577 7389 11580
rect 7423 11577 7435 11611
rect 7377 11571 7435 11577
rect 7466 11568 7472 11620
rect 7524 11608 7530 11620
rect 7806 11611 7864 11617
rect 7806 11608 7818 11611
rect 7524 11580 7818 11608
rect 7524 11568 7530 11580
rect 7806 11577 7818 11580
rect 7852 11577 7864 11611
rect 7806 11571 7864 11577
rect 4614 11540 4620 11552
rect 3099 11512 3280 11540
rect 4575 11512 4620 11540
rect 3099 11509 3111 11512
rect 3053 11503 3111 11509
rect 4614 11500 4620 11512
rect 4672 11500 4678 11552
rect 5261 11543 5319 11549
rect 5261 11509 5273 11543
rect 5307 11540 5319 11543
rect 5350 11540 5356 11552
rect 5307 11512 5356 11540
rect 5307 11509 5319 11512
rect 5261 11503 5319 11509
rect 5350 11500 5356 11512
rect 5408 11500 5414 11552
rect 6454 11500 6460 11552
rect 6512 11540 6518 11552
rect 6549 11543 6607 11549
rect 6549 11540 6561 11543
rect 6512 11512 6561 11540
rect 6512 11500 6518 11512
rect 6549 11509 6561 11512
rect 6595 11540 6607 11543
rect 6730 11540 6736 11552
rect 6595 11512 6736 11540
rect 6595 11509 6607 11512
rect 6549 11503 6607 11509
rect 6730 11500 6736 11512
rect 6788 11500 6794 11552
rect 7006 11540 7012 11552
rect 6967 11512 7012 11540
rect 7006 11500 7012 11512
rect 7064 11500 7070 11552
rect 9766 11540 9772 11552
rect 9727 11512 9772 11540
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 10042 11540 10048 11552
rect 10003 11512 10048 11540
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 10134 11500 10140 11552
rect 10192 11540 10198 11552
rect 10505 11543 10563 11549
rect 10505 11540 10517 11543
rect 10192 11512 10517 11540
rect 10192 11500 10198 11512
rect 10505 11509 10517 11512
rect 10551 11509 10563 11543
rect 10505 11503 10563 11509
rect 11149 11543 11207 11549
rect 11149 11509 11161 11543
rect 11195 11540 11207 11543
rect 12158 11540 12164 11552
rect 11195 11512 12164 11540
rect 11195 11509 11207 11512
rect 11149 11503 11207 11509
rect 12158 11500 12164 11512
rect 12216 11500 12222 11552
rect 12437 11543 12495 11549
rect 12437 11509 12449 11543
rect 12483 11540 12495 11543
rect 12710 11540 12716 11552
rect 12483 11512 12716 11540
rect 12483 11509 12495 11512
rect 12437 11503 12495 11509
rect 12710 11500 12716 11512
rect 12768 11500 12774 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 2869 11339 2927 11345
rect 2869 11305 2881 11339
rect 2915 11336 2927 11339
rect 3326 11336 3332 11348
rect 2915 11308 3332 11336
rect 2915 11305 2927 11308
rect 2869 11299 2927 11305
rect 3326 11296 3332 11308
rect 3384 11296 3390 11348
rect 3694 11296 3700 11348
rect 3752 11336 3758 11348
rect 4249 11339 4307 11345
rect 4249 11336 4261 11339
rect 3752 11308 4261 11336
rect 3752 11296 3758 11308
rect 4249 11305 4261 11308
rect 4295 11305 4307 11339
rect 4249 11299 4307 11305
rect 4985 11339 5043 11345
rect 4985 11305 4997 11339
rect 5031 11336 5043 11339
rect 5442 11336 5448 11348
rect 5031 11308 5448 11336
rect 5031 11305 5043 11308
rect 4985 11299 5043 11305
rect 5442 11296 5448 11308
rect 5500 11336 5506 11348
rect 6733 11339 6791 11345
rect 6733 11336 6745 11339
rect 5500 11308 6745 11336
rect 5500 11296 5506 11308
rect 6733 11305 6745 11308
rect 6779 11336 6791 11339
rect 7006 11336 7012 11348
rect 6779 11308 7012 11336
rect 6779 11305 6791 11308
rect 6733 11299 6791 11305
rect 7006 11296 7012 11308
rect 7064 11296 7070 11348
rect 8294 11296 8300 11348
rect 8352 11336 8358 11348
rect 8573 11339 8631 11345
rect 8573 11336 8585 11339
rect 8352 11308 8585 11336
rect 8352 11296 8358 11308
rect 8573 11305 8585 11308
rect 8619 11336 8631 11339
rect 9401 11339 9459 11345
rect 9401 11336 9413 11339
rect 8619 11308 9413 11336
rect 8619 11305 8631 11308
rect 8573 11299 8631 11305
rect 9401 11305 9413 11308
rect 9447 11305 9459 11339
rect 9401 11299 9459 11305
rect 1756 11271 1814 11277
rect 1756 11237 1768 11271
rect 1802 11268 1814 11271
rect 2038 11268 2044 11280
rect 1802 11240 2044 11268
rect 1802 11237 1814 11240
rect 1756 11231 1814 11237
rect 2038 11228 2044 11240
rect 2096 11228 2102 11280
rect 5534 11228 5540 11280
rect 5592 11277 5598 11280
rect 11146 11277 11152 11280
rect 5592 11271 5656 11277
rect 5592 11237 5610 11271
rect 5644 11237 5656 11271
rect 11140 11268 11152 11277
rect 11107 11240 11152 11268
rect 5592 11231 5656 11237
rect 11140 11231 11152 11240
rect 5592 11228 5598 11231
rect 11146 11228 11152 11231
rect 11204 11228 11210 11280
rect 3878 11160 3884 11212
rect 3936 11200 3942 11212
rect 4065 11203 4123 11209
rect 4065 11200 4077 11203
rect 3936 11172 4077 11200
rect 3936 11160 3942 11172
rect 4065 11169 4077 11172
rect 4111 11169 4123 11203
rect 4065 11163 4123 11169
rect 8202 11160 8208 11212
rect 8260 11200 8266 11212
rect 8389 11203 8447 11209
rect 8389 11200 8401 11203
rect 8260 11172 8401 11200
rect 8260 11160 8266 11172
rect 8389 11169 8401 11172
rect 8435 11200 8447 11203
rect 9677 11203 9735 11209
rect 9677 11200 9689 11203
rect 8435 11172 9689 11200
rect 8435 11169 8447 11172
rect 8389 11163 8447 11169
rect 9677 11169 9689 11172
rect 9723 11169 9735 11203
rect 16206 11200 16212 11212
rect 16167 11172 16212 11200
rect 9677 11163 9735 11169
rect 16206 11160 16212 11172
rect 16264 11160 16270 11212
rect 1486 11132 1492 11144
rect 1447 11104 1492 11132
rect 1486 11092 1492 11104
rect 1544 11092 1550 11144
rect 5258 11092 5264 11144
rect 5316 11132 5322 11144
rect 5353 11135 5411 11141
rect 5353 11132 5365 11135
rect 5316 11104 5365 11132
rect 5316 11092 5322 11104
rect 5353 11101 5365 11104
rect 5399 11101 5411 11135
rect 5353 11095 5411 11101
rect 8570 11092 8576 11144
rect 8628 11132 8634 11144
rect 8665 11135 8723 11141
rect 8665 11132 8677 11135
rect 8628 11104 8677 11132
rect 8628 11092 8634 11104
rect 8665 11101 8677 11104
rect 8711 11101 8723 11135
rect 9030 11132 9036 11144
rect 8991 11104 9036 11132
rect 8665 11095 8723 11101
rect 9030 11092 9036 11104
rect 9088 11092 9094 11144
rect 9766 11092 9772 11144
rect 9824 11132 9830 11144
rect 10873 11135 10931 11141
rect 10873 11132 10885 11135
rect 9824 11104 10885 11132
rect 9824 11092 9830 11104
rect 10873 11101 10885 11104
rect 10919 11101 10931 11135
rect 13354 11132 13360 11144
rect 13315 11104 13360 11132
rect 10873 11095 10931 11101
rect 13354 11092 13360 11104
rect 13412 11092 13418 11144
rect 16482 11132 16488 11144
rect 16443 11104 16488 11132
rect 16482 11092 16488 11104
rect 16540 11092 16546 11144
rect 3881 11067 3939 11073
rect 3881 11033 3893 11067
rect 3927 11064 3939 11067
rect 4614 11064 4620 11076
rect 3927 11036 4620 11064
rect 3927 11033 3939 11036
rect 3881 11027 3939 11033
rect 4614 11024 4620 11036
rect 4672 11024 4678 11076
rect 8110 11064 8116 11076
rect 8071 11036 8116 11064
rect 8110 11024 8116 11036
rect 8168 11024 8174 11076
rect 9674 11024 9680 11076
rect 9732 11064 9738 11076
rect 10137 11067 10195 11073
rect 10137 11064 10149 11067
rect 9732 11036 10149 11064
rect 9732 11024 9738 11036
rect 10137 11033 10149 11036
rect 10183 11033 10195 11067
rect 10137 11027 10195 11033
rect 12342 11024 12348 11076
rect 12400 11064 12406 11076
rect 15562 11064 15568 11076
rect 12400 11036 15568 11064
rect 12400 11024 12406 11036
rect 15562 11024 15568 11036
rect 15620 11024 15626 11076
rect 3510 10996 3516 11008
rect 3471 10968 3516 10996
rect 3510 10956 3516 10968
rect 3568 10956 3574 11008
rect 7466 10956 7472 11008
rect 7524 10996 7530 11008
rect 7561 10999 7619 11005
rect 7561 10996 7573 10999
rect 7524 10968 7573 10996
rect 7524 10956 7530 10968
rect 7561 10965 7573 10968
rect 7607 10965 7619 10999
rect 7561 10959 7619 10965
rect 12066 10956 12072 11008
rect 12124 10996 12130 11008
rect 12253 10999 12311 11005
rect 12253 10996 12265 10999
rect 12124 10968 12265 10996
rect 12124 10956 12130 10968
rect 12253 10965 12265 10968
rect 12299 10965 12311 10999
rect 12253 10959 12311 10965
rect 12897 10999 12955 11005
rect 12897 10965 12909 10999
rect 12943 10996 12955 10999
rect 12986 10996 12992 11008
rect 12943 10968 12992 10996
rect 12943 10965 12955 10968
rect 12897 10959 12955 10965
rect 12986 10956 12992 10968
rect 13044 10956 13050 11008
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1762 10752 1768 10804
rect 1820 10792 1826 10804
rect 2038 10792 2044 10804
rect 1820 10764 2044 10792
rect 1820 10752 1826 10764
rect 2038 10752 2044 10764
rect 2096 10752 2102 10804
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 5629 10795 5687 10801
rect 5629 10792 5641 10795
rect 5592 10764 5641 10792
rect 5592 10752 5598 10764
rect 5629 10761 5641 10764
rect 5675 10761 5687 10795
rect 6638 10792 6644 10804
rect 6599 10764 6644 10792
rect 5629 10755 5687 10761
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 8113 10795 8171 10801
rect 8113 10761 8125 10795
rect 8159 10792 8171 10795
rect 8202 10792 8208 10804
rect 8159 10764 8208 10792
rect 8159 10761 8171 10764
rect 8113 10755 8171 10761
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 8570 10752 8576 10804
rect 8628 10792 8634 10804
rect 10045 10795 10103 10801
rect 10045 10792 10057 10795
rect 8628 10764 10057 10792
rect 8628 10752 8634 10764
rect 10045 10761 10057 10764
rect 10091 10792 10103 10795
rect 10134 10792 10140 10804
rect 10091 10764 10140 10792
rect 10091 10761 10103 10764
rect 10045 10755 10103 10761
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 6656 10656 6684 10752
rect 6917 10727 6975 10733
rect 6917 10693 6929 10727
rect 6963 10724 6975 10727
rect 8662 10724 8668 10736
rect 6963 10696 8668 10724
rect 6963 10693 6975 10696
rect 6917 10687 6975 10693
rect 8662 10684 8668 10696
rect 8720 10684 8726 10736
rect 12526 10724 12532 10736
rect 12487 10696 12532 10724
rect 12526 10684 12532 10696
rect 12584 10684 12590 10736
rect 16206 10724 16212 10736
rect 16167 10696 16212 10724
rect 16206 10684 16212 10696
rect 16264 10684 16270 10736
rect 7285 10659 7343 10665
rect 7285 10656 7297 10659
rect 6656 10628 7297 10656
rect 7285 10625 7297 10628
rect 7331 10625 7343 10659
rect 7285 10619 7343 10625
rect 1486 10548 1492 10600
rect 1544 10588 1550 10600
rect 1765 10591 1823 10597
rect 1765 10588 1777 10591
rect 1544 10560 1777 10588
rect 1544 10548 1550 10560
rect 1765 10557 1777 10560
rect 1811 10588 1823 10591
rect 2774 10588 2780 10600
rect 1811 10560 2780 10588
rect 1811 10557 1823 10560
rect 1765 10551 1823 10557
rect 2774 10548 2780 10560
rect 2832 10588 2838 10600
rect 8938 10597 8944 10600
rect 4249 10591 4307 10597
rect 2832 10560 3832 10588
rect 2832 10548 2838 10560
rect 2032 10523 2090 10529
rect 2032 10489 2044 10523
rect 2078 10520 2090 10523
rect 2314 10520 2320 10532
rect 2078 10492 2320 10520
rect 2078 10489 2090 10492
rect 2032 10483 2090 10489
rect 2314 10480 2320 10492
rect 2372 10480 2378 10532
rect 3804 10529 3832 10560
rect 4249 10557 4261 10591
rect 4295 10588 4307 10591
rect 8665 10591 8723 10597
rect 8665 10588 8677 10591
rect 4295 10560 4329 10588
rect 8496 10560 8677 10588
rect 4295 10557 4307 10560
rect 4249 10551 4307 10557
rect 3789 10523 3847 10529
rect 3789 10489 3801 10523
rect 3835 10520 3847 10523
rect 4264 10520 4292 10551
rect 4516 10523 4574 10529
rect 3835 10492 4476 10520
rect 3835 10489 3847 10492
rect 3789 10483 3847 10489
rect 1670 10452 1676 10464
rect 1631 10424 1676 10452
rect 1670 10412 1676 10424
rect 1728 10412 1734 10464
rect 3142 10452 3148 10464
rect 3103 10424 3148 10452
rect 3142 10412 3148 10424
rect 3200 10412 3206 10464
rect 3878 10412 3884 10464
rect 3936 10452 3942 10464
rect 4157 10455 4215 10461
rect 4157 10452 4169 10455
rect 3936 10424 4169 10452
rect 3936 10412 3942 10424
rect 4157 10421 4169 10424
rect 4203 10452 4215 10455
rect 4338 10452 4344 10464
rect 4203 10424 4344 10452
rect 4203 10421 4215 10424
rect 4157 10415 4215 10421
rect 4338 10412 4344 10424
rect 4396 10412 4402 10464
rect 4448 10452 4476 10492
rect 4516 10489 4528 10523
rect 4562 10520 4574 10523
rect 4614 10520 4620 10532
rect 4562 10492 4620 10520
rect 4562 10489 4574 10492
rect 4516 10483 4574 10489
rect 4614 10480 4620 10492
rect 4672 10520 4678 10532
rect 5074 10520 5080 10532
rect 4672 10492 5080 10520
rect 4672 10480 4678 10492
rect 5074 10480 5080 10492
rect 5132 10480 5138 10532
rect 7466 10520 7472 10532
rect 7427 10492 7472 10520
rect 7466 10480 7472 10492
rect 7524 10480 7530 10532
rect 8496 10520 8524 10560
rect 8665 10557 8677 10560
rect 8711 10557 8723 10591
rect 8932 10588 8944 10597
rect 8899 10560 8944 10588
rect 8665 10551 8723 10557
rect 8932 10551 8944 10560
rect 8938 10548 8944 10551
rect 8996 10548 9002 10600
rect 11885 10591 11943 10597
rect 11885 10557 11897 10591
rect 11931 10588 11943 10591
rect 12066 10588 12072 10600
rect 11931 10560 12072 10588
rect 11931 10557 11943 10560
rect 11885 10551 11943 10557
rect 12066 10548 12072 10560
rect 12124 10588 12130 10600
rect 13081 10591 13139 10597
rect 13081 10588 13093 10591
rect 12124 10560 13093 10588
rect 12124 10548 12130 10560
rect 13081 10557 13093 10560
rect 13127 10557 13139 10591
rect 16666 10588 16672 10600
rect 16627 10560 16672 10588
rect 13081 10551 13139 10557
rect 16666 10548 16672 10560
rect 16724 10588 16730 10600
rect 17405 10591 17463 10597
rect 17405 10588 17417 10591
rect 16724 10560 17417 10588
rect 16724 10548 16730 10560
rect 17405 10557 17417 10560
rect 17451 10557 17463 10591
rect 17405 10551 17463 10557
rect 9766 10520 9772 10532
rect 8496 10492 9772 10520
rect 8496 10464 8524 10492
rect 9766 10480 9772 10492
rect 9824 10520 9830 10532
rect 10873 10523 10931 10529
rect 10873 10520 10885 10523
rect 9824 10492 10885 10520
rect 9824 10480 9830 10492
rect 10873 10489 10885 10492
rect 10919 10489 10931 10523
rect 10873 10483 10931 10489
rect 11241 10523 11299 10529
rect 11241 10489 11253 10523
rect 11287 10520 11299 10523
rect 12161 10523 12219 10529
rect 12161 10520 12173 10523
rect 11287 10492 12173 10520
rect 11287 10489 11299 10492
rect 11241 10483 11299 10489
rect 12161 10489 12173 10492
rect 12207 10520 12219 10523
rect 12805 10523 12863 10529
rect 12805 10520 12817 10523
rect 12207 10492 12817 10520
rect 12207 10489 12219 10492
rect 12161 10483 12219 10489
rect 12805 10489 12817 10492
rect 12851 10489 12863 10523
rect 16942 10520 16948 10532
rect 16903 10492 16948 10520
rect 12805 10483 12863 10489
rect 16942 10480 16948 10492
rect 17000 10480 17006 10532
rect 5258 10452 5264 10464
rect 4448 10424 5264 10452
rect 5258 10412 5264 10424
rect 5316 10452 5322 10464
rect 6273 10455 6331 10461
rect 6273 10452 6285 10455
rect 5316 10424 6285 10452
rect 5316 10412 5322 10424
rect 6273 10421 6285 10424
rect 6319 10452 6331 10455
rect 6730 10452 6736 10464
rect 6319 10424 6736 10452
rect 6319 10421 6331 10424
rect 6273 10415 6331 10421
rect 6730 10412 6736 10424
rect 6788 10412 6794 10464
rect 7374 10452 7380 10464
rect 7335 10424 7380 10452
rect 7374 10412 7380 10424
rect 7432 10412 7438 10464
rect 8478 10452 8484 10464
rect 8439 10424 8484 10452
rect 8478 10412 8484 10424
rect 8536 10412 8542 10464
rect 8662 10412 8668 10464
rect 8720 10452 8726 10464
rect 9398 10452 9404 10464
rect 8720 10424 9404 10452
rect 8720 10412 8726 10424
rect 9398 10412 9404 10424
rect 9456 10412 9462 10464
rect 12986 10452 12992 10464
rect 12947 10424 12992 10452
rect 12986 10412 12992 10424
rect 13044 10412 13050 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 3053 10251 3111 10257
rect 3053 10248 3065 10251
rect 2832 10220 3065 10248
rect 2832 10208 2838 10220
rect 3053 10217 3065 10220
rect 3099 10217 3111 10251
rect 3053 10211 3111 10217
rect 3142 10208 3148 10260
rect 3200 10248 3206 10260
rect 3789 10251 3847 10257
rect 3789 10248 3801 10251
rect 3200 10220 3801 10248
rect 3200 10208 3206 10220
rect 3789 10217 3801 10220
rect 3835 10217 3847 10251
rect 5445 10251 5503 10257
rect 3789 10211 3847 10217
rect 4531 10220 5028 10248
rect 1762 10140 1768 10192
rect 1820 10180 1826 10192
rect 2225 10183 2283 10189
rect 2225 10180 2237 10183
rect 1820 10152 2237 10180
rect 1820 10140 1826 10152
rect 2225 10149 2237 10152
rect 2271 10149 2283 10183
rect 2225 10143 2283 10149
rect 566 10072 572 10124
rect 624 10112 630 10124
rect 4531 10112 4559 10220
rect 4614 10140 4620 10192
rect 4672 10180 4678 10192
rect 4893 10183 4951 10189
rect 4893 10180 4905 10183
rect 4672 10152 4905 10180
rect 4672 10140 4678 10152
rect 4893 10149 4905 10152
rect 4939 10149 4951 10183
rect 5000 10180 5028 10220
rect 5445 10217 5457 10251
rect 5491 10248 5503 10251
rect 5534 10248 5540 10260
rect 5491 10220 5540 10248
rect 5491 10217 5503 10220
rect 5445 10211 5503 10217
rect 5534 10208 5540 10220
rect 5592 10208 5598 10260
rect 6362 10248 6368 10260
rect 5644 10220 6368 10248
rect 5644 10180 5672 10220
rect 6362 10208 6368 10220
rect 6420 10208 6426 10260
rect 7009 10251 7067 10257
rect 7009 10217 7021 10251
rect 7055 10248 7067 10251
rect 7466 10248 7472 10260
rect 7055 10220 7472 10248
rect 7055 10217 7067 10220
rect 7009 10211 7067 10217
rect 7466 10208 7472 10220
rect 7524 10208 7530 10260
rect 8021 10251 8079 10257
rect 8021 10217 8033 10251
rect 8067 10248 8079 10251
rect 8110 10248 8116 10260
rect 8067 10220 8116 10248
rect 8067 10217 8079 10220
rect 8021 10211 8079 10217
rect 8110 10208 8116 10220
rect 8168 10208 8174 10260
rect 8570 10248 8576 10260
rect 8531 10220 8576 10248
rect 8570 10208 8576 10220
rect 8628 10208 8634 10260
rect 8938 10248 8944 10260
rect 8899 10220 8944 10248
rect 8938 10208 8944 10220
rect 8996 10208 9002 10260
rect 9493 10251 9551 10257
rect 9493 10217 9505 10251
rect 9539 10248 9551 10251
rect 10965 10251 11023 10257
rect 10965 10248 10977 10251
rect 9539 10220 10977 10248
rect 9539 10217 9551 10220
rect 9493 10211 9551 10217
rect 6270 10180 6276 10192
rect 5000 10152 5672 10180
rect 6231 10152 6276 10180
rect 4893 10143 4951 10149
rect 6270 10140 6276 10152
rect 6328 10140 6334 10192
rect 6454 10180 6460 10192
rect 6415 10152 6460 10180
rect 6454 10140 6460 10152
rect 6512 10140 6518 10192
rect 9674 10140 9680 10192
rect 9732 10180 9738 10192
rect 10137 10183 10195 10189
rect 10137 10180 10149 10183
rect 9732 10152 10149 10180
rect 9732 10140 9738 10152
rect 10137 10149 10149 10152
rect 10183 10149 10195 10183
rect 10137 10143 10195 10149
rect 10226 10140 10232 10192
rect 10284 10180 10290 10192
rect 10428 10189 10456 10220
rect 10965 10217 10977 10220
rect 11011 10248 11023 10251
rect 11146 10248 11152 10260
rect 11011 10220 11152 10248
rect 11011 10217 11023 10220
rect 10965 10211 11023 10217
rect 11146 10208 11152 10220
rect 11204 10208 11210 10260
rect 12066 10189 12072 10192
rect 10321 10183 10379 10189
rect 10321 10180 10333 10183
rect 10284 10152 10333 10180
rect 10284 10140 10290 10152
rect 10321 10149 10333 10152
rect 10367 10149 10379 10183
rect 10321 10143 10379 10149
rect 10413 10183 10471 10189
rect 10413 10149 10425 10183
rect 10459 10149 10471 10183
rect 12060 10180 12072 10189
rect 12027 10152 12072 10180
rect 10413 10143 10471 10149
rect 12060 10143 12072 10152
rect 12066 10140 12072 10143
rect 12124 10140 12130 10192
rect 624 10084 4559 10112
rect 4709 10115 4767 10121
rect 624 10072 630 10084
rect 4709 10081 4721 10115
rect 4755 10112 4767 10115
rect 5166 10112 5172 10124
rect 4755 10084 5172 10112
rect 4755 10081 4767 10084
rect 4709 10075 4767 10081
rect 5166 10072 5172 10084
rect 5224 10072 5230 10124
rect 5813 10115 5871 10121
rect 5813 10081 5825 10115
rect 5859 10112 5871 10115
rect 6549 10115 6607 10121
rect 6549 10112 6561 10115
rect 5859 10084 6561 10112
rect 5859 10081 5871 10084
rect 5813 10075 5871 10081
rect 6549 10081 6561 10084
rect 6595 10112 6607 10115
rect 6822 10112 6828 10124
rect 6595 10084 6828 10112
rect 6595 10081 6607 10084
rect 6549 10075 6607 10081
rect 6822 10072 6828 10084
rect 6880 10072 6886 10124
rect 7377 10115 7435 10121
rect 7377 10081 7389 10115
rect 7423 10112 7435 10115
rect 8113 10115 8171 10121
rect 8113 10112 8125 10115
rect 7423 10084 8125 10112
rect 7423 10081 7435 10084
rect 7377 10075 7435 10081
rect 8113 10081 8125 10084
rect 8159 10112 8171 10115
rect 8294 10112 8300 10124
rect 8159 10084 8300 10112
rect 8159 10081 8171 10084
rect 8113 10075 8171 10081
rect 8294 10072 8300 10084
rect 8352 10072 8358 10124
rect 2130 10044 2136 10056
rect 2091 10016 2136 10044
rect 2130 10004 2136 10016
rect 2188 10004 2194 10056
rect 2314 10044 2320 10056
rect 2227 10016 2320 10044
rect 2314 10004 2320 10016
rect 2372 10044 2378 10056
rect 4985 10047 5043 10053
rect 2372 10016 3556 10044
rect 2372 10004 2378 10016
rect 1765 9979 1823 9985
rect 1765 9945 1777 9979
rect 1811 9976 1823 9979
rect 1946 9976 1952 9988
rect 1811 9948 1952 9976
rect 1811 9945 1823 9948
rect 1765 9939 1823 9945
rect 1946 9936 1952 9948
rect 2004 9936 2010 9988
rect 3528 9920 3556 10016
rect 4985 10013 4997 10047
rect 5031 10044 5043 10047
rect 5074 10044 5080 10056
rect 5031 10016 5080 10044
rect 5031 10013 5043 10016
rect 4985 10007 5043 10013
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 8018 10044 8024 10056
rect 7979 10016 8024 10044
rect 8018 10004 8024 10016
rect 8076 10004 8082 10056
rect 11514 10004 11520 10056
rect 11572 10044 11578 10056
rect 11793 10047 11851 10053
rect 11793 10044 11805 10047
rect 11572 10016 11805 10044
rect 11572 10004 11578 10016
rect 11793 10013 11805 10016
rect 11839 10013 11851 10047
rect 15286 10044 15292 10056
rect 15247 10016 15292 10044
rect 11793 10007 11851 10013
rect 15286 10004 15292 10016
rect 15344 10004 15350 10056
rect 4433 9979 4491 9985
rect 4433 9945 4445 9979
rect 4479 9976 4491 9979
rect 4890 9976 4896 9988
rect 4479 9948 4896 9976
rect 4479 9945 4491 9948
rect 4433 9939 4491 9945
rect 4890 9936 4896 9948
rect 4948 9936 4954 9988
rect 7558 9976 7564 9988
rect 7519 9948 7564 9976
rect 7558 9936 7564 9948
rect 7616 9936 7622 9988
rect 9858 9976 9864 9988
rect 9819 9948 9864 9976
rect 9858 9936 9864 9948
rect 9916 9936 9922 9988
rect 3510 9908 3516 9920
rect 3471 9880 3516 9908
rect 3510 9868 3516 9880
rect 3568 9868 3574 9920
rect 5997 9911 6055 9917
rect 5997 9877 6009 9911
rect 6043 9908 6055 9911
rect 8110 9908 8116 9920
rect 6043 9880 8116 9908
rect 6043 9877 6055 9880
rect 5997 9871 6055 9877
rect 8110 9868 8116 9880
rect 8168 9868 8174 9920
rect 11146 9868 11152 9920
rect 11204 9908 11210 9920
rect 11241 9911 11299 9917
rect 11241 9908 11253 9911
rect 11204 9880 11253 9908
rect 11204 9868 11210 9880
rect 11241 9877 11253 9880
rect 11287 9877 11299 9911
rect 11241 9871 11299 9877
rect 12986 9868 12992 9920
rect 13044 9908 13050 9920
rect 13173 9911 13231 9917
rect 13173 9908 13185 9911
rect 13044 9880 13185 9908
rect 13044 9868 13050 9880
rect 13173 9877 13185 9880
rect 13219 9908 13231 9911
rect 13725 9911 13783 9917
rect 13725 9908 13737 9911
rect 13219 9880 13737 9908
rect 13219 9877 13231 9880
rect 13173 9871 13231 9877
rect 13725 9877 13737 9880
rect 13771 9877 13783 9911
rect 13725 9871 13783 9877
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 4614 9704 4620 9716
rect 4080 9676 4620 9704
rect 2590 9636 2596 9648
rect 2551 9608 2596 9636
rect 2590 9596 2596 9608
rect 2648 9596 2654 9648
rect 3881 9639 3939 9645
rect 3881 9605 3893 9639
rect 3927 9636 3939 9639
rect 4080 9636 4108 9676
rect 4614 9664 4620 9676
rect 4672 9664 4678 9716
rect 5445 9707 5503 9713
rect 5445 9673 5457 9707
rect 5491 9704 5503 9707
rect 5534 9704 5540 9716
rect 5491 9676 5540 9704
rect 5491 9673 5503 9676
rect 5445 9667 5503 9673
rect 4430 9636 4436 9648
rect 3927 9608 4108 9636
rect 4391 9608 4436 9636
rect 3927 9605 3939 9608
rect 3881 9599 3939 9605
rect 4430 9596 4436 9608
rect 4488 9596 4494 9648
rect 3970 9528 3976 9580
rect 4028 9568 4034 9580
rect 4338 9568 4344 9580
rect 4028 9540 4344 9568
rect 4028 9528 4034 9540
rect 4338 9528 4344 9540
rect 4396 9528 4402 9580
rect 4985 9571 5043 9577
rect 4985 9537 4997 9571
rect 5031 9568 5043 9571
rect 5460 9568 5488 9667
rect 5534 9664 5540 9676
rect 5592 9664 5598 9716
rect 6270 9704 6276 9716
rect 6231 9676 6276 9704
rect 6270 9664 6276 9676
rect 6328 9664 6334 9716
rect 7837 9707 7895 9713
rect 7837 9673 7849 9707
rect 7883 9704 7895 9707
rect 8018 9704 8024 9716
rect 7883 9676 8024 9704
rect 7883 9673 7895 9676
rect 7837 9667 7895 9673
rect 8018 9664 8024 9676
rect 8076 9664 8082 9716
rect 8478 9704 8484 9716
rect 8312 9676 8484 9704
rect 6730 9596 6736 9648
rect 6788 9636 6794 9648
rect 8113 9639 8171 9645
rect 8113 9636 8125 9639
rect 6788 9608 8125 9636
rect 6788 9596 6794 9608
rect 8113 9605 8125 9608
rect 8159 9636 8171 9639
rect 8312 9636 8340 9676
rect 8478 9664 8484 9676
rect 8536 9664 8542 9716
rect 12066 9664 12072 9716
rect 12124 9704 12130 9716
rect 12161 9707 12219 9713
rect 12161 9704 12173 9707
rect 12124 9676 12173 9704
rect 12124 9664 12130 9676
rect 12161 9673 12173 9676
rect 12207 9673 12219 9707
rect 12161 9667 12219 9673
rect 8159 9608 8340 9636
rect 8159 9605 8171 9608
rect 8113 9599 8171 9605
rect 5031 9540 5488 9568
rect 5031 9537 5043 9540
rect 4985 9531 5043 9537
rect 5534 9528 5540 9580
rect 5592 9568 5598 9580
rect 5905 9571 5963 9577
rect 5905 9568 5917 9571
rect 5592 9540 5917 9568
rect 5592 9528 5598 9540
rect 5905 9537 5917 9540
rect 5951 9568 5963 9571
rect 6454 9568 6460 9580
rect 5951 9540 6460 9568
rect 5951 9537 5963 9540
rect 5905 9531 5963 9537
rect 6454 9528 6460 9540
rect 6512 9528 6518 9580
rect 8312 9577 8340 9608
rect 9674 9596 9680 9648
rect 9732 9636 9738 9648
rect 10873 9639 10931 9645
rect 10873 9636 10885 9639
rect 9732 9608 10885 9636
rect 9732 9596 9738 9608
rect 10873 9605 10885 9608
rect 10919 9605 10931 9639
rect 10873 9599 10931 9605
rect 16390 9596 16396 9648
rect 16448 9636 16454 9648
rect 17862 9636 17868 9648
rect 16448 9608 17868 9636
rect 16448 9596 16454 9608
rect 17862 9596 17868 9608
rect 17920 9596 17926 9648
rect 8297 9571 8355 9577
rect 8297 9537 8309 9571
rect 8343 9537 8355 9571
rect 10226 9568 10232 9580
rect 10187 9540 10232 9568
rect 8297 9531 8355 9537
rect 10226 9528 10232 9540
rect 10284 9568 10290 9580
rect 11606 9568 11612 9580
rect 10284 9540 11612 9568
rect 10284 9528 10290 9540
rect 11606 9528 11612 9540
rect 11664 9528 11670 9580
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 1670 9500 1676 9512
rect 1443 9472 1676 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1670 9460 1676 9472
rect 1728 9500 1734 9512
rect 2406 9500 2412 9512
rect 1728 9472 2412 9500
rect 1728 9460 1734 9472
rect 2406 9460 2412 9472
rect 2464 9460 2470 9512
rect 2866 9500 2872 9512
rect 2827 9472 2872 9500
rect 2866 9460 2872 9472
rect 2924 9460 2930 9512
rect 4706 9500 4712 9512
rect 4667 9472 4712 9500
rect 4706 9460 4712 9472
rect 4764 9460 4770 9512
rect 6825 9503 6883 9509
rect 6825 9469 6837 9503
rect 6871 9500 6883 9503
rect 7469 9503 7527 9509
rect 7469 9500 7481 9503
rect 6871 9472 7481 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 7469 9469 7481 9472
rect 7515 9500 7527 9503
rect 8110 9500 8116 9512
rect 7515 9472 8116 9500
rect 7515 9469 7527 9472
rect 7469 9463 7527 9469
rect 8110 9460 8116 9472
rect 8168 9460 8174 9512
rect 8386 9460 8392 9512
rect 8444 9500 8450 9512
rect 8553 9503 8611 9509
rect 8553 9500 8565 9503
rect 8444 9472 8565 9500
rect 8444 9460 8450 9472
rect 8553 9469 8565 9472
rect 8599 9469 8611 9503
rect 8553 9463 8611 9469
rect 11514 9460 11520 9512
rect 11572 9500 11578 9512
rect 11885 9503 11943 9509
rect 11885 9500 11897 9503
rect 11572 9472 11897 9500
rect 11572 9460 11578 9472
rect 11885 9469 11897 9472
rect 11931 9500 11943 9503
rect 12713 9503 12771 9509
rect 12713 9500 12725 9503
rect 11931 9472 12725 9500
rect 11931 9469 11943 9472
rect 11885 9463 11943 9469
rect 12713 9469 12725 9472
rect 12759 9500 12771 9503
rect 12802 9500 12808 9512
rect 12759 9472 12808 9500
rect 12759 9469 12771 9472
rect 12713 9463 12771 9469
rect 12802 9460 12808 9472
rect 12860 9460 12866 9512
rect 12986 9509 12992 9512
rect 12980 9500 12992 9509
rect 12912 9472 12992 9500
rect 3142 9432 3148 9444
rect 3103 9404 3148 9432
rect 3142 9392 3148 9404
rect 3200 9392 3206 9444
rect 4246 9432 4252 9444
rect 3712 9404 4252 9432
rect 1486 9324 1492 9376
rect 1544 9364 1550 9376
rect 1581 9367 1639 9373
rect 1581 9364 1593 9367
rect 1544 9336 1593 9364
rect 1544 9324 1550 9336
rect 1581 9333 1593 9336
rect 1627 9333 1639 9367
rect 1581 9327 1639 9333
rect 1762 9324 1768 9376
rect 1820 9364 1826 9376
rect 1946 9364 1952 9376
rect 1820 9336 1952 9364
rect 1820 9324 1826 9336
rect 1946 9324 1952 9336
rect 2004 9324 2010 9376
rect 2130 9324 2136 9376
rect 2188 9364 2194 9376
rect 2409 9367 2467 9373
rect 2409 9364 2421 9367
rect 2188 9336 2421 9364
rect 2188 9324 2194 9336
rect 2409 9333 2421 9336
rect 2455 9364 2467 9367
rect 2682 9364 2688 9376
rect 2455 9336 2688 9364
rect 2455 9333 2467 9336
rect 2409 9327 2467 9333
rect 2682 9324 2688 9336
rect 2740 9324 2746 9376
rect 3050 9364 3056 9376
rect 3011 9336 3056 9364
rect 3050 9324 3056 9336
rect 3108 9364 3114 9376
rect 3712 9364 3740 9404
rect 4246 9392 4252 9404
rect 4304 9392 4310 9444
rect 4890 9432 4896 9444
rect 4851 9404 4896 9432
rect 4890 9392 4896 9404
rect 4948 9392 4954 9444
rect 9766 9392 9772 9444
rect 9824 9432 9830 9444
rect 10689 9435 10747 9441
rect 10689 9432 10701 9435
rect 9824 9404 10701 9432
rect 9824 9392 9830 9404
rect 10689 9401 10701 9404
rect 10735 9432 10747 9435
rect 11149 9435 11207 9441
rect 11149 9432 11161 9435
rect 10735 9404 11161 9432
rect 10735 9401 10747 9404
rect 10689 9395 10747 9401
rect 11149 9401 11161 9404
rect 11195 9401 11207 9435
rect 11149 9395 11207 9401
rect 11238 9392 11244 9444
rect 11296 9432 11302 9444
rect 11425 9435 11483 9441
rect 11425 9432 11437 9435
rect 11296 9404 11437 9432
rect 11296 9392 11302 9404
rect 11425 9401 11437 9404
rect 11471 9401 11483 9435
rect 11425 9395 11483 9401
rect 11974 9392 11980 9444
rect 12032 9432 12038 9444
rect 12912 9432 12940 9472
rect 12980 9463 12992 9472
rect 12986 9460 12992 9463
rect 13044 9460 13050 9512
rect 18046 9500 18052 9512
rect 18007 9472 18052 9500
rect 18046 9460 18052 9472
rect 18104 9500 18110 9512
rect 18785 9503 18843 9509
rect 18785 9500 18797 9503
rect 18104 9472 18797 9500
rect 18104 9460 18110 9472
rect 18785 9469 18797 9472
rect 18831 9469 18843 9503
rect 18785 9463 18843 9469
rect 18322 9432 18328 9444
rect 12032 9404 12940 9432
rect 18283 9404 18328 9432
rect 12032 9392 12038 9404
rect 18322 9392 18328 9404
rect 18380 9392 18386 9444
rect 3108 9336 3740 9364
rect 3108 9324 3114 9336
rect 3786 9324 3792 9376
rect 3844 9364 3850 9376
rect 4157 9367 4215 9373
rect 4157 9364 4169 9367
rect 3844 9336 4169 9364
rect 3844 9324 3850 9336
rect 4157 9333 4169 9336
rect 4203 9364 4215 9367
rect 5166 9364 5172 9376
rect 4203 9336 5172 9364
rect 4203 9333 4215 9336
rect 4157 9327 4215 9333
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 7009 9367 7067 9373
rect 7009 9333 7021 9367
rect 7055 9364 7067 9367
rect 7190 9364 7196 9376
rect 7055 9336 7196 9364
rect 7055 9333 7067 9336
rect 7009 9327 7067 9333
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 9490 9324 9496 9376
rect 9548 9364 9554 9376
rect 9677 9367 9735 9373
rect 9677 9364 9689 9367
rect 9548 9336 9689 9364
rect 9548 9324 9554 9336
rect 9677 9333 9689 9336
rect 9723 9333 9735 9367
rect 11330 9364 11336 9376
rect 11291 9336 11336 9364
rect 9677 9327 9735 9333
rect 11330 9324 11336 9336
rect 11388 9324 11394 9376
rect 14090 9364 14096 9376
rect 14051 9336 14096 9364
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 15197 9367 15255 9373
rect 15197 9333 15209 9367
rect 15243 9364 15255 9367
rect 15562 9364 15568 9376
rect 15243 9336 15568 9364
rect 15243 9333 15255 9336
rect 15197 9327 15255 9333
rect 15562 9324 15568 9336
rect 15620 9324 15626 9376
rect 16666 9324 16672 9376
rect 16724 9364 16730 9376
rect 18690 9364 18696 9376
rect 16724 9336 18696 9364
rect 16724 9324 16730 9336
rect 18690 9324 18696 9336
rect 18748 9324 18754 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 1946 9120 1952 9172
rect 2004 9160 2010 9172
rect 2130 9160 2136 9172
rect 2004 9132 2136 9160
rect 2004 9120 2010 9132
rect 2130 9120 2136 9132
rect 2188 9120 2194 9172
rect 2869 9163 2927 9169
rect 2869 9129 2881 9163
rect 2915 9160 2927 9163
rect 3510 9160 3516 9172
rect 2915 9132 3516 9160
rect 2915 9129 2927 9132
rect 2869 9123 2927 9129
rect 3510 9120 3516 9132
rect 3568 9160 3574 9172
rect 5074 9160 5080 9172
rect 3568 9132 3924 9160
rect 5035 9132 5080 9160
rect 3568 9120 3574 9132
rect 3326 9052 3332 9104
rect 3384 9092 3390 9104
rect 3602 9092 3608 9104
rect 3384 9064 3608 9092
rect 3384 9052 3390 9064
rect 3602 9052 3608 9064
rect 3660 9052 3666 9104
rect 1756 9027 1814 9033
rect 1756 8993 1768 9027
rect 1802 9024 1814 9027
rect 3142 9024 3148 9036
rect 1802 8996 3148 9024
rect 1802 8993 1814 8996
rect 1756 8987 1814 8993
rect 3142 8984 3148 8996
rect 3200 9024 3206 9036
rect 3896 9033 3924 9132
rect 5074 9120 5080 9132
rect 5132 9120 5138 9172
rect 5534 9160 5540 9172
rect 5495 9132 5540 9160
rect 5534 9120 5540 9132
rect 5592 9120 5598 9172
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 8481 9163 8539 9169
rect 8481 9160 8493 9163
rect 8352 9132 8493 9160
rect 8352 9120 8358 9132
rect 8481 9129 8493 9132
rect 8527 9160 8539 9163
rect 9033 9163 9091 9169
rect 9033 9160 9045 9163
rect 8527 9132 9045 9160
rect 8527 9129 8539 9132
rect 8481 9123 8539 9129
rect 9033 9129 9045 9132
rect 9079 9129 9091 9163
rect 9398 9160 9404 9172
rect 9359 9132 9404 9160
rect 9033 9123 9091 9129
rect 9398 9120 9404 9132
rect 9456 9120 9462 9172
rect 11415 9163 11473 9169
rect 11415 9129 11427 9163
rect 11461 9160 11473 9163
rect 13449 9163 13507 9169
rect 13449 9160 13461 9163
rect 11461 9132 13461 9160
rect 11461 9129 11473 9132
rect 11415 9123 11473 9129
rect 13449 9129 13461 9132
rect 13495 9160 13507 9163
rect 14277 9163 14335 9169
rect 14277 9160 14289 9163
rect 13495 9132 14289 9160
rect 13495 9129 13507 9132
rect 13449 9123 13507 9129
rect 14277 9129 14289 9132
rect 14323 9129 14335 9163
rect 14277 9123 14335 9129
rect 14826 9120 14832 9172
rect 14884 9160 14890 9172
rect 15841 9163 15899 9169
rect 15841 9160 15853 9163
rect 14884 9132 15853 9160
rect 14884 9120 14890 9132
rect 15841 9129 15853 9132
rect 15887 9160 15899 9163
rect 16666 9160 16672 9172
rect 15887 9132 16672 9160
rect 15887 9129 15899 9132
rect 15841 9123 15899 9129
rect 16666 9120 16672 9132
rect 16724 9120 16730 9172
rect 4617 9095 4675 9101
rect 4617 9061 4629 9095
rect 4663 9092 4675 9095
rect 5350 9092 5356 9104
rect 4663 9064 5356 9092
rect 4663 9061 4675 9064
rect 4617 9055 4675 9061
rect 5350 9052 5356 9064
rect 5408 9052 5414 9104
rect 6914 9052 6920 9104
rect 6972 9092 6978 9104
rect 7346 9095 7404 9101
rect 7346 9092 7358 9095
rect 6972 9064 7358 9092
rect 6972 9052 6978 9064
rect 7346 9061 7358 9064
rect 7392 9092 7404 9095
rect 8202 9092 8208 9104
rect 7392 9064 8208 9092
rect 7392 9061 7404 9064
rect 7346 9055 7404 9061
rect 8202 9052 8208 9064
rect 8260 9052 8266 9104
rect 8754 9052 8760 9104
rect 8812 9092 8818 9104
rect 10045 9095 10103 9101
rect 10045 9092 10057 9095
rect 8812 9064 10057 9092
rect 8812 9052 8818 9064
rect 10045 9061 10057 9064
rect 10091 9061 10103 9095
rect 10045 9055 10103 9061
rect 10229 9095 10287 9101
rect 10229 9061 10241 9095
rect 10275 9092 10287 9095
rect 11698 9092 11704 9104
rect 10275 9064 10456 9092
rect 11659 9064 11704 9092
rect 10275 9061 10287 9064
rect 10229 9055 10287 9061
rect 3881 9027 3939 9033
rect 3200 8996 3556 9024
rect 3200 8984 3206 8996
rect 1489 8959 1547 8965
rect 1489 8925 1501 8959
rect 1535 8925 1547 8959
rect 1489 8919 1547 8925
rect 1504 8820 1532 8919
rect 1762 8820 1768 8832
rect 1504 8792 1768 8820
rect 1762 8780 1768 8792
rect 1820 8780 1826 8832
rect 3528 8829 3556 8996
rect 3881 8993 3893 9027
rect 3927 9024 3939 9027
rect 4709 9027 4767 9033
rect 4709 9024 4721 9027
rect 3927 8996 4721 9024
rect 3927 8993 3939 8996
rect 3881 8987 3939 8993
rect 4709 8993 4721 8996
rect 4755 8993 4767 9027
rect 4709 8987 4767 8993
rect 5629 9027 5687 9033
rect 5629 8993 5641 9027
rect 5675 9024 5687 9027
rect 6086 9024 6092 9036
rect 5675 8996 6092 9024
rect 5675 8993 5687 8996
rect 5629 8987 5687 8993
rect 6086 8984 6092 8996
rect 6144 8984 6150 9036
rect 9490 8984 9496 9036
rect 9548 9024 9554 9036
rect 10321 9027 10379 9033
rect 10321 9024 10333 9027
rect 9548 8996 10333 9024
rect 9548 8984 9554 8996
rect 10321 8993 10333 8996
rect 10367 8993 10379 9027
rect 10321 8987 10379 8993
rect 4522 8956 4528 8968
rect 4483 8928 4528 8956
rect 4522 8916 4528 8928
rect 4580 8916 4586 8968
rect 7101 8959 7159 8965
rect 7101 8956 7113 8959
rect 6840 8928 7113 8956
rect 4154 8888 4160 8900
rect 4115 8860 4160 8888
rect 4154 8848 4160 8860
rect 4212 8848 4218 8900
rect 6840 8832 6868 8928
rect 7101 8925 7113 8928
rect 7147 8925 7159 8959
rect 7101 8919 7159 8925
rect 9122 8916 9128 8968
rect 9180 8956 9186 8968
rect 10428 8956 10456 9064
rect 11698 9052 11704 9064
rect 11756 9052 11762 9104
rect 11882 9092 11888 9104
rect 11843 9064 11888 9092
rect 11882 9052 11888 9064
rect 11940 9052 11946 9104
rect 13265 9095 13323 9101
rect 13265 9061 13277 9095
rect 13311 9092 13323 9095
rect 13354 9092 13360 9104
rect 13311 9064 13360 9092
rect 13311 9061 13323 9064
rect 13265 9055 13323 9061
rect 13354 9052 13360 9064
rect 13412 9052 13418 9104
rect 15286 9052 15292 9104
rect 15344 9092 15350 9104
rect 15654 9092 15660 9104
rect 15344 9064 15660 9092
rect 15344 9052 15350 9064
rect 15654 9052 15660 9064
rect 15712 9052 15718 9104
rect 12437 9027 12495 9033
rect 12437 8993 12449 9027
rect 12483 9024 12495 9027
rect 13541 9027 13599 9033
rect 13541 9024 13553 9027
rect 12483 8996 13553 9024
rect 12483 8993 12495 8996
rect 12437 8987 12495 8993
rect 13541 8993 13553 8996
rect 13587 9024 13599 9027
rect 13909 9027 13967 9033
rect 13909 9024 13921 9027
rect 13587 8996 13921 9024
rect 13587 8993 13599 8996
rect 13541 8987 13599 8993
rect 13909 8993 13921 8996
rect 13955 9024 13967 9027
rect 14090 9024 14096 9036
rect 13955 8996 14096 9024
rect 13955 8993 13967 8996
rect 13909 8987 13967 8993
rect 14090 8984 14096 8996
rect 14148 8984 14154 9036
rect 18322 9024 18328 9036
rect 18283 8996 18328 9024
rect 18322 8984 18328 8996
rect 18380 8984 18386 9036
rect 11974 8956 11980 8968
rect 9180 8928 10456 8956
rect 11935 8928 11980 8956
rect 9180 8916 9186 8928
rect 11974 8916 11980 8928
rect 12032 8916 12038 8968
rect 15930 8956 15936 8968
rect 15891 8928 15936 8956
rect 15930 8916 15936 8928
rect 15988 8916 15994 8968
rect 16853 8959 16911 8965
rect 16853 8925 16865 8959
rect 16899 8956 16911 8959
rect 17770 8956 17776 8968
rect 16899 8928 17776 8956
rect 16899 8925 16911 8928
rect 16853 8919 16911 8925
rect 17770 8916 17776 8928
rect 17828 8916 17834 8968
rect 9858 8848 9864 8900
rect 9916 8888 9922 8900
rect 10873 8891 10931 8897
rect 10873 8888 10885 8891
rect 9916 8860 10885 8888
rect 9916 8848 9922 8860
rect 10873 8857 10885 8860
rect 10919 8888 10931 8891
rect 11330 8888 11336 8900
rect 10919 8860 11336 8888
rect 10919 8857 10931 8860
rect 10873 8851 10931 8857
rect 11330 8848 11336 8860
rect 11388 8888 11394 8900
rect 12250 8888 12256 8900
rect 11388 8860 12256 8888
rect 11388 8848 11394 8860
rect 12250 8848 12256 8860
rect 12308 8848 12314 8900
rect 12802 8888 12808 8900
rect 12715 8860 12808 8888
rect 12802 8848 12808 8860
rect 12860 8888 12866 8900
rect 13538 8888 13544 8900
rect 12860 8860 13544 8888
rect 12860 8848 12866 8860
rect 13538 8848 13544 8860
rect 13596 8848 13602 8900
rect 3513 8823 3571 8829
rect 3513 8789 3525 8823
rect 3559 8820 3571 8823
rect 3602 8820 3608 8832
rect 3559 8792 3608 8820
rect 3559 8789 3571 8792
rect 3513 8783 3571 8789
rect 3602 8780 3608 8792
rect 3660 8780 3666 8832
rect 5813 8823 5871 8829
rect 5813 8789 5825 8823
rect 5859 8820 5871 8823
rect 6362 8820 6368 8832
rect 5859 8792 6368 8820
rect 5859 8789 5871 8792
rect 5813 8783 5871 8789
rect 6362 8780 6368 8792
rect 6420 8780 6426 8832
rect 6549 8823 6607 8829
rect 6549 8789 6561 8823
rect 6595 8820 6607 8823
rect 6638 8820 6644 8832
rect 6595 8792 6644 8820
rect 6595 8789 6607 8792
rect 6549 8783 6607 8789
rect 6638 8780 6644 8792
rect 6696 8780 6702 8832
rect 6822 8820 6828 8832
rect 6783 8792 6828 8820
rect 6822 8780 6828 8792
rect 6880 8780 6886 8832
rect 9766 8820 9772 8832
rect 9727 8792 9772 8820
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 11238 8820 11244 8832
rect 11199 8792 11244 8820
rect 11238 8780 11244 8792
rect 11296 8780 11302 8832
rect 12986 8820 12992 8832
rect 12947 8792 12992 8820
rect 12986 8780 12992 8792
rect 13044 8780 13050 8832
rect 15378 8820 15384 8832
rect 15339 8792 15384 8820
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 18509 8823 18567 8829
rect 18509 8789 18521 8823
rect 18555 8820 18567 8823
rect 19150 8820 19156 8832
rect 18555 8792 19156 8820
rect 18555 8789 18567 8792
rect 18509 8783 18567 8789
rect 19150 8780 19156 8792
rect 19208 8780 19214 8832
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1765 8619 1823 8625
rect 1765 8585 1777 8619
rect 1811 8616 1823 8619
rect 2866 8616 2872 8628
rect 1811 8588 2872 8616
rect 1811 8585 1823 8588
rect 1765 8579 1823 8585
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 8202 8616 8208 8628
rect 8163 8588 8208 8616
rect 8202 8576 8208 8588
rect 8260 8576 8266 8628
rect 8754 8616 8760 8628
rect 8715 8588 8760 8616
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 9122 8616 9128 8628
rect 9083 8588 9128 8616
rect 9122 8576 9128 8588
rect 9180 8576 9186 8628
rect 11698 8616 11704 8628
rect 11659 8588 11704 8616
rect 11698 8576 11704 8588
rect 11756 8576 11762 8628
rect 12618 8616 12624 8628
rect 12579 8588 12624 8616
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 15654 8616 15660 8628
rect 15615 8588 15660 8616
rect 15654 8576 15660 8588
rect 15712 8576 15718 8628
rect 15930 8576 15936 8628
rect 15988 8616 15994 8628
rect 16025 8619 16083 8625
rect 16025 8616 16037 8619
rect 15988 8588 16037 8616
rect 15988 8576 15994 8588
rect 16025 8585 16037 8588
rect 16071 8585 16083 8619
rect 16666 8616 16672 8628
rect 16627 8588 16672 8616
rect 16025 8579 16083 8585
rect 16666 8576 16672 8588
rect 16724 8576 16730 8628
rect 18322 8616 18328 8628
rect 18283 8588 18328 8616
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 4522 8508 4528 8560
rect 4580 8548 4586 8560
rect 5537 8551 5595 8557
rect 5537 8548 5549 8551
rect 4580 8520 5549 8548
rect 4580 8508 4586 8520
rect 5537 8517 5549 8520
rect 5583 8517 5595 8551
rect 5537 8511 5595 8517
rect 8478 8508 8484 8560
rect 8536 8548 8542 8560
rect 9140 8548 9168 8576
rect 8536 8520 9168 8548
rect 12253 8551 12311 8557
rect 8536 8508 8542 8520
rect 12253 8517 12265 8551
rect 12299 8548 12311 8551
rect 13354 8548 13360 8560
rect 12299 8520 13360 8548
rect 12299 8517 12311 8520
rect 12253 8511 12311 8517
rect 13354 8508 13360 8520
rect 13412 8508 13418 8560
rect 1394 8440 1400 8492
rect 1452 8480 1458 8492
rect 2225 8483 2283 8489
rect 2225 8480 2237 8483
rect 1452 8452 2237 8480
rect 1452 8440 1458 8452
rect 2225 8449 2237 8452
rect 2271 8480 2283 8483
rect 2685 8483 2743 8489
rect 2685 8480 2697 8483
rect 2271 8452 2697 8480
rect 2271 8449 2283 8452
rect 2225 8443 2283 8449
rect 2685 8449 2697 8452
rect 2731 8449 2743 8483
rect 2685 8443 2743 8449
rect 1762 8372 1768 8424
rect 1820 8412 1826 8424
rect 3053 8415 3111 8421
rect 3053 8412 3065 8415
rect 1820 8384 3065 8412
rect 1820 8372 1826 8384
rect 3053 8381 3065 8384
rect 3099 8412 3111 8415
rect 3237 8415 3295 8421
rect 3237 8412 3249 8415
rect 3099 8384 3249 8412
rect 3099 8381 3111 8384
rect 3053 8375 3111 8381
rect 3237 8381 3249 8384
rect 3283 8381 3295 8415
rect 3237 8375 3295 8381
rect 5534 8372 5540 8424
rect 5592 8412 5598 8424
rect 5721 8415 5779 8421
rect 5721 8412 5733 8415
rect 5592 8384 5733 8412
rect 5592 8372 5598 8384
rect 5721 8381 5733 8384
rect 5767 8381 5779 8415
rect 6822 8412 6828 8424
rect 5721 8375 5779 8381
rect 6564 8384 6828 8412
rect 2222 8344 2228 8356
rect 2183 8316 2228 8344
rect 2222 8304 2228 8316
rect 2280 8304 2286 8356
rect 2317 8347 2375 8353
rect 2317 8313 2329 8347
rect 2363 8344 2375 8347
rect 2498 8344 2504 8356
rect 2363 8316 2504 8344
rect 2363 8313 2375 8316
rect 2317 8307 2375 8313
rect 2498 8304 2504 8316
rect 2556 8304 2562 8356
rect 3510 8353 3516 8356
rect 3504 8344 3516 8353
rect 3471 8316 3516 8344
rect 3504 8307 3516 8316
rect 3510 8304 3516 8307
rect 3568 8304 3574 8356
rect 5261 8347 5319 8353
rect 5261 8313 5273 8347
rect 5307 8344 5319 8347
rect 5350 8344 5356 8356
rect 5307 8316 5356 8344
rect 5307 8313 5319 8316
rect 5261 8307 5319 8313
rect 5350 8304 5356 8316
rect 5408 8304 5414 8356
rect 6086 8304 6092 8356
rect 6144 8344 6150 8356
rect 6181 8347 6239 8353
rect 6181 8344 6193 8347
rect 6144 8316 6193 8344
rect 6144 8304 6150 8316
rect 6181 8313 6193 8316
rect 6227 8313 6239 8347
rect 6181 8307 6239 8313
rect 6564 8288 6592 8384
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 9306 8412 9312 8424
rect 9267 8384 9312 8412
rect 9306 8372 9312 8384
rect 9364 8372 9370 8424
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8381 12495 8415
rect 12437 8375 12495 8381
rect 13725 8415 13783 8421
rect 13725 8381 13737 8415
rect 13771 8381 13783 8415
rect 13725 8375 13783 8381
rect 6638 8304 6644 8356
rect 6696 8344 6702 8356
rect 7092 8347 7150 8353
rect 7092 8344 7104 8347
rect 6696 8316 7104 8344
rect 6696 8304 6702 8316
rect 7092 8313 7104 8316
rect 7138 8344 7150 8347
rect 7282 8344 7288 8356
rect 7138 8316 7288 8344
rect 7138 8313 7150 8316
rect 7092 8307 7150 8313
rect 7282 8304 7288 8316
rect 7340 8304 7346 8356
rect 9030 8304 9036 8356
rect 9088 8344 9094 8356
rect 9490 8344 9496 8356
rect 9088 8316 9496 8344
rect 9088 8304 9094 8316
rect 9490 8304 9496 8316
rect 9548 8353 9554 8356
rect 9548 8347 9612 8353
rect 9548 8313 9566 8347
rect 9600 8313 9612 8347
rect 9548 8307 9612 8313
rect 11425 8347 11483 8353
rect 11425 8313 11437 8347
rect 11471 8344 11483 8347
rect 11882 8344 11888 8356
rect 11471 8316 11888 8344
rect 11471 8313 11483 8316
rect 11425 8307 11483 8313
rect 9548 8304 9554 8307
rect 11882 8304 11888 8316
rect 11940 8304 11946 8356
rect 12452 8344 12480 8375
rect 13081 8347 13139 8353
rect 13081 8344 13093 8347
rect 12452 8316 13093 8344
rect 13081 8313 13093 8316
rect 13127 8344 13139 8347
rect 13630 8344 13636 8356
rect 13127 8316 13636 8344
rect 13127 8313 13139 8316
rect 13081 8307 13139 8313
rect 13630 8304 13636 8316
rect 13688 8304 13694 8356
rect 4430 8236 4436 8288
rect 4488 8276 4494 8288
rect 4617 8279 4675 8285
rect 4617 8276 4629 8279
rect 4488 8248 4629 8276
rect 4488 8236 4494 8248
rect 4617 8245 4629 8248
rect 4663 8245 4675 8279
rect 6546 8276 6552 8288
rect 6507 8248 6552 8276
rect 4617 8239 4675 8245
rect 6546 8236 6552 8248
rect 6604 8236 6610 8288
rect 10689 8279 10747 8285
rect 10689 8245 10701 8279
rect 10735 8276 10747 8279
rect 10870 8276 10876 8288
rect 10735 8248 10876 8276
rect 10735 8245 10747 8248
rect 10689 8239 10747 8245
rect 10870 8236 10876 8248
rect 10928 8236 10934 8288
rect 13538 8276 13544 8288
rect 13499 8248 13544 8276
rect 13538 8236 13544 8248
rect 13596 8276 13602 8288
rect 13740 8276 13768 8375
rect 13992 8347 14050 8353
rect 13992 8313 14004 8347
rect 14038 8344 14050 8347
rect 14090 8344 14096 8356
rect 14038 8316 14096 8344
rect 14038 8313 14050 8316
rect 13992 8307 14050 8313
rect 14090 8304 14096 8316
rect 14148 8304 14154 8356
rect 16206 8344 16212 8356
rect 16167 8316 16212 8344
rect 16206 8304 16212 8316
rect 16264 8304 16270 8356
rect 13596 8248 13768 8276
rect 13596 8236 13602 8248
rect 14734 8236 14740 8288
rect 14792 8276 14798 8288
rect 15105 8279 15163 8285
rect 15105 8276 15117 8279
rect 14792 8248 15117 8276
rect 14792 8236 14798 8248
rect 15105 8245 15117 8248
rect 15151 8245 15163 8279
rect 15105 8239 15163 8245
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1394 8072 1400 8084
rect 1355 8044 1400 8072
rect 1394 8032 1400 8044
rect 1452 8032 1458 8084
rect 1762 8032 1768 8084
rect 1820 8072 1826 8084
rect 1857 8075 1915 8081
rect 1857 8072 1869 8075
rect 1820 8044 1869 8072
rect 1820 8032 1826 8044
rect 1857 8041 1869 8044
rect 1903 8041 1915 8075
rect 1857 8035 1915 8041
rect 2317 8075 2375 8081
rect 2317 8041 2329 8075
rect 2363 8072 2375 8075
rect 3602 8072 3608 8084
rect 2363 8044 3608 8072
rect 2363 8041 2375 8044
rect 2317 8035 2375 8041
rect 3602 8032 3608 8044
rect 3660 8032 3666 8084
rect 3786 8032 3792 8084
rect 3844 8032 3850 8084
rect 8294 8072 8300 8084
rect 8255 8044 8300 8072
rect 8294 8032 8300 8044
rect 8352 8032 8358 8084
rect 11425 8075 11483 8081
rect 11425 8041 11437 8075
rect 11471 8072 11483 8075
rect 11974 8072 11980 8084
rect 11471 8044 11980 8072
rect 11471 8041 11483 8044
rect 11425 8035 11483 8041
rect 11974 8032 11980 8044
rect 12032 8032 12038 8084
rect 13814 8072 13820 8084
rect 13775 8044 13820 8072
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 15930 8032 15936 8084
rect 15988 8072 15994 8084
rect 16669 8075 16727 8081
rect 16669 8072 16681 8075
rect 15988 8044 16681 8072
rect 15988 8032 15994 8044
rect 16669 8041 16681 8044
rect 16715 8041 16727 8075
rect 16669 8035 16727 8041
rect 2961 8007 3019 8013
rect 2961 7973 2973 8007
rect 3007 8004 3019 8007
rect 3804 8004 3832 8032
rect 4338 8004 4344 8016
rect 3007 7976 4344 8004
rect 3007 7973 3019 7976
rect 2961 7967 3019 7973
rect 2314 7896 2320 7948
rect 2372 7936 2378 7948
rect 2976 7936 3004 7967
rect 4338 7964 4344 7976
rect 4396 7964 4402 8016
rect 4614 8004 4620 8016
rect 4575 7976 4620 8004
rect 4614 7964 4620 7976
rect 4672 7964 4678 8016
rect 6546 8004 6552 8016
rect 5920 7976 6552 8004
rect 2372 7908 3004 7936
rect 3053 7939 3111 7945
rect 2372 7896 2378 7908
rect 3053 7905 3065 7939
rect 3099 7936 3111 7939
rect 3510 7936 3516 7948
rect 3099 7908 3516 7936
rect 3099 7905 3111 7908
rect 3053 7899 3111 7905
rect 3510 7896 3516 7908
rect 3568 7896 3574 7948
rect 3786 7896 3792 7948
rect 3844 7936 3850 7948
rect 4430 7936 4436 7948
rect 3844 7908 4436 7936
rect 3844 7896 3850 7908
rect 4430 7896 4436 7908
rect 4488 7936 4494 7948
rect 5920 7945 5948 7976
rect 6546 7964 6552 7976
rect 6604 7964 6610 8016
rect 9674 7964 9680 8016
rect 9732 8004 9738 8016
rect 10045 8007 10103 8013
rect 10045 8004 10057 8007
rect 9732 7976 10057 8004
rect 9732 7964 9738 7976
rect 10045 7973 10057 7976
rect 10091 8004 10103 8007
rect 10134 8004 10140 8016
rect 10091 7976 10140 8004
rect 10091 7973 10103 7976
rect 10045 7967 10103 7973
rect 10134 7964 10140 7976
rect 10192 7964 10198 8016
rect 10229 8007 10287 8013
rect 10229 7973 10241 8007
rect 10275 7973 10287 8007
rect 10229 7967 10287 7973
rect 5077 7939 5135 7945
rect 5077 7936 5089 7939
rect 4488 7908 5089 7936
rect 4488 7896 4494 7908
rect 5077 7905 5089 7908
rect 5123 7905 5135 7939
rect 5077 7899 5135 7905
rect 5905 7939 5963 7945
rect 5905 7905 5917 7939
rect 5951 7905 5963 7939
rect 5905 7899 5963 7905
rect 6172 7939 6230 7945
rect 6172 7905 6184 7939
rect 6218 7936 6230 7939
rect 6638 7936 6644 7948
rect 6218 7908 6644 7936
rect 6218 7905 6230 7908
rect 6172 7899 6230 7905
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 8386 7936 8392 7948
rect 8347 7908 8392 7936
rect 8386 7896 8392 7908
rect 8444 7896 8450 7948
rect 9766 7896 9772 7948
rect 9824 7936 9830 7948
rect 10244 7936 10272 7967
rect 10318 7964 10324 8016
rect 10376 8004 10382 8016
rect 10870 8004 10876 8016
rect 10376 7976 10876 8004
rect 10376 7964 10382 7976
rect 10870 7964 10876 7976
rect 10928 7964 10934 8016
rect 14734 7964 14740 8016
rect 14792 8004 14798 8016
rect 15534 8007 15592 8013
rect 15534 8004 15546 8007
rect 14792 7976 15546 8004
rect 14792 7964 14798 7976
rect 15534 7973 15546 7976
rect 15580 7973 15592 8007
rect 15534 7967 15592 7973
rect 11784 7939 11842 7945
rect 9824 7908 10916 7936
rect 9824 7896 9830 7908
rect 10888 7880 10916 7908
rect 11784 7905 11796 7939
rect 11830 7936 11842 7939
rect 12342 7936 12348 7948
rect 11830 7908 12348 7936
rect 11830 7905 11842 7908
rect 11784 7899 11842 7905
rect 12342 7896 12348 7908
rect 12400 7896 12406 7948
rect 13538 7896 13544 7948
rect 13596 7936 13602 7948
rect 15289 7939 15347 7945
rect 15289 7936 15301 7939
rect 13596 7908 15301 7936
rect 13596 7896 13602 7908
rect 15289 7905 15301 7908
rect 15335 7936 15347 7939
rect 16022 7936 16028 7948
rect 15335 7908 16028 7936
rect 15335 7905 15347 7908
rect 15289 7899 15347 7905
rect 16022 7896 16028 7908
rect 16080 7896 16086 7948
rect 18322 7936 18328 7948
rect 18283 7908 18328 7936
rect 18322 7896 18328 7908
rect 18380 7896 18386 7948
rect 20898 7936 20904 7948
rect 20859 7908 20904 7936
rect 20898 7896 20904 7908
rect 20956 7896 20962 7948
rect 2222 7828 2228 7880
rect 2280 7828 2286 7880
rect 2961 7871 3019 7877
rect 2961 7837 2973 7871
rect 3007 7868 3019 7871
rect 3234 7868 3240 7880
rect 3007 7840 3240 7868
rect 3007 7837 3019 7840
rect 2961 7831 3019 7837
rect 3234 7828 3240 7840
rect 3292 7828 3298 7880
rect 4522 7868 4528 7880
rect 4483 7840 4528 7868
rect 4522 7828 4528 7840
rect 4580 7828 4586 7880
rect 4706 7868 4712 7880
rect 4667 7840 4712 7868
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 10870 7828 10876 7880
rect 10928 7828 10934 7880
rect 11514 7868 11520 7880
rect 11475 7840 11520 7868
rect 11514 7828 11520 7840
rect 11572 7828 11578 7880
rect 14001 7871 14059 7877
rect 14001 7837 14013 7871
rect 14047 7868 14059 7871
rect 14366 7868 14372 7880
rect 14047 7840 14372 7868
rect 14047 7837 14059 7840
rect 14001 7831 14059 7837
rect 14366 7828 14372 7840
rect 14424 7828 14430 7880
rect 18601 7871 18659 7877
rect 18601 7837 18613 7871
rect 18647 7868 18659 7871
rect 19334 7868 19340 7880
rect 18647 7840 19340 7868
rect 18647 7837 18659 7840
rect 18601 7831 18659 7837
rect 19334 7828 19340 7840
rect 19392 7828 19398 7880
rect 21177 7871 21235 7877
rect 21177 7837 21189 7871
rect 21223 7868 21235 7871
rect 22002 7868 22008 7880
rect 21223 7840 22008 7868
rect 21223 7837 21235 7840
rect 21177 7831 21235 7837
rect 22002 7828 22008 7840
rect 22060 7828 22066 7880
rect 2240 7800 2268 7828
rect 2501 7803 2559 7809
rect 2501 7800 2513 7803
rect 2240 7772 2513 7800
rect 2501 7769 2513 7772
rect 2547 7769 2559 7803
rect 3510 7800 3516 7812
rect 3423 7772 3516 7800
rect 2501 7763 2559 7769
rect 3510 7760 3516 7772
rect 3568 7800 3574 7812
rect 4724 7800 4752 7828
rect 3568 7772 4752 7800
rect 3568 7760 3574 7772
rect 7006 7760 7012 7812
rect 7064 7800 7070 7812
rect 8573 7803 8631 7809
rect 8573 7800 8585 7803
rect 7064 7772 8585 7800
rect 7064 7760 7070 7772
rect 8573 7769 8585 7772
rect 8619 7769 8631 7803
rect 9766 7800 9772 7812
rect 9727 7772 9772 7800
rect 8573 7763 8631 7769
rect 9766 7760 9772 7772
rect 9824 7760 9830 7812
rect 2590 7692 2596 7744
rect 2648 7732 2654 7744
rect 2958 7732 2964 7744
rect 2648 7704 2964 7732
rect 2648 7692 2654 7704
rect 2958 7692 2964 7704
rect 3016 7692 3022 7744
rect 3786 7732 3792 7744
rect 3747 7704 3792 7732
rect 3786 7692 3792 7704
rect 3844 7692 3850 7744
rect 4062 7692 4068 7744
rect 4120 7732 4126 7744
rect 4157 7735 4215 7741
rect 4157 7732 4169 7735
rect 4120 7704 4169 7732
rect 4120 7692 4126 7704
rect 4157 7701 4169 7704
rect 4203 7701 4215 7735
rect 4157 7695 4215 7701
rect 5813 7735 5871 7741
rect 5813 7701 5825 7735
rect 5859 7732 5871 7735
rect 6914 7732 6920 7744
rect 5859 7704 6920 7732
rect 5859 7701 5871 7704
rect 5813 7695 5871 7701
rect 6914 7692 6920 7704
rect 6972 7692 6978 7744
rect 7282 7732 7288 7744
rect 7243 7704 7288 7732
rect 7282 7692 7288 7704
rect 7340 7692 7346 7744
rect 7929 7735 7987 7741
rect 7929 7701 7941 7735
rect 7975 7732 7987 7735
rect 8018 7732 8024 7744
rect 7975 7704 8024 7732
rect 7975 7701 7987 7704
rect 7929 7695 7987 7701
rect 8018 7692 8024 7704
rect 8076 7692 8082 7744
rect 9030 7732 9036 7744
rect 8991 7704 9036 7732
rect 9030 7692 9036 7704
rect 9088 7692 9094 7744
rect 9306 7732 9312 7744
rect 9267 7704 9312 7732
rect 9306 7692 9312 7704
rect 9364 7692 9370 7744
rect 10781 7735 10839 7741
rect 10781 7701 10793 7735
rect 10827 7732 10839 7735
rect 11330 7732 11336 7744
rect 10827 7704 11336 7732
rect 10827 7701 10839 7704
rect 10781 7695 10839 7701
rect 11330 7692 11336 7704
rect 11388 7692 11394 7744
rect 12894 7732 12900 7744
rect 12855 7704 12900 7732
rect 12894 7692 12900 7704
rect 12952 7692 12958 7744
rect 14458 7732 14464 7744
rect 14419 7704 14464 7732
rect 14458 7692 14464 7704
rect 14516 7692 14522 7744
rect 18138 7732 18144 7744
rect 18099 7704 18144 7732
rect 18138 7692 18144 7704
rect 18196 7692 18202 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 2314 7528 2320 7540
rect 2275 7500 2320 7528
rect 2314 7488 2320 7500
rect 2372 7488 2378 7540
rect 3602 7488 3608 7540
rect 3660 7528 3666 7540
rect 3789 7531 3847 7537
rect 3789 7528 3801 7531
rect 3660 7500 3801 7528
rect 3660 7488 3666 7500
rect 3789 7497 3801 7500
rect 3835 7497 3847 7531
rect 3789 7491 3847 7497
rect 4433 7531 4491 7537
rect 4433 7497 4445 7531
rect 4479 7528 4491 7531
rect 4522 7528 4528 7540
rect 4479 7500 4528 7528
rect 4479 7497 4491 7500
rect 4433 7491 4491 7497
rect 4522 7488 4528 7500
rect 4580 7488 4586 7540
rect 4614 7488 4620 7540
rect 4672 7528 4678 7540
rect 4801 7531 4859 7537
rect 4801 7528 4813 7531
rect 4672 7500 4813 7528
rect 4672 7488 4678 7500
rect 4801 7497 4813 7500
rect 4847 7528 4859 7531
rect 6638 7528 6644 7540
rect 4847 7500 5488 7528
rect 6599 7500 6644 7528
rect 4847 7497 4859 7500
rect 4801 7491 4859 7497
rect 5258 7460 5264 7472
rect 5219 7432 5264 7460
rect 5258 7420 5264 7432
rect 5316 7420 5322 7472
rect 5460 7460 5488 7500
rect 6638 7488 6644 7500
rect 6696 7488 6702 7540
rect 7193 7531 7251 7537
rect 7193 7497 7205 7531
rect 7239 7528 7251 7531
rect 7926 7528 7932 7540
rect 7239 7500 7932 7528
rect 7239 7497 7251 7500
rect 7193 7491 7251 7497
rect 7208 7460 7236 7491
rect 7926 7488 7932 7500
rect 7984 7488 7990 7540
rect 10134 7528 10140 7540
rect 10095 7500 10140 7528
rect 10134 7488 10140 7500
rect 10192 7488 10198 7540
rect 12618 7528 12624 7540
rect 12579 7500 12624 7528
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 13817 7531 13875 7537
rect 13817 7497 13829 7531
rect 13863 7528 13875 7531
rect 14826 7528 14832 7540
rect 13863 7500 14832 7528
rect 13863 7497 13875 7500
rect 13817 7491 13875 7497
rect 14826 7488 14832 7500
rect 14884 7488 14890 7540
rect 20898 7528 20904 7540
rect 20859 7500 20904 7528
rect 20898 7488 20904 7500
rect 20956 7488 20962 7540
rect 7742 7460 7748 7472
rect 5460 7432 7236 7460
rect 7703 7432 7748 7460
rect 7742 7420 7748 7432
rect 7800 7420 7806 7472
rect 9125 7463 9183 7469
rect 9125 7429 9137 7463
rect 9171 7460 9183 7463
rect 9766 7460 9772 7472
rect 9171 7432 9772 7460
rect 9171 7429 9183 7432
rect 9125 7423 9183 7429
rect 9766 7420 9772 7432
rect 9824 7460 9830 7472
rect 10318 7460 10324 7472
rect 9824 7432 10324 7460
rect 9824 7420 9830 7432
rect 10318 7420 10324 7432
rect 10376 7420 10382 7472
rect 10781 7463 10839 7469
rect 10781 7429 10793 7463
rect 10827 7460 10839 7463
rect 10962 7460 10968 7472
rect 10827 7432 10968 7460
rect 10827 7429 10839 7432
rect 10781 7423 10839 7429
rect 10962 7420 10968 7432
rect 11020 7420 11026 7472
rect 1762 7352 1768 7404
rect 1820 7392 1826 7404
rect 2314 7392 2320 7404
rect 1820 7364 2320 7392
rect 1820 7352 1826 7364
rect 2314 7352 2320 7364
rect 2372 7392 2378 7404
rect 2409 7395 2467 7401
rect 2409 7392 2421 7395
rect 2372 7364 2421 7392
rect 2372 7352 2378 7364
rect 2409 7361 2421 7364
rect 2455 7361 2467 7395
rect 5718 7392 5724 7404
rect 5679 7364 5724 7392
rect 2409 7355 2467 7361
rect 5718 7352 5724 7364
rect 5776 7352 5782 7404
rect 7558 7392 7564 7404
rect 7471 7364 7564 7392
rect 7558 7352 7564 7364
rect 7616 7392 7622 7404
rect 8113 7395 8171 7401
rect 8113 7392 8125 7395
rect 7616 7364 8125 7392
rect 7616 7352 7622 7364
rect 8113 7361 8125 7364
rect 8159 7392 8171 7395
rect 8478 7392 8484 7404
rect 8159 7364 8484 7392
rect 8159 7361 8171 7364
rect 8113 7355 8171 7361
rect 8478 7352 8484 7364
rect 8536 7352 8542 7404
rect 10042 7352 10048 7404
rect 10100 7392 10106 7404
rect 10505 7395 10563 7401
rect 10505 7392 10517 7395
rect 10100 7364 10517 7392
rect 10100 7352 10106 7364
rect 10505 7361 10517 7364
rect 10551 7361 10563 7395
rect 11330 7392 11336 7404
rect 11291 7364 11336 7392
rect 10505 7355 10563 7361
rect 2498 7284 2504 7336
rect 2556 7324 2562 7336
rect 2665 7327 2723 7333
rect 2665 7324 2677 7327
rect 2556 7296 2677 7324
rect 2556 7284 2562 7296
rect 2665 7293 2677 7296
rect 2711 7324 2723 7327
rect 3050 7324 3056 7336
rect 2711 7296 3056 7324
rect 2711 7293 2723 7296
rect 2665 7287 2723 7293
rect 3050 7284 3056 7296
rect 3108 7284 3114 7336
rect 6178 7324 6184 7336
rect 5644 7296 6184 7324
rect 1394 7188 1400 7200
rect 1355 7160 1400 7188
rect 1394 7148 1400 7160
rect 1452 7148 1458 7200
rect 1949 7191 2007 7197
rect 1949 7157 1961 7191
rect 1995 7188 2007 7191
rect 3234 7188 3240 7200
rect 1995 7160 3240 7188
rect 1995 7157 2007 7160
rect 1949 7151 2007 7157
rect 3234 7148 3240 7160
rect 3292 7148 3298 7200
rect 5644 7188 5672 7296
rect 6178 7284 6184 7296
rect 6236 7284 6242 7336
rect 8202 7284 8208 7336
rect 8260 7324 8266 7336
rect 8665 7327 8723 7333
rect 8665 7324 8677 7327
rect 8260 7296 8677 7324
rect 8260 7284 8266 7296
rect 8665 7293 8677 7296
rect 8711 7293 8723 7327
rect 8665 7287 8723 7293
rect 9122 7284 9128 7336
rect 9180 7324 9186 7336
rect 9217 7327 9275 7333
rect 9217 7324 9229 7327
rect 9180 7296 9229 7324
rect 9180 7284 9186 7296
rect 9217 7293 9229 7296
rect 9263 7324 9275 7327
rect 9769 7327 9827 7333
rect 9769 7324 9781 7327
rect 9263 7296 9781 7324
rect 9263 7293 9275 7296
rect 9217 7287 9275 7293
rect 9769 7293 9781 7296
rect 9815 7293 9827 7327
rect 9769 7287 9827 7293
rect 5810 7256 5816 7268
rect 5771 7228 5816 7256
rect 5810 7216 5816 7228
rect 5868 7256 5874 7268
rect 7282 7256 7288 7268
rect 5868 7228 7288 7256
rect 5868 7216 5874 7228
rect 7282 7216 7288 7228
rect 7340 7216 7346 7268
rect 8018 7216 8024 7268
rect 8076 7256 8082 7268
rect 8297 7259 8355 7265
rect 8297 7256 8309 7259
rect 8076 7228 8309 7256
rect 8076 7216 8082 7228
rect 8297 7225 8309 7228
rect 8343 7256 8355 7259
rect 9490 7256 9496 7268
rect 8343 7228 9496 7256
rect 8343 7225 8355 7228
rect 8297 7219 8355 7225
rect 9490 7216 9496 7228
rect 9548 7216 9554 7268
rect 10520 7256 10548 7355
rect 11330 7352 11336 7364
rect 11388 7352 11394 7404
rect 13265 7395 13323 7401
rect 13265 7361 13277 7395
rect 13311 7392 13323 7395
rect 14369 7395 14427 7401
rect 14369 7392 14381 7395
rect 13311 7364 14381 7392
rect 13311 7361 13323 7364
rect 13265 7355 13323 7361
rect 14369 7361 14381 7364
rect 14415 7392 14427 7395
rect 14734 7392 14740 7404
rect 14415 7364 14740 7392
rect 14415 7361 14427 7364
rect 14369 7355 14427 7361
rect 14734 7352 14740 7364
rect 14792 7392 14798 7404
rect 15010 7392 15016 7404
rect 14792 7364 15016 7392
rect 14792 7352 14798 7364
rect 15010 7352 15016 7364
rect 15068 7352 15074 7404
rect 17865 7395 17923 7401
rect 17865 7361 17877 7395
rect 17911 7392 17923 7395
rect 18046 7392 18052 7404
rect 17911 7364 18052 7392
rect 17911 7361 17923 7364
rect 17865 7355 17923 7361
rect 10686 7284 10692 7336
rect 10744 7324 10750 7336
rect 11057 7327 11115 7333
rect 11057 7324 11069 7327
rect 10744 7296 11069 7324
rect 10744 7284 10750 7296
rect 11057 7293 11069 7296
rect 11103 7293 11115 7327
rect 11057 7287 11115 7293
rect 12434 7284 12440 7336
rect 12492 7324 12498 7336
rect 14458 7324 14464 7336
rect 12492 7296 14464 7324
rect 12492 7284 12498 7296
rect 14458 7284 14464 7296
rect 14516 7284 14522 7336
rect 14921 7327 14979 7333
rect 14921 7293 14933 7327
rect 14967 7324 14979 7327
rect 15381 7327 15439 7333
rect 15381 7324 15393 7327
rect 14967 7296 15393 7324
rect 14967 7293 14979 7296
rect 14921 7287 14979 7293
rect 15381 7293 15393 7296
rect 15427 7324 15439 7327
rect 15473 7327 15531 7333
rect 15473 7324 15485 7327
rect 15427 7296 15485 7324
rect 15427 7293 15439 7296
rect 15381 7287 15439 7293
rect 15473 7293 15485 7296
rect 15519 7324 15531 7327
rect 16022 7324 16028 7336
rect 15519 7296 16028 7324
rect 15519 7293 15531 7296
rect 15473 7287 15531 7293
rect 16022 7284 16028 7296
rect 16080 7324 16086 7336
rect 16080 7296 16436 7324
rect 16080 7284 16086 7296
rect 16408 7268 16436 7296
rect 11241 7259 11299 7265
rect 11241 7256 11253 7259
rect 10520 7228 11253 7256
rect 11241 7225 11253 7228
rect 11287 7256 11299 7259
rect 11606 7256 11612 7268
rect 11287 7228 11612 7256
rect 11287 7225 11299 7228
rect 11241 7219 11299 7225
rect 11606 7216 11612 7228
rect 11664 7216 11670 7268
rect 13814 7216 13820 7268
rect 13872 7256 13878 7268
rect 14093 7259 14151 7265
rect 14093 7256 14105 7259
rect 13872 7228 14105 7256
rect 13872 7216 13878 7228
rect 14093 7225 14105 7228
rect 14139 7225 14151 7259
rect 14093 7219 14151 7225
rect 15740 7259 15798 7265
rect 15740 7225 15752 7259
rect 15786 7256 15798 7259
rect 15930 7256 15936 7268
rect 15786 7228 15936 7256
rect 15786 7225 15798 7228
rect 15740 7219 15798 7225
rect 15930 7216 15936 7228
rect 15988 7216 15994 7268
rect 16390 7216 16396 7268
rect 16448 7256 16454 7268
rect 17880 7256 17908 7355
rect 18046 7352 18052 7364
rect 18104 7352 18110 7404
rect 18138 7284 18144 7336
rect 18196 7324 18202 7336
rect 18305 7327 18363 7333
rect 18305 7324 18317 7327
rect 18196 7296 18317 7324
rect 18196 7284 18202 7296
rect 18305 7293 18317 7296
rect 18351 7293 18363 7327
rect 21358 7324 21364 7336
rect 21319 7296 21364 7324
rect 18305 7287 18363 7293
rect 21358 7284 21364 7296
rect 21416 7324 21422 7336
rect 22097 7327 22155 7333
rect 22097 7324 22109 7327
rect 21416 7296 22109 7324
rect 21416 7284 21422 7296
rect 22097 7293 22109 7296
rect 22143 7293 22155 7327
rect 22097 7287 22155 7293
rect 21634 7256 21640 7268
rect 16448 7228 17908 7256
rect 21595 7228 21640 7256
rect 16448 7216 16454 7228
rect 21634 7216 21640 7228
rect 21692 7216 21698 7268
rect 5721 7191 5779 7197
rect 5721 7188 5733 7191
rect 5644 7160 5733 7188
rect 5721 7157 5733 7160
rect 5767 7157 5779 7191
rect 5721 7151 5779 7157
rect 6273 7191 6331 7197
rect 6273 7157 6285 7191
rect 6319 7188 6331 7191
rect 6546 7188 6552 7200
rect 6319 7160 6552 7188
rect 6319 7157 6331 7160
rect 6273 7151 6331 7157
rect 6546 7148 6552 7160
rect 6604 7148 6610 7200
rect 7926 7148 7932 7200
rect 7984 7188 7990 7200
rect 8205 7191 8263 7197
rect 8205 7188 8217 7191
rect 7984 7160 8217 7188
rect 7984 7148 7990 7160
rect 8205 7157 8217 7160
rect 8251 7157 8263 7191
rect 8205 7151 8263 7157
rect 8754 7148 8760 7200
rect 8812 7188 8818 7200
rect 9401 7191 9459 7197
rect 9401 7188 9413 7191
rect 8812 7160 9413 7188
rect 8812 7148 8818 7160
rect 9401 7157 9413 7160
rect 9447 7157 9459 7191
rect 9401 7151 9459 7157
rect 11514 7148 11520 7200
rect 11572 7188 11578 7200
rect 11701 7191 11759 7197
rect 11701 7188 11713 7191
rect 11572 7160 11713 7188
rect 11572 7148 11578 7160
rect 11701 7157 11713 7160
rect 11747 7157 11759 7191
rect 11701 7151 11759 7157
rect 12161 7191 12219 7197
rect 12161 7157 12173 7191
rect 12207 7188 12219 7191
rect 12342 7188 12348 7200
rect 12207 7160 12348 7188
rect 12207 7157 12219 7160
rect 12161 7151 12219 7157
rect 12342 7148 12348 7160
rect 12400 7188 12406 7200
rect 12618 7188 12624 7200
rect 12400 7160 12624 7188
rect 12400 7148 12406 7160
rect 12618 7148 12624 7160
rect 12676 7148 12682 7200
rect 13538 7188 13544 7200
rect 13499 7160 13544 7188
rect 13538 7148 13544 7160
rect 13596 7188 13602 7200
rect 14182 7188 14188 7200
rect 13596 7160 14188 7188
rect 13596 7148 13602 7160
rect 14182 7148 14188 7160
rect 14240 7188 14246 7200
rect 14277 7191 14335 7197
rect 14277 7188 14289 7191
rect 14240 7160 14289 7188
rect 14240 7148 14246 7160
rect 14277 7157 14289 7160
rect 14323 7157 14335 7191
rect 16850 7188 16856 7200
rect 16811 7160 16856 7188
rect 14277 7151 14335 7157
rect 16850 7148 16856 7160
rect 16908 7148 16914 7200
rect 19426 7188 19432 7200
rect 19387 7160 19432 7188
rect 19426 7148 19432 7160
rect 19484 7148 19490 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 2314 6984 2320 6996
rect 2275 6956 2320 6984
rect 2314 6944 2320 6956
rect 2372 6944 2378 6996
rect 3513 6987 3571 6993
rect 3513 6953 3525 6987
rect 3559 6984 3571 6987
rect 3881 6987 3939 6993
rect 3881 6984 3893 6987
rect 3559 6956 3893 6984
rect 3559 6953 3571 6956
rect 3513 6947 3571 6953
rect 3881 6953 3893 6956
rect 3927 6984 3939 6987
rect 4246 6984 4252 6996
rect 3927 6956 4252 6984
rect 3927 6953 3939 6956
rect 3881 6947 3939 6953
rect 4246 6944 4252 6956
rect 4304 6984 4310 6996
rect 6638 6984 6644 6996
rect 4304 6956 4752 6984
rect 4304 6944 4310 6956
rect 4724 6928 4752 6956
rect 6288 6956 6644 6984
rect 2682 6876 2688 6928
rect 2740 6916 2746 6928
rect 2961 6919 3019 6925
rect 2740 6888 2912 6916
rect 2740 6876 2746 6888
rect 2884 6792 2912 6888
rect 2961 6885 2973 6919
rect 3007 6916 3019 6919
rect 4062 6916 4068 6928
rect 3007 6888 4068 6916
rect 3007 6885 3019 6888
rect 2961 6879 3019 6885
rect 4062 6876 4068 6888
rect 4120 6876 4126 6928
rect 4617 6919 4675 6925
rect 4617 6885 4629 6919
rect 4663 6885 4675 6919
rect 4617 6879 4675 6885
rect 4430 6848 4436 6860
rect 4391 6820 4436 6848
rect 4430 6808 4436 6820
rect 4488 6808 4494 6860
rect 4632 6848 4660 6879
rect 4706 6876 4712 6928
rect 4764 6916 4770 6928
rect 5810 6916 5816 6928
rect 4764 6888 4809 6916
rect 5460 6888 5816 6916
rect 4764 6876 4770 6888
rect 5261 6851 5319 6857
rect 4632 6820 4752 6848
rect 4724 6792 4752 6820
rect 5261 6817 5273 6851
rect 5307 6848 5319 6851
rect 5460 6848 5488 6888
rect 5810 6876 5816 6888
rect 5868 6876 5874 6928
rect 6288 6925 6316 6956
rect 6638 6944 6644 6956
rect 6696 6944 6702 6996
rect 7742 6984 7748 6996
rect 7655 6956 7748 6984
rect 7742 6944 7748 6956
rect 7800 6984 7806 6996
rect 8205 6987 8263 6993
rect 8205 6984 8217 6987
rect 7800 6956 8217 6984
rect 7800 6944 7806 6956
rect 8205 6953 8217 6956
rect 8251 6953 8263 6987
rect 8205 6947 8263 6953
rect 9030 6944 9036 6996
rect 9088 6984 9094 6996
rect 9309 6987 9367 6993
rect 9309 6984 9321 6987
rect 9088 6956 9321 6984
rect 9088 6944 9094 6956
rect 9309 6953 9321 6956
rect 9355 6953 9367 6987
rect 9309 6947 9367 6953
rect 9858 6944 9864 6996
rect 9916 6984 9922 6996
rect 10229 6987 10287 6993
rect 10229 6984 10241 6987
rect 9916 6956 10241 6984
rect 9916 6944 9922 6956
rect 10229 6953 10241 6956
rect 10275 6984 10287 6987
rect 13541 6987 13599 6993
rect 13541 6984 13553 6987
rect 10275 6956 13553 6984
rect 10275 6953 10287 6956
rect 10229 6947 10287 6953
rect 13541 6953 13553 6956
rect 13587 6953 13599 6987
rect 13906 6984 13912 6996
rect 13867 6956 13912 6984
rect 13541 6947 13599 6953
rect 13906 6944 13912 6956
rect 13964 6944 13970 6996
rect 15010 6984 15016 6996
rect 14971 6956 15016 6984
rect 15010 6944 15016 6956
rect 15068 6944 15074 6996
rect 15930 6984 15936 6996
rect 15891 6956 15936 6984
rect 15930 6944 15936 6956
rect 15988 6944 15994 6996
rect 18322 6984 18328 6996
rect 18283 6956 18328 6984
rect 18322 6944 18328 6956
rect 18380 6944 18386 6996
rect 6181 6919 6239 6925
rect 6181 6885 6193 6919
rect 6227 6885 6239 6919
rect 6181 6879 6239 6885
rect 6273 6919 6331 6925
rect 6273 6885 6285 6919
rect 6319 6885 6331 6919
rect 6273 6879 6331 6885
rect 5307 6820 5488 6848
rect 5307 6817 5319 6820
rect 5261 6811 5319 6817
rect 5994 6808 6000 6860
rect 6052 6848 6058 6860
rect 6196 6848 6224 6879
rect 7374 6876 7380 6928
rect 7432 6916 7438 6928
rect 7834 6916 7840 6928
rect 7432 6888 7840 6916
rect 7432 6876 7438 6888
rect 7834 6876 7840 6888
rect 7892 6876 7898 6928
rect 11330 6876 11336 6928
rect 11388 6916 11394 6928
rect 11486 6919 11544 6925
rect 11486 6916 11498 6919
rect 11388 6888 11498 6916
rect 11388 6876 11394 6888
rect 11486 6885 11498 6888
rect 11532 6885 11544 6919
rect 16660 6919 16718 6925
rect 16660 6916 16672 6919
rect 11486 6879 11544 6885
rect 16592 6888 16672 6916
rect 6052 6820 6224 6848
rect 6052 6808 6058 6820
rect 7650 6808 7656 6860
rect 7708 6848 7714 6860
rect 8941 6851 8999 6857
rect 8941 6848 8953 6851
rect 7708 6820 8953 6848
rect 7708 6808 7714 6820
rect 8941 6817 8953 6820
rect 8987 6817 8999 6851
rect 10042 6848 10048 6860
rect 10003 6820 10048 6848
rect 8941 6811 8999 6817
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 10686 6848 10692 6860
rect 10647 6820 10692 6848
rect 10686 6808 10692 6820
rect 10744 6808 10750 6860
rect 13170 6848 13176 6860
rect 13131 6820 13176 6848
rect 13170 6808 13176 6820
rect 13228 6808 13234 6860
rect 13722 6848 13728 6860
rect 13683 6820 13728 6848
rect 13722 6808 13728 6820
rect 13780 6808 13786 6860
rect 14826 6808 14832 6860
rect 14884 6848 14890 6860
rect 15289 6851 15347 6857
rect 15289 6848 15301 6851
rect 14884 6820 15301 6848
rect 14884 6808 14890 6820
rect 15289 6817 15301 6820
rect 15335 6817 15347 6851
rect 16298 6848 16304 6860
rect 16211 6820 16304 6848
rect 15289 6811 15347 6817
rect 16298 6808 16304 6820
rect 16356 6848 16362 6860
rect 16592 6848 16620 6888
rect 16660 6885 16672 6888
rect 16706 6916 16718 6919
rect 16850 6916 16856 6928
rect 16706 6888 16856 6916
rect 16706 6885 16718 6888
rect 16660 6879 16718 6885
rect 16850 6876 16856 6888
rect 16908 6876 16914 6928
rect 16356 6820 16620 6848
rect 16356 6808 16362 6820
rect 19334 6808 19340 6860
rect 19392 6848 19398 6860
rect 19429 6851 19487 6857
rect 19429 6848 19441 6851
rect 19392 6820 19441 6848
rect 19392 6808 19398 6820
rect 19429 6817 19441 6820
rect 19475 6817 19487 6851
rect 19429 6811 19487 6817
rect 1394 6780 1400 6792
rect 1355 6752 1400 6780
rect 1394 6740 1400 6752
rect 1452 6740 1458 6792
rect 2866 6740 2872 6792
rect 2924 6740 2930 6792
rect 2961 6783 3019 6789
rect 2961 6749 2973 6783
rect 3007 6749 3019 6783
rect 2961 6743 3019 6749
rect 2976 6712 3004 6743
rect 3050 6740 3056 6792
rect 3108 6780 3114 6792
rect 3786 6780 3792 6792
rect 3108 6752 3792 6780
rect 3108 6740 3114 6752
rect 3786 6740 3792 6752
rect 3844 6740 3850 6792
rect 4706 6740 4712 6792
rect 4764 6740 4770 6792
rect 5166 6740 5172 6792
rect 5224 6780 5230 6792
rect 6089 6783 6147 6789
rect 6089 6780 6101 6783
rect 5224 6752 6101 6780
rect 5224 6740 5230 6752
rect 6089 6749 6101 6752
rect 6135 6749 6147 6783
rect 7742 6780 7748 6792
rect 7703 6752 7748 6780
rect 6089 6743 6147 6749
rect 7742 6740 7748 6752
rect 7800 6740 7806 6792
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6780 7895 6783
rect 8386 6780 8392 6792
rect 7883 6752 8392 6780
rect 7883 6749 7895 6752
rect 7837 6743 7895 6749
rect 8386 6740 8392 6752
rect 8444 6740 8450 6792
rect 10134 6740 10140 6792
rect 10192 6780 10198 6792
rect 10321 6783 10379 6789
rect 10321 6780 10333 6783
rect 10192 6752 10333 6780
rect 10192 6740 10198 6752
rect 10321 6749 10333 6752
rect 10367 6749 10379 6783
rect 11054 6780 11060 6792
rect 11015 6752 11060 6780
rect 10321 6743 10379 6749
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 11241 6783 11299 6789
rect 11241 6749 11253 6783
rect 11287 6749 11299 6783
rect 16390 6780 16396 6792
rect 16351 6752 16396 6780
rect 11241 6743 11299 6749
rect 4154 6712 4160 6724
rect 2976 6684 4160 6712
rect 4154 6672 4160 6684
rect 4212 6672 4218 6724
rect 5718 6712 5724 6724
rect 5679 6684 5724 6712
rect 5718 6672 5724 6684
rect 5776 6672 5782 6724
rect 7760 6712 7788 6740
rect 8573 6715 8631 6721
rect 8573 6712 8585 6715
rect 7760 6684 8585 6712
rect 8573 6681 8585 6684
rect 8619 6681 8631 6715
rect 8573 6675 8631 6681
rect 9306 6672 9312 6724
rect 9364 6712 9370 6724
rect 11256 6712 11284 6743
rect 16390 6740 16396 6752
rect 16448 6740 16454 6792
rect 15470 6712 15476 6724
rect 9364 6684 11284 6712
rect 15431 6684 15476 6712
rect 9364 6672 9370 6684
rect 1946 6644 1952 6656
rect 1907 6616 1952 6644
rect 1946 6604 1952 6616
rect 2004 6604 2010 6656
rect 2501 6647 2559 6653
rect 2501 6613 2513 6647
rect 2547 6644 2559 6647
rect 2958 6644 2964 6656
rect 2547 6616 2964 6644
rect 2547 6613 2559 6616
rect 2501 6607 2559 6613
rect 2958 6604 2964 6616
rect 3016 6604 3022 6656
rect 7098 6644 7104 6656
rect 7059 6616 7104 6644
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 7285 6647 7343 6653
rect 7285 6613 7297 6647
rect 7331 6644 7343 6647
rect 7374 6644 7380 6656
rect 7331 6616 7380 6644
rect 7331 6613 7343 6616
rect 7285 6607 7343 6613
rect 7374 6604 7380 6616
rect 7432 6644 7438 6656
rect 8202 6644 8208 6656
rect 7432 6616 8208 6644
rect 7432 6604 7438 6616
rect 8202 6604 8208 6616
rect 8260 6604 8266 6656
rect 9769 6647 9827 6653
rect 9769 6613 9781 6647
rect 9815 6644 9827 6647
rect 10686 6644 10692 6656
rect 9815 6616 10692 6644
rect 9815 6613 9827 6616
rect 9769 6607 9827 6613
rect 10686 6604 10692 6616
rect 10744 6604 10750 6656
rect 11256 6644 11284 6684
rect 15470 6672 15476 6684
rect 15528 6672 15534 6724
rect 17773 6715 17831 6721
rect 17773 6681 17785 6715
rect 17819 6712 17831 6715
rect 18138 6712 18144 6724
rect 17819 6684 18144 6712
rect 17819 6681 17831 6684
rect 17773 6675 17831 6681
rect 18138 6672 18144 6684
rect 18196 6672 18202 6724
rect 11514 6644 11520 6656
rect 11256 6616 11520 6644
rect 11514 6604 11520 6616
rect 11572 6604 11578 6656
rect 12618 6644 12624 6656
rect 12531 6616 12624 6644
rect 12618 6604 12624 6616
rect 12676 6644 12682 6656
rect 13078 6644 13084 6656
rect 12676 6616 13084 6644
rect 12676 6604 12682 6616
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 14274 6644 14280 6656
rect 14235 6616 14280 6644
rect 14274 6604 14280 6616
rect 14332 6604 14338 6656
rect 14642 6644 14648 6656
rect 14603 6616 14648 6644
rect 14642 6604 14648 6616
rect 14700 6604 14706 6656
rect 19613 6647 19671 6653
rect 19613 6613 19625 6647
rect 19659 6644 19671 6647
rect 20622 6644 20628 6656
rect 19659 6616 20628 6644
rect 19659 6613 19671 6616
rect 19613 6607 19671 6613
rect 20622 6604 20628 6616
rect 20680 6604 20686 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 2314 6400 2320 6452
rect 2372 6440 2378 6452
rect 2685 6443 2743 6449
rect 2685 6440 2697 6443
rect 2372 6412 2697 6440
rect 2372 6400 2378 6412
rect 2685 6409 2697 6412
rect 2731 6440 2743 6443
rect 4246 6440 4252 6452
rect 2731 6412 2912 6440
rect 4207 6412 4252 6440
rect 2731 6409 2743 6412
rect 2685 6403 2743 6409
rect 2884 6313 2912 6412
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 5166 6440 5172 6452
rect 5127 6412 5172 6440
rect 5166 6400 5172 6412
rect 5224 6400 5230 6452
rect 5994 6440 6000 6452
rect 5955 6412 6000 6440
rect 5994 6400 6000 6412
rect 6052 6400 6058 6452
rect 9306 6440 9312 6452
rect 7024 6412 9312 6440
rect 2869 6307 2927 6313
rect 2869 6273 2881 6307
rect 2915 6273 2927 6307
rect 2869 6267 2927 6273
rect 1578 6236 1584 6248
rect 1539 6208 1584 6236
rect 1578 6196 1584 6208
rect 1636 6236 1642 6248
rect 2498 6236 2504 6248
rect 1636 6208 2504 6236
rect 1636 6196 1642 6208
rect 2498 6196 2504 6208
rect 2556 6196 2562 6248
rect 5350 6236 5356 6248
rect 5311 6208 5356 6236
rect 5350 6196 5356 6208
rect 5408 6196 5414 6248
rect 7024 6245 7052 6412
rect 9306 6400 9312 6412
rect 9364 6400 9370 6452
rect 11330 6400 11336 6452
rect 11388 6440 11394 6452
rect 11793 6443 11851 6449
rect 11793 6440 11805 6443
rect 11388 6412 11805 6440
rect 11388 6400 11394 6412
rect 11793 6409 11805 6412
rect 11839 6409 11851 6443
rect 11793 6403 11851 6409
rect 12713 6443 12771 6449
rect 12713 6409 12725 6443
rect 12759 6440 12771 6443
rect 12802 6440 12808 6452
rect 12759 6412 12808 6440
rect 12759 6409 12771 6412
rect 12713 6403 12771 6409
rect 12802 6400 12808 6412
rect 12860 6440 12866 6452
rect 13446 6440 13452 6452
rect 12860 6412 13452 6440
rect 12860 6400 12866 6412
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 15197 6443 15255 6449
rect 15197 6409 15209 6443
rect 15243 6440 15255 6443
rect 15378 6440 15384 6452
rect 15243 6412 15384 6440
rect 15243 6409 15255 6412
rect 15197 6403 15255 6409
rect 15378 6400 15384 6412
rect 15436 6400 15442 6452
rect 16390 6400 16396 6452
rect 16448 6440 16454 6452
rect 16669 6443 16727 6449
rect 16669 6440 16681 6443
rect 16448 6412 16681 6440
rect 16448 6400 16454 6412
rect 16669 6409 16681 6412
rect 16715 6409 16727 6443
rect 17770 6440 17776 6452
rect 17731 6412 17776 6440
rect 16669 6403 16727 6409
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 19334 6400 19340 6452
rect 19392 6440 19398 6452
rect 19429 6443 19487 6449
rect 19429 6440 19441 6443
rect 19392 6412 19441 6440
rect 19392 6400 19398 6412
rect 19429 6409 19441 6412
rect 19475 6409 19487 6443
rect 19429 6403 19487 6409
rect 9324 6304 9352 6400
rect 14185 6375 14243 6381
rect 14185 6341 14197 6375
rect 14231 6372 14243 6375
rect 15286 6372 15292 6384
rect 14231 6344 15292 6372
rect 14231 6341 14243 6344
rect 14185 6335 14243 6341
rect 15286 6332 15292 6344
rect 15344 6332 15350 6384
rect 9493 6307 9551 6313
rect 9493 6304 9505 6307
rect 9324 6276 9505 6304
rect 9493 6273 9505 6276
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 12253 6307 12311 6313
rect 12253 6273 12265 6307
rect 12299 6304 12311 6307
rect 15396 6304 15424 6400
rect 15749 6375 15807 6381
rect 15749 6341 15761 6375
rect 15795 6372 15807 6375
rect 17405 6375 17463 6381
rect 17405 6372 17417 6375
rect 15795 6344 17417 6372
rect 15795 6341 15807 6344
rect 15749 6335 15807 6341
rect 17405 6341 17417 6344
rect 17451 6341 17463 6375
rect 18138 6372 18144 6384
rect 18099 6344 18144 6372
rect 17405 6335 17463 6341
rect 16117 6307 16175 6313
rect 16117 6304 16129 6307
rect 12299 6276 12940 6304
rect 15396 6276 16129 6304
rect 12299 6273 12311 6276
rect 12253 6267 12311 6273
rect 7282 6245 7288 6248
rect 7009 6239 7067 6245
rect 7009 6236 7021 6239
rect 6564 6208 7021 6236
rect 1857 6171 1915 6177
rect 1857 6137 1869 6171
rect 1903 6168 1915 6171
rect 2958 6168 2964 6180
rect 1903 6140 2964 6168
rect 1903 6137 1915 6140
rect 1857 6131 1915 6137
rect 2958 6128 2964 6140
rect 3016 6128 3022 6180
rect 3142 6177 3148 6180
rect 3136 6168 3148 6177
rect 3103 6140 3148 6168
rect 3136 6131 3148 6140
rect 3142 6128 3148 6131
rect 3200 6128 3206 6180
rect 2409 6103 2467 6109
rect 2409 6069 2421 6103
rect 2455 6100 2467 6103
rect 3151 6100 3179 6128
rect 6564 6112 6592 6208
rect 7009 6205 7021 6208
rect 7055 6205 7067 6239
rect 7276 6236 7288 6245
rect 7195 6208 7288 6236
rect 7009 6199 7067 6205
rect 7276 6199 7288 6208
rect 7340 6236 7346 6248
rect 8018 6236 8024 6248
rect 7340 6208 8024 6236
rect 7282 6196 7288 6199
rect 7340 6196 7346 6208
rect 8018 6196 8024 6208
rect 8076 6196 8082 6248
rect 9766 6245 9772 6248
rect 9760 6236 9772 6245
rect 9727 6208 9772 6236
rect 9760 6199 9772 6208
rect 9766 6196 9772 6199
rect 9824 6196 9830 6248
rect 11514 6236 11520 6248
rect 11427 6208 11520 6236
rect 11514 6196 11520 6208
rect 11572 6236 11578 6248
rect 12526 6236 12532 6248
rect 11572 6208 12532 6236
rect 11572 6196 11578 6208
rect 12526 6196 12532 6208
rect 12584 6236 12590 6248
rect 12802 6236 12808 6248
rect 12584 6208 12808 6236
rect 12584 6196 12590 6208
rect 12802 6196 12808 6208
rect 12860 6196 12866 6248
rect 12912 6236 12940 6276
rect 16117 6273 16129 6276
rect 16163 6273 16175 6307
rect 16298 6304 16304 6316
rect 16259 6276 16304 6304
rect 16117 6267 16175 6273
rect 16298 6264 16304 6276
rect 16356 6304 16362 6316
rect 17037 6307 17095 6313
rect 17037 6304 17049 6307
rect 16356 6276 17049 6304
rect 16356 6264 16362 6276
rect 17037 6273 17049 6276
rect 17083 6273 17095 6307
rect 17037 6267 17095 6273
rect 13061 6239 13119 6245
rect 13061 6236 13073 6239
rect 12912 6208 13073 6236
rect 13061 6205 13073 6208
rect 13107 6236 13119 6239
rect 13538 6236 13544 6248
rect 13107 6208 13544 6236
rect 13107 6205 13119 6208
rect 13061 6199 13119 6205
rect 13538 6196 13544 6208
rect 13596 6196 13602 6248
rect 17420 6236 17448 6335
rect 18138 6332 18144 6344
rect 18196 6332 18202 6384
rect 25498 6372 25504 6384
rect 25459 6344 25504 6372
rect 25498 6332 25504 6344
rect 25556 6332 25562 6384
rect 18230 6264 18236 6316
rect 18288 6304 18294 6316
rect 18693 6307 18751 6313
rect 18693 6304 18705 6307
rect 18288 6276 18705 6304
rect 18288 6264 18294 6276
rect 18693 6273 18705 6276
rect 18739 6273 18751 6307
rect 18693 6267 18751 6273
rect 24029 6307 24087 6313
rect 24029 6273 24041 6307
rect 24075 6304 24087 6307
rect 24075 6276 24256 6304
rect 24075 6273 24087 6276
rect 24029 6267 24087 6273
rect 17420 6208 18644 6236
rect 17770 6128 17776 6180
rect 17828 6168 17834 6180
rect 18616 6177 18644 6208
rect 19426 6196 19432 6248
rect 19484 6236 19490 6248
rect 19613 6239 19671 6245
rect 19613 6236 19625 6239
rect 19484 6208 19625 6236
rect 19484 6196 19490 6208
rect 19613 6205 19625 6208
rect 19659 6236 19671 6239
rect 20349 6239 20407 6245
rect 20349 6236 20361 6239
rect 19659 6208 20361 6236
rect 19659 6205 19671 6208
rect 19613 6199 19671 6205
rect 20349 6205 20361 6208
rect 20395 6205 20407 6239
rect 24118 6236 24124 6248
rect 24079 6208 24124 6236
rect 20349 6199 20407 6205
rect 24118 6196 24124 6208
rect 24176 6196 24182 6248
rect 24228 6236 24256 6276
rect 24388 6239 24446 6245
rect 24388 6236 24400 6239
rect 24228 6208 24400 6236
rect 24388 6205 24400 6208
rect 24434 6236 24446 6239
rect 24762 6236 24768 6248
rect 24434 6208 24768 6236
rect 24434 6205 24446 6208
rect 24388 6199 24446 6205
rect 24762 6196 24768 6208
rect 24820 6196 24826 6248
rect 18417 6171 18475 6177
rect 18417 6168 18429 6171
rect 17828 6140 18429 6168
rect 17828 6128 17834 6140
rect 18417 6137 18429 6140
rect 18463 6137 18475 6171
rect 18417 6131 18475 6137
rect 18601 6171 18659 6177
rect 18601 6137 18613 6171
rect 18647 6137 18659 6171
rect 18601 6131 18659 6137
rect 19889 6171 19947 6177
rect 19889 6137 19901 6171
rect 19935 6168 19947 6171
rect 20898 6168 20904 6180
rect 19935 6140 20904 6168
rect 19935 6137 19947 6140
rect 19889 6131 19947 6137
rect 20898 6128 20904 6140
rect 20956 6128 20962 6180
rect 2455 6072 3179 6100
rect 2455 6069 2467 6072
rect 2409 6063 2467 6069
rect 4706 6060 4712 6112
rect 4764 6100 4770 6112
rect 4801 6103 4859 6109
rect 4801 6100 4813 6103
rect 4764 6072 4813 6100
rect 4764 6060 4770 6072
rect 4801 6069 4813 6072
rect 4847 6069 4859 6103
rect 4801 6063 4859 6069
rect 5537 6103 5595 6109
rect 5537 6069 5549 6103
rect 5583 6100 5595 6103
rect 5994 6100 6000 6112
rect 5583 6072 6000 6100
rect 5583 6069 5595 6072
rect 5537 6063 5595 6069
rect 5994 6060 6000 6072
rect 6052 6060 6058 6112
rect 6546 6100 6552 6112
rect 6507 6072 6552 6100
rect 6546 6060 6552 6072
rect 6604 6060 6610 6112
rect 8386 6100 8392 6112
rect 8347 6072 8392 6100
rect 8386 6060 8392 6072
rect 8444 6100 8450 6112
rect 8941 6103 8999 6109
rect 8941 6100 8953 6103
rect 8444 6072 8953 6100
rect 8444 6060 8450 6072
rect 8941 6069 8953 6072
rect 8987 6069 8999 6103
rect 10870 6100 10876 6112
rect 10831 6072 10876 6100
rect 8941 6063 8999 6069
rect 10870 6060 10876 6072
rect 10928 6060 10934 6112
rect 14274 6060 14280 6112
rect 14332 6100 14338 6112
rect 14737 6103 14795 6109
rect 14737 6100 14749 6103
rect 14332 6072 14749 6100
rect 14332 6060 14338 6072
rect 14737 6069 14749 6072
rect 14783 6100 14795 6103
rect 14826 6100 14832 6112
rect 14783 6072 14832 6100
rect 14783 6069 14795 6072
rect 14737 6063 14795 6069
rect 14826 6060 14832 6072
rect 14884 6060 14890 6112
rect 15378 6060 15384 6112
rect 15436 6100 15442 6112
rect 15473 6103 15531 6109
rect 15473 6100 15485 6103
rect 15436 6072 15485 6100
rect 15436 6060 15442 6072
rect 15473 6069 15485 6072
rect 15519 6100 15531 6103
rect 16209 6103 16267 6109
rect 16209 6100 16221 6103
rect 15519 6072 16221 6100
rect 15519 6069 15531 6072
rect 15473 6063 15531 6069
rect 16209 6069 16221 6072
rect 16255 6069 16267 6103
rect 16209 6063 16267 6069
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1949 5899 2007 5905
rect 1949 5865 1961 5899
rect 1995 5896 2007 5899
rect 2038 5896 2044 5908
rect 1995 5868 2044 5896
rect 1995 5865 2007 5868
rect 1949 5859 2007 5865
rect 2038 5856 2044 5868
rect 2096 5856 2102 5908
rect 2314 5856 2320 5908
rect 2372 5896 2378 5908
rect 2409 5899 2467 5905
rect 2409 5896 2421 5899
rect 2372 5868 2421 5896
rect 2372 5856 2378 5868
rect 2409 5865 2421 5868
rect 2455 5865 2467 5899
rect 2409 5859 2467 5865
rect 3881 5899 3939 5905
rect 3881 5865 3893 5899
rect 3927 5896 3939 5899
rect 4246 5896 4252 5908
rect 3927 5868 4252 5896
rect 3927 5865 3939 5868
rect 3881 5859 3939 5865
rect 4246 5856 4252 5868
rect 4304 5856 4310 5908
rect 6822 5856 6828 5908
rect 6880 5896 6886 5908
rect 7098 5896 7104 5908
rect 6880 5868 7104 5896
rect 6880 5856 6886 5868
rect 7098 5856 7104 5868
rect 7156 5896 7162 5908
rect 8941 5899 8999 5905
rect 8941 5896 8953 5899
rect 7156 5868 8953 5896
rect 7156 5856 7162 5868
rect 8941 5865 8953 5868
rect 8987 5865 8999 5899
rect 8941 5859 8999 5865
rect 9766 5856 9772 5908
rect 9824 5896 9830 5908
rect 9861 5899 9919 5905
rect 9861 5896 9873 5899
rect 9824 5868 9873 5896
rect 9824 5856 9830 5868
rect 9861 5865 9873 5868
rect 9907 5865 9919 5899
rect 9861 5859 9919 5865
rect 10134 5856 10140 5908
rect 10192 5896 10198 5908
rect 10229 5899 10287 5905
rect 10229 5896 10241 5899
rect 10192 5868 10241 5896
rect 10192 5856 10198 5868
rect 10229 5865 10241 5868
rect 10275 5865 10287 5899
rect 10229 5859 10287 5865
rect 11514 5856 11520 5908
rect 11572 5896 11578 5908
rect 17221 5899 17279 5905
rect 17221 5896 17233 5899
rect 11572 5868 17233 5896
rect 11572 5856 11578 5868
rect 17221 5865 17233 5868
rect 17267 5865 17279 5899
rect 17221 5859 17279 5865
rect 18141 5899 18199 5905
rect 18141 5865 18153 5899
rect 18187 5896 18199 5899
rect 18230 5896 18236 5908
rect 18187 5868 18236 5896
rect 18187 5865 18199 5868
rect 18141 5859 18199 5865
rect 18230 5856 18236 5868
rect 18288 5856 18294 5908
rect 24118 5896 24124 5908
rect 24079 5868 24124 5896
rect 24118 5856 24124 5868
rect 24176 5856 24182 5908
rect 1394 5788 1400 5840
rect 1452 5828 1458 5840
rect 1765 5831 1823 5837
rect 1765 5828 1777 5831
rect 1452 5800 1777 5828
rect 1452 5788 1458 5800
rect 1765 5797 1777 5800
rect 1811 5828 1823 5831
rect 2777 5831 2835 5837
rect 2777 5828 2789 5831
rect 1811 5800 2789 5828
rect 1811 5797 1823 5800
rect 1765 5791 1823 5797
rect 2777 5797 2789 5800
rect 2823 5797 2835 5831
rect 2958 5828 2964 5840
rect 2919 5800 2964 5828
rect 2777 5791 2835 5797
rect 2958 5788 2964 5800
rect 3016 5788 3022 5840
rect 7006 5828 7012 5840
rect 3151 5800 7012 5828
rect 1302 5720 1308 5772
rect 1360 5760 1366 5772
rect 3151 5760 3179 5800
rect 7006 5788 7012 5800
rect 7064 5788 7070 5840
rect 7558 5828 7564 5840
rect 7519 5800 7564 5828
rect 7558 5788 7564 5800
rect 7616 5788 7622 5840
rect 7650 5788 7656 5840
rect 7708 5828 7714 5840
rect 7745 5831 7803 5837
rect 7745 5828 7757 5831
rect 7708 5800 7757 5828
rect 7708 5788 7714 5800
rect 7745 5797 7757 5800
rect 7791 5797 7803 5831
rect 10680 5831 10738 5837
rect 7745 5791 7803 5797
rect 10060 5800 10548 5828
rect 10060 5772 10088 5800
rect 1360 5732 3179 5760
rect 1360 5720 1366 5732
rect 4154 5720 4160 5772
rect 4212 5760 4218 5772
rect 4965 5763 5023 5769
rect 4965 5760 4977 5763
rect 4212 5732 4977 5760
rect 4212 5720 4218 5732
rect 4965 5729 4977 5732
rect 5011 5760 5023 5763
rect 5442 5760 5448 5772
rect 5011 5732 5448 5760
rect 5011 5729 5023 5732
rect 4965 5723 5023 5729
rect 5442 5720 5448 5732
rect 5500 5720 5506 5772
rect 6730 5720 6736 5772
rect 6788 5760 6794 5772
rect 7837 5763 7895 5769
rect 7837 5760 7849 5763
rect 6788 5732 7849 5760
rect 6788 5720 6794 5732
rect 7837 5729 7849 5732
rect 7883 5760 7895 5763
rect 8386 5760 8392 5772
rect 7883 5732 8392 5760
rect 7883 5729 7895 5732
rect 7837 5723 7895 5729
rect 8386 5720 8392 5732
rect 8444 5720 8450 5772
rect 9306 5720 9312 5772
rect 9364 5760 9370 5772
rect 10042 5760 10048 5772
rect 9364 5732 10048 5760
rect 9364 5720 9370 5732
rect 10042 5720 10048 5732
rect 10100 5720 10106 5772
rect 10420 5763 10478 5769
rect 10420 5729 10432 5763
rect 10466 5760 10478 5763
rect 10520 5760 10548 5800
rect 10680 5797 10692 5831
rect 10726 5828 10738 5831
rect 10870 5828 10876 5840
rect 10726 5800 10876 5828
rect 10726 5797 10738 5800
rect 10680 5791 10738 5797
rect 10870 5788 10876 5800
rect 10928 5828 10934 5840
rect 11054 5828 11060 5840
rect 10928 5800 11060 5828
rect 10928 5788 10934 5800
rect 11054 5788 11060 5800
rect 11112 5788 11118 5840
rect 12066 5788 12072 5840
rect 12124 5828 12130 5840
rect 13449 5831 13507 5837
rect 13449 5828 13461 5831
rect 12124 5800 13461 5828
rect 12124 5788 12130 5800
rect 13449 5797 13461 5800
rect 13495 5797 13507 5831
rect 13449 5791 13507 5797
rect 13538 5788 13544 5840
rect 13596 5828 13602 5840
rect 13814 5828 13820 5840
rect 13596 5800 13820 5828
rect 13596 5788 13602 5800
rect 13814 5788 13820 5800
rect 13872 5828 13878 5840
rect 14277 5831 14335 5837
rect 14277 5828 14289 5831
rect 13872 5800 14289 5828
rect 13872 5788 13878 5800
rect 14277 5797 14289 5800
rect 14323 5797 14335 5831
rect 14277 5791 14335 5797
rect 15286 5788 15292 5840
rect 15344 5828 15350 5840
rect 15534 5831 15592 5837
rect 15534 5828 15546 5831
rect 15344 5800 15546 5828
rect 15344 5788 15350 5800
rect 15534 5797 15546 5800
rect 15580 5797 15592 5831
rect 15534 5791 15592 5797
rect 13262 5760 13268 5772
rect 10466 5732 10548 5760
rect 13223 5732 13268 5760
rect 10466 5729 10478 5732
rect 10420 5723 10478 5729
rect 13262 5720 13268 5732
rect 13320 5760 13326 5772
rect 13906 5760 13912 5772
rect 13320 5732 13912 5760
rect 13320 5720 13326 5732
rect 13906 5720 13912 5732
rect 13964 5720 13970 5772
rect 15930 5760 15936 5772
rect 15304 5732 15936 5760
rect 1946 5652 1952 5704
rect 2004 5692 2010 5704
rect 2041 5695 2099 5701
rect 2041 5692 2053 5695
rect 2004 5664 2053 5692
rect 2004 5652 2010 5664
rect 2041 5661 2053 5664
rect 2087 5692 2099 5695
rect 2087 5664 2912 5692
rect 2087 5661 2099 5664
rect 2041 5655 2099 5661
rect 1489 5627 1547 5633
rect 1489 5593 1501 5627
rect 1535 5624 1547 5627
rect 2682 5624 2688 5636
rect 1535 5596 2688 5624
rect 1535 5593 1547 5596
rect 1489 5587 1547 5593
rect 2682 5584 2688 5596
rect 2740 5584 2746 5636
rect 2884 5624 2912 5664
rect 4246 5652 4252 5704
rect 4304 5692 4310 5704
rect 4709 5695 4767 5701
rect 4709 5692 4721 5695
rect 4304 5664 4721 5692
rect 4304 5652 4310 5664
rect 4709 5661 4721 5664
rect 4755 5661 4767 5695
rect 4709 5655 4767 5661
rect 7101 5695 7159 5701
rect 7101 5661 7113 5695
rect 7147 5692 7159 5695
rect 7190 5692 7196 5704
rect 7147 5664 7196 5692
rect 7147 5661 7159 5664
rect 7101 5655 7159 5661
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 14826 5652 14832 5704
rect 14884 5692 14890 5704
rect 15304 5701 15332 5732
rect 15930 5720 15936 5732
rect 15988 5760 15994 5772
rect 16390 5760 16396 5772
rect 15988 5732 16396 5760
rect 15988 5720 15994 5732
rect 16390 5720 16396 5732
rect 16448 5720 16454 5772
rect 18138 5720 18144 5772
rect 18196 5760 18202 5772
rect 18509 5763 18567 5769
rect 18509 5760 18521 5763
rect 18196 5732 18521 5760
rect 18196 5720 18202 5732
rect 18509 5729 18521 5732
rect 18555 5760 18567 5763
rect 18966 5760 18972 5772
rect 18555 5732 18972 5760
rect 18555 5729 18567 5732
rect 18509 5723 18567 5729
rect 18966 5720 18972 5732
rect 19024 5720 19030 5772
rect 20898 5760 20904 5772
rect 20859 5732 20904 5760
rect 20898 5720 20904 5732
rect 20956 5720 20962 5772
rect 15289 5695 15347 5701
rect 15289 5692 15301 5695
rect 14884 5664 15301 5692
rect 14884 5652 14890 5664
rect 15289 5661 15301 5664
rect 15335 5661 15347 5695
rect 17586 5692 17592 5704
rect 17547 5664 17592 5692
rect 15289 5655 15347 5661
rect 17586 5652 17592 5664
rect 17644 5652 17650 5704
rect 18782 5692 18788 5704
rect 18743 5664 18788 5692
rect 18782 5652 18788 5664
rect 18840 5652 18846 5704
rect 19794 5692 19800 5704
rect 19755 5664 19800 5692
rect 19794 5652 19800 5664
rect 19852 5652 19858 5704
rect 3513 5627 3571 5633
rect 3513 5624 3525 5627
rect 2884 5596 3525 5624
rect 3513 5593 3525 5596
rect 3559 5624 3571 5627
rect 4062 5624 4068 5636
rect 3559 5596 4068 5624
rect 3559 5593 3571 5596
rect 3513 5587 3571 5593
rect 4062 5584 4068 5596
rect 4120 5584 4126 5636
rect 6914 5584 6920 5636
rect 6972 5624 6978 5636
rect 7285 5627 7343 5633
rect 7285 5624 7297 5627
rect 6972 5596 7297 5624
rect 6972 5584 6978 5596
rect 7285 5593 7297 5596
rect 7331 5593 7343 5627
rect 7285 5587 7343 5593
rect 11974 5584 11980 5636
rect 12032 5624 12038 5636
rect 13722 5624 13728 5636
rect 12032 5596 13728 5624
rect 12032 5584 12038 5596
rect 13722 5584 13728 5596
rect 13780 5624 13786 5636
rect 13909 5627 13967 5633
rect 13909 5624 13921 5627
rect 13780 5596 13921 5624
rect 13780 5584 13786 5596
rect 13909 5593 13921 5596
rect 13955 5593 13967 5627
rect 13909 5587 13967 5593
rect 3878 5516 3884 5568
rect 3936 5556 3942 5568
rect 4249 5559 4307 5565
rect 4249 5556 4261 5559
rect 3936 5528 4261 5556
rect 3936 5516 3942 5528
rect 4249 5525 4261 5528
rect 4295 5556 4307 5559
rect 4430 5556 4436 5568
rect 4295 5528 4436 5556
rect 4295 5525 4307 5528
rect 4249 5519 4307 5525
rect 4430 5516 4436 5528
rect 4488 5516 4494 5568
rect 5350 5516 5356 5568
rect 5408 5556 5414 5568
rect 6089 5559 6147 5565
rect 6089 5556 6101 5559
rect 5408 5528 6101 5556
rect 5408 5516 5414 5528
rect 6089 5525 6101 5528
rect 6135 5525 6147 5559
rect 6730 5556 6736 5568
rect 6691 5528 6736 5556
rect 6089 5519 6147 5525
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 8297 5559 8355 5565
rect 8297 5525 8309 5559
rect 8343 5556 8355 5559
rect 8478 5556 8484 5568
rect 8343 5528 8484 5556
rect 8343 5525 8355 5528
rect 8297 5519 8355 5525
rect 8478 5516 8484 5528
rect 8536 5556 8542 5568
rect 8573 5559 8631 5565
rect 8573 5556 8585 5559
rect 8536 5528 8585 5556
rect 8536 5516 8542 5528
rect 8573 5525 8585 5528
rect 8619 5525 8631 5559
rect 9398 5556 9404 5568
rect 9359 5528 9404 5556
rect 8573 5519 8631 5525
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 11146 5516 11152 5568
rect 11204 5556 11210 5568
rect 11793 5559 11851 5565
rect 11793 5556 11805 5559
rect 11204 5528 11805 5556
rect 11204 5516 11210 5528
rect 11793 5525 11805 5528
rect 11839 5556 11851 5559
rect 12437 5559 12495 5565
rect 12437 5556 12449 5559
rect 11839 5528 12449 5556
rect 11839 5525 11851 5528
rect 11793 5519 11851 5525
rect 12437 5525 12449 5528
rect 12483 5556 12495 5559
rect 12618 5556 12624 5568
rect 12483 5528 12624 5556
rect 12483 5525 12495 5528
rect 12437 5519 12495 5525
rect 12618 5516 12624 5528
rect 12676 5516 12682 5568
rect 12989 5559 13047 5565
rect 12989 5525 13001 5559
rect 13035 5556 13047 5559
rect 13446 5556 13452 5568
rect 13035 5528 13452 5556
rect 13035 5525 13047 5528
rect 12989 5519 13047 5525
rect 13446 5516 13452 5528
rect 13504 5516 13510 5568
rect 15013 5559 15071 5565
rect 15013 5525 15025 5559
rect 15059 5556 15071 5559
rect 15470 5556 15476 5568
rect 15059 5528 15476 5556
rect 15059 5525 15071 5528
rect 15013 5519 15071 5525
rect 15470 5516 15476 5528
rect 15528 5556 15534 5568
rect 16669 5559 16727 5565
rect 16669 5556 16681 5559
rect 15528 5528 16681 5556
rect 15528 5516 15534 5528
rect 16669 5525 16681 5528
rect 16715 5525 16727 5559
rect 21082 5556 21088 5568
rect 21043 5528 21088 5556
rect 16669 5519 16727 5525
rect 21082 5516 21088 5528
rect 21140 5516 21146 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 1673 5355 1731 5361
rect 1673 5321 1685 5355
rect 1719 5352 1731 5355
rect 2038 5352 2044 5364
rect 1719 5324 2044 5352
rect 1719 5321 1731 5324
rect 1673 5315 1731 5321
rect 2038 5312 2044 5324
rect 2096 5312 2102 5364
rect 3142 5312 3148 5364
rect 3200 5352 3206 5364
rect 3237 5355 3295 5361
rect 3237 5352 3249 5355
rect 3200 5324 3249 5352
rect 3200 5312 3206 5324
rect 3237 5321 3249 5324
rect 3283 5321 3295 5355
rect 3237 5315 3295 5321
rect 3973 5355 4031 5361
rect 3973 5321 3985 5355
rect 4019 5352 4031 5355
rect 4154 5352 4160 5364
rect 4019 5324 4160 5352
rect 4019 5321 4031 5324
rect 3973 5315 4031 5321
rect 4154 5312 4160 5324
rect 4212 5312 4218 5364
rect 4614 5352 4620 5364
rect 4575 5324 4620 5352
rect 4614 5312 4620 5324
rect 4672 5352 4678 5364
rect 6273 5355 6331 5361
rect 6273 5352 6285 5355
rect 4672 5324 5672 5352
rect 4672 5312 4678 5324
rect 4338 5244 4344 5296
rect 4396 5284 4402 5296
rect 4985 5287 5043 5293
rect 4985 5284 4997 5287
rect 4396 5256 4997 5284
rect 4396 5244 4402 5256
rect 4985 5253 4997 5256
rect 5031 5253 5043 5287
rect 5258 5284 5264 5296
rect 5219 5256 5264 5284
rect 4985 5247 5043 5253
rect 1857 5151 1915 5157
rect 1857 5117 1869 5151
rect 1903 5148 1915 5151
rect 1903 5120 2360 5148
rect 1903 5117 1915 5120
rect 1857 5111 1915 5117
rect 2332 5092 2360 5120
rect 2038 5040 2044 5092
rect 2096 5089 2102 5092
rect 2096 5083 2160 5089
rect 2096 5049 2114 5083
rect 2148 5049 2160 5083
rect 2096 5043 2160 5049
rect 2096 5040 2102 5043
rect 2314 5040 2320 5092
rect 2372 5080 2378 5092
rect 4154 5080 4160 5092
rect 2372 5052 4160 5080
rect 2372 5040 2378 5052
rect 4154 5040 4160 5052
rect 4212 5080 4218 5092
rect 4249 5083 4307 5089
rect 4249 5080 4261 5083
rect 4212 5052 4261 5080
rect 4212 5040 4218 5052
rect 4249 5049 4261 5052
rect 4295 5049 4307 5083
rect 5000 5080 5028 5247
rect 5258 5244 5264 5256
rect 5316 5244 5322 5296
rect 5644 5225 5672 5324
rect 5828 5324 6285 5352
rect 5828 5225 5856 5324
rect 6273 5321 6285 5324
rect 6319 5352 6331 5355
rect 7282 5352 7288 5364
rect 6319 5324 7288 5352
rect 6319 5321 6331 5324
rect 6273 5315 6331 5321
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 10042 5312 10048 5364
rect 10100 5352 10106 5364
rect 10597 5355 10655 5361
rect 10597 5352 10609 5355
rect 10100 5324 10609 5352
rect 10100 5312 10106 5324
rect 10597 5321 10609 5324
rect 10643 5321 10655 5355
rect 10597 5315 10655 5321
rect 10778 5312 10784 5364
rect 10836 5312 10842 5364
rect 11054 5352 11060 5364
rect 11015 5324 11060 5352
rect 11054 5312 11060 5324
rect 11112 5352 11118 5364
rect 11701 5355 11759 5361
rect 11701 5352 11713 5355
rect 11112 5324 11713 5352
rect 11112 5312 11118 5324
rect 11701 5321 11713 5324
rect 11747 5352 11759 5355
rect 11882 5352 11888 5364
rect 11747 5324 11888 5352
rect 11747 5321 11759 5324
rect 11701 5315 11759 5321
rect 11882 5312 11888 5324
rect 11940 5312 11946 5364
rect 13814 5352 13820 5364
rect 13775 5324 13820 5352
rect 13814 5312 13820 5324
rect 13872 5312 13878 5364
rect 13906 5312 13912 5364
rect 13964 5352 13970 5364
rect 14369 5355 14427 5361
rect 14369 5352 14381 5355
rect 13964 5324 14381 5352
rect 13964 5312 13970 5324
rect 14369 5321 14381 5324
rect 14415 5321 14427 5355
rect 14826 5352 14832 5364
rect 14787 5324 14832 5352
rect 14369 5315 14427 5321
rect 14826 5312 14832 5324
rect 14884 5312 14890 5364
rect 16390 5312 16396 5364
rect 16448 5352 16454 5364
rect 16853 5355 16911 5361
rect 16853 5352 16865 5355
rect 16448 5324 16865 5352
rect 16448 5312 16454 5324
rect 16853 5321 16865 5324
rect 16899 5321 16911 5355
rect 18966 5352 18972 5364
rect 18927 5324 18972 5352
rect 16853 5315 16911 5321
rect 18966 5312 18972 5324
rect 19024 5312 19030 5364
rect 20898 5312 20904 5364
rect 20956 5352 20962 5364
rect 21177 5355 21235 5361
rect 21177 5352 21189 5355
rect 20956 5324 21189 5352
rect 20956 5312 20962 5324
rect 21177 5321 21189 5324
rect 21223 5321 21235 5355
rect 21177 5315 21235 5321
rect 9674 5284 9680 5296
rect 9635 5256 9680 5284
rect 9674 5244 9680 5256
rect 9732 5244 9738 5296
rect 5629 5219 5687 5225
rect 5629 5185 5641 5219
rect 5675 5185 5687 5219
rect 5629 5179 5687 5185
rect 5813 5219 5871 5225
rect 5813 5185 5825 5219
rect 5859 5185 5871 5219
rect 5813 5179 5871 5185
rect 6546 5176 6552 5228
rect 6604 5216 6610 5228
rect 7101 5219 7159 5225
rect 7101 5216 7113 5219
rect 6604 5188 7113 5216
rect 6604 5176 6610 5188
rect 7101 5185 7113 5188
rect 7147 5185 7159 5219
rect 7101 5179 7159 5185
rect 10796 5160 10824 5312
rect 11514 5176 11520 5228
rect 11572 5176 11578 5228
rect 14844 5216 14872 5312
rect 14921 5219 14979 5225
rect 14921 5216 14933 5219
rect 14844 5188 14933 5216
rect 14921 5185 14933 5188
rect 14967 5185 14979 5219
rect 14921 5179 14979 5185
rect 9493 5151 9551 5157
rect 9493 5117 9505 5151
rect 9539 5148 9551 5151
rect 10229 5151 10287 5157
rect 10229 5148 10241 5151
rect 9539 5120 10241 5148
rect 9539 5117 9551 5120
rect 9493 5111 9551 5117
rect 10229 5117 10241 5120
rect 10275 5148 10287 5151
rect 10686 5148 10692 5160
rect 10275 5120 10692 5148
rect 10275 5117 10287 5120
rect 10229 5111 10287 5117
rect 10686 5108 10692 5120
rect 10744 5108 10750 5160
rect 10778 5108 10784 5160
rect 10836 5108 10842 5160
rect 11149 5151 11207 5157
rect 11149 5117 11161 5151
rect 11195 5148 11207 5151
rect 11238 5148 11244 5160
rect 11195 5120 11244 5148
rect 11195 5117 11207 5120
rect 11149 5111 11207 5117
rect 11238 5108 11244 5120
rect 11296 5108 11302 5160
rect 5721 5083 5779 5089
rect 5721 5080 5733 5083
rect 5000 5052 5733 5080
rect 4249 5043 4307 5049
rect 5721 5049 5733 5052
rect 5767 5049 5779 5083
rect 5721 5043 5779 5049
rect 4264 5012 4292 5043
rect 6730 5040 6736 5092
rect 6788 5080 6794 5092
rect 7346 5083 7404 5089
rect 7346 5080 7358 5083
rect 6788 5052 7358 5080
rect 6788 5040 6794 5052
rect 7346 5049 7358 5052
rect 7392 5049 7404 5083
rect 9953 5083 10011 5089
rect 9953 5080 9965 5083
rect 7346 5043 7404 5049
rect 9048 5052 9965 5080
rect 9048 5024 9076 5052
rect 9953 5049 9965 5052
rect 9999 5049 10011 5083
rect 10134 5080 10140 5092
rect 10047 5052 10140 5080
rect 9953 5043 10011 5049
rect 10134 5040 10140 5052
rect 10192 5080 10198 5092
rect 11532 5080 11560 5176
rect 12342 5108 12348 5160
rect 12400 5148 12406 5160
rect 12437 5151 12495 5157
rect 12437 5148 12449 5151
rect 12400 5120 12449 5148
rect 12400 5108 12406 5120
rect 12437 5117 12449 5120
rect 12483 5117 12495 5151
rect 12693 5151 12751 5157
rect 12693 5148 12705 5151
rect 12437 5111 12495 5117
rect 12636 5120 12705 5148
rect 10192 5052 11560 5080
rect 10192 5040 10198 5052
rect 12636 5024 12664 5120
rect 12693 5117 12705 5120
rect 12739 5117 12751 5151
rect 12693 5111 12751 5117
rect 15188 5151 15246 5157
rect 15188 5117 15200 5151
rect 15234 5148 15246 5151
rect 15470 5148 15476 5160
rect 15234 5120 15476 5148
rect 15234 5117 15246 5120
rect 15188 5111 15246 5117
rect 15470 5108 15476 5120
rect 15528 5108 15534 5160
rect 17586 5148 17592 5160
rect 17547 5120 17592 5148
rect 17586 5108 17592 5120
rect 17644 5108 17650 5160
rect 18049 5151 18107 5157
rect 18049 5117 18061 5151
rect 18095 5148 18107 5151
rect 18322 5148 18328 5160
rect 18095 5120 18328 5148
rect 18095 5117 18107 5120
rect 18049 5111 18107 5117
rect 18322 5108 18328 5120
rect 18380 5148 18386 5160
rect 18601 5151 18659 5157
rect 18601 5148 18613 5151
rect 18380 5120 18613 5148
rect 18380 5108 18386 5120
rect 18601 5117 18613 5120
rect 18647 5117 18659 5151
rect 18601 5111 18659 5117
rect 18690 5108 18696 5160
rect 18748 5148 18754 5160
rect 19153 5151 19211 5157
rect 19153 5148 19165 5151
rect 18748 5120 19165 5148
rect 18748 5108 18754 5120
rect 19153 5117 19165 5120
rect 19199 5148 19211 5151
rect 19705 5151 19763 5157
rect 19705 5148 19717 5151
rect 19199 5120 19717 5148
rect 19199 5117 19211 5120
rect 19153 5111 19211 5117
rect 19705 5117 19717 5120
rect 19751 5117 19763 5151
rect 20254 5148 20260 5160
rect 20215 5120 20260 5148
rect 19705 5111 19763 5117
rect 20254 5108 20260 5120
rect 20312 5148 20318 5160
rect 20809 5151 20867 5157
rect 20809 5148 20821 5151
rect 20312 5120 20821 5148
rect 20312 5108 20318 5120
rect 20809 5117 20821 5120
rect 20855 5117 20867 5151
rect 21358 5148 21364 5160
rect 21319 5120 21364 5148
rect 20809 5111 20867 5117
rect 21358 5108 21364 5120
rect 21416 5148 21422 5160
rect 21913 5151 21971 5157
rect 21913 5148 21925 5151
rect 21416 5120 21925 5148
rect 21416 5108 21422 5120
rect 21913 5117 21925 5120
rect 21959 5117 21971 5151
rect 21913 5111 21971 5117
rect 22094 5108 22100 5160
rect 22152 5148 22158 5160
rect 22465 5151 22523 5157
rect 22465 5148 22477 5151
rect 22152 5120 22477 5148
rect 22152 5108 22158 5120
rect 22465 5117 22477 5120
rect 22511 5148 22523 5151
rect 23017 5151 23075 5157
rect 23017 5148 23029 5151
rect 22511 5120 23029 5148
rect 22511 5117 22523 5120
rect 22465 5111 22523 5117
rect 23017 5117 23029 5120
rect 23063 5117 23075 5151
rect 23017 5111 23075 5117
rect 22002 5080 22008 5092
rect 21560 5052 22008 5080
rect 6546 5012 6552 5024
rect 4264 4984 6552 5012
rect 6546 4972 6552 4984
rect 6604 4972 6610 5024
rect 7466 4972 7472 5024
rect 7524 5012 7530 5024
rect 8481 5015 8539 5021
rect 8481 5012 8493 5015
rect 7524 4984 8493 5012
rect 7524 4972 7530 4984
rect 8481 4981 8493 4984
rect 8527 4981 8539 5015
rect 9030 5012 9036 5024
rect 8991 4984 9036 5012
rect 8481 4975 8539 4981
rect 9030 4972 9036 4984
rect 9088 4972 9094 5024
rect 11333 5015 11391 5021
rect 11333 4981 11345 5015
rect 11379 5012 11391 5015
rect 11422 5012 11428 5024
rect 11379 4984 11428 5012
rect 11379 4981 11391 4984
rect 11333 4975 11391 4981
rect 11422 4972 11428 4984
rect 11480 4972 11486 5024
rect 12066 4972 12072 5024
rect 12124 5012 12130 5024
rect 12161 5015 12219 5021
rect 12161 5012 12173 5015
rect 12124 4984 12173 5012
rect 12124 4972 12130 4984
rect 12161 4981 12173 4984
rect 12207 4981 12219 5015
rect 12161 4975 12219 4981
rect 12618 4972 12624 5024
rect 12676 4972 12682 5024
rect 16206 4972 16212 5024
rect 16264 5012 16270 5024
rect 16301 5015 16359 5021
rect 16301 5012 16313 5015
rect 16264 4984 16313 5012
rect 16264 4972 16270 4984
rect 16301 4981 16313 4984
rect 16347 4981 16359 5015
rect 17218 5012 17224 5024
rect 17179 4984 17224 5012
rect 16301 4975 16359 4981
rect 17218 4972 17224 4984
rect 17276 4972 17282 5024
rect 18230 5012 18236 5024
rect 18191 4984 18236 5012
rect 18230 4972 18236 4984
rect 18288 4972 18294 5024
rect 19242 4972 19248 5024
rect 19300 5012 19306 5024
rect 19337 5015 19395 5021
rect 19337 5012 19349 5015
rect 19300 4984 19349 5012
rect 19300 4972 19306 4984
rect 19337 4981 19349 4984
rect 19383 4981 19395 5015
rect 19337 4975 19395 4981
rect 20070 4972 20076 5024
rect 20128 5012 20134 5024
rect 21560 5021 21588 5052
rect 22002 5040 22008 5052
rect 22060 5040 22066 5092
rect 20441 5015 20499 5021
rect 20441 5012 20453 5015
rect 20128 4984 20453 5012
rect 20128 4972 20134 4984
rect 20441 4981 20453 4984
rect 20487 4981 20499 5015
rect 20441 4975 20499 4981
rect 21545 5015 21603 5021
rect 21545 4981 21557 5015
rect 21591 4981 21603 5015
rect 21545 4975 21603 4981
rect 22649 5015 22707 5021
rect 22649 4981 22661 5015
rect 22695 5012 22707 5015
rect 23566 5012 23572 5024
rect 22695 4984 23572 5012
rect 22695 4981 22707 4984
rect 22649 4975 22707 4981
rect 23566 4972 23572 4984
rect 23624 4972 23630 5024
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1394 4808 1400 4820
rect 1355 4780 1400 4808
rect 1394 4768 1400 4780
rect 1452 4768 1458 4820
rect 3786 4808 3792 4820
rect 3747 4780 3792 4808
rect 3786 4768 3792 4780
rect 3844 4768 3850 4820
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 5445 4811 5503 4817
rect 5445 4808 5457 4811
rect 4120 4780 5457 4808
rect 4120 4768 4126 4780
rect 5445 4777 5457 4780
rect 5491 4777 5503 4811
rect 6730 4808 6736 4820
rect 6691 4780 6736 4808
rect 5445 4771 5503 4777
rect 6730 4768 6736 4780
rect 6788 4768 6794 4820
rect 7374 4808 7380 4820
rect 7335 4780 7380 4808
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 7558 4768 7564 4820
rect 7616 4808 7622 4820
rect 7837 4811 7895 4817
rect 7837 4808 7849 4811
rect 7616 4780 7849 4808
rect 7616 4768 7622 4780
rect 7837 4777 7849 4780
rect 7883 4777 7895 4811
rect 8570 4808 8576 4820
rect 8531 4780 8576 4808
rect 7837 4771 7895 4777
rect 8570 4768 8576 4780
rect 8628 4768 8634 4820
rect 9490 4768 9496 4820
rect 9548 4808 9554 4820
rect 9858 4808 9864 4820
rect 9548 4780 9864 4808
rect 9548 4768 9554 4780
rect 9858 4768 9864 4780
rect 9916 4768 9922 4820
rect 10873 4811 10931 4817
rect 10873 4777 10885 4811
rect 10919 4808 10931 4811
rect 11146 4808 11152 4820
rect 10919 4780 11152 4808
rect 10919 4777 10931 4780
rect 10873 4771 10931 4777
rect 11146 4768 11152 4780
rect 11204 4768 11210 4820
rect 11698 4768 11704 4820
rect 11756 4808 11762 4820
rect 11793 4811 11851 4817
rect 11793 4808 11805 4811
rect 11756 4780 11805 4808
rect 11756 4768 11762 4780
rect 11793 4777 11805 4780
rect 11839 4777 11851 4811
rect 12526 4808 12532 4820
rect 12487 4780 12532 4808
rect 11793 4771 11851 4777
rect 12526 4768 12532 4780
rect 12584 4768 12590 4820
rect 14369 4811 14427 4817
rect 14369 4808 14381 4811
rect 13556 4780 14381 4808
rect 2961 4743 3019 4749
rect 2961 4709 2973 4743
rect 3007 4740 3019 4743
rect 3050 4740 3056 4752
rect 3007 4712 3056 4740
rect 3007 4709 3019 4712
rect 2961 4703 3019 4709
rect 3050 4700 3056 4712
rect 3108 4700 3114 4752
rect 3513 4743 3571 4749
rect 3513 4709 3525 4743
rect 3559 4740 3571 4743
rect 4332 4743 4390 4749
rect 4332 4740 4344 4743
rect 3559 4712 4344 4740
rect 3559 4709 3571 4712
rect 3513 4703 3571 4709
rect 4332 4709 4344 4712
rect 4378 4740 4390 4743
rect 5350 4740 5356 4752
rect 4378 4712 5356 4740
rect 4378 4709 4390 4712
rect 4332 4703 4390 4709
rect 2866 4604 2872 4616
rect 2827 4576 2872 4604
rect 2866 4564 2872 4576
rect 2924 4564 2930 4616
rect 2958 4564 2964 4616
rect 3016 4604 3022 4616
rect 3053 4607 3111 4613
rect 3053 4604 3065 4607
rect 3016 4576 3065 4604
rect 3016 4564 3022 4576
rect 3053 4573 3065 4576
rect 3099 4604 3111 4607
rect 3528 4604 3556 4703
rect 5350 4700 5356 4712
rect 5408 4700 5414 4752
rect 6914 4700 6920 4752
rect 6972 4740 6978 4752
rect 7193 4743 7251 4749
rect 7193 4740 7205 4743
rect 6972 4712 7205 4740
rect 6972 4700 6978 4712
rect 7193 4709 7205 4712
rect 7239 4709 7251 4743
rect 7466 4740 7472 4752
rect 7427 4712 7472 4740
rect 7193 4703 7251 4709
rect 7466 4700 7472 4712
rect 7524 4700 7530 4752
rect 10226 4740 10232 4752
rect 10187 4712 10232 4740
rect 10226 4700 10232 4712
rect 10284 4700 10290 4752
rect 11330 4700 11336 4752
rect 11388 4740 11394 4752
rect 11609 4743 11667 4749
rect 11609 4740 11621 4743
rect 11388 4712 11621 4740
rect 11388 4700 11394 4712
rect 11609 4709 11621 4712
rect 11655 4709 11667 4743
rect 11609 4703 11667 4709
rect 11882 4700 11888 4752
rect 11940 4740 11946 4752
rect 13446 4740 13452 4752
rect 11940 4712 11985 4740
rect 13407 4712 13452 4740
rect 11940 4700 11946 4712
rect 13446 4700 13452 4712
rect 13504 4700 13510 4752
rect 13556 4749 13584 4780
rect 14369 4777 14381 4780
rect 14415 4808 14427 4811
rect 15102 4808 15108 4820
rect 14415 4780 15108 4808
rect 14415 4777 14427 4780
rect 14369 4771 14427 4777
rect 15102 4768 15108 4780
rect 15160 4768 15166 4820
rect 15746 4808 15752 4820
rect 15707 4780 15752 4808
rect 15746 4768 15752 4780
rect 15804 4768 15810 4820
rect 15838 4768 15844 4820
rect 15896 4808 15902 4820
rect 17862 4808 17868 4820
rect 15896 4780 17868 4808
rect 15896 4768 15902 4780
rect 17862 4768 17868 4780
rect 17920 4768 17926 4820
rect 13541 4743 13599 4749
rect 13541 4709 13553 4743
rect 13587 4709 13599 4743
rect 18230 4740 18236 4752
rect 18191 4712 18236 4740
rect 13541 4703 13599 4709
rect 18230 4700 18236 4712
rect 18288 4700 18294 4752
rect 18598 4700 18604 4752
rect 18656 4740 18662 4752
rect 18969 4743 19027 4749
rect 18969 4740 18981 4743
rect 18656 4712 18981 4740
rect 18656 4700 18662 4712
rect 18969 4709 18981 4712
rect 19015 4709 19027 4743
rect 18969 4703 19027 4709
rect 4065 4675 4123 4681
rect 4065 4641 4077 4675
rect 4111 4672 4123 4675
rect 4154 4672 4160 4684
rect 4111 4644 4160 4672
rect 4111 4641 4123 4644
rect 4065 4635 4123 4641
rect 4154 4632 4160 4644
rect 4212 4632 4218 4684
rect 8386 4672 8392 4684
rect 8347 4644 8392 4672
rect 8386 4632 8392 4644
rect 8444 4632 8450 4684
rect 10045 4675 10103 4681
rect 10045 4641 10057 4675
rect 10091 4672 10103 4675
rect 10410 4672 10416 4684
rect 10091 4644 10416 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 10410 4632 10416 4644
rect 10468 4632 10474 4684
rect 15930 4672 15936 4684
rect 15891 4644 15936 4672
rect 15930 4632 15936 4644
rect 15988 4632 15994 4684
rect 16206 4681 16212 4684
rect 16200 4672 16212 4681
rect 16119 4644 16212 4672
rect 16200 4635 16212 4644
rect 16264 4672 16270 4684
rect 20901 4675 20959 4681
rect 16264 4644 19104 4672
rect 16206 4632 16212 4635
rect 16264 4632 16270 4644
rect 19076 4616 19104 4644
rect 20901 4641 20913 4675
rect 20947 4672 20959 4675
rect 20990 4672 20996 4684
rect 20947 4644 20996 4672
rect 20947 4641 20959 4644
rect 20901 4635 20959 4641
rect 20990 4632 20996 4644
rect 21048 4632 21054 4684
rect 22462 4672 22468 4684
rect 22423 4644 22468 4672
rect 22462 4632 22468 4644
rect 22520 4632 22526 4684
rect 22741 4675 22799 4681
rect 22741 4641 22753 4675
rect 22787 4672 22799 4675
rect 23750 4672 23756 4684
rect 22787 4644 23756 4672
rect 22787 4641 22799 4644
rect 22741 4635 22799 4641
rect 23750 4632 23756 4644
rect 23808 4632 23814 4684
rect 3099 4576 3556 4604
rect 10321 4607 10379 4613
rect 3099 4573 3111 4576
rect 3053 4567 3111 4573
rect 10321 4573 10333 4607
rect 10367 4573 10379 4607
rect 13354 4604 13360 4616
rect 13315 4576 13360 4604
rect 10321 4567 10379 4573
rect 2774 4536 2780 4548
rect 2332 4508 2780 4536
rect 2332 4480 2360 4508
rect 2774 4496 2780 4508
rect 2832 4496 2838 4548
rect 9398 4536 9404 4548
rect 8312 4508 9404 4536
rect 8312 4480 8340 4508
rect 9398 4496 9404 4508
rect 9456 4536 9462 4548
rect 10336 4536 10364 4567
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 14642 4604 14648 4616
rect 14603 4576 14648 4604
rect 14642 4564 14648 4576
rect 14700 4564 14706 4616
rect 18874 4604 18880 4616
rect 18835 4576 18880 4604
rect 18874 4564 18880 4576
rect 18932 4564 18938 4616
rect 19058 4604 19064 4616
rect 19019 4576 19064 4604
rect 19058 4564 19064 4576
rect 19116 4564 19122 4616
rect 9456 4508 10364 4536
rect 12989 4539 13047 4545
rect 9456 4496 9462 4508
rect 12989 4505 13001 4539
rect 13035 4536 13047 4539
rect 13722 4536 13728 4548
rect 13035 4508 13728 4536
rect 13035 4505 13047 4508
rect 12989 4499 13047 4505
rect 13722 4496 13728 4508
rect 13780 4496 13786 4548
rect 2133 4471 2191 4477
rect 2133 4437 2145 4471
rect 2179 4468 2191 4471
rect 2314 4468 2320 4480
rect 2179 4440 2320 4468
rect 2179 4437 2191 4440
rect 2133 4431 2191 4437
rect 2314 4428 2320 4440
rect 2372 4428 2378 4480
rect 2501 4471 2559 4477
rect 2501 4437 2513 4471
rect 2547 4468 2559 4471
rect 2590 4468 2596 4480
rect 2547 4440 2596 4468
rect 2547 4437 2559 4440
rect 2501 4431 2559 4437
rect 2590 4428 2596 4440
rect 2648 4428 2654 4480
rect 5994 4468 6000 4480
rect 5955 4440 6000 4468
rect 5994 4428 6000 4440
rect 6052 4428 6058 4480
rect 6914 4468 6920 4480
rect 6875 4440 6920 4468
rect 6914 4428 6920 4440
rect 6972 4428 6978 4480
rect 8294 4468 8300 4480
rect 8255 4440 8300 4468
rect 8294 4428 8300 4440
rect 8352 4428 8358 4480
rect 9309 4471 9367 4477
rect 9309 4437 9321 4471
rect 9355 4468 9367 4471
rect 9582 4468 9588 4480
rect 9355 4440 9588 4468
rect 9355 4437 9367 4440
rect 9309 4431 9367 4437
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 9769 4471 9827 4477
rect 9769 4437 9781 4471
rect 9815 4468 9827 4471
rect 10134 4468 10140 4480
rect 9815 4440 10140 4468
rect 9815 4437 9827 4440
rect 9769 4431 9827 4437
rect 10134 4428 10140 4440
rect 10192 4428 10198 4480
rect 11330 4468 11336 4480
rect 11291 4440 11336 4468
rect 11330 4428 11336 4440
rect 11388 4428 11394 4480
rect 13078 4428 13084 4480
rect 13136 4468 13142 4480
rect 13909 4471 13967 4477
rect 13909 4468 13921 4471
rect 13136 4440 13921 4468
rect 13136 4428 13142 4440
rect 13909 4437 13921 4440
rect 13955 4437 13967 4471
rect 17310 4468 17316 4480
rect 17271 4440 17316 4468
rect 13909 4431 13967 4437
rect 17310 4428 17316 4440
rect 17368 4428 17374 4480
rect 18506 4468 18512 4480
rect 18467 4440 18512 4468
rect 18506 4428 18512 4440
rect 18564 4428 18570 4480
rect 20898 4428 20904 4480
rect 20956 4468 20962 4480
rect 21085 4471 21143 4477
rect 21085 4468 21097 4471
rect 20956 4440 21097 4468
rect 20956 4428 20962 4440
rect 21085 4437 21097 4440
rect 21131 4437 21143 4471
rect 21085 4431 21143 4437
rect 23937 4471 23995 4477
rect 23937 4437 23949 4471
rect 23983 4468 23995 4471
rect 25406 4468 25412 4480
rect 23983 4440 25412 4468
rect 23983 4437 23995 4440
rect 23937 4431 23995 4437
rect 25406 4428 25412 4440
rect 25464 4428 25470 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 6178 4264 6184 4276
rect 2884 4236 6184 4264
rect 2884 4208 2912 4236
rect 6178 4224 6184 4236
rect 6236 4224 6242 4276
rect 7101 4267 7159 4273
rect 7101 4233 7113 4267
rect 7147 4264 7159 4267
rect 7466 4264 7472 4276
rect 7147 4236 7472 4264
rect 7147 4233 7159 4236
rect 7101 4227 7159 4233
rect 7466 4224 7472 4236
rect 7524 4224 7530 4276
rect 7742 4264 7748 4276
rect 7703 4236 7748 4264
rect 7742 4224 7748 4236
rect 7800 4224 7806 4276
rect 9306 4264 9312 4276
rect 9267 4236 9312 4264
rect 9306 4224 9312 4236
rect 9364 4224 9370 4276
rect 10045 4267 10103 4273
rect 10045 4233 10057 4267
rect 10091 4264 10103 4267
rect 10410 4264 10416 4276
rect 10091 4236 10416 4264
rect 10091 4233 10103 4236
rect 10045 4227 10103 4233
rect 10410 4224 10416 4236
rect 10468 4224 10474 4276
rect 10689 4267 10747 4273
rect 10689 4233 10701 4267
rect 10735 4264 10747 4267
rect 11238 4264 11244 4276
rect 10735 4236 11244 4264
rect 10735 4233 10747 4236
rect 10689 4227 10747 4233
rect 11238 4224 11244 4236
rect 11296 4224 11302 4276
rect 11698 4224 11704 4276
rect 11756 4264 11762 4276
rect 11793 4267 11851 4273
rect 11793 4264 11805 4267
rect 11756 4236 11805 4264
rect 11756 4224 11762 4236
rect 11793 4233 11805 4236
rect 11839 4233 11851 4267
rect 11793 4227 11851 4233
rect 12529 4267 12587 4273
rect 12529 4233 12541 4267
rect 12575 4264 12587 4267
rect 12802 4264 12808 4276
rect 12575 4236 12808 4264
rect 12575 4233 12587 4236
rect 12529 4227 12587 4233
rect 12802 4224 12808 4236
rect 12860 4224 12866 4276
rect 13354 4224 13360 4276
rect 13412 4264 13418 4276
rect 13449 4267 13507 4273
rect 13449 4264 13461 4267
rect 13412 4236 13461 4264
rect 13412 4224 13418 4236
rect 13449 4233 13461 4236
rect 13495 4233 13507 4267
rect 13449 4227 13507 4233
rect 15930 4224 15936 4276
rect 15988 4264 15994 4276
rect 16758 4264 16764 4276
rect 15988 4236 16764 4264
rect 15988 4224 15994 4236
rect 16758 4224 16764 4236
rect 16816 4224 16822 4276
rect 18874 4264 18880 4276
rect 18835 4236 18880 4264
rect 18874 4224 18880 4236
rect 18932 4224 18938 4276
rect 19058 4224 19064 4276
rect 19116 4264 19122 4276
rect 19153 4267 19211 4273
rect 19153 4264 19165 4267
rect 19116 4236 19165 4264
rect 19116 4224 19122 4236
rect 19153 4233 19165 4236
rect 19199 4233 19211 4267
rect 19153 4227 19211 4233
rect 22462 4224 22468 4276
rect 22520 4264 22526 4276
rect 22833 4267 22891 4273
rect 22833 4264 22845 4267
rect 22520 4236 22845 4264
rect 22520 4224 22526 4236
rect 22833 4233 22845 4236
rect 22879 4233 22891 4267
rect 22833 4227 22891 4233
rect 23750 4224 23756 4276
rect 23808 4264 23814 4276
rect 24581 4267 24639 4273
rect 24581 4264 24593 4267
rect 23808 4236 24593 4264
rect 23808 4224 23814 4236
rect 24581 4233 24593 4236
rect 24627 4233 24639 4267
rect 24581 4227 24639 4233
rect 2866 4196 2872 4208
rect 2608 4168 2872 4196
rect 1765 4131 1823 4137
rect 1765 4097 1777 4131
rect 1811 4128 1823 4131
rect 2608 4128 2636 4168
rect 2866 4156 2872 4168
rect 2924 4156 2930 4208
rect 3050 4196 3056 4208
rect 3011 4168 3056 4196
rect 3050 4156 3056 4168
rect 3108 4156 3114 4208
rect 7282 4156 7288 4208
rect 7340 4196 7346 4208
rect 8018 4196 8024 4208
rect 7340 4168 8024 4196
rect 7340 4156 7346 4168
rect 8018 4156 8024 4168
rect 8076 4196 8082 4208
rect 8076 4168 8340 4196
rect 8076 4156 8082 4168
rect 1811 4100 2636 4128
rect 2685 4131 2743 4137
rect 1811 4097 1823 4100
rect 1765 4091 1823 4097
rect 2685 4097 2697 4131
rect 2731 4128 2743 4131
rect 2958 4128 2964 4140
rect 2731 4100 2964 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4128 4307 4131
rect 6181 4131 6239 4137
rect 6181 4128 6193 4131
rect 4295 4100 6193 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 6181 4097 6193 4100
rect 6227 4128 6239 4131
rect 6549 4131 6607 4137
rect 6549 4128 6561 4131
rect 6227 4100 6561 4128
rect 6227 4097 6239 4100
rect 6181 4091 6239 4097
rect 6549 4097 6561 4100
rect 6595 4128 6607 4131
rect 7098 4128 7104 4140
rect 6595 4100 7104 4128
rect 6595 4097 6607 4100
rect 6549 4091 6607 4097
rect 7098 4088 7104 4100
rect 7156 4088 7162 4140
rect 7374 4088 7380 4140
rect 7432 4128 7438 4140
rect 8312 4137 8340 4168
rect 9582 4156 9588 4208
rect 9640 4156 9646 4208
rect 10870 4196 10876 4208
rect 10831 4168 10876 4196
rect 10870 4156 10876 4168
rect 10928 4156 10934 4208
rect 15470 4196 15476 4208
rect 15212 4168 15476 4196
rect 7469 4131 7527 4137
rect 7469 4128 7481 4131
rect 7432 4100 7481 4128
rect 7432 4088 7438 4100
rect 7469 4097 7481 4100
rect 7515 4097 7527 4131
rect 7469 4091 7527 4097
rect 8297 4131 8355 4137
rect 8297 4097 8309 4131
rect 8343 4097 8355 4131
rect 9600 4128 9628 4156
rect 9861 4131 9919 4137
rect 9861 4128 9873 4131
rect 9600 4100 9873 4128
rect 8297 4091 8355 4097
rect 9861 4097 9873 4100
rect 9907 4128 9919 4131
rect 10042 4128 10048 4140
rect 9907 4100 10048 4128
rect 9907 4097 9919 4100
rect 9861 4091 9919 4097
rect 1670 4020 1676 4072
rect 1728 4060 1734 4072
rect 5077 4063 5135 4069
rect 1728 4032 2636 4060
rect 1728 4020 1734 4032
rect 2314 3952 2320 4004
rect 2372 3992 2378 4004
rect 2608 4001 2636 4032
rect 5077 4029 5089 4063
rect 5123 4060 5135 4063
rect 5534 4060 5540 4072
rect 5123 4032 5540 4060
rect 5123 4029 5135 4032
rect 5077 4023 5135 4029
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 7484 4060 7512 4091
rect 10042 4088 10048 4100
rect 10100 4088 10106 4140
rect 11146 4088 11152 4140
rect 11204 4128 11210 4140
rect 11425 4131 11483 4137
rect 11425 4128 11437 4131
rect 11204 4100 11437 4128
rect 11204 4088 11210 4100
rect 11425 4097 11437 4100
rect 11471 4097 11483 4131
rect 12158 4128 12164 4140
rect 12119 4100 12164 4128
rect 11425 4091 11483 4097
rect 12158 4088 12164 4100
rect 12216 4128 12222 4140
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 12216 4100 12909 4128
rect 12216 4088 12222 4100
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 13078 4128 13084 4140
rect 13039 4100 13084 4128
rect 12897 4091 12955 4097
rect 13078 4088 13084 4100
rect 13136 4088 13142 4140
rect 13909 4131 13967 4137
rect 13909 4097 13921 4131
rect 13955 4128 13967 4131
rect 14182 4128 14188 4140
rect 13955 4100 14188 4128
rect 13955 4097 13967 4100
rect 13909 4091 13967 4097
rect 7484 4032 8248 4060
rect 2409 3995 2467 4001
rect 2409 3992 2421 3995
rect 2372 3964 2421 3992
rect 2372 3952 2378 3964
rect 2409 3961 2421 3964
rect 2455 3961 2467 3995
rect 2409 3955 2467 3961
rect 2593 3995 2651 4001
rect 2593 3961 2605 3995
rect 2639 3961 2651 3995
rect 2593 3955 2651 3961
rect 2774 3952 2780 4004
rect 2832 3992 2838 4004
rect 3513 3995 3571 4001
rect 3513 3992 3525 3995
rect 2832 3964 3525 3992
rect 2832 3952 2838 3964
rect 3513 3961 3525 3964
rect 3559 3992 3571 3995
rect 3973 3995 4031 4001
rect 3973 3992 3985 3995
rect 3559 3964 3985 3992
rect 3559 3961 3571 3964
rect 3513 3955 3571 3961
rect 3973 3961 3985 3964
rect 4019 3961 4031 3995
rect 3973 3955 4031 3961
rect 4062 3952 4068 4004
rect 4120 3992 4126 4004
rect 4157 3995 4215 4001
rect 4157 3992 4169 3995
rect 4120 3964 4169 3992
rect 4120 3952 4126 3964
rect 4157 3961 4169 3964
rect 4203 3992 4215 3995
rect 4798 3992 4804 4004
rect 4203 3964 4804 3992
rect 4203 3961 4215 3964
rect 4157 3955 4215 3961
rect 4798 3952 4804 3964
rect 4856 3952 4862 4004
rect 5810 3992 5816 4004
rect 5771 3964 5816 3992
rect 5810 3952 5816 3964
rect 5868 3952 5874 4004
rect 7650 3952 7656 4004
rect 7708 3992 7714 4004
rect 8220 4001 8248 4032
rect 9766 4020 9772 4072
rect 9824 4060 9830 4072
rect 10134 4060 10140 4072
rect 9824 4032 10140 4060
rect 9824 4020 9830 4032
rect 10134 4020 10140 4032
rect 10192 4020 10198 4072
rect 8021 3995 8079 4001
rect 8021 3992 8033 3995
rect 7708 3964 8033 3992
rect 7708 3952 7714 3964
rect 8021 3961 8033 3964
rect 8067 3961 8079 3995
rect 8021 3955 8079 3961
rect 8205 3995 8263 4001
rect 8205 3961 8217 3995
rect 8251 3961 8263 3995
rect 8205 3955 8263 3961
rect 8386 3952 8392 4004
rect 8444 3992 8450 4004
rect 8757 3995 8815 4001
rect 8757 3992 8769 3995
rect 8444 3964 8769 3992
rect 8444 3952 8450 3964
rect 8757 3961 8769 3964
rect 8803 3992 8815 3995
rect 9214 3992 9220 4004
rect 8803 3964 9220 3992
rect 8803 3961 8815 3964
rect 8757 3955 8815 3961
rect 9214 3952 9220 3964
rect 9272 3952 9278 4004
rect 9398 3952 9404 4004
rect 9456 3992 9462 4004
rect 9585 3995 9643 4001
rect 9585 3992 9597 3995
rect 9456 3964 9597 3992
rect 9456 3952 9462 3964
rect 9585 3961 9597 3964
rect 9631 3992 9643 3995
rect 10045 3995 10103 4001
rect 10045 3992 10057 3995
rect 9631 3964 10057 3992
rect 9631 3961 9643 3964
rect 9585 3955 9643 3961
rect 10045 3961 10057 3964
rect 10091 3961 10103 3995
rect 10045 3955 10103 3961
rect 10226 3952 10232 4004
rect 10284 3992 10290 4004
rect 10321 3995 10379 4001
rect 10321 3992 10333 3995
rect 10284 3964 10333 3992
rect 10284 3952 10290 3964
rect 10321 3961 10333 3964
rect 10367 3992 10379 3995
rect 10870 3992 10876 4004
rect 10367 3964 10876 3992
rect 10367 3961 10379 3964
rect 10321 3955 10379 3961
rect 10870 3952 10876 3964
rect 10928 3952 10934 4004
rect 11149 3995 11207 4001
rect 11149 3961 11161 3995
rect 11195 3961 11207 3995
rect 11330 3992 11336 4004
rect 11291 3964 11336 3992
rect 11149 3955 11207 3961
rect 1394 3884 1400 3936
rect 1452 3924 1458 3936
rect 1765 3927 1823 3933
rect 1765 3924 1777 3927
rect 1452 3896 1777 3924
rect 1452 3884 1458 3896
rect 1765 3893 1777 3896
rect 1811 3924 1823 3927
rect 1857 3927 1915 3933
rect 1857 3924 1869 3927
rect 1811 3896 1869 3924
rect 1811 3893 1823 3896
rect 1765 3887 1823 3893
rect 1857 3893 1869 3896
rect 1903 3893 1915 3927
rect 1857 3887 1915 3893
rect 2123 3927 2181 3933
rect 2123 3893 2135 3927
rect 2169 3924 2181 3927
rect 2866 3924 2872 3936
rect 2169 3896 2872 3924
rect 2169 3893 2181 3896
rect 2123 3887 2181 3893
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 3694 3933 3700 3936
rect 3687 3927 3700 3933
rect 3687 3893 3699 3927
rect 3752 3924 3758 3936
rect 4709 3927 4767 3933
rect 3752 3896 3787 3924
rect 3687 3887 3700 3893
rect 3694 3884 3700 3887
rect 3752 3884 3758 3896
rect 4709 3893 4721 3927
rect 4755 3924 4767 3927
rect 5074 3924 5080 3936
rect 4755 3896 5080 3924
rect 4755 3893 4767 3896
rect 4709 3887 4767 3893
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 5258 3933 5264 3936
rect 5251 3927 5264 3933
rect 5251 3924 5263 3927
rect 5219 3896 5263 3924
rect 5251 3893 5263 3896
rect 5251 3887 5264 3893
rect 5258 3884 5264 3887
rect 5316 3884 5322 3936
rect 5718 3924 5724 3936
rect 5679 3896 5724 3924
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 9125 3927 9183 3933
rect 9125 3893 9137 3927
rect 9171 3924 9183 3927
rect 9766 3924 9772 3936
rect 9171 3896 9772 3924
rect 9171 3893 9183 3896
rect 9125 3887 9183 3893
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 11054 3884 11060 3936
rect 11112 3924 11118 3936
rect 11164 3924 11192 3955
rect 11330 3952 11336 3964
rect 11388 3952 11394 4004
rect 12986 3992 12992 4004
rect 12947 3964 12992 3992
rect 12986 3952 12992 3964
rect 13044 3952 13050 4004
rect 13924 3992 13952 4091
rect 14182 4088 14188 4100
rect 14240 4088 14246 4140
rect 14458 4088 14464 4140
rect 14516 4128 14522 4140
rect 14645 4131 14703 4137
rect 14645 4128 14657 4131
rect 14516 4100 14657 4128
rect 14516 4088 14522 4100
rect 14645 4097 14657 4100
rect 14691 4128 14703 4131
rect 15212 4128 15240 4168
rect 15470 4156 15476 4168
rect 15528 4156 15534 4208
rect 15841 4199 15899 4205
rect 15841 4165 15853 4199
rect 15887 4165 15899 4199
rect 15841 4159 15899 4165
rect 14691 4100 15240 4128
rect 15856 4128 15884 4159
rect 16942 4128 16948 4140
rect 15856 4100 16948 4128
rect 14691 4097 14703 4100
rect 14645 4091 14703 4097
rect 16942 4088 16948 4100
rect 17000 4088 17006 4140
rect 17770 4128 17776 4140
rect 17731 4100 17776 4128
rect 17770 4088 17776 4100
rect 17828 4088 17834 4140
rect 18322 4128 18328 4140
rect 18283 4100 18328 4128
rect 18322 4088 18328 4100
rect 18380 4088 18386 4140
rect 13998 4020 14004 4072
rect 14056 4060 14062 4072
rect 14369 4063 14427 4069
rect 14369 4060 14381 4063
rect 14056 4032 14381 4060
rect 14056 4020 14062 4032
rect 14369 4029 14381 4032
rect 14415 4029 14427 4063
rect 14369 4023 14427 4029
rect 15746 4020 15752 4072
rect 15804 4060 15810 4072
rect 16117 4063 16175 4069
rect 16117 4060 16129 4063
rect 15804 4032 16129 4060
rect 15804 4020 15810 4032
rect 16117 4029 16129 4032
rect 16163 4029 16175 4063
rect 17126 4060 17132 4072
rect 17087 4032 17132 4060
rect 16117 4023 16175 4029
rect 17126 4020 17132 4032
rect 17184 4020 17190 4072
rect 17788 4060 17816 4088
rect 18049 4063 18107 4069
rect 18049 4060 18061 4063
rect 17788 4032 18061 4060
rect 18049 4029 18061 4032
rect 18095 4029 18107 4063
rect 19334 4060 19340 4072
rect 19295 4032 19340 4060
rect 18049 4023 18107 4029
rect 19334 4020 19340 4032
rect 19392 4060 19398 4072
rect 19889 4063 19947 4069
rect 19889 4060 19901 4063
rect 19392 4032 19901 4060
rect 19392 4020 19398 4032
rect 19889 4029 19901 4032
rect 19935 4029 19947 4063
rect 19889 4023 19947 4029
rect 20254 4020 20260 4072
rect 20312 4060 20318 4072
rect 20441 4063 20499 4069
rect 20441 4060 20453 4063
rect 20312 4032 20453 4060
rect 20312 4020 20318 4032
rect 20441 4029 20453 4032
rect 20487 4029 20499 4063
rect 21726 4060 21732 4072
rect 21687 4032 21732 4060
rect 20441 4023 20499 4029
rect 21726 4020 21732 4032
rect 21784 4060 21790 4072
rect 22465 4063 22523 4069
rect 22465 4060 22477 4063
rect 21784 4032 22477 4060
rect 21784 4020 21790 4032
rect 22465 4029 22477 4032
rect 22511 4029 22523 4063
rect 23658 4060 23664 4072
rect 23619 4032 23664 4060
rect 22465 4023 22523 4029
rect 23658 4020 23664 4032
rect 23716 4060 23722 4072
rect 24213 4063 24271 4069
rect 24213 4060 24225 4063
rect 23716 4032 24225 4060
rect 23716 4020 23722 4032
rect 24213 4029 24225 4032
rect 24259 4029 24271 4063
rect 24762 4060 24768 4072
rect 24723 4032 24768 4060
rect 24213 4023 24271 4029
rect 24762 4020 24768 4032
rect 24820 4060 24826 4072
rect 25317 4063 25375 4069
rect 25317 4060 25329 4063
rect 24820 4032 25329 4060
rect 24820 4020 24826 4032
rect 25317 4029 25329 4032
rect 25363 4029 25375 4063
rect 25317 4023 25375 4029
rect 14553 3995 14611 4001
rect 14553 3992 14565 3995
rect 13924 3964 14565 3992
rect 14553 3961 14565 3964
rect 14599 3961 14611 3995
rect 14553 3955 14611 3961
rect 15289 3995 15347 4001
rect 15289 3961 15301 3995
rect 15335 3992 15347 3995
rect 15930 3992 15936 4004
rect 15335 3964 15936 3992
rect 15335 3961 15347 3964
rect 15289 3955 15347 3961
rect 15930 3952 15936 3964
rect 15988 3992 15994 4004
rect 16393 3995 16451 4001
rect 16393 3992 16405 3995
rect 15988 3964 16405 3992
rect 15988 3952 15994 3964
rect 16393 3961 16405 3964
rect 16439 3992 16451 3995
rect 17310 3992 17316 4004
rect 16439 3964 17316 3992
rect 16439 3961 16451 3964
rect 16393 3955 16451 3961
rect 17310 3952 17316 3964
rect 17368 3952 17374 4004
rect 18690 3952 18696 4004
rect 18748 3992 18754 4004
rect 22002 3992 22008 4004
rect 18748 3964 20668 3992
rect 21963 3964 22008 3992
rect 18748 3952 18754 3964
rect 12710 3924 12716 3936
rect 11112 3896 12716 3924
rect 11112 3884 11118 3896
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 14083 3927 14141 3933
rect 14083 3893 14095 3927
rect 14129 3924 14141 3927
rect 14182 3924 14188 3936
rect 14129 3896 14188 3924
rect 14129 3893 14141 3896
rect 14083 3887 14141 3893
rect 14182 3884 14188 3896
rect 14240 3884 14246 3936
rect 14642 3884 14648 3936
rect 14700 3924 14706 3936
rect 15378 3924 15384 3936
rect 14700 3896 15384 3924
rect 14700 3884 14706 3896
rect 15378 3884 15384 3896
rect 15436 3924 15442 3936
rect 15565 3927 15623 3933
rect 15565 3924 15577 3927
rect 15436 3896 15577 3924
rect 15436 3884 15442 3896
rect 15565 3893 15577 3896
rect 15611 3924 15623 3927
rect 16301 3927 16359 3933
rect 16301 3924 16313 3927
rect 15611 3896 16313 3924
rect 15611 3893 15623 3896
rect 15565 3887 15623 3893
rect 16301 3893 16313 3896
rect 16347 3893 16359 3927
rect 19518 3924 19524 3936
rect 19479 3896 19524 3924
rect 16301 3887 16359 3893
rect 19518 3884 19524 3896
rect 19576 3884 19582 3936
rect 20254 3924 20260 3936
rect 20215 3896 20260 3924
rect 20254 3884 20260 3896
rect 20312 3884 20318 3936
rect 20640 3933 20668 3964
rect 22002 3952 22008 3964
rect 22060 3952 22066 4004
rect 20625 3927 20683 3933
rect 20625 3893 20637 3927
rect 20671 3893 20683 3927
rect 20990 3924 20996 3936
rect 20951 3896 20996 3924
rect 20625 3887 20683 3893
rect 20990 3884 20996 3896
rect 21048 3884 21054 3936
rect 23845 3927 23903 3933
rect 23845 3893 23857 3927
rect 23891 3924 23903 3927
rect 24118 3924 24124 3936
rect 23891 3896 24124 3924
rect 23891 3893 23903 3896
rect 23845 3887 23903 3893
rect 24118 3884 24124 3896
rect 24176 3884 24182 3936
rect 24949 3927 25007 3933
rect 24949 3893 24961 3927
rect 24995 3924 25007 3927
rect 25958 3924 25964 3936
rect 24995 3896 25964 3924
rect 24995 3893 25007 3896
rect 24949 3887 25007 3893
rect 25958 3884 25964 3896
rect 26016 3884 26022 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1670 3680 1676 3732
rect 1728 3720 1734 3732
rect 2041 3723 2099 3729
rect 2041 3720 2053 3723
rect 1728 3692 2053 3720
rect 1728 3680 1734 3692
rect 2041 3689 2053 3692
rect 2087 3720 2099 3723
rect 2406 3720 2412 3732
rect 2087 3692 2412 3720
rect 2087 3689 2099 3692
rect 2041 3683 2099 3689
rect 2406 3680 2412 3692
rect 2464 3680 2470 3732
rect 2590 3680 2596 3732
rect 2648 3720 2654 3732
rect 2648 3692 3004 3720
rect 2648 3680 2654 3692
rect 2976 3664 3004 3692
rect 3050 3680 3056 3732
rect 3108 3720 3114 3732
rect 3421 3723 3479 3729
rect 3421 3720 3433 3723
rect 3108 3692 3433 3720
rect 3108 3680 3114 3692
rect 3421 3689 3433 3692
rect 3467 3720 3479 3723
rect 3789 3723 3847 3729
rect 3789 3720 3801 3723
rect 3467 3692 3801 3720
rect 3467 3689 3479 3692
rect 3421 3683 3479 3689
rect 3789 3689 3801 3692
rect 3835 3689 3847 3723
rect 7098 3720 7104 3732
rect 3789 3683 3847 3689
rect 4448 3692 6408 3720
rect 7059 3692 7104 3720
rect 2958 3652 2964 3664
rect 2919 3624 2964 3652
rect 2958 3612 2964 3624
rect 3016 3612 3022 3664
rect 3234 3612 3240 3664
rect 3292 3652 3298 3664
rect 4448 3661 4476 3692
rect 4433 3655 4491 3661
rect 4433 3652 4445 3655
rect 3292 3624 4445 3652
rect 3292 3612 3298 3624
rect 4433 3621 4445 3624
rect 4479 3621 4491 3655
rect 4614 3652 4620 3664
rect 4575 3624 4620 3652
rect 4433 3615 4491 3621
rect 4614 3612 4620 3624
rect 4672 3612 4678 3664
rect 5537 3655 5595 3661
rect 5537 3621 5549 3655
rect 5583 3652 5595 3655
rect 5810 3652 5816 3664
rect 5583 3624 5816 3652
rect 5583 3621 5595 3624
rect 5537 3615 5595 3621
rect 5810 3612 5816 3624
rect 5868 3652 5874 3664
rect 6270 3652 6276 3664
rect 5868 3624 6276 3652
rect 5868 3612 5874 3624
rect 6270 3612 6276 3624
rect 6328 3612 6334 3664
rect 6380 3652 6408 3692
rect 7098 3680 7104 3692
rect 7156 3680 7162 3732
rect 8018 3720 8024 3732
rect 7979 3692 8024 3720
rect 8018 3680 8024 3692
rect 8076 3680 8082 3732
rect 9217 3723 9275 3729
rect 9217 3720 9229 3723
rect 8312 3692 9229 3720
rect 8312 3652 8340 3692
rect 9217 3689 9229 3692
rect 9263 3720 9275 3723
rect 9398 3720 9404 3732
rect 9263 3692 9404 3720
rect 9263 3689 9275 3692
rect 9217 3683 9275 3689
rect 9398 3680 9404 3692
rect 9456 3720 9462 3732
rect 10413 3723 10471 3729
rect 10413 3720 10425 3723
rect 9456 3692 10425 3720
rect 9456 3680 9462 3692
rect 10413 3689 10425 3692
rect 10459 3689 10471 3723
rect 10413 3683 10471 3689
rect 10873 3723 10931 3729
rect 10873 3689 10885 3723
rect 10919 3720 10931 3723
rect 11054 3720 11060 3732
rect 10919 3692 11060 3720
rect 10919 3689 10931 3692
rect 10873 3683 10931 3689
rect 11054 3680 11060 3692
rect 11112 3680 11118 3732
rect 11790 3720 11796 3732
rect 11532 3692 11796 3720
rect 6380 3624 8340 3652
rect 8481 3655 8539 3661
rect 8481 3621 8493 3655
rect 8527 3652 8539 3655
rect 8662 3652 8668 3664
rect 8527 3624 8668 3652
rect 8527 3621 8539 3624
rect 8481 3615 8539 3621
rect 8662 3612 8668 3624
rect 8720 3612 8726 3664
rect 9858 3612 9864 3664
rect 9916 3612 9922 3664
rect 9953 3655 10011 3661
rect 9953 3621 9965 3655
rect 9999 3652 10011 3655
rect 10134 3652 10140 3664
rect 9999 3624 10140 3652
rect 9999 3621 10011 3624
rect 9953 3615 10011 3621
rect 10134 3612 10140 3624
rect 10192 3612 10198 3664
rect 11532 3661 11560 3692
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 12526 3720 12532 3732
rect 12487 3692 12532 3720
rect 12526 3680 12532 3692
rect 12584 3680 12590 3732
rect 13262 3720 13268 3732
rect 13223 3692 13268 3720
rect 13262 3680 13268 3692
rect 13320 3680 13326 3732
rect 13998 3720 14004 3732
rect 13959 3692 14004 3720
rect 13998 3680 14004 3692
rect 14056 3680 14062 3732
rect 14458 3720 14464 3732
rect 14419 3692 14464 3720
rect 14458 3680 14464 3692
rect 14516 3680 14522 3732
rect 16117 3723 16175 3729
rect 16117 3689 16129 3723
rect 16163 3720 16175 3723
rect 16206 3720 16212 3732
rect 16163 3692 16212 3720
rect 16163 3689 16175 3692
rect 16117 3683 16175 3689
rect 16206 3680 16212 3692
rect 16264 3680 16270 3732
rect 16298 3680 16304 3732
rect 16356 3720 16362 3732
rect 16393 3723 16451 3729
rect 16393 3720 16405 3723
rect 16356 3692 16405 3720
rect 16356 3680 16362 3692
rect 16393 3689 16405 3692
rect 16439 3689 16451 3723
rect 16393 3683 16451 3689
rect 16942 3680 16948 3732
rect 17000 3720 17006 3732
rect 19061 3723 19119 3729
rect 19061 3720 19073 3723
rect 17000 3692 19073 3720
rect 17000 3680 17006 3692
rect 19061 3689 19073 3692
rect 19107 3689 19119 3723
rect 19061 3683 19119 3689
rect 19426 3680 19432 3732
rect 19484 3720 19490 3732
rect 19797 3723 19855 3729
rect 19797 3720 19809 3723
rect 19484 3692 19809 3720
rect 19484 3680 19490 3692
rect 19797 3689 19809 3692
rect 19843 3689 19855 3723
rect 19978 3720 19984 3732
rect 19939 3692 19984 3720
rect 19797 3683 19855 3689
rect 19978 3680 19984 3692
rect 20036 3680 20042 3732
rect 11517 3655 11575 3661
rect 11517 3621 11529 3655
rect 11563 3621 11575 3655
rect 11517 3615 11575 3621
rect 11606 3612 11612 3664
rect 11664 3652 11670 3664
rect 11701 3655 11759 3661
rect 11701 3652 11713 3655
rect 11664 3624 11713 3652
rect 11664 3612 11670 3624
rect 11701 3621 11713 3624
rect 11747 3621 11759 3655
rect 14734 3652 14740 3664
rect 14695 3624 14740 3652
rect 11701 3615 11759 3621
rect 14734 3612 14740 3624
rect 14792 3612 14798 3664
rect 17028 3655 17086 3661
rect 17028 3621 17040 3655
rect 17074 3652 17086 3655
rect 17310 3652 17316 3664
rect 17074 3624 17316 3652
rect 17074 3621 17086 3624
rect 17028 3615 17086 3621
rect 17310 3612 17316 3624
rect 17368 3612 17374 3664
rect 18506 3612 18512 3664
rect 18564 3652 18570 3664
rect 18693 3655 18751 3661
rect 18693 3652 18705 3655
rect 18564 3624 18705 3652
rect 18564 3612 18570 3624
rect 18693 3621 18705 3624
rect 18739 3621 18751 3655
rect 18693 3615 18751 3621
rect 23017 3655 23075 3661
rect 23017 3621 23029 3655
rect 23063 3652 23075 3655
rect 24762 3652 24768 3664
rect 23063 3624 24768 3652
rect 23063 3621 23075 3624
rect 23017 3615 23075 3621
rect 24762 3612 24768 3624
rect 24820 3612 24826 3664
rect 2774 3544 2780 3596
rect 2832 3584 2838 3596
rect 3053 3587 3111 3593
rect 3053 3584 3065 3587
rect 2832 3556 3065 3584
rect 2832 3544 2838 3556
rect 3053 3553 3065 3556
rect 3099 3553 3111 3587
rect 3053 3547 3111 3553
rect 5626 3544 5632 3596
rect 5684 3584 5690 3596
rect 5988 3587 6046 3593
rect 5988 3584 6000 3587
rect 5684 3556 6000 3584
rect 5684 3544 5690 3556
rect 5988 3553 6000 3556
rect 6034 3584 6046 3587
rect 6822 3584 6828 3596
rect 6034 3556 6828 3584
rect 6034 3553 6046 3556
rect 5988 3547 6046 3553
rect 6822 3544 6828 3556
rect 6880 3544 6886 3596
rect 8202 3584 8208 3596
rect 8163 3556 8208 3584
rect 8202 3544 8208 3556
rect 8260 3544 8266 3596
rect 9677 3587 9735 3593
rect 9677 3553 9689 3587
rect 9723 3584 9735 3587
rect 9876 3584 9904 3612
rect 9723 3556 9904 3584
rect 13081 3587 13139 3593
rect 9723 3553 9735 3556
rect 9677 3547 9735 3553
rect 13081 3553 13093 3587
rect 13127 3584 13139 3587
rect 14366 3584 14372 3596
rect 13127 3556 14372 3584
rect 13127 3553 13139 3556
rect 13081 3547 13139 3553
rect 14366 3544 14372 3556
rect 14424 3544 14430 3596
rect 15289 3587 15347 3593
rect 15289 3553 15301 3587
rect 15335 3584 15347 3587
rect 15838 3584 15844 3596
rect 15335 3556 15844 3584
rect 15335 3553 15347 3556
rect 15289 3547 15347 3553
rect 15838 3544 15844 3556
rect 15896 3544 15902 3596
rect 16758 3584 16764 3596
rect 16719 3556 16764 3584
rect 16758 3544 16764 3556
rect 16816 3544 16822 3596
rect 18414 3544 18420 3596
rect 18472 3584 18478 3596
rect 19245 3587 19303 3593
rect 19245 3584 19257 3587
rect 18472 3556 19257 3584
rect 18472 3544 18478 3556
rect 19245 3553 19257 3556
rect 19291 3584 19303 3587
rect 19978 3584 19984 3596
rect 19291 3556 19984 3584
rect 19291 3553 19303 3556
rect 19245 3547 19303 3553
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 20714 3544 20720 3596
rect 20772 3584 20778 3596
rect 20901 3587 20959 3593
rect 20901 3584 20913 3587
rect 20772 3556 20913 3584
rect 20772 3544 20778 3556
rect 20901 3553 20913 3556
rect 20947 3584 20959 3587
rect 21634 3584 21640 3596
rect 20947 3556 21640 3584
rect 20947 3553 20959 3556
rect 20901 3547 20959 3553
rect 21634 3544 21640 3556
rect 21692 3544 21698 3596
rect 22738 3584 22744 3596
rect 22699 3556 22744 3584
rect 22738 3544 22744 3556
rect 22796 3544 22802 3596
rect 24026 3584 24032 3596
rect 23987 3556 24032 3584
rect 24026 3544 24032 3556
rect 24084 3544 24090 3596
rect 25130 3584 25136 3596
rect 25091 3556 25136 3584
rect 25130 3544 25136 3556
rect 25188 3544 25194 3596
rect 1397 3519 1455 3525
rect 1397 3485 1409 3519
rect 1443 3516 1455 3519
rect 2222 3516 2228 3528
rect 1443 3488 2228 3516
rect 1443 3485 1455 3488
rect 1397 3479 1455 3485
rect 2222 3476 2228 3488
rect 2280 3476 2286 3528
rect 2958 3516 2964 3528
rect 2919 3488 2964 3516
rect 2958 3476 2964 3488
rect 3016 3476 3022 3528
rect 4706 3516 4712 3528
rect 4667 3488 4712 3516
rect 4706 3476 4712 3488
rect 4764 3476 4770 3528
rect 5074 3476 5080 3528
rect 5132 3516 5138 3528
rect 5721 3519 5779 3525
rect 5721 3516 5733 3519
rect 5132 3488 5733 3516
rect 5132 3476 5138 3488
rect 5721 3485 5733 3488
rect 5767 3485 5779 3519
rect 11790 3516 11796 3528
rect 11751 3488 11796 3516
rect 5721 3479 5779 3485
rect 11790 3476 11796 3488
rect 11848 3516 11854 3528
rect 12710 3516 12716 3528
rect 11848 3488 12716 3516
rect 11848 3476 11854 3488
rect 12710 3476 12716 3488
rect 12768 3476 12774 3528
rect 13354 3516 13360 3528
rect 13315 3488 13360 3516
rect 13354 3476 13360 3488
rect 13412 3476 13418 3528
rect 15562 3516 15568 3528
rect 15523 3488 15568 3516
rect 15562 3476 15568 3488
rect 15620 3476 15626 3528
rect 20806 3476 20812 3528
rect 20864 3516 20870 3528
rect 20990 3516 20996 3528
rect 20864 3488 20996 3516
rect 20864 3476 20870 3488
rect 20990 3476 20996 3488
rect 21048 3476 21054 3528
rect 2498 3448 2504 3460
rect 2459 3420 2504 3448
rect 2498 3408 2504 3420
rect 2556 3408 2562 3460
rect 3050 3408 3056 3460
rect 3108 3448 3114 3460
rect 3878 3448 3884 3460
rect 3108 3420 3884 3448
rect 3108 3408 3114 3420
rect 3878 3408 3884 3420
rect 3936 3448 3942 3460
rect 11241 3451 11299 3457
rect 3936 3420 5764 3448
rect 3936 3408 3942 3420
rect 4154 3380 4160 3392
rect 4115 3352 4160 3380
rect 4154 3340 4160 3352
rect 4212 3340 4218 3392
rect 5074 3380 5080 3392
rect 5035 3352 5080 3380
rect 5074 3340 5080 3352
rect 5132 3340 5138 3392
rect 5736 3380 5764 3420
rect 11241 3417 11253 3451
rect 11287 3448 11299 3451
rect 13262 3448 13268 3460
rect 11287 3420 13268 3448
rect 11287 3417 11299 3420
rect 11241 3411 11299 3417
rect 13262 3408 13268 3420
rect 13320 3408 13326 3460
rect 19429 3451 19487 3457
rect 19429 3417 19441 3451
rect 19475 3448 19487 3451
rect 19981 3451 20039 3457
rect 19981 3448 19993 3451
rect 19475 3420 19993 3448
rect 19475 3417 19487 3420
rect 19429 3411 19487 3417
rect 19981 3417 19993 3420
rect 20027 3417 20039 3451
rect 19981 3411 20039 3417
rect 7650 3380 7656 3392
rect 5736 3352 7656 3380
rect 7650 3340 7656 3352
rect 7708 3380 7714 3392
rect 9582 3380 9588 3392
rect 7708 3352 9588 3380
rect 7708 3340 7714 3352
rect 9582 3340 9588 3352
rect 9640 3340 9646 3392
rect 12802 3380 12808 3392
rect 12763 3352 12808 3380
rect 12802 3340 12808 3352
rect 12860 3340 12866 3392
rect 17954 3340 17960 3392
rect 18012 3380 18018 3392
rect 18141 3383 18199 3389
rect 18141 3380 18153 3383
rect 18012 3352 18153 3380
rect 18012 3340 18018 3352
rect 18141 3349 18153 3352
rect 18187 3349 18199 3383
rect 20162 3380 20168 3392
rect 20123 3352 20168 3380
rect 18141 3343 18199 3349
rect 20162 3340 20168 3352
rect 20220 3340 20226 3392
rect 20806 3340 20812 3392
rect 20864 3380 20870 3392
rect 21085 3383 21143 3389
rect 21085 3380 21097 3383
rect 20864 3352 21097 3380
rect 20864 3340 20870 3352
rect 21085 3349 21097 3352
rect 21131 3349 21143 3383
rect 21085 3343 21143 3349
rect 23198 3340 23204 3392
rect 23256 3380 23262 3392
rect 24213 3383 24271 3389
rect 24213 3380 24225 3383
rect 23256 3352 24225 3380
rect 23256 3340 23262 3352
rect 24213 3349 24225 3352
rect 24259 3349 24271 3383
rect 24213 3343 24271 3349
rect 24946 3340 24952 3392
rect 25004 3380 25010 3392
rect 25317 3383 25375 3389
rect 25317 3380 25329 3383
rect 25004 3352 25329 3380
rect 25004 3340 25010 3352
rect 25317 3349 25329 3352
rect 25363 3349 25375 3383
rect 25317 3343 25375 3349
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 2777 3179 2835 3185
rect 2777 3145 2789 3179
rect 2823 3176 2835 3179
rect 4062 3176 4068 3188
rect 2823 3148 4068 3176
rect 2823 3145 2835 3148
rect 2777 3139 2835 3145
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 5629 3179 5687 3185
rect 5629 3176 5641 3179
rect 5592 3148 5641 3176
rect 5592 3136 5598 3148
rect 5629 3145 5641 3148
rect 5675 3145 5687 3179
rect 9122 3176 9128 3188
rect 9083 3148 9128 3176
rect 5629 3139 5687 3145
rect 9122 3136 9128 3148
rect 9180 3136 9186 3188
rect 10686 3136 10692 3188
rect 10744 3176 10750 3188
rect 10962 3176 10968 3188
rect 10744 3148 10968 3176
rect 10744 3136 10750 3148
rect 10962 3136 10968 3148
rect 11020 3136 11026 3188
rect 11606 3176 11612 3188
rect 11567 3148 11612 3176
rect 11606 3136 11612 3148
rect 11664 3136 11670 3188
rect 11882 3176 11888 3188
rect 11843 3148 11888 3176
rect 11882 3136 11888 3148
rect 11940 3136 11946 3188
rect 13354 3136 13360 3188
rect 13412 3176 13418 3188
rect 13814 3176 13820 3188
rect 13412 3148 13820 3176
rect 13412 3136 13418 3148
rect 13814 3136 13820 3148
rect 13872 3136 13878 3188
rect 14366 3176 14372 3188
rect 14327 3148 14372 3176
rect 14366 3136 14372 3148
rect 14424 3136 14430 3188
rect 15930 3176 15936 3188
rect 15891 3148 15936 3176
rect 15930 3136 15936 3148
rect 15988 3136 15994 3188
rect 16482 3176 16488 3188
rect 16443 3148 16488 3176
rect 16482 3136 16488 3148
rect 16540 3136 16546 3188
rect 16758 3136 16764 3188
rect 16816 3176 16822 3188
rect 17405 3179 17463 3185
rect 17405 3176 17417 3179
rect 16816 3148 17417 3176
rect 16816 3136 16822 3148
rect 17405 3145 17417 3148
rect 17451 3176 17463 3179
rect 17773 3179 17831 3185
rect 17773 3176 17785 3179
rect 17451 3148 17785 3176
rect 17451 3145 17463 3148
rect 17405 3139 17463 3145
rect 17773 3145 17785 3148
rect 17819 3145 17831 3179
rect 19978 3176 19984 3188
rect 19939 3148 19984 3176
rect 17773 3139 17831 3145
rect 3234 3108 3240 3120
rect 3160 3080 3240 3108
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3040 1731 3043
rect 2130 3040 2136 3052
rect 1719 3012 2136 3040
rect 1719 3009 1731 3012
rect 1673 3003 1731 3009
rect 2130 3000 2136 3012
rect 2188 3000 2194 3052
rect 2866 3000 2872 3052
rect 2924 3040 2930 3052
rect 3160 3049 3188 3080
rect 3234 3068 3240 3080
rect 3292 3108 3298 3120
rect 3697 3111 3755 3117
rect 3697 3108 3709 3111
rect 3292 3080 3709 3108
rect 3292 3068 3298 3080
rect 3697 3077 3709 3080
rect 3743 3077 3755 3111
rect 3697 3071 3755 3077
rect 3145 3043 3203 3049
rect 3145 3040 3157 3043
rect 2924 3012 3157 3040
rect 2924 3000 2930 3012
rect 3145 3009 3157 3012
rect 3191 3009 3203 3043
rect 3326 3040 3332 3052
rect 3287 3012 3332 3040
rect 3145 3003 3203 3009
rect 3326 3000 3332 3012
rect 3384 3000 3390 3052
rect 14734 3000 14740 3052
rect 14792 3040 14798 3052
rect 15378 3040 15384 3052
rect 14792 3012 15148 3040
rect 15339 3012 15384 3040
rect 14792 3000 14798 3012
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2972 1455 2975
rect 3694 2972 3700 2984
rect 1443 2944 3700 2972
rect 1443 2941 1455 2944
rect 1397 2935 1455 2941
rect 3694 2932 3700 2944
rect 3752 2932 3758 2984
rect 3970 2932 3976 2984
rect 4028 2972 4034 2984
rect 4249 2975 4307 2981
rect 4249 2972 4261 2975
rect 4028 2944 4261 2972
rect 4028 2932 4034 2944
rect 4249 2941 4261 2944
rect 4295 2972 4307 2975
rect 5074 2972 5080 2984
rect 4295 2944 5080 2972
rect 4295 2941 4307 2944
rect 4249 2935 4307 2941
rect 5074 2932 5080 2944
rect 5132 2972 5138 2984
rect 6181 2975 6239 2981
rect 6181 2972 6193 2975
rect 5132 2944 6193 2972
rect 5132 2932 5138 2944
rect 6181 2941 6193 2944
rect 6227 2972 6239 2975
rect 6549 2975 6607 2981
rect 6549 2972 6561 2975
rect 6227 2944 6561 2972
rect 6227 2941 6239 2944
rect 6181 2935 6239 2941
rect 6549 2941 6561 2944
rect 6595 2972 6607 2975
rect 6730 2972 6736 2984
rect 6595 2944 6736 2972
rect 6595 2941 6607 2944
rect 6549 2935 6607 2941
rect 6730 2932 6736 2944
rect 6788 2972 6794 2984
rect 7374 2981 7380 2984
rect 7101 2975 7159 2981
rect 7101 2972 7113 2975
rect 6788 2944 7113 2972
rect 6788 2932 6794 2944
rect 7101 2941 7113 2944
rect 7147 2941 7159 2975
rect 7368 2972 7380 2981
rect 7101 2935 7159 2941
rect 7208 2944 7380 2972
rect 2225 2907 2283 2913
rect 2225 2873 2237 2907
rect 2271 2904 2283 2907
rect 2866 2904 2872 2916
rect 2271 2876 2872 2904
rect 2271 2873 2283 2876
rect 2225 2867 2283 2873
rect 2866 2864 2872 2876
rect 2924 2864 2930 2916
rect 4516 2907 4574 2913
rect 4516 2873 4528 2907
rect 4562 2904 4574 2907
rect 5442 2904 5448 2916
rect 4562 2876 5448 2904
rect 4562 2873 4574 2876
rect 4516 2867 4574 2873
rect 5442 2864 5448 2876
rect 5500 2864 5506 2916
rect 6270 2864 6276 2916
rect 6328 2904 6334 2916
rect 7208 2904 7236 2944
rect 7368 2935 7380 2944
rect 7374 2932 7380 2935
rect 7432 2932 7438 2984
rect 9490 2972 9496 2984
rect 9403 2944 9496 2972
rect 9490 2932 9496 2944
rect 9548 2972 9554 2984
rect 9585 2975 9643 2981
rect 9585 2972 9597 2975
rect 9548 2944 9597 2972
rect 9548 2932 9554 2944
rect 9585 2941 9597 2944
rect 9631 2941 9643 2975
rect 9585 2935 9643 2941
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2972 12495 2975
rect 12526 2972 12532 2984
rect 12483 2944 12532 2972
rect 12483 2941 12495 2944
rect 12437 2935 12495 2941
rect 12526 2932 12532 2944
rect 12584 2932 12590 2984
rect 12710 2981 12716 2984
rect 12704 2972 12716 2981
rect 12623 2944 12716 2972
rect 12704 2935 12716 2944
rect 12768 2972 12774 2984
rect 14826 2972 14832 2984
rect 12768 2944 14832 2972
rect 12710 2932 12716 2935
rect 12768 2932 12774 2944
rect 14826 2932 14832 2944
rect 14884 2932 14890 2984
rect 15120 2981 15148 3012
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 16301 3043 16359 3049
rect 16301 3009 16313 3043
rect 16347 3040 16359 3043
rect 16945 3043 17003 3049
rect 16945 3040 16957 3043
rect 16347 3012 16957 3040
rect 16347 3009 16359 3012
rect 16301 3003 16359 3009
rect 16945 3009 16957 3012
rect 16991 3040 17003 3043
rect 17678 3040 17684 3052
rect 16991 3012 17684 3040
rect 16991 3009 17003 3012
rect 16945 3003 17003 3009
rect 17678 3000 17684 3012
rect 17736 3000 17742 3052
rect 17788 3040 17816 3139
rect 19978 3136 19984 3148
rect 20036 3136 20042 3188
rect 21634 3176 21640 3188
rect 21595 3148 21640 3176
rect 21634 3136 21640 3148
rect 21692 3136 21698 3188
rect 22738 3176 22744 3188
rect 22699 3148 22744 3176
rect 22738 3136 22744 3148
rect 22796 3136 22802 3188
rect 23474 3176 23480 3188
rect 23435 3148 23480 3176
rect 23474 3136 23480 3148
rect 23532 3136 23538 3188
rect 25130 3136 25136 3188
rect 25188 3176 25194 3188
rect 25501 3179 25559 3185
rect 25501 3176 25513 3179
rect 25188 3148 25513 3176
rect 25188 3136 25194 3148
rect 25501 3145 25513 3148
rect 25547 3145 25559 3179
rect 25501 3139 25559 3145
rect 18049 3043 18107 3049
rect 18049 3040 18061 3043
rect 17788 3012 18061 3040
rect 18049 3009 18061 3012
rect 18095 3009 18107 3043
rect 18049 3003 18107 3009
rect 19978 3000 19984 3052
rect 20036 3040 20042 3052
rect 20438 3040 20444 3052
rect 20036 3012 20444 3040
rect 20036 3000 20042 3012
rect 20438 3000 20444 3012
rect 20496 3000 20502 3052
rect 15105 2975 15163 2981
rect 15105 2941 15117 2975
rect 15151 2941 15163 2975
rect 15105 2935 15163 2941
rect 9830 2907 9888 2913
rect 9830 2904 9842 2907
rect 6328 2876 7236 2904
rect 9692 2876 9842 2904
rect 6328 2864 6334 2876
rect 2593 2839 2651 2845
rect 2593 2805 2605 2839
rect 2639 2836 2651 2839
rect 3234 2836 3240 2848
rect 2639 2808 3240 2836
rect 2639 2805 2651 2808
rect 2593 2799 2651 2805
rect 3234 2796 3240 2808
rect 3292 2796 3298 2848
rect 4157 2839 4215 2845
rect 4157 2805 4169 2839
rect 4203 2836 4215 2839
rect 4614 2836 4620 2848
rect 4203 2808 4620 2836
rect 4203 2805 4215 2808
rect 4157 2799 4215 2805
rect 4614 2796 4620 2808
rect 4672 2836 4678 2848
rect 5258 2836 5264 2848
rect 4672 2808 5264 2836
rect 4672 2796 4678 2808
rect 5258 2796 5264 2808
rect 5316 2796 5322 2848
rect 8478 2836 8484 2848
rect 8439 2808 8484 2836
rect 8478 2796 8484 2808
rect 8536 2796 8542 2848
rect 9582 2796 9588 2848
rect 9640 2836 9646 2848
rect 9692 2836 9720 2876
rect 9830 2873 9842 2876
rect 9876 2873 9888 2907
rect 9830 2867 9888 2873
rect 9640 2808 9720 2836
rect 15120 2836 15148 2935
rect 16574 2932 16580 2984
rect 16632 2972 16638 2984
rect 17037 2975 17095 2981
rect 17037 2972 17049 2975
rect 16632 2944 17049 2972
rect 16632 2932 16638 2944
rect 17037 2941 17049 2944
rect 17083 2972 17095 2975
rect 17954 2972 17960 2984
rect 17083 2944 17960 2972
rect 17083 2941 17095 2944
rect 17037 2935 17095 2941
rect 17954 2932 17960 2944
rect 18012 2932 18018 2984
rect 20530 2972 20536 2984
rect 20491 2944 20536 2972
rect 20530 2932 20536 2944
rect 20588 2972 20594 2984
rect 21269 2975 21327 2981
rect 21269 2972 21281 2975
rect 20588 2944 21281 2972
rect 20588 2932 20594 2944
rect 21269 2941 21281 2944
rect 21315 2941 21327 2975
rect 21818 2972 21824 2984
rect 21779 2944 21824 2972
rect 21269 2935 21327 2941
rect 21818 2932 21824 2944
rect 21876 2972 21882 2984
rect 22373 2975 22431 2981
rect 22373 2972 22385 2975
rect 21876 2944 22385 2972
rect 21876 2932 21882 2944
rect 22373 2941 22385 2944
rect 22419 2941 22431 2975
rect 22373 2935 22431 2941
rect 23474 2932 23480 2984
rect 23532 2972 23538 2984
rect 23661 2975 23719 2981
rect 23661 2972 23673 2975
rect 23532 2944 23673 2972
rect 23532 2932 23538 2944
rect 23661 2941 23673 2944
rect 23707 2941 23719 2975
rect 24026 2972 24032 2984
rect 23661 2935 23719 2941
rect 23768 2944 24032 2972
rect 16942 2904 16948 2916
rect 16903 2876 16948 2904
rect 16942 2864 16948 2876
rect 17000 2864 17006 2916
rect 17972 2904 18000 2932
rect 18294 2907 18352 2913
rect 18294 2904 18306 2907
rect 17972 2876 18306 2904
rect 18294 2873 18306 2876
rect 18340 2873 18352 2907
rect 20349 2907 20407 2913
rect 20349 2904 20361 2907
rect 18294 2867 18352 2873
rect 18984 2876 20361 2904
rect 18984 2836 19012 2876
rect 20349 2873 20361 2876
rect 20395 2873 20407 2907
rect 20349 2867 20407 2873
rect 20809 2907 20867 2913
rect 20809 2873 20821 2907
rect 20855 2904 20867 2907
rect 23768 2904 23796 2944
rect 24026 2932 24032 2944
rect 24084 2972 24090 2984
rect 24397 2975 24455 2981
rect 24397 2972 24409 2975
rect 24084 2944 24409 2972
rect 24084 2932 24090 2944
rect 24397 2941 24409 2944
rect 24443 2941 24455 2975
rect 24397 2935 24455 2941
rect 24762 2932 24768 2984
rect 24820 2972 24826 2984
rect 24857 2975 24915 2981
rect 24857 2972 24869 2975
rect 24820 2944 24869 2972
rect 24820 2932 24826 2944
rect 24857 2941 24869 2944
rect 24903 2972 24915 2975
rect 24949 2975 25007 2981
rect 24949 2972 24961 2975
rect 24903 2944 24961 2972
rect 24903 2941 24915 2944
rect 24857 2935 24915 2941
rect 24949 2941 24961 2944
rect 24995 2941 25007 2975
rect 24949 2935 25007 2941
rect 20855 2876 23796 2904
rect 23937 2907 23995 2913
rect 20855 2873 20867 2876
rect 20809 2867 20867 2873
rect 23937 2873 23949 2907
rect 23983 2904 23995 2907
rect 25038 2904 25044 2916
rect 23983 2876 25044 2904
rect 23983 2873 23995 2876
rect 23937 2867 23995 2873
rect 25038 2864 25044 2876
rect 25096 2864 25102 2916
rect 19426 2836 19432 2848
rect 15120 2808 19012 2836
rect 19387 2808 19432 2836
rect 9640 2796 9646 2808
rect 19426 2796 19432 2808
rect 19484 2796 19490 2848
rect 22002 2836 22008 2848
rect 21963 2808 22008 2836
rect 22002 2796 22008 2808
rect 22060 2796 22066 2848
rect 25130 2836 25136 2848
rect 25091 2808 25136 2836
rect 25130 2796 25136 2808
rect 25188 2796 25194 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 2222 2632 2228 2644
rect 2183 2604 2228 2632
rect 2222 2592 2228 2604
rect 2280 2632 2286 2644
rect 3237 2635 3295 2641
rect 2280 2604 2820 2632
rect 2280 2592 2286 2604
rect 1397 2567 1455 2573
rect 1397 2533 1409 2567
rect 1443 2564 1455 2567
rect 2682 2564 2688 2576
rect 1443 2536 2688 2564
rect 1443 2533 1455 2536
rect 1397 2527 1455 2533
rect 2682 2524 2688 2536
rect 2740 2524 2746 2576
rect 2792 2573 2820 2604
rect 3237 2601 3249 2635
rect 3283 2632 3295 2635
rect 3513 2635 3571 2641
rect 3513 2632 3525 2635
rect 3283 2604 3525 2632
rect 3283 2601 3295 2604
rect 3237 2595 3295 2601
rect 3513 2601 3525 2604
rect 3559 2632 3571 2635
rect 5442 2632 5448 2644
rect 3559 2604 5448 2632
rect 3559 2601 3571 2604
rect 3513 2595 3571 2601
rect 5442 2592 5448 2604
rect 5500 2632 5506 2644
rect 5994 2632 6000 2644
rect 5500 2604 6000 2632
rect 5500 2592 5506 2604
rect 5994 2592 6000 2604
rect 6052 2592 6058 2644
rect 6270 2632 6276 2644
rect 6231 2604 6276 2632
rect 6270 2592 6276 2604
rect 6328 2592 6334 2644
rect 6730 2632 6736 2644
rect 6691 2604 6736 2632
rect 6730 2592 6736 2604
rect 6788 2592 6794 2644
rect 8294 2592 8300 2644
rect 8352 2632 8358 2644
rect 8573 2635 8631 2641
rect 8573 2632 8585 2635
rect 8352 2604 8585 2632
rect 8352 2592 8358 2604
rect 8573 2601 8585 2604
rect 8619 2632 8631 2635
rect 9582 2632 9588 2644
rect 8619 2604 9588 2632
rect 8619 2601 8631 2604
rect 8573 2595 8631 2601
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 11146 2632 11152 2644
rect 11107 2604 11152 2632
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 12437 2635 12495 2641
rect 12437 2601 12449 2635
rect 12483 2632 12495 2635
rect 12526 2632 12532 2644
rect 12483 2604 12532 2632
rect 12483 2601 12495 2604
rect 12437 2595 12495 2601
rect 12526 2592 12532 2604
rect 12584 2592 12590 2644
rect 13998 2632 14004 2644
rect 13959 2604 14004 2632
rect 13998 2592 14004 2604
rect 14056 2592 14062 2644
rect 16485 2635 16543 2641
rect 16485 2601 16497 2635
rect 16531 2632 16543 2635
rect 16574 2632 16580 2644
rect 16531 2604 16580 2632
rect 16531 2601 16543 2604
rect 16485 2595 16543 2601
rect 16574 2592 16580 2604
rect 16632 2592 16638 2644
rect 17954 2592 17960 2644
rect 18012 2632 18018 2644
rect 18049 2635 18107 2641
rect 18049 2632 18061 2635
rect 18012 2604 18061 2632
rect 18012 2592 18018 2604
rect 18049 2601 18061 2604
rect 18095 2601 18107 2635
rect 18049 2595 18107 2601
rect 19797 2635 19855 2641
rect 19797 2601 19809 2635
rect 19843 2632 19855 2635
rect 19978 2632 19984 2644
rect 19843 2604 19984 2632
rect 19843 2601 19855 2604
rect 19797 2595 19855 2601
rect 19978 2592 19984 2604
rect 20036 2592 20042 2644
rect 20990 2592 20996 2644
rect 21048 2632 21054 2644
rect 21361 2635 21419 2641
rect 21361 2632 21373 2635
rect 21048 2604 21373 2632
rect 21048 2592 21054 2604
rect 21361 2601 21373 2604
rect 21407 2601 21419 2635
rect 21361 2595 21419 2601
rect 2777 2567 2835 2573
rect 2777 2533 2789 2567
rect 2823 2533 2835 2567
rect 2777 2527 2835 2533
rect 2961 2567 3019 2573
rect 2961 2533 2973 2567
rect 3007 2564 3019 2567
rect 4062 2564 4068 2576
rect 3007 2536 4068 2564
rect 3007 2533 3019 2536
rect 2961 2527 3019 2533
rect 4062 2524 4068 2536
rect 4120 2524 4126 2576
rect 4332 2567 4390 2573
rect 4332 2533 4344 2567
rect 4378 2564 4390 2567
rect 4706 2564 4712 2576
rect 4378 2536 4712 2564
rect 4378 2533 4390 2536
rect 4332 2527 4390 2533
rect 4706 2524 4712 2536
rect 4764 2524 4770 2576
rect 3053 2499 3111 2505
rect 3053 2465 3065 2499
rect 3099 2496 3111 2499
rect 3237 2499 3295 2505
rect 3237 2496 3249 2499
rect 3099 2468 3249 2496
rect 3099 2465 3111 2468
rect 3053 2459 3111 2465
rect 3237 2465 3249 2468
rect 3283 2465 3295 2499
rect 6748 2496 6776 2592
rect 7098 2524 7104 2576
rect 7156 2564 7162 2576
rect 10042 2573 10048 2576
rect 7438 2567 7496 2573
rect 7438 2564 7450 2567
rect 7156 2536 7450 2564
rect 7156 2524 7162 2536
rect 7438 2533 7450 2536
rect 7484 2533 7496 2567
rect 7438 2527 7496 2533
rect 9217 2567 9275 2573
rect 9217 2533 9229 2567
rect 9263 2564 9275 2567
rect 10036 2564 10048 2573
rect 9263 2536 10048 2564
rect 9263 2533 9275 2536
rect 9217 2527 9275 2533
rect 10036 2527 10048 2536
rect 10042 2524 10048 2527
rect 10100 2524 10106 2576
rect 12069 2567 12127 2573
rect 12069 2533 12081 2567
rect 12115 2564 12127 2567
rect 12866 2567 12924 2573
rect 12866 2564 12878 2567
rect 12115 2536 12878 2564
rect 12115 2533 12127 2536
rect 12069 2527 12127 2533
rect 12866 2533 12878 2536
rect 12912 2564 12924 2567
rect 13814 2564 13820 2576
rect 12912 2536 13820 2564
rect 12912 2533 12924 2536
rect 12866 2527 12924 2533
rect 13814 2524 13820 2536
rect 13872 2564 13878 2576
rect 14553 2567 14611 2573
rect 14553 2564 14565 2567
rect 13872 2536 14565 2564
rect 13872 2524 13878 2536
rect 14553 2533 14565 2536
rect 14599 2533 14611 2567
rect 17034 2564 17040 2576
rect 16995 2536 17040 2564
rect 14553 2527 14611 2533
rect 17034 2524 17040 2536
rect 17092 2524 17098 2576
rect 18598 2564 18604 2576
rect 18559 2536 18604 2564
rect 18598 2524 18604 2536
rect 18656 2524 18662 2576
rect 24305 2567 24363 2573
rect 24305 2533 24317 2567
rect 24351 2564 24363 2567
rect 24762 2564 24768 2576
rect 24351 2536 24768 2564
rect 24351 2533 24363 2536
rect 24305 2527 24363 2533
rect 24762 2524 24768 2536
rect 24820 2524 24826 2576
rect 7193 2499 7251 2505
rect 7193 2496 7205 2499
rect 6748 2468 7205 2496
rect 3237 2459 3295 2465
rect 7193 2465 7205 2468
rect 7239 2496 7251 2499
rect 9490 2496 9496 2508
rect 7239 2468 9496 2496
rect 7239 2465 7251 2468
rect 7193 2459 7251 2465
rect 9490 2456 9496 2468
rect 9548 2496 9554 2508
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 9548 2468 9781 2496
rect 9548 2456 9554 2468
rect 9769 2465 9781 2468
rect 9815 2496 9827 2499
rect 12526 2496 12532 2508
rect 9815 2468 12532 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 12526 2456 12532 2468
rect 12584 2496 12590 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12584 2468 12633 2496
rect 12584 2456 12590 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 15470 2496 15476 2508
rect 12621 2459 12679 2465
rect 12728 2468 15476 2496
rect 1949 2431 2007 2437
rect 1949 2397 1961 2431
rect 1995 2428 2007 2431
rect 2038 2428 2044 2440
rect 1995 2400 2044 2428
rect 1995 2397 2007 2400
rect 1949 2391 2007 2397
rect 2038 2388 2044 2400
rect 2096 2428 2102 2440
rect 2682 2428 2688 2440
rect 2096 2400 2688 2428
rect 2096 2388 2102 2400
rect 2682 2388 2688 2400
rect 2740 2388 2746 2440
rect 3881 2431 3939 2437
rect 3881 2397 3893 2431
rect 3927 2428 3939 2431
rect 3970 2428 3976 2440
rect 3927 2400 3976 2428
rect 3927 2397 3939 2400
rect 3881 2391 3939 2397
rect 3970 2388 3976 2400
rect 4028 2428 4034 2440
rect 4065 2431 4123 2437
rect 4065 2428 4077 2431
rect 4028 2400 4077 2428
rect 4028 2388 4034 2400
rect 4065 2397 4077 2400
rect 4111 2397 4123 2431
rect 4065 2391 4123 2397
rect 11514 2388 11520 2440
rect 11572 2428 11578 2440
rect 12728 2428 12756 2468
rect 15470 2456 15476 2468
rect 15528 2456 15534 2508
rect 16758 2496 16764 2508
rect 16719 2468 16764 2496
rect 16758 2456 16764 2468
rect 16816 2496 16822 2508
rect 17497 2499 17555 2505
rect 17497 2496 17509 2499
rect 16816 2468 17509 2496
rect 16816 2456 16822 2468
rect 17497 2465 17509 2468
rect 17543 2465 17555 2499
rect 17497 2459 17555 2465
rect 18230 2456 18236 2508
rect 18288 2496 18294 2508
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 18288 2468 18337 2496
rect 18288 2456 18294 2468
rect 18325 2465 18337 2468
rect 18371 2496 18383 2499
rect 19061 2499 19119 2505
rect 19061 2496 19073 2499
rect 18371 2468 19073 2496
rect 18371 2465 18383 2468
rect 18325 2459 18383 2465
rect 19061 2465 19073 2468
rect 19107 2465 19119 2499
rect 19610 2496 19616 2508
rect 19571 2468 19616 2496
rect 19061 2459 19119 2465
rect 19610 2456 19616 2468
rect 19668 2496 19674 2508
rect 20165 2499 20223 2505
rect 20165 2496 20177 2499
rect 19668 2468 20177 2496
rect 19668 2456 19674 2468
rect 20165 2465 20177 2468
rect 20211 2465 20223 2499
rect 21174 2496 21180 2508
rect 21135 2468 21180 2496
rect 20165 2459 20223 2465
rect 21174 2456 21180 2468
rect 21232 2496 21238 2508
rect 21729 2499 21787 2505
rect 21729 2496 21741 2499
rect 21232 2468 21741 2496
rect 21232 2456 21238 2468
rect 21729 2465 21741 2468
rect 21775 2465 21787 2499
rect 22278 2496 22284 2508
rect 22239 2468 22284 2496
rect 21729 2459 21787 2465
rect 22278 2456 22284 2468
rect 22336 2496 22342 2508
rect 22833 2499 22891 2505
rect 22833 2496 22845 2499
rect 22336 2468 22845 2496
rect 22336 2456 22342 2468
rect 22833 2465 22845 2468
rect 22879 2465 22891 2499
rect 24026 2496 24032 2508
rect 23987 2468 24032 2496
rect 22833 2459 22891 2465
rect 24026 2456 24032 2468
rect 24084 2496 24090 2508
rect 24857 2499 24915 2505
rect 24857 2496 24869 2499
rect 24084 2468 24869 2496
rect 24084 2456 24090 2468
rect 24857 2465 24869 2468
rect 24903 2465 24915 2499
rect 24857 2459 24915 2465
rect 25038 2456 25044 2508
rect 25096 2496 25102 2508
rect 25317 2499 25375 2505
rect 25317 2496 25329 2499
rect 25096 2468 25329 2496
rect 25096 2456 25102 2468
rect 25317 2465 25329 2468
rect 25363 2496 25375 2499
rect 25869 2499 25927 2505
rect 25869 2496 25881 2499
rect 25363 2468 25881 2496
rect 25363 2465 25375 2468
rect 25317 2459 25375 2465
rect 25869 2465 25881 2468
rect 25915 2465 25927 2499
rect 25869 2459 25927 2465
rect 15746 2428 15752 2440
rect 11572 2400 12756 2428
rect 15707 2400 15752 2428
rect 11572 2388 11578 2400
rect 15746 2388 15752 2400
rect 15804 2388 15810 2440
rect 20530 2428 20536 2440
rect 20491 2400 20536 2428
rect 20530 2388 20536 2400
rect 20588 2388 20594 2440
rect 1578 2320 1584 2372
rect 1636 2360 1642 2372
rect 2501 2363 2559 2369
rect 2501 2360 2513 2363
rect 1636 2332 2513 2360
rect 1636 2320 1642 2332
rect 2501 2329 2513 2332
rect 2547 2329 2559 2363
rect 2501 2323 2559 2329
rect 25501 2363 25559 2369
rect 25501 2329 25513 2363
rect 25547 2360 25559 2363
rect 26510 2360 26516 2372
rect 25547 2332 26516 2360
rect 25547 2329 25559 2332
rect 25501 2323 25559 2329
rect 26510 2320 26516 2332
rect 26568 2320 26574 2372
rect 14642 2252 14648 2304
rect 14700 2292 14706 2304
rect 14921 2295 14979 2301
rect 14921 2292 14933 2295
rect 14700 2264 14933 2292
rect 14700 2252 14706 2264
rect 14921 2261 14933 2264
rect 14967 2261 14979 2295
rect 19426 2292 19432 2304
rect 19387 2264 19432 2292
rect 14921 2255 14979 2261
rect 19426 2252 19432 2264
rect 19484 2252 19490 2304
rect 22462 2292 22468 2304
rect 22423 2264 22468 2292
rect 22462 2252 22468 2264
rect 22520 2252 22526 2304
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 9674 2048 9680 2100
rect 9732 2088 9738 2100
rect 15378 2088 15384 2100
rect 9732 2060 15384 2088
rect 9732 2048 9738 2060
rect 15378 2048 15384 2060
rect 15436 2048 15442 2100
rect 16666 2048 16672 2100
rect 16724 2088 16730 2100
rect 20714 2088 20720 2100
rect 16724 2060 20720 2088
rect 16724 2048 16730 2060
rect 20714 2048 20720 2060
rect 20772 2048 20778 2100
rect 14826 1096 14832 1148
rect 14884 1136 14890 1148
rect 15654 1136 15660 1148
rect 14884 1108 15660 1136
rect 14884 1096 14890 1108
rect 15654 1096 15660 1108
rect 15712 1096 15718 1148
rect 9030 660 9036 672
rect 6932 632 9036 660
rect 6932 604 6960 632
rect 9030 620 9036 632
rect 9088 620 9094 672
rect 6914 552 6920 604
rect 6972 552 6978 604
rect 7558 552 7564 604
rect 7616 592 7622 604
rect 7834 592 7840 604
rect 7616 564 7840 592
rect 7616 552 7622 564
rect 7834 552 7840 564
rect 7892 552 7898 604
rect 12250 552 12256 604
rect 12308 592 12314 604
rect 15930 592 15936 604
rect 12308 564 15936 592
rect 12308 552 12314 564
rect 15930 552 15936 564
rect 15988 552 15994 604
<< via1 >>
rect 2964 26256 3016 26308
rect 15752 26256 15804 26308
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 3424 24896 3476 24948
rect 13268 24896 13320 24948
rect 3516 24828 3568 24880
rect 14004 24828 14056 24880
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2412 14356 2464 14408
rect 1400 14220 1452 14272
rect 1952 14263 2004 14272
rect 1952 14229 1961 14263
rect 1961 14229 1995 14263
rect 1995 14229 2004 14263
rect 1952 14220 2004 14229
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 2044 14059 2096 14068
rect 2044 14025 2053 14059
rect 2053 14025 2087 14059
rect 2087 14025 2096 14059
rect 2044 14016 2096 14025
rect 2872 13880 2924 13932
rect 2044 13812 2096 13864
rect 2228 13812 2280 13864
rect 2136 13744 2188 13796
rect 1584 13719 1636 13728
rect 1584 13685 1593 13719
rect 1593 13685 1627 13719
rect 1627 13685 1636 13719
rect 1584 13676 1636 13685
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 7840 13515 7892 13524
rect 7840 13481 7849 13515
rect 7849 13481 7883 13515
rect 7883 13481 7892 13515
rect 7840 13472 7892 13481
rect 2596 13336 2648 13388
rect 4988 13336 5040 13388
rect 4160 13268 4212 13320
rect 2504 13200 2556 13252
rect 2964 13200 3016 13252
rect 1860 13132 1912 13184
rect 2320 13175 2372 13184
rect 2320 13141 2329 13175
rect 2329 13141 2363 13175
rect 2363 13141 2372 13175
rect 2320 13132 2372 13141
rect 2688 13175 2740 13184
rect 2688 13141 2697 13175
rect 2697 13141 2731 13175
rect 2731 13141 2740 13175
rect 2688 13132 2740 13141
rect 3424 13175 3476 13184
rect 3424 13141 3433 13175
rect 3433 13141 3467 13175
rect 3467 13141 3476 13175
rect 3424 13132 3476 13141
rect 4804 13132 4856 13184
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 2596 12971 2648 12980
rect 2596 12937 2605 12971
rect 2605 12937 2639 12971
rect 2639 12937 2648 12971
rect 2596 12928 2648 12937
rect 3700 12971 3752 12980
rect 3700 12937 3709 12971
rect 3709 12937 3743 12971
rect 3743 12937 3752 12971
rect 3700 12928 3752 12937
rect 6092 12928 6144 12980
rect 4712 12860 4764 12912
rect 8300 12860 8352 12912
rect 2136 12835 2188 12844
rect 2136 12801 2145 12835
rect 2145 12801 2179 12835
rect 2179 12801 2188 12835
rect 2136 12792 2188 12801
rect 2320 12792 2372 12844
rect 2780 12792 2832 12844
rect 5448 12792 5500 12844
rect 8944 12724 8996 12776
rect 2044 12656 2096 12708
rect 3424 12656 3476 12708
rect 3700 12656 3752 12708
rect 4620 12656 4672 12708
rect 7840 12656 7892 12708
rect 3056 12631 3108 12640
rect 3056 12597 3065 12631
rect 3065 12597 3099 12631
rect 3099 12597 3108 12631
rect 3056 12588 3108 12597
rect 4896 12631 4948 12640
rect 4896 12597 4905 12631
rect 4905 12597 4939 12631
rect 4939 12597 4948 12631
rect 4896 12588 4948 12597
rect 6644 12588 6696 12640
rect 9128 12588 9180 12640
rect 9588 12588 9640 12640
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1952 12384 2004 12436
rect 2412 12384 2464 12436
rect 2780 12384 2832 12436
rect 3332 12384 3384 12436
rect 3148 12316 3200 12368
rect 3608 12316 3660 12368
rect 3884 12316 3936 12368
rect 5264 12359 5316 12368
rect 5264 12325 5273 12359
rect 5273 12325 5307 12359
rect 5307 12325 5316 12359
rect 5264 12316 5316 12325
rect 5356 12316 5408 12368
rect 5908 12359 5960 12368
rect 5908 12325 5917 12359
rect 5917 12325 5951 12359
rect 5951 12325 5960 12359
rect 5908 12316 5960 12325
rect 10140 12316 10192 12368
rect 1400 12248 1452 12300
rect 2320 12248 2372 12300
rect 2044 12112 2096 12164
rect 4620 12180 4672 12232
rect 5448 12180 5500 12232
rect 6460 12223 6512 12232
rect 6460 12189 6469 12223
rect 6469 12189 6503 12223
rect 6503 12189 6512 12223
rect 6460 12180 6512 12189
rect 9772 12223 9824 12232
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 3148 12044 3200 12096
rect 4068 12044 4120 12096
rect 4252 12044 4304 12096
rect 4988 12087 5040 12096
rect 4988 12053 4997 12087
rect 4997 12053 5031 12087
rect 5031 12053 5040 12087
rect 4988 12044 5040 12053
rect 7472 12044 7524 12096
rect 11152 12087 11204 12096
rect 11152 12053 11161 12087
rect 11161 12053 11195 12087
rect 11195 12053 11204 12087
rect 11152 12044 11204 12053
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 2136 11840 2188 11892
rect 5264 11840 5316 11892
rect 8944 11883 8996 11892
rect 8944 11849 8953 11883
rect 8953 11849 8987 11883
rect 8987 11849 8996 11883
rect 8944 11840 8996 11849
rect 11244 11840 11296 11892
rect 16396 11840 16448 11892
rect 2412 11704 2464 11756
rect 5540 11704 5592 11756
rect 2044 11611 2096 11620
rect 2044 11577 2053 11611
rect 2053 11577 2087 11611
rect 2087 11577 2096 11611
rect 2044 11568 2096 11577
rect 3148 11568 3200 11620
rect 1492 11500 1544 11552
rect 2780 11500 2832 11552
rect 3332 11636 3384 11688
rect 7472 11568 7524 11620
rect 4620 11543 4672 11552
rect 4620 11509 4629 11543
rect 4629 11509 4663 11543
rect 4663 11509 4672 11543
rect 4620 11500 4672 11509
rect 5356 11500 5408 11552
rect 6460 11500 6512 11552
rect 6736 11500 6788 11552
rect 7012 11543 7064 11552
rect 7012 11509 7021 11543
rect 7021 11509 7055 11543
rect 7055 11509 7064 11543
rect 7012 11500 7064 11509
rect 9772 11543 9824 11552
rect 9772 11509 9781 11543
rect 9781 11509 9815 11543
rect 9815 11509 9824 11543
rect 9772 11500 9824 11509
rect 10048 11543 10100 11552
rect 10048 11509 10057 11543
rect 10057 11509 10091 11543
rect 10091 11509 10100 11543
rect 10048 11500 10100 11509
rect 10140 11500 10192 11552
rect 12164 11500 12216 11552
rect 12716 11500 12768 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 3332 11296 3384 11348
rect 3700 11296 3752 11348
rect 5448 11296 5500 11348
rect 7012 11296 7064 11348
rect 8300 11296 8352 11348
rect 2044 11228 2096 11280
rect 5540 11228 5592 11280
rect 11152 11271 11204 11280
rect 11152 11237 11186 11271
rect 11186 11237 11204 11271
rect 11152 11228 11204 11237
rect 3884 11160 3936 11212
rect 8208 11160 8260 11212
rect 16212 11203 16264 11212
rect 16212 11169 16221 11203
rect 16221 11169 16255 11203
rect 16255 11169 16264 11203
rect 16212 11160 16264 11169
rect 1492 11135 1544 11144
rect 1492 11101 1501 11135
rect 1501 11101 1535 11135
rect 1535 11101 1544 11135
rect 1492 11092 1544 11101
rect 5264 11092 5316 11144
rect 8576 11092 8628 11144
rect 9036 11135 9088 11144
rect 9036 11101 9045 11135
rect 9045 11101 9079 11135
rect 9079 11101 9088 11135
rect 9036 11092 9088 11101
rect 9772 11092 9824 11144
rect 13360 11135 13412 11144
rect 13360 11101 13369 11135
rect 13369 11101 13403 11135
rect 13403 11101 13412 11135
rect 13360 11092 13412 11101
rect 16488 11135 16540 11144
rect 16488 11101 16497 11135
rect 16497 11101 16531 11135
rect 16531 11101 16540 11135
rect 16488 11092 16540 11101
rect 4620 11024 4672 11076
rect 8116 11067 8168 11076
rect 8116 11033 8125 11067
rect 8125 11033 8159 11067
rect 8159 11033 8168 11067
rect 8116 11024 8168 11033
rect 9680 11024 9732 11076
rect 12348 11024 12400 11076
rect 15568 11024 15620 11076
rect 3516 10999 3568 11008
rect 3516 10965 3525 10999
rect 3525 10965 3559 10999
rect 3559 10965 3568 10999
rect 3516 10956 3568 10965
rect 7472 10956 7524 11008
rect 12072 10956 12124 11008
rect 12992 10956 13044 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1768 10752 1820 10804
rect 2044 10752 2096 10804
rect 5540 10752 5592 10804
rect 6644 10795 6696 10804
rect 6644 10761 6653 10795
rect 6653 10761 6687 10795
rect 6687 10761 6696 10795
rect 6644 10752 6696 10761
rect 8208 10752 8260 10804
rect 8576 10752 8628 10804
rect 10140 10752 10192 10804
rect 8668 10684 8720 10736
rect 12532 10727 12584 10736
rect 12532 10693 12541 10727
rect 12541 10693 12575 10727
rect 12575 10693 12584 10727
rect 12532 10684 12584 10693
rect 16212 10727 16264 10736
rect 16212 10693 16221 10727
rect 16221 10693 16255 10727
rect 16255 10693 16264 10727
rect 16212 10684 16264 10693
rect 1492 10548 1544 10600
rect 2780 10548 2832 10600
rect 2320 10480 2372 10532
rect 1676 10455 1728 10464
rect 1676 10421 1685 10455
rect 1685 10421 1719 10455
rect 1719 10421 1728 10455
rect 1676 10412 1728 10421
rect 3148 10455 3200 10464
rect 3148 10421 3157 10455
rect 3157 10421 3191 10455
rect 3191 10421 3200 10455
rect 3148 10412 3200 10421
rect 3884 10412 3936 10464
rect 4344 10412 4396 10464
rect 4620 10480 4672 10532
rect 5080 10480 5132 10532
rect 7472 10523 7524 10532
rect 7472 10489 7481 10523
rect 7481 10489 7515 10523
rect 7515 10489 7524 10523
rect 7472 10480 7524 10489
rect 8944 10591 8996 10600
rect 8944 10557 8978 10591
rect 8978 10557 8996 10591
rect 8944 10548 8996 10557
rect 12072 10548 12124 10600
rect 16672 10591 16724 10600
rect 16672 10557 16681 10591
rect 16681 10557 16715 10591
rect 16715 10557 16724 10591
rect 16672 10548 16724 10557
rect 9772 10480 9824 10532
rect 16948 10523 17000 10532
rect 16948 10489 16957 10523
rect 16957 10489 16991 10523
rect 16991 10489 17000 10523
rect 16948 10480 17000 10489
rect 5264 10412 5316 10464
rect 6736 10412 6788 10464
rect 7380 10455 7432 10464
rect 7380 10421 7389 10455
rect 7389 10421 7423 10455
rect 7423 10421 7432 10455
rect 7380 10412 7432 10421
rect 8484 10455 8536 10464
rect 8484 10421 8493 10455
rect 8493 10421 8527 10455
rect 8527 10421 8536 10455
rect 8484 10412 8536 10421
rect 8668 10412 8720 10464
rect 9404 10412 9456 10464
rect 12992 10455 13044 10464
rect 12992 10421 13001 10455
rect 13001 10421 13035 10455
rect 13035 10421 13044 10455
rect 12992 10412 13044 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2780 10251 2832 10260
rect 2780 10217 2789 10251
rect 2789 10217 2823 10251
rect 2823 10217 2832 10251
rect 2780 10208 2832 10217
rect 3148 10208 3200 10260
rect 1768 10140 1820 10192
rect 572 10072 624 10124
rect 4620 10140 4672 10192
rect 5540 10208 5592 10260
rect 6368 10208 6420 10260
rect 7472 10208 7524 10260
rect 8116 10208 8168 10260
rect 8576 10251 8628 10260
rect 8576 10217 8585 10251
rect 8585 10217 8619 10251
rect 8619 10217 8628 10251
rect 8576 10208 8628 10217
rect 8944 10251 8996 10260
rect 8944 10217 8953 10251
rect 8953 10217 8987 10251
rect 8987 10217 8996 10251
rect 8944 10208 8996 10217
rect 6276 10183 6328 10192
rect 6276 10149 6285 10183
rect 6285 10149 6319 10183
rect 6319 10149 6328 10183
rect 6276 10140 6328 10149
rect 6460 10183 6512 10192
rect 6460 10149 6469 10183
rect 6469 10149 6503 10183
rect 6503 10149 6512 10183
rect 6460 10140 6512 10149
rect 9680 10140 9732 10192
rect 10232 10140 10284 10192
rect 11152 10208 11204 10260
rect 12072 10183 12124 10192
rect 12072 10149 12106 10183
rect 12106 10149 12124 10183
rect 12072 10140 12124 10149
rect 5172 10072 5224 10124
rect 6828 10072 6880 10124
rect 8300 10072 8352 10124
rect 2136 10047 2188 10056
rect 2136 10013 2145 10047
rect 2145 10013 2179 10047
rect 2179 10013 2188 10047
rect 2136 10004 2188 10013
rect 2320 10047 2372 10056
rect 2320 10013 2329 10047
rect 2329 10013 2363 10047
rect 2363 10013 2372 10047
rect 2320 10004 2372 10013
rect 1952 9936 2004 9988
rect 5080 10004 5132 10056
rect 8024 10047 8076 10056
rect 8024 10013 8033 10047
rect 8033 10013 8067 10047
rect 8067 10013 8076 10047
rect 8024 10004 8076 10013
rect 11520 10004 11572 10056
rect 15292 10047 15344 10056
rect 15292 10013 15301 10047
rect 15301 10013 15335 10047
rect 15335 10013 15344 10047
rect 15292 10004 15344 10013
rect 4896 9936 4948 9988
rect 7564 9979 7616 9988
rect 7564 9945 7573 9979
rect 7573 9945 7607 9979
rect 7607 9945 7616 9979
rect 7564 9936 7616 9945
rect 9864 9979 9916 9988
rect 9864 9945 9873 9979
rect 9873 9945 9907 9979
rect 9907 9945 9916 9979
rect 9864 9936 9916 9945
rect 3516 9911 3568 9920
rect 3516 9877 3525 9911
rect 3525 9877 3559 9911
rect 3559 9877 3568 9911
rect 3516 9868 3568 9877
rect 8116 9868 8168 9920
rect 11152 9868 11204 9920
rect 12992 9868 13044 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 2596 9639 2648 9648
rect 2596 9605 2605 9639
rect 2605 9605 2639 9639
rect 2639 9605 2648 9639
rect 2596 9596 2648 9605
rect 4620 9664 4672 9716
rect 4436 9639 4488 9648
rect 4436 9605 4445 9639
rect 4445 9605 4479 9639
rect 4479 9605 4488 9639
rect 4436 9596 4488 9605
rect 3976 9528 4028 9580
rect 4344 9528 4396 9580
rect 5540 9664 5592 9716
rect 6276 9707 6328 9716
rect 6276 9673 6285 9707
rect 6285 9673 6319 9707
rect 6319 9673 6328 9707
rect 6276 9664 6328 9673
rect 8024 9664 8076 9716
rect 6736 9596 6788 9648
rect 8484 9664 8536 9716
rect 12072 9664 12124 9716
rect 5540 9528 5592 9580
rect 6460 9528 6512 9580
rect 9680 9596 9732 9648
rect 16396 9596 16448 9648
rect 17868 9596 17920 9648
rect 10232 9571 10284 9580
rect 10232 9537 10241 9571
rect 10241 9537 10275 9571
rect 10275 9537 10284 9571
rect 10232 9528 10284 9537
rect 11612 9528 11664 9580
rect 1676 9460 1728 9512
rect 2412 9460 2464 9512
rect 2872 9503 2924 9512
rect 2872 9469 2881 9503
rect 2881 9469 2915 9503
rect 2915 9469 2924 9503
rect 2872 9460 2924 9469
rect 4712 9503 4764 9512
rect 4712 9469 4721 9503
rect 4721 9469 4755 9503
rect 4755 9469 4764 9503
rect 4712 9460 4764 9469
rect 8116 9460 8168 9512
rect 8392 9460 8444 9512
rect 11520 9460 11572 9512
rect 12808 9460 12860 9512
rect 12992 9503 13044 9512
rect 3148 9435 3200 9444
rect 3148 9401 3157 9435
rect 3157 9401 3191 9435
rect 3191 9401 3200 9435
rect 3148 9392 3200 9401
rect 1492 9324 1544 9376
rect 1768 9324 1820 9376
rect 1952 9367 2004 9376
rect 1952 9333 1961 9367
rect 1961 9333 1995 9367
rect 1995 9333 2004 9367
rect 1952 9324 2004 9333
rect 2136 9324 2188 9376
rect 2688 9324 2740 9376
rect 3056 9367 3108 9376
rect 3056 9333 3065 9367
rect 3065 9333 3099 9367
rect 3099 9333 3108 9367
rect 4252 9392 4304 9444
rect 4896 9435 4948 9444
rect 4896 9401 4905 9435
rect 4905 9401 4939 9435
rect 4939 9401 4948 9435
rect 4896 9392 4948 9401
rect 9772 9392 9824 9444
rect 11244 9392 11296 9444
rect 11980 9392 12032 9444
rect 12992 9469 13026 9503
rect 13026 9469 13044 9503
rect 12992 9460 13044 9469
rect 18052 9503 18104 9512
rect 18052 9469 18061 9503
rect 18061 9469 18095 9503
rect 18095 9469 18104 9503
rect 18052 9460 18104 9469
rect 18328 9435 18380 9444
rect 18328 9401 18337 9435
rect 18337 9401 18371 9435
rect 18371 9401 18380 9435
rect 18328 9392 18380 9401
rect 3056 9324 3108 9333
rect 3792 9324 3844 9376
rect 5172 9324 5224 9376
rect 7196 9324 7248 9376
rect 9496 9324 9548 9376
rect 11336 9367 11388 9376
rect 11336 9333 11345 9367
rect 11345 9333 11379 9367
rect 11379 9333 11388 9367
rect 11336 9324 11388 9333
rect 14096 9367 14148 9376
rect 14096 9333 14105 9367
rect 14105 9333 14139 9367
rect 14139 9333 14148 9367
rect 14096 9324 14148 9333
rect 15568 9324 15620 9376
rect 16672 9324 16724 9376
rect 18696 9324 18748 9376
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 1952 9120 2004 9172
rect 2136 9120 2188 9172
rect 3516 9120 3568 9172
rect 5080 9163 5132 9172
rect 3332 9052 3384 9104
rect 3608 9052 3660 9104
rect 3148 8984 3200 9036
rect 5080 9129 5089 9163
rect 5089 9129 5123 9163
rect 5123 9129 5132 9163
rect 5080 9120 5132 9129
rect 5540 9163 5592 9172
rect 5540 9129 5549 9163
rect 5549 9129 5583 9163
rect 5583 9129 5592 9163
rect 5540 9120 5592 9129
rect 8300 9120 8352 9172
rect 9404 9163 9456 9172
rect 9404 9129 9413 9163
rect 9413 9129 9447 9163
rect 9447 9129 9456 9163
rect 9404 9120 9456 9129
rect 14832 9120 14884 9172
rect 16672 9120 16724 9172
rect 5356 9052 5408 9104
rect 6920 9052 6972 9104
rect 8208 9052 8260 9104
rect 8760 9052 8812 9104
rect 11704 9095 11756 9104
rect 1768 8780 1820 8832
rect 6092 8984 6144 9036
rect 9496 8984 9548 9036
rect 4528 8959 4580 8968
rect 4528 8925 4537 8959
rect 4537 8925 4571 8959
rect 4571 8925 4580 8959
rect 4528 8916 4580 8925
rect 4160 8891 4212 8900
rect 4160 8857 4169 8891
rect 4169 8857 4203 8891
rect 4203 8857 4212 8891
rect 4160 8848 4212 8857
rect 9128 8916 9180 8968
rect 11704 9061 11713 9095
rect 11713 9061 11747 9095
rect 11747 9061 11756 9095
rect 11704 9052 11756 9061
rect 11888 9095 11940 9104
rect 11888 9061 11897 9095
rect 11897 9061 11931 9095
rect 11931 9061 11940 9095
rect 11888 9052 11940 9061
rect 13360 9052 13412 9104
rect 15292 9052 15344 9104
rect 15660 9095 15712 9104
rect 15660 9061 15669 9095
rect 15669 9061 15703 9095
rect 15703 9061 15712 9095
rect 15660 9052 15712 9061
rect 14096 8984 14148 9036
rect 18328 9027 18380 9036
rect 18328 8993 18337 9027
rect 18337 8993 18371 9027
rect 18371 8993 18380 9027
rect 18328 8984 18380 8993
rect 11980 8959 12032 8968
rect 11980 8925 11989 8959
rect 11989 8925 12023 8959
rect 12023 8925 12032 8959
rect 11980 8916 12032 8925
rect 15936 8959 15988 8968
rect 15936 8925 15945 8959
rect 15945 8925 15979 8959
rect 15979 8925 15988 8959
rect 15936 8916 15988 8925
rect 17776 8916 17828 8968
rect 9864 8848 9916 8900
rect 11336 8848 11388 8900
rect 12256 8848 12308 8900
rect 12808 8891 12860 8900
rect 12808 8857 12817 8891
rect 12817 8857 12851 8891
rect 12851 8857 12860 8891
rect 12808 8848 12860 8857
rect 13544 8848 13596 8900
rect 3608 8780 3660 8832
rect 6368 8780 6420 8832
rect 6644 8780 6696 8832
rect 6828 8823 6880 8832
rect 6828 8789 6837 8823
rect 6837 8789 6871 8823
rect 6871 8789 6880 8823
rect 6828 8780 6880 8789
rect 9772 8823 9824 8832
rect 9772 8789 9781 8823
rect 9781 8789 9815 8823
rect 9815 8789 9824 8823
rect 9772 8780 9824 8789
rect 11244 8823 11296 8832
rect 11244 8789 11253 8823
rect 11253 8789 11287 8823
rect 11287 8789 11296 8823
rect 11244 8780 11296 8789
rect 12992 8823 13044 8832
rect 12992 8789 13001 8823
rect 13001 8789 13035 8823
rect 13035 8789 13044 8823
rect 12992 8780 13044 8789
rect 15384 8823 15436 8832
rect 15384 8789 15393 8823
rect 15393 8789 15427 8823
rect 15427 8789 15436 8823
rect 15384 8780 15436 8789
rect 19156 8780 19208 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 2872 8576 2924 8628
rect 8208 8619 8260 8628
rect 8208 8585 8217 8619
rect 8217 8585 8251 8619
rect 8251 8585 8260 8619
rect 8208 8576 8260 8585
rect 8760 8619 8812 8628
rect 8760 8585 8769 8619
rect 8769 8585 8803 8619
rect 8803 8585 8812 8619
rect 8760 8576 8812 8585
rect 9128 8619 9180 8628
rect 9128 8585 9137 8619
rect 9137 8585 9171 8619
rect 9171 8585 9180 8619
rect 9128 8576 9180 8585
rect 11704 8619 11756 8628
rect 11704 8585 11713 8619
rect 11713 8585 11747 8619
rect 11747 8585 11756 8619
rect 11704 8576 11756 8585
rect 12624 8619 12676 8628
rect 12624 8585 12633 8619
rect 12633 8585 12667 8619
rect 12667 8585 12676 8619
rect 12624 8576 12676 8585
rect 15660 8619 15712 8628
rect 15660 8585 15669 8619
rect 15669 8585 15703 8619
rect 15703 8585 15712 8619
rect 15660 8576 15712 8585
rect 15936 8576 15988 8628
rect 16672 8619 16724 8628
rect 16672 8585 16681 8619
rect 16681 8585 16715 8619
rect 16715 8585 16724 8619
rect 16672 8576 16724 8585
rect 18328 8619 18380 8628
rect 18328 8585 18337 8619
rect 18337 8585 18371 8619
rect 18371 8585 18380 8619
rect 18328 8576 18380 8585
rect 4528 8508 4580 8560
rect 8484 8508 8536 8560
rect 13360 8508 13412 8560
rect 1400 8440 1452 8492
rect 1768 8372 1820 8424
rect 5540 8372 5592 8424
rect 6828 8415 6880 8424
rect 2228 8347 2280 8356
rect 2228 8313 2237 8347
rect 2237 8313 2271 8347
rect 2271 8313 2280 8347
rect 2228 8304 2280 8313
rect 2504 8304 2556 8356
rect 3516 8347 3568 8356
rect 3516 8313 3550 8347
rect 3550 8313 3568 8347
rect 3516 8304 3568 8313
rect 5356 8304 5408 8356
rect 6092 8304 6144 8356
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 9312 8415 9364 8424
rect 9312 8381 9321 8415
rect 9321 8381 9355 8415
rect 9355 8381 9364 8415
rect 9312 8372 9364 8381
rect 6644 8304 6696 8356
rect 7288 8304 7340 8356
rect 9036 8304 9088 8356
rect 9496 8304 9548 8356
rect 11888 8304 11940 8356
rect 13636 8304 13688 8356
rect 4436 8236 4488 8288
rect 6552 8279 6604 8288
rect 6552 8245 6561 8279
rect 6561 8245 6595 8279
rect 6595 8245 6604 8279
rect 6552 8236 6604 8245
rect 10876 8236 10928 8288
rect 13544 8279 13596 8288
rect 13544 8245 13553 8279
rect 13553 8245 13587 8279
rect 13587 8245 13596 8279
rect 14096 8304 14148 8356
rect 16212 8347 16264 8356
rect 16212 8313 16221 8347
rect 16221 8313 16255 8347
rect 16255 8313 16264 8347
rect 16212 8304 16264 8313
rect 13544 8236 13596 8245
rect 14740 8236 14792 8288
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1400 8075 1452 8084
rect 1400 8041 1409 8075
rect 1409 8041 1443 8075
rect 1443 8041 1452 8075
rect 1400 8032 1452 8041
rect 1768 8032 1820 8084
rect 3608 8032 3660 8084
rect 3792 8032 3844 8084
rect 8300 8075 8352 8084
rect 8300 8041 8309 8075
rect 8309 8041 8343 8075
rect 8343 8041 8352 8075
rect 8300 8032 8352 8041
rect 11980 8032 12032 8084
rect 13820 8075 13872 8084
rect 13820 8041 13829 8075
rect 13829 8041 13863 8075
rect 13863 8041 13872 8075
rect 13820 8032 13872 8041
rect 15936 8032 15988 8084
rect 2320 7896 2372 7948
rect 4344 7964 4396 8016
rect 4620 8007 4672 8016
rect 4620 7973 4629 8007
rect 4629 7973 4663 8007
rect 4663 7973 4672 8007
rect 4620 7964 4672 7973
rect 3516 7896 3568 7948
rect 3792 7896 3844 7948
rect 4436 7896 4488 7948
rect 6552 7964 6604 8016
rect 9680 7964 9732 8016
rect 10140 7964 10192 8016
rect 6644 7896 6696 7948
rect 8392 7939 8444 7948
rect 8392 7905 8401 7939
rect 8401 7905 8435 7939
rect 8435 7905 8444 7939
rect 8392 7896 8444 7905
rect 9772 7896 9824 7948
rect 10324 8007 10376 8016
rect 10324 7973 10333 8007
rect 10333 7973 10367 8007
rect 10367 7973 10376 8007
rect 10324 7964 10376 7973
rect 10876 7964 10928 8016
rect 14740 7964 14792 8016
rect 12348 7896 12400 7948
rect 13544 7896 13596 7948
rect 16028 7896 16080 7948
rect 18328 7939 18380 7948
rect 18328 7905 18337 7939
rect 18337 7905 18371 7939
rect 18371 7905 18380 7939
rect 18328 7896 18380 7905
rect 20904 7939 20956 7948
rect 20904 7905 20913 7939
rect 20913 7905 20947 7939
rect 20947 7905 20956 7939
rect 20904 7896 20956 7905
rect 2228 7828 2280 7880
rect 3240 7828 3292 7880
rect 4528 7871 4580 7880
rect 4528 7837 4537 7871
rect 4537 7837 4571 7871
rect 4571 7837 4580 7871
rect 4528 7828 4580 7837
rect 4712 7871 4764 7880
rect 4712 7837 4721 7871
rect 4721 7837 4755 7871
rect 4755 7837 4764 7871
rect 4712 7828 4764 7837
rect 10876 7828 10928 7880
rect 11520 7871 11572 7880
rect 11520 7837 11529 7871
rect 11529 7837 11563 7871
rect 11563 7837 11572 7871
rect 11520 7828 11572 7837
rect 14372 7828 14424 7880
rect 19340 7828 19392 7880
rect 22008 7828 22060 7880
rect 3516 7803 3568 7812
rect 3516 7769 3525 7803
rect 3525 7769 3559 7803
rect 3559 7769 3568 7803
rect 3516 7760 3568 7769
rect 7012 7760 7064 7812
rect 9772 7803 9824 7812
rect 9772 7769 9781 7803
rect 9781 7769 9815 7803
rect 9815 7769 9824 7803
rect 9772 7760 9824 7769
rect 2596 7692 2648 7744
rect 2964 7692 3016 7744
rect 3792 7735 3844 7744
rect 3792 7701 3801 7735
rect 3801 7701 3835 7735
rect 3835 7701 3844 7735
rect 3792 7692 3844 7701
rect 4068 7692 4120 7744
rect 6920 7692 6972 7744
rect 7288 7735 7340 7744
rect 7288 7701 7297 7735
rect 7297 7701 7331 7735
rect 7331 7701 7340 7735
rect 7288 7692 7340 7701
rect 8024 7692 8076 7744
rect 9036 7735 9088 7744
rect 9036 7701 9045 7735
rect 9045 7701 9079 7735
rect 9079 7701 9088 7735
rect 9036 7692 9088 7701
rect 9312 7735 9364 7744
rect 9312 7701 9321 7735
rect 9321 7701 9355 7735
rect 9355 7701 9364 7735
rect 9312 7692 9364 7701
rect 11336 7692 11388 7744
rect 12900 7735 12952 7744
rect 12900 7701 12909 7735
rect 12909 7701 12943 7735
rect 12943 7701 12952 7735
rect 12900 7692 12952 7701
rect 14464 7735 14516 7744
rect 14464 7701 14473 7735
rect 14473 7701 14507 7735
rect 14507 7701 14516 7735
rect 14464 7692 14516 7701
rect 18144 7735 18196 7744
rect 18144 7701 18153 7735
rect 18153 7701 18187 7735
rect 18187 7701 18196 7735
rect 18144 7692 18196 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 2320 7531 2372 7540
rect 2320 7497 2329 7531
rect 2329 7497 2363 7531
rect 2363 7497 2372 7531
rect 2320 7488 2372 7497
rect 3608 7488 3660 7540
rect 4528 7488 4580 7540
rect 4620 7488 4672 7540
rect 6644 7531 6696 7540
rect 5264 7463 5316 7472
rect 5264 7429 5273 7463
rect 5273 7429 5307 7463
rect 5307 7429 5316 7463
rect 5264 7420 5316 7429
rect 6644 7497 6653 7531
rect 6653 7497 6687 7531
rect 6687 7497 6696 7531
rect 6644 7488 6696 7497
rect 7932 7488 7984 7540
rect 10140 7531 10192 7540
rect 10140 7497 10149 7531
rect 10149 7497 10183 7531
rect 10183 7497 10192 7531
rect 10140 7488 10192 7497
rect 12624 7531 12676 7540
rect 12624 7497 12633 7531
rect 12633 7497 12667 7531
rect 12667 7497 12676 7531
rect 12624 7488 12676 7497
rect 14832 7488 14884 7540
rect 20904 7531 20956 7540
rect 20904 7497 20913 7531
rect 20913 7497 20947 7531
rect 20947 7497 20956 7531
rect 20904 7488 20956 7497
rect 7748 7463 7800 7472
rect 7748 7429 7757 7463
rect 7757 7429 7791 7463
rect 7791 7429 7800 7463
rect 7748 7420 7800 7429
rect 9772 7420 9824 7472
rect 10324 7420 10376 7472
rect 10968 7420 11020 7472
rect 1768 7352 1820 7404
rect 2320 7352 2372 7404
rect 5724 7395 5776 7404
rect 5724 7361 5733 7395
rect 5733 7361 5767 7395
rect 5767 7361 5776 7395
rect 5724 7352 5776 7361
rect 7564 7395 7616 7404
rect 7564 7361 7573 7395
rect 7573 7361 7607 7395
rect 7607 7361 7616 7395
rect 7564 7352 7616 7361
rect 8484 7352 8536 7404
rect 10048 7352 10100 7404
rect 11336 7395 11388 7404
rect 2504 7284 2556 7336
rect 3056 7284 3108 7336
rect 1400 7191 1452 7200
rect 1400 7157 1409 7191
rect 1409 7157 1443 7191
rect 1443 7157 1452 7191
rect 1400 7148 1452 7157
rect 3240 7148 3292 7200
rect 6184 7284 6236 7336
rect 8208 7284 8260 7336
rect 9128 7284 9180 7336
rect 5816 7259 5868 7268
rect 5816 7225 5825 7259
rect 5825 7225 5859 7259
rect 5859 7225 5868 7259
rect 5816 7216 5868 7225
rect 7288 7216 7340 7268
rect 8024 7216 8076 7268
rect 9496 7216 9548 7268
rect 11336 7361 11345 7395
rect 11345 7361 11379 7395
rect 11379 7361 11388 7395
rect 11336 7352 11388 7361
rect 14740 7352 14792 7404
rect 15016 7352 15068 7404
rect 18052 7395 18104 7404
rect 10692 7284 10744 7336
rect 12440 7327 12492 7336
rect 12440 7293 12449 7327
rect 12449 7293 12483 7327
rect 12483 7293 12492 7327
rect 12440 7284 12492 7293
rect 14464 7284 14516 7336
rect 16028 7284 16080 7336
rect 11612 7216 11664 7268
rect 13820 7216 13872 7268
rect 15936 7216 15988 7268
rect 16396 7216 16448 7268
rect 18052 7361 18061 7395
rect 18061 7361 18095 7395
rect 18095 7361 18104 7395
rect 18052 7352 18104 7361
rect 18144 7284 18196 7336
rect 21364 7327 21416 7336
rect 21364 7293 21373 7327
rect 21373 7293 21407 7327
rect 21407 7293 21416 7327
rect 21364 7284 21416 7293
rect 21640 7259 21692 7268
rect 21640 7225 21649 7259
rect 21649 7225 21683 7259
rect 21683 7225 21692 7259
rect 21640 7216 21692 7225
rect 6552 7148 6604 7200
rect 7932 7148 7984 7200
rect 8760 7148 8812 7200
rect 11520 7148 11572 7200
rect 12348 7148 12400 7200
rect 12624 7148 12676 7200
rect 13544 7191 13596 7200
rect 13544 7157 13553 7191
rect 13553 7157 13587 7191
rect 13587 7157 13596 7191
rect 13544 7148 13596 7157
rect 14188 7148 14240 7200
rect 16856 7191 16908 7200
rect 16856 7157 16865 7191
rect 16865 7157 16899 7191
rect 16899 7157 16908 7191
rect 16856 7148 16908 7157
rect 19432 7191 19484 7200
rect 19432 7157 19441 7191
rect 19441 7157 19475 7191
rect 19475 7157 19484 7191
rect 19432 7148 19484 7157
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 2320 6987 2372 6996
rect 2320 6953 2329 6987
rect 2329 6953 2363 6987
rect 2363 6953 2372 6987
rect 2320 6944 2372 6953
rect 4252 6944 4304 6996
rect 6644 6987 6696 6996
rect 2688 6876 2740 6928
rect 4068 6876 4120 6928
rect 4436 6851 4488 6860
rect 4436 6817 4445 6851
rect 4445 6817 4479 6851
rect 4479 6817 4488 6851
rect 4436 6808 4488 6817
rect 4712 6919 4764 6928
rect 4712 6885 4721 6919
rect 4721 6885 4755 6919
rect 4755 6885 4764 6919
rect 4712 6876 4764 6885
rect 5816 6876 5868 6928
rect 6644 6953 6653 6987
rect 6653 6953 6687 6987
rect 6687 6953 6696 6987
rect 6644 6944 6696 6953
rect 7748 6987 7800 6996
rect 7748 6953 7757 6987
rect 7757 6953 7791 6987
rect 7791 6953 7800 6987
rect 7748 6944 7800 6953
rect 9036 6944 9088 6996
rect 9864 6944 9916 6996
rect 13912 6987 13964 6996
rect 13912 6953 13921 6987
rect 13921 6953 13955 6987
rect 13955 6953 13964 6987
rect 13912 6944 13964 6953
rect 15016 6987 15068 6996
rect 15016 6953 15025 6987
rect 15025 6953 15059 6987
rect 15059 6953 15068 6987
rect 15016 6944 15068 6953
rect 15936 6987 15988 6996
rect 15936 6953 15945 6987
rect 15945 6953 15979 6987
rect 15979 6953 15988 6987
rect 15936 6944 15988 6953
rect 18328 6987 18380 6996
rect 18328 6953 18337 6987
rect 18337 6953 18371 6987
rect 18371 6953 18380 6987
rect 18328 6944 18380 6953
rect 6000 6808 6052 6860
rect 7380 6876 7432 6928
rect 7840 6876 7892 6928
rect 11336 6876 11388 6928
rect 7656 6808 7708 6860
rect 10048 6851 10100 6860
rect 10048 6817 10057 6851
rect 10057 6817 10091 6851
rect 10091 6817 10100 6851
rect 10048 6808 10100 6817
rect 10692 6851 10744 6860
rect 10692 6817 10701 6851
rect 10701 6817 10735 6851
rect 10735 6817 10744 6851
rect 10692 6808 10744 6817
rect 13176 6851 13228 6860
rect 13176 6817 13185 6851
rect 13185 6817 13219 6851
rect 13219 6817 13228 6851
rect 13176 6808 13228 6817
rect 13728 6851 13780 6860
rect 13728 6817 13737 6851
rect 13737 6817 13771 6851
rect 13771 6817 13780 6851
rect 13728 6808 13780 6817
rect 14832 6808 14884 6860
rect 16304 6851 16356 6860
rect 16304 6817 16313 6851
rect 16313 6817 16347 6851
rect 16347 6817 16356 6851
rect 16856 6876 16908 6928
rect 16304 6808 16356 6817
rect 19340 6808 19392 6860
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 2872 6740 2924 6792
rect 3056 6783 3108 6792
rect 3056 6749 3065 6783
rect 3065 6749 3099 6783
rect 3099 6749 3108 6783
rect 3056 6740 3108 6749
rect 3792 6740 3844 6792
rect 4712 6740 4764 6792
rect 5172 6740 5224 6792
rect 7748 6783 7800 6792
rect 7748 6749 7757 6783
rect 7757 6749 7791 6783
rect 7791 6749 7800 6783
rect 7748 6740 7800 6749
rect 8392 6740 8444 6792
rect 10140 6740 10192 6792
rect 11060 6783 11112 6792
rect 11060 6749 11069 6783
rect 11069 6749 11103 6783
rect 11103 6749 11112 6783
rect 11060 6740 11112 6749
rect 16396 6783 16448 6792
rect 4160 6715 4212 6724
rect 4160 6681 4169 6715
rect 4169 6681 4203 6715
rect 4203 6681 4212 6715
rect 4160 6672 4212 6681
rect 5724 6715 5776 6724
rect 5724 6681 5733 6715
rect 5733 6681 5767 6715
rect 5767 6681 5776 6715
rect 5724 6672 5776 6681
rect 9312 6672 9364 6724
rect 16396 6749 16405 6783
rect 16405 6749 16439 6783
rect 16439 6749 16448 6783
rect 16396 6740 16448 6749
rect 15476 6715 15528 6724
rect 1952 6647 2004 6656
rect 1952 6613 1961 6647
rect 1961 6613 1995 6647
rect 1995 6613 2004 6647
rect 1952 6604 2004 6613
rect 2964 6604 3016 6656
rect 7104 6647 7156 6656
rect 7104 6613 7113 6647
rect 7113 6613 7147 6647
rect 7147 6613 7156 6647
rect 7104 6604 7156 6613
rect 7380 6604 7432 6656
rect 8208 6604 8260 6656
rect 10692 6604 10744 6656
rect 15476 6681 15485 6715
rect 15485 6681 15519 6715
rect 15519 6681 15528 6715
rect 15476 6672 15528 6681
rect 18144 6672 18196 6724
rect 11520 6604 11572 6656
rect 12624 6647 12676 6656
rect 12624 6613 12633 6647
rect 12633 6613 12667 6647
rect 12667 6613 12676 6647
rect 12624 6604 12676 6613
rect 13084 6604 13136 6656
rect 14280 6647 14332 6656
rect 14280 6613 14289 6647
rect 14289 6613 14323 6647
rect 14323 6613 14332 6647
rect 14280 6604 14332 6613
rect 14648 6647 14700 6656
rect 14648 6613 14657 6647
rect 14657 6613 14691 6647
rect 14691 6613 14700 6647
rect 14648 6604 14700 6613
rect 20628 6604 20680 6656
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 2320 6400 2372 6452
rect 4252 6443 4304 6452
rect 4252 6409 4261 6443
rect 4261 6409 4295 6443
rect 4295 6409 4304 6443
rect 4252 6400 4304 6409
rect 5172 6443 5224 6452
rect 5172 6409 5181 6443
rect 5181 6409 5215 6443
rect 5215 6409 5224 6443
rect 5172 6400 5224 6409
rect 6000 6443 6052 6452
rect 6000 6409 6009 6443
rect 6009 6409 6043 6443
rect 6043 6409 6052 6443
rect 6000 6400 6052 6409
rect 9312 6443 9364 6452
rect 1584 6239 1636 6248
rect 1584 6205 1593 6239
rect 1593 6205 1627 6239
rect 1627 6205 1636 6239
rect 1584 6196 1636 6205
rect 2504 6196 2556 6248
rect 5356 6239 5408 6248
rect 5356 6205 5365 6239
rect 5365 6205 5399 6239
rect 5399 6205 5408 6239
rect 5356 6196 5408 6205
rect 9312 6409 9321 6443
rect 9321 6409 9355 6443
rect 9355 6409 9364 6443
rect 9312 6400 9364 6409
rect 11336 6400 11388 6452
rect 12808 6400 12860 6452
rect 13452 6400 13504 6452
rect 15384 6400 15436 6452
rect 16396 6400 16448 6452
rect 17776 6443 17828 6452
rect 17776 6409 17785 6443
rect 17785 6409 17819 6443
rect 17819 6409 17828 6443
rect 17776 6400 17828 6409
rect 19340 6400 19392 6452
rect 15292 6332 15344 6384
rect 18144 6375 18196 6384
rect 2964 6128 3016 6180
rect 3148 6171 3200 6180
rect 3148 6137 3182 6171
rect 3182 6137 3200 6171
rect 3148 6128 3200 6137
rect 7288 6239 7340 6248
rect 7288 6205 7322 6239
rect 7322 6205 7340 6239
rect 7288 6196 7340 6205
rect 8024 6196 8076 6248
rect 9772 6239 9824 6248
rect 9772 6205 9806 6239
rect 9806 6205 9824 6239
rect 9772 6196 9824 6205
rect 11520 6239 11572 6248
rect 11520 6205 11529 6239
rect 11529 6205 11563 6239
rect 11563 6205 11572 6239
rect 11520 6196 11572 6205
rect 12532 6196 12584 6248
rect 12808 6239 12860 6248
rect 12808 6205 12817 6239
rect 12817 6205 12851 6239
rect 12851 6205 12860 6239
rect 12808 6196 12860 6205
rect 16304 6307 16356 6316
rect 16304 6273 16313 6307
rect 16313 6273 16347 6307
rect 16347 6273 16356 6307
rect 16304 6264 16356 6273
rect 13544 6196 13596 6248
rect 18144 6341 18153 6375
rect 18153 6341 18187 6375
rect 18187 6341 18196 6375
rect 18144 6332 18196 6341
rect 25504 6375 25556 6384
rect 25504 6341 25513 6375
rect 25513 6341 25547 6375
rect 25547 6341 25556 6375
rect 25504 6332 25556 6341
rect 18236 6264 18288 6316
rect 17776 6128 17828 6180
rect 19432 6196 19484 6248
rect 24124 6239 24176 6248
rect 24124 6205 24133 6239
rect 24133 6205 24167 6239
rect 24167 6205 24176 6239
rect 24124 6196 24176 6205
rect 24768 6196 24820 6248
rect 20904 6128 20956 6180
rect 4712 6060 4764 6112
rect 6000 6060 6052 6112
rect 6552 6103 6604 6112
rect 6552 6069 6561 6103
rect 6561 6069 6595 6103
rect 6595 6069 6604 6103
rect 6552 6060 6604 6069
rect 8392 6103 8444 6112
rect 8392 6069 8401 6103
rect 8401 6069 8435 6103
rect 8435 6069 8444 6103
rect 8392 6060 8444 6069
rect 10876 6103 10928 6112
rect 10876 6069 10885 6103
rect 10885 6069 10919 6103
rect 10919 6069 10928 6103
rect 10876 6060 10928 6069
rect 14280 6060 14332 6112
rect 14832 6060 14884 6112
rect 15384 6060 15436 6112
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 2044 5856 2096 5908
rect 2320 5856 2372 5908
rect 4252 5856 4304 5908
rect 6828 5856 6880 5908
rect 7104 5856 7156 5908
rect 9772 5856 9824 5908
rect 10140 5856 10192 5908
rect 11520 5856 11572 5908
rect 18236 5856 18288 5908
rect 24124 5899 24176 5908
rect 24124 5865 24133 5899
rect 24133 5865 24167 5899
rect 24167 5865 24176 5899
rect 24124 5856 24176 5865
rect 1400 5788 1452 5840
rect 2964 5831 3016 5840
rect 2964 5797 2973 5831
rect 2973 5797 3007 5831
rect 3007 5797 3016 5831
rect 2964 5788 3016 5797
rect 1308 5720 1360 5772
rect 7012 5788 7064 5840
rect 7564 5831 7616 5840
rect 7564 5797 7573 5831
rect 7573 5797 7607 5831
rect 7607 5797 7616 5831
rect 7564 5788 7616 5797
rect 7656 5788 7708 5840
rect 4160 5720 4212 5772
rect 5448 5720 5500 5772
rect 6736 5720 6788 5772
rect 8392 5720 8444 5772
rect 9312 5720 9364 5772
rect 10048 5720 10100 5772
rect 10876 5788 10928 5840
rect 11060 5788 11112 5840
rect 12072 5788 12124 5840
rect 13544 5831 13596 5840
rect 13544 5797 13553 5831
rect 13553 5797 13587 5831
rect 13587 5797 13596 5831
rect 13544 5788 13596 5797
rect 13820 5788 13872 5840
rect 15292 5788 15344 5840
rect 13268 5763 13320 5772
rect 13268 5729 13277 5763
rect 13277 5729 13311 5763
rect 13311 5729 13320 5763
rect 13268 5720 13320 5729
rect 13912 5720 13964 5772
rect 1952 5652 2004 5704
rect 2688 5584 2740 5636
rect 4252 5652 4304 5704
rect 7196 5652 7248 5704
rect 14832 5652 14884 5704
rect 15936 5720 15988 5772
rect 16396 5720 16448 5772
rect 18144 5720 18196 5772
rect 18972 5720 19024 5772
rect 20904 5763 20956 5772
rect 20904 5729 20913 5763
rect 20913 5729 20947 5763
rect 20947 5729 20956 5763
rect 20904 5720 20956 5729
rect 17592 5695 17644 5704
rect 17592 5661 17601 5695
rect 17601 5661 17635 5695
rect 17635 5661 17644 5695
rect 17592 5652 17644 5661
rect 18788 5695 18840 5704
rect 18788 5661 18797 5695
rect 18797 5661 18831 5695
rect 18831 5661 18840 5695
rect 18788 5652 18840 5661
rect 19800 5695 19852 5704
rect 19800 5661 19809 5695
rect 19809 5661 19843 5695
rect 19843 5661 19852 5695
rect 19800 5652 19852 5661
rect 4068 5584 4120 5636
rect 6920 5584 6972 5636
rect 11980 5584 12032 5636
rect 13728 5584 13780 5636
rect 3884 5516 3936 5568
rect 4436 5516 4488 5568
rect 5356 5516 5408 5568
rect 6736 5559 6788 5568
rect 6736 5525 6745 5559
rect 6745 5525 6779 5559
rect 6779 5525 6788 5559
rect 6736 5516 6788 5525
rect 8484 5516 8536 5568
rect 9404 5559 9456 5568
rect 9404 5525 9413 5559
rect 9413 5525 9447 5559
rect 9447 5525 9456 5559
rect 9404 5516 9456 5525
rect 11152 5516 11204 5568
rect 12624 5516 12676 5568
rect 13452 5516 13504 5568
rect 15476 5516 15528 5568
rect 21088 5559 21140 5568
rect 21088 5525 21097 5559
rect 21097 5525 21131 5559
rect 21131 5525 21140 5559
rect 21088 5516 21140 5525
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 2044 5312 2096 5364
rect 3148 5312 3200 5364
rect 4160 5312 4212 5364
rect 4620 5355 4672 5364
rect 4620 5321 4629 5355
rect 4629 5321 4663 5355
rect 4663 5321 4672 5355
rect 4620 5312 4672 5321
rect 4344 5244 4396 5296
rect 5264 5287 5316 5296
rect 2044 5040 2096 5092
rect 2320 5040 2372 5092
rect 4160 5040 4212 5092
rect 5264 5253 5273 5287
rect 5273 5253 5307 5287
rect 5307 5253 5316 5287
rect 5264 5244 5316 5253
rect 7288 5312 7340 5364
rect 10048 5312 10100 5364
rect 10784 5312 10836 5364
rect 11060 5355 11112 5364
rect 11060 5321 11069 5355
rect 11069 5321 11103 5355
rect 11103 5321 11112 5355
rect 11060 5312 11112 5321
rect 11888 5312 11940 5364
rect 13820 5355 13872 5364
rect 13820 5321 13829 5355
rect 13829 5321 13863 5355
rect 13863 5321 13872 5355
rect 13820 5312 13872 5321
rect 13912 5312 13964 5364
rect 14832 5355 14884 5364
rect 14832 5321 14841 5355
rect 14841 5321 14875 5355
rect 14875 5321 14884 5355
rect 14832 5312 14884 5321
rect 16396 5312 16448 5364
rect 18972 5355 19024 5364
rect 18972 5321 18981 5355
rect 18981 5321 19015 5355
rect 19015 5321 19024 5355
rect 18972 5312 19024 5321
rect 20904 5312 20956 5364
rect 9680 5287 9732 5296
rect 9680 5253 9689 5287
rect 9689 5253 9723 5287
rect 9723 5253 9732 5287
rect 9680 5244 9732 5253
rect 6552 5176 6604 5228
rect 11520 5176 11572 5228
rect 10692 5108 10744 5160
rect 10784 5108 10836 5160
rect 11244 5108 11296 5160
rect 6736 5040 6788 5092
rect 10140 5083 10192 5092
rect 10140 5049 10149 5083
rect 10149 5049 10183 5083
rect 10183 5049 10192 5083
rect 12348 5108 12400 5160
rect 10140 5040 10192 5049
rect 15476 5108 15528 5160
rect 17592 5151 17644 5160
rect 17592 5117 17601 5151
rect 17601 5117 17635 5151
rect 17635 5117 17644 5151
rect 17592 5108 17644 5117
rect 18328 5108 18380 5160
rect 18696 5108 18748 5160
rect 20260 5151 20312 5160
rect 20260 5117 20269 5151
rect 20269 5117 20303 5151
rect 20303 5117 20312 5151
rect 20260 5108 20312 5117
rect 21364 5151 21416 5160
rect 21364 5117 21373 5151
rect 21373 5117 21407 5151
rect 21407 5117 21416 5151
rect 21364 5108 21416 5117
rect 22100 5108 22152 5160
rect 6552 5015 6604 5024
rect 6552 4981 6561 5015
rect 6561 4981 6595 5015
rect 6595 4981 6604 5015
rect 6552 4972 6604 4981
rect 7472 4972 7524 5024
rect 9036 5015 9088 5024
rect 9036 4981 9045 5015
rect 9045 4981 9079 5015
rect 9079 4981 9088 5015
rect 9036 4972 9088 4981
rect 11428 4972 11480 5024
rect 12072 4972 12124 5024
rect 12624 4972 12676 5024
rect 16212 4972 16264 5024
rect 17224 5015 17276 5024
rect 17224 4981 17233 5015
rect 17233 4981 17267 5015
rect 17267 4981 17276 5015
rect 17224 4972 17276 4981
rect 18236 5015 18288 5024
rect 18236 4981 18245 5015
rect 18245 4981 18279 5015
rect 18279 4981 18288 5015
rect 18236 4972 18288 4981
rect 19248 4972 19300 5024
rect 20076 4972 20128 5024
rect 22008 5040 22060 5092
rect 23572 4972 23624 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1400 4811 1452 4820
rect 1400 4777 1409 4811
rect 1409 4777 1443 4811
rect 1443 4777 1452 4811
rect 1400 4768 1452 4777
rect 3792 4811 3844 4820
rect 3792 4777 3801 4811
rect 3801 4777 3835 4811
rect 3835 4777 3844 4811
rect 3792 4768 3844 4777
rect 4068 4768 4120 4820
rect 6736 4811 6788 4820
rect 6736 4777 6745 4811
rect 6745 4777 6779 4811
rect 6779 4777 6788 4811
rect 6736 4768 6788 4777
rect 7380 4811 7432 4820
rect 7380 4777 7389 4811
rect 7389 4777 7423 4811
rect 7423 4777 7432 4811
rect 7380 4768 7432 4777
rect 7564 4768 7616 4820
rect 8576 4811 8628 4820
rect 8576 4777 8585 4811
rect 8585 4777 8619 4811
rect 8619 4777 8628 4811
rect 8576 4768 8628 4777
rect 9496 4768 9548 4820
rect 9864 4768 9916 4820
rect 11152 4768 11204 4820
rect 11704 4768 11756 4820
rect 12532 4811 12584 4820
rect 12532 4777 12541 4811
rect 12541 4777 12575 4811
rect 12575 4777 12584 4811
rect 12532 4768 12584 4777
rect 3056 4700 3108 4752
rect 2872 4607 2924 4616
rect 2872 4573 2881 4607
rect 2881 4573 2915 4607
rect 2915 4573 2924 4607
rect 2872 4564 2924 4573
rect 2964 4564 3016 4616
rect 5356 4700 5408 4752
rect 6920 4700 6972 4752
rect 7472 4743 7524 4752
rect 7472 4709 7481 4743
rect 7481 4709 7515 4743
rect 7515 4709 7524 4743
rect 7472 4700 7524 4709
rect 10232 4743 10284 4752
rect 10232 4709 10241 4743
rect 10241 4709 10275 4743
rect 10275 4709 10284 4743
rect 10232 4700 10284 4709
rect 11336 4700 11388 4752
rect 11888 4743 11940 4752
rect 11888 4709 11897 4743
rect 11897 4709 11931 4743
rect 11931 4709 11940 4743
rect 13452 4743 13504 4752
rect 11888 4700 11940 4709
rect 13452 4709 13461 4743
rect 13461 4709 13495 4743
rect 13495 4709 13504 4743
rect 13452 4700 13504 4709
rect 15108 4811 15160 4820
rect 15108 4777 15117 4811
rect 15117 4777 15151 4811
rect 15151 4777 15160 4811
rect 15108 4768 15160 4777
rect 15752 4811 15804 4820
rect 15752 4777 15761 4811
rect 15761 4777 15795 4811
rect 15795 4777 15804 4811
rect 15752 4768 15804 4777
rect 15844 4768 15896 4820
rect 17868 4811 17920 4820
rect 17868 4777 17877 4811
rect 17877 4777 17911 4811
rect 17911 4777 17920 4811
rect 17868 4768 17920 4777
rect 18236 4743 18288 4752
rect 18236 4709 18245 4743
rect 18245 4709 18279 4743
rect 18279 4709 18288 4743
rect 18236 4700 18288 4709
rect 18604 4700 18656 4752
rect 4160 4632 4212 4684
rect 8392 4675 8444 4684
rect 8392 4641 8401 4675
rect 8401 4641 8435 4675
rect 8435 4641 8444 4675
rect 8392 4632 8444 4641
rect 10416 4632 10468 4684
rect 15936 4675 15988 4684
rect 15936 4641 15945 4675
rect 15945 4641 15979 4675
rect 15979 4641 15988 4675
rect 15936 4632 15988 4641
rect 16212 4675 16264 4684
rect 16212 4641 16246 4675
rect 16246 4641 16264 4675
rect 16212 4632 16264 4641
rect 20996 4632 21048 4684
rect 22468 4675 22520 4684
rect 22468 4641 22477 4675
rect 22477 4641 22511 4675
rect 22511 4641 22520 4675
rect 22468 4632 22520 4641
rect 23756 4675 23808 4684
rect 23756 4641 23765 4675
rect 23765 4641 23799 4675
rect 23799 4641 23808 4675
rect 23756 4632 23808 4641
rect 13360 4607 13412 4616
rect 2780 4496 2832 4548
rect 9404 4496 9456 4548
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 14648 4607 14700 4616
rect 14648 4573 14657 4607
rect 14657 4573 14691 4607
rect 14691 4573 14700 4607
rect 14648 4564 14700 4573
rect 18880 4607 18932 4616
rect 18880 4573 18889 4607
rect 18889 4573 18923 4607
rect 18923 4573 18932 4607
rect 18880 4564 18932 4573
rect 19064 4607 19116 4616
rect 19064 4573 19073 4607
rect 19073 4573 19107 4607
rect 19107 4573 19116 4607
rect 19064 4564 19116 4573
rect 13728 4496 13780 4548
rect 2320 4428 2372 4480
rect 2596 4428 2648 4480
rect 6000 4471 6052 4480
rect 6000 4437 6009 4471
rect 6009 4437 6043 4471
rect 6043 4437 6052 4471
rect 6000 4428 6052 4437
rect 6920 4471 6972 4480
rect 6920 4437 6929 4471
rect 6929 4437 6963 4471
rect 6963 4437 6972 4471
rect 6920 4428 6972 4437
rect 8300 4471 8352 4480
rect 8300 4437 8309 4471
rect 8309 4437 8343 4471
rect 8343 4437 8352 4471
rect 8300 4428 8352 4437
rect 9588 4428 9640 4480
rect 10140 4428 10192 4480
rect 11336 4471 11388 4480
rect 11336 4437 11345 4471
rect 11345 4437 11379 4471
rect 11379 4437 11388 4471
rect 11336 4428 11388 4437
rect 13084 4428 13136 4480
rect 17316 4471 17368 4480
rect 17316 4437 17325 4471
rect 17325 4437 17359 4471
rect 17359 4437 17368 4471
rect 17316 4428 17368 4437
rect 18512 4471 18564 4480
rect 18512 4437 18521 4471
rect 18521 4437 18555 4471
rect 18555 4437 18564 4471
rect 18512 4428 18564 4437
rect 20904 4428 20956 4480
rect 25412 4428 25464 4480
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 6184 4224 6236 4276
rect 7472 4224 7524 4276
rect 7748 4267 7800 4276
rect 7748 4233 7757 4267
rect 7757 4233 7791 4267
rect 7791 4233 7800 4267
rect 7748 4224 7800 4233
rect 9312 4267 9364 4276
rect 9312 4233 9321 4267
rect 9321 4233 9355 4267
rect 9355 4233 9364 4267
rect 9312 4224 9364 4233
rect 10416 4224 10468 4276
rect 11244 4224 11296 4276
rect 11704 4224 11756 4276
rect 12808 4224 12860 4276
rect 13360 4224 13412 4276
rect 15936 4224 15988 4276
rect 16764 4267 16816 4276
rect 16764 4233 16773 4267
rect 16773 4233 16807 4267
rect 16807 4233 16816 4267
rect 16764 4224 16816 4233
rect 18880 4267 18932 4276
rect 18880 4233 18889 4267
rect 18889 4233 18923 4267
rect 18923 4233 18932 4267
rect 18880 4224 18932 4233
rect 19064 4224 19116 4276
rect 22468 4224 22520 4276
rect 23756 4224 23808 4276
rect 2872 4156 2924 4208
rect 3056 4199 3108 4208
rect 3056 4165 3065 4199
rect 3065 4165 3099 4199
rect 3099 4165 3108 4199
rect 3056 4156 3108 4165
rect 7288 4156 7340 4208
rect 8024 4156 8076 4208
rect 2964 4088 3016 4140
rect 7104 4088 7156 4140
rect 7380 4088 7432 4140
rect 9588 4156 9640 4208
rect 10876 4199 10928 4208
rect 10876 4165 10885 4199
rect 10885 4165 10919 4199
rect 10919 4165 10928 4199
rect 10876 4156 10928 4165
rect 1676 4020 1728 4072
rect 2320 3952 2372 4004
rect 5540 4063 5592 4072
rect 5540 4029 5549 4063
rect 5549 4029 5583 4063
rect 5583 4029 5592 4063
rect 5540 4020 5592 4029
rect 10048 4088 10100 4140
rect 11152 4088 11204 4140
rect 12164 4131 12216 4140
rect 12164 4097 12173 4131
rect 12173 4097 12207 4131
rect 12207 4097 12216 4131
rect 12164 4088 12216 4097
rect 13084 4131 13136 4140
rect 13084 4097 13093 4131
rect 13093 4097 13127 4131
rect 13127 4097 13136 4131
rect 13084 4088 13136 4097
rect 2780 3952 2832 4004
rect 4068 3952 4120 4004
rect 4804 3952 4856 4004
rect 5816 3995 5868 4004
rect 5816 3961 5825 3995
rect 5825 3961 5859 3995
rect 5859 3961 5868 3995
rect 5816 3952 5868 3961
rect 7656 3952 7708 4004
rect 9772 4020 9824 4072
rect 10140 4020 10192 4072
rect 8392 3952 8444 4004
rect 9220 3952 9272 4004
rect 9404 3952 9456 4004
rect 10232 3952 10284 4004
rect 10876 3952 10928 4004
rect 11336 3995 11388 4004
rect 1400 3884 1452 3936
rect 2872 3884 2924 3936
rect 3700 3927 3752 3936
rect 3700 3893 3733 3927
rect 3733 3893 3752 3927
rect 3700 3884 3752 3893
rect 5080 3884 5132 3936
rect 5264 3927 5316 3936
rect 5264 3893 5297 3927
rect 5297 3893 5316 3927
rect 5264 3884 5316 3893
rect 5724 3927 5776 3936
rect 5724 3893 5733 3927
rect 5733 3893 5767 3927
rect 5767 3893 5776 3927
rect 5724 3884 5776 3893
rect 9772 3927 9824 3936
rect 9772 3893 9781 3927
rect 9781 3893 9815 3927
rect 9815 3893 9824 3927
rect 9772 3884 9824 3893
rect 11060 3884 11112 3936
rect 11336 3961 11345 3995
rect 11345 3961 11379 3995
rect 11379 3961 11388 3995
rect 11336 3952 11388 3961
rect 12992 3995 13044 4004
rect 12992 3961 13001 3995
rect 13001 3961 13035 3995
rect 13035 3961 13044 3995
rect 12992 3952 13044 3961
rect 14188 4088 14240 4140
rect 14464 4088 14516 4140
rect 15476 4156 15528 4208
rect 16948 4088 17000 4140
rect 17776 4131 17828 4140
rect 17776 4097 17785 4131
rect 17785 4097 17819 4131
rect 17819 4097 17828 4131
rect 17776 4088 17828 4097
rect 18328 4131 18380 4140
rect 18328 4097 18337 4131
rect 18337 4097 18371 4131
rect 18371 4097 18380 4131
rect 18328 4088 18380 4097
rect 14004 4020 14056 4072
rect 15752 4020 15804 4072
rect 17132 4063 17184 4072
rect 17132 4029 17141 4063
rect 17141 4029 17175 4063
rect 17175 4029 17184 4063
rect 17132 4020 17184 4029
rect 19340 4063 19392 4072
rect 19340 4029 19349 4063
rect 19349 4029 19383 4063
rect 19383 4029 19392 4063
rect 19340 4020 19392 4029
rect 20260 4020 20312 4072
rect 21732 4063 21784 4072
rect 21732 4029 21741 4063
rect 21741 4029 21775 4063
rect 21775 4029 21784 4063
rect 21732 4020 21784 4029
rect 23664 4063 23716 4072
rect 23664 4029 23673 4063
rect 23673 4029 23707 4063
rect 23707 4029 23716 4063
rect 23664 4020 23716 4029
rect 24768 4063 24820 4072
rect 24768 4029 24777 4063
rect 24777 4029 24811 4063
rect 24811 4029 24820 4063
rect 24768 4020 24820 4029
rect 15936 3952 15988 4004
rect 17316 3952 17368 4004
rect 18696 3952 18748 4004
rect 22008 3995 22060 4004
rect 12716 3884 12768 3936
rect 14188 3884 14240 3936
rect 14648 3884 14700 3936
rect 15384 3884 15436 3936
rect 19524 3927 19576 3936
rect 19524 3893 19533 3927
rect 19533 3893 19567 3927
rect 19567 3893 19576 3927
rect 19524 3884 19576 3893
rect 20260 3927 20312 3936
rect 20260 3893 20269 3927
rect 20269 3893 20303 3927
rect 20303 3893 20312 3927
rect 20260 3884 20312 3893
rect 22008 3961 22017 3995
rect 22017 3961 22051 3995
rect 22051 3961 22060 3995
rect 22008 3952 22060 3961
rect 20996 3927 21048 3936
rect 20996 3893 21005 3927
rect 21005 3893 21039 3927
rect 21039 3893 21048 3927
rect 20996 3884 21048 3893
rect 24124 3884 24176 3936
rect 25964 3884 26016 3936
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1676 3680 1728 3732
rect 2412 3680 2464 3732
rect 2596 3680 2648 3732
rect 3056 3680 3108 3732
rect 7104 3723 7156 3732
rect 2964 3655 3016 3664
rect 2964 3621 2973 3655
rect 2973 3621 3007 3655
rect 3007 3621 3016 3655
rect 2964 3612 3016 3621
rect 3240 3612 3292 3664
rect 4620 3655 4672 3664
rect 4620 3621 4629 3655
rect 4629 3621 4663 3655
rect 4663 3621 4672 3655
rect 4620 3612 4672 3621
rect 5816 3612 5868 3664
rect 6276 3612 6328 3664
rect 7104 3689 7113 3723
rect 7113 3689 7147 3723
rect 7147 3689 7156 3723
rect 7104 3680 7156 3689
rect 8024 3723 8076 3732
rect 8024 3689 8033 3723
rect 8033 3689 8067 3723
rect 8067 3689 8076 3723
rect 8024 3680 8076 3689
rect 9404 3680 9456 3732
rect 11060 3680 11112 3732
rect 8668 3612 8720 3664
rect 9864 3612 9916 3664
rect 10140 3612 10192 3664
rect 11796 3680 11848 3732
rect 12532 3723 12584 3732
rect 12532 3689 12541 3723
rect 12541 3689 12575 3723
rect 12575 3689 12584 3723
rect 12532 3680 12584 3689
rect 13268 3723 13320 3732
rect 13268 3689 13277 3723
rect 13277 3689 13311 3723
rect 13311 3689 13320 3723
rect 13268 3680 13320 3689
rect 14004 3723 14056 3732
rect 14004 3689 14013 3723
rect 14013 3689 14047 3723
rect 14047 3689 14056 3723
rect 14004 3680 14056 3689
rect 14464 3723 14516 3732
rect 14464 3689 14473 3723
rect 14473 3689 14507 3723
rect 14507 3689 14516 3723
rect 14464 3680 14516 3689
rect 16212 3680 16264 3732
rect 16304 3680 16356 3732
rect 16948 3680 17000 3732
rect 19432 3680 19484 3732
rect 19984 3723 20036 3732
rect 19984 3689 19993 3723
rect 19993 3689 20027 3723
rect 20027 3689 20036 3723
rect 19984 3680 20036 3689
rect 11612 3612 11664 3664
rect 14740 3655 14792 3664
rect 14740 3621 14749 3655
rect 14749 3621 14783 3655
rect 14783 3621 14792 3655
rect 14740 3612 14792 3621
rect 17316 3612 17368 3664
rect 18512 3612 18564 3664
rect 24768 3612 24820 3664
rect 2780 3544 2832 3596
rect 5632 3544 5684 3596
rect 6828 3544 6880 3596
rect 8208 3587 8260 3596
rect 8208 3553 8217 3587
rect 8217 3553 8251 3587
rect 8251 3553 8260 3587
rect 8208 3544 8260 3553
rect 14372 3544 14424 3596
rect 15844 3544 15896 3596
rect 16764 3587 16816 3596
rect 16764 3553 16773 3587
rect 16773 3553 16807 3587
rect 16807 3553 16816 3587
rect 16764 3544 16816 3553
rect 18420 3544 18472 3596
rect 19984 3544 20036 3596
rect 20720 3544 20772 3596
rect 21640 3544 21692 3596
rect 22744 3587 22796 3596
rect 22744 3553 22753 3587
rect 22753 3553 22787 3587
rect 22787 3553 22796 3587
rect 22744 3544 22796 3553
rect 24032 3587 24084 3596
rect 24032 3553 24041 3587
rect 24041 3553 24075 3587
rect 24075 3553 24084 3587
rect 24032 3544 24084 3553
rect 25136 3587 25188 3596
rect 25136 3553 25145 3587
rect 25145 3553 25179 3587
rect 25179 3553 25188 3587
rect 25136 3544 25188 3553
rect 2228 3476 2280 3528
rect 2964 3519 3016 3528
rect 2964 3485 2973 3519
rect 2973 3485 3007 3519
rect 3007 3485 3016 3519
rect 2964 3476 3016 3485
rect 4712 3519 4764 3528
rect 4712 3485 4721 3519
rect 4721 3485 4755 3519
rect 4755 3485 4764 3519
rect 4712 3476 4764 3485
rect 5080 3476 5132 3528
rect 11796 3519 11848 3528
rect 11796 3485 11805 3519
rect 11805 3485 11839 3519
rect 11839 3485 11848 3519
rect 11796 3476 11848 3485
rect 12716 3476 12768 3528
rect 13360 3519 13412 3528
rect 13360 3485 13369 3519
rect 13369 3485 13403 3519
rect 13403 3485 13412 3519
rect 13360 3476 13412 3485
rect 15568 3519 15620 3528
rect 15568 3485 15577 3519
rect 15577 3485 15611 3519
rect 15611 3485 15620 3519
rect 15568 3476 15620 3485
rect 20812 3476 20864 3528
rect 20996 3476 21048 3528
rect 2504 3451 2556 3460
rect 2504 3417 2513 3451
rect 2513 3417 2547 3451
rect 2547 3417 2556 3451
rect 2504 3408 2556 3417
rect 3056 3408 3108 3460
rect 3884 3408 3936 3460
rect 4160 3383 4212 3392
rect 4160 3349 4169 3383
rect 4169 3349 4203 3383
rect 4203 3349 4212 3383
rect 4160 3340 4212 3349
rect 5080 3383 5132 3392
rect 5080 3349 5089 3383
rect 5089 3349 5123 3383
rect 5123 3349 5132 3383
rect 5080 3340 5132 3349
rect 13268 3408 13320 3460
rect 7656 3383 7708 3392
rect 7656 3349 7665 3383
rect 7665 3349 7699 3383
rect 7699 3349 7708 3383
rect 7656 3340 7708 3349
rect 9588 3340 9640 3392
rect 12808 3383 12860 3392
rect 12808 3349 12817 3383
rect 12817 3349 12851 3383
rect 12851 3349 12860 3383
rect 12808 3340 12860 3349
rect 17960 3340 18012 3392
rect 20168 3383 20220 3392
rect 20168 3349 20177 3383
rect 20177 3349 20211 3383
rect 20211 3349 20220 3383
rect 20168 3340 20220 3349
rect 20812 3340 20864 3392
rect 23204 3340 23256 3392
rect 24952 3340 25004 3392
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 4068 3136 4120 3188
rect 5540 3136 5592 3188
rect 9128 3179 9180 3188
rect 9128 3145 9137 3179
rect 9137 3145 9171 3179
rect 9171 3145 9180 3179
rect 9128 3136 9180 3145
rect 10692 3136 10744 3188
rect 10968 3179 11020 3188
rect 10968 3145 10977 3179
rect 10977 3145 11011 3179
rect 11011 3145 11020 3179
rect 10968 3136 11020 3145
rect 11612 3179 11664 3188
rect 11612 3145 11621 3179
rect 11621 3145 11655 3179
rect 11655 3145 11664 3179
rect 11612 3136 11664 3145
rect 11888 3179 11940 3188
rect 11888 3145 11897 3179
rect 11897 3145 11931 3179
rect 11931 3145 11940 3179
rect 11888 3136 11940 3145
rect 13360 3136 13412 3188
rect 13820 3179 13872 3188
rect 13820 3145 13829 3179
rect 13829 3145 13863 3179
rect 13863 3145 13872 3179
rect 13820 3136 13872 3145
rect 14372 3179 14424 3188
rect 14372 3145 14381 3179
rect 14381 3145 14415 3179
rect 14415 3145 14424 3179
rect 14372 3136 14424 3145
rect 15936 3179 15988 3188
rect 15936 3145 15945 3179
rect 15945 3145 15979 3179
rect 15979 3145 15988 3179
rect 15936 3136 15988 3145
rect 16488 3179 16540 3188
rect 16488 3145 16497 3179
rect 16497 3145 16531 3179
rect 16531 3145 16540 3179
rect 16488 3136 16540 3145
rect 16764 3136 16816 3188
rect 19984 3179 20036 3188
rect 2136 3000 2188 3052
rect 2872 3000 2924 3052
rect 3240 3068 3292 3120
rect 3332 3043 3384 3052
rect 3332 3009 3341 3043
rect 3341 3009 3375 3043
rect 3375 3009 3384 3043
rect 3332 3000 3384 3009
rect 14740 3000 14792 3052
rect 15384 3043 15436 3052
rect 3700 2932 3752 2984
rect 3976 2932 4028 2984
rect 5080 2932 5132 2984
rect 6736 2932 6788 2984
rect 7380 2975 7432 2984
rect 2872 2864 2924 2916
rect 5448 2864 5500 2916
rect 6276 2864 6328 2916
rect 7380 2941 7414 2975
rect 7414 2941 7432 2975
rect 7380 2932 7432 2941
rect 9496 2975 9548 2984
rect 9496 2941 9505 2975
rect 9505 2941 9539 2975
rect 9539 2941 9548 2975
rect 9496 2932 9548 2941
rect 12532 2932 12584 2984
rect 12716 2975 12768 2984
rect 12716 2941 12750 2975
rect 12750 2941 12768 2975
rect 14832 2975 14884 2984
rect 12716 2932 12768 2941
rect 14832 2941 14841 2975
rect 14841 2941 14875 2975
rect 14875 2941 14884 2975
rect 14832 2932 14884 2941
rect 15384 3009 15393 3043
rect 15393 3009 15427 3043
rect 15427 3009 15436 3043
rect 15384 3000 15436 3009
rect 17684 3000 17736 3052
rect 19984 3145 19993 3179
rect 19993 3145 20027 3179
rect 20027 3145 20036 3179
rect 19984 3136 20036 3145
rect 21640 3179 21692 3188
rect 21640 3145 21649 3179
rect 21649 3145 21683 3179
rect 21683 3145 21692 3179
rect 21640 3136 21692 3145
rect 22744 3179 22796 3188
rect 22744 3145 22753 3179
rect 22753 3145 22787 3179
rect 22787 3145 22796 3179
rect 22744 3136 22796 3145
rect 23480 3179 23532 3188
rect 23480 3145 23489 3179
rect 23489 3145 23523 3179
rect 23523 3145 23532 3179
rect 23480 3136 23532 3145
rect 25136 3136 25188 3188
rect 19984 3000 20036 3052
rect 20444 3000 20496 3052
rect 3240 2839 3292 2848
rect 3240 2805 3249 2839
rect 3249 2805 3283 2839
rect 3283 2805 3292 2839
rect 3240 2796 3292 2805
rect 4620 2796 4672 2848
rect 5264 2796 5316 2848
rect 8484 2839 8536 2848
rect 8484 2805 8493 2839
rect 8493 2805 8527 2839
rect 8527 2805 8536 2839
rect 8484 2796 8536 2805
rect 9588 2796 9640 2848
rect 16580 2932 16632 2984
rect 17960 2932 18012 2984
rect 20536 2975 20588 2984
rect 20536 2941 20545 2975
rect 20545 2941 20579 2975
rect 20579 2941 20588 2975
rect 20536 2932 20588 2941
rect 21824 2975 21876 2984
rect 21824 2941 21833 2975
rect 21833 2941 21867 2975
rect 21867 2941 21876 2975
rect 21824 2932 21876 2941
rect 23480 2932 23532 2984
rect 16948 2907 17000 2916
rect 16948 2873 16957 2907
rect 16957 2873 16991 2907
rect 16991 2873 17000 2907
rect 16948 2864 17000 2873
rect 24032 2932 24084 2984
rect 24768 2932 24820 2984
rect 25044 2864 25096 2916
rect 19432 2839 19484 2848
rect 19432 2805 19441 2839
rect 19441 2805 19475 2839
rect 19475 2805 19484 2839
rect 19432 2796 19484 2805
rect 22008 2839 22060 2848
rect 22008 2805 22017 2839
rect 22017 2805 22051 2839
rect 22051 2805 22060 2839
rect 22008 2796 22060 2805
rect 25136 2839 25188 2848
rect 25136 2805 25145 2839
rect 25145 2805 25179 2839
rect 25179 2805 25188 2839
rect 25136 2796 25188 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 2228 2635 2280 2644
rect 2228 2601 2237 2635
rect 2237 2601 2271 2635
rect 2271 2601 2280 2635
rect 2228 2592 2280 2601
rect 2688 2524 2740 2576
rect 5448 2635 5500 2644
rect 5448 2601 5457 2635
rect 5457 2601 5491 2635
rect 5491 2601 5500 2635
rect 5448 2592 5500 2601
rect 6000 2592 6052 2644
rect 6276 2635 6328 2644
rect 6276 2601 6285 2635
rect 6285 2601 6319 2635
rect 6319 2601 6328 2635
rect 6276 2592 6328 2601
rect 6736 2635 6788 2644
rect 6736 2601 6745 2635
rect 6745 2601 6779 2635
rect 6779 2601 6788 2635
rect 6736 2592 6788 2601
rect 8300 2592 8352 2644
rect 9588 2592 9640 2644
rect 11152 2635 11204 2644
rect 11152 2601 11161 2635
rect 11161 2601 11195 2635
rect 11195 2601 11204 2635
rect 11152 2592 11204 2601
rect 12532 2592 12584 2644
rect 14004 2635 14056 2644
rect 14004 2601 14013 2635
rect 14013 2601 14047 2635
rect 14047 2601 14056 2635
rect 14004 2592 14056 2601
rect 16580 2592 16632 2644
rect 17960 2592 18012 2644
rect 19984 2592 20036 2644
rect 20996 2592 21048 2644
rect 4068 2524 4120 2576
rect 4712 2524 4764 2576
rect 7104 2524 7156 2576
rect 10048 2567 10100 2576
rect 10048 2533 10082 2567
rect 10082 2533 10100 2567
rect 10048 2524 10100 2533
rect 13820 2524 13872 2576
rect 17040 2567 17092 2576
rect 17040 2533 17049 2567
rect 17049 2533 17083 2567
rect 17083 2533 17092 2567
rect 17040 2524 17092 2533
rect 18604 2567 18656 2576
rect 18604 2533 18613 2567
rect 18613 2533 18647 2567
rect 18647 2533 18656 2567
rect 18604 2524 18656 2533
rect 24768 2524 24820 2576
rect 9496 2499 9548 2508
rect 9496 2465 9505 2499
rect 9505 2465 9539 2499
rect 9539 2465 9548 2499
rect 9496 2456 9548 2465
rect 12532 2456 12584 2508
rect 15476 2499 15528 2508
rect 2044 2388 2096 2440
rect 2688 2388 2740 2440
rect 3976 2388 4028 2440
rect 11520 2388 11572 2440
rect 15476 2465 15485 2499
rect 15485 2465 15519 2499
rect 15519 2465 15528 2499
rect 15476 2456 15528 2465
rect 16764 2499 16816 2508
rect 16764 2465 16773 2499
rect 16773 2465 16807 2499
rect 16807 2465 16816 2499
rect 16764 2456 16816 2465
rect 18236 2456 18288 2508
rect 19616 2499 19668 2508
rect 19616 2465 19625 2499
rect 19625 2465 19659 2499
rect 19659 2465 19668 2499
rect 19616 2456 19668 2465
rect 21180 2499 21232 2508
rect 21180 2465 21189 2499
rect 21189 2465 21223 2499
rect 21223 2465 21232 2499
rect 21180 2456 21232 2465
rect 22284 2499 22336 2508
rect 22284 2465 22293 2499
rect 22293 2465 22327 2499
rect 22327 2465 22336 2499
rect 22284 2456 22336 2465
rect 24032 2499 24084 2508
rect 24032 2465 24041 2499
rect 24041 2465 24075 2499
rect 24075 2465 24084 2499
rect 24032 2456 24084 2465
rect 25044 2456 25096 2508
rect 15752 2431 15804 2440
rect 15752 2397 15761 2431
rect 15761 2397 15795 2431
rect 15795 2397 15804 2431
rect 15752 2388 15804 2397
rect 20536 2431 20588 2440
rect 20536 2397 20545 2431
rect 20545 2397 20579 2431
rect 20579 2397 20588 2431
rect 20536 2388 20588 2397
rect 1584 2320 1636 2372
rect 26516 2320 26568 2372
rect 14648 2252 14700 2304
rect 19432 2295 19484 2304
rect 19432 2261 19441 2295
rect 19441 2261 19475 2295
rect 19475 2261 19484 2295
rect 19432 2252 19484 2261
rect 22468 2295 22520 2304
rect 22468 2261 22477 2295
rect 22477 2261 22511 2295
rect 22511 2261 22520 2295
rect 22468 2252 22520 2261
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 9680 2048 9732 2100
rect 15384 2048 15436 2100
rect 16672 2048 16724 2100
rect 20720 2048 20772 2100
rect 14832 1096 14884 1148
rect 15660 1096 15712 1148
rect 9036 620 9088 672
rect 6920 552 6972 604
rect 7564 552 7616 604
rect 7840 552 7892 604
rect 12256 552 12308 604
rect 15936 552 15988 604
<< metal2 >>
rect 3146 27568 3202 27577
rect 3146 27503 3202 27512
rect 2962 26888 3018 26897
rect 2962 26823 3018 26832
rect 2976 26314 3004 26823
rect 2964 26308 3016 26314
rect 2964 26250 3016 26256
rect 570 24848 626 24857
rect 570 24783 626 24792
rect 584 23769 612 24783
rect 570 23760 626 23769
rect 570 23695 626 23704
rect 1490 16688 1546 16697
rect 1490 16623 1546 16632
rect 1400 14272 1452 14278
rect 1400 14214 1452 14220
rect 1412 12306 1440 14214
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 1504 11558 1532 16623
rect 1766 15328 1822 15337
rect 1766 15263 1822 15272
rect 1584 13728 1636 13734
rect 1584 13670 1636 13676
rect 1492 11552 1544 11558
rect 1492 11494 1544 11500
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1504 10606 1532 11086
rect 1492 10600 1544 10606
rect 1492 10542 1544 10548
rect 572 10124 624 10130
rect 572 10066 624 10072
rect 584 9897 612 10066
rect 570 9888 626 9897
rect 570 9823 626 9832
rect 1492 9376 1544 9382
rect 1492 9318 1544 9324
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 8090 1440 8434
rect 1400 8084 1452 8090
rect 1400 8026 1452 8032
rect 846 7304 902 7313
rect 846 7239 902 7248
rect 294 4176 350 4185
rect 294 4111 350 4120
rect 308 480 336 4111
rect 860 480 888 7239
rect 1400 7200 1452 7206
rect 1400 7142 1452 7148
rect 1412 6905 1440 7142
rect 1398 6896 1454 6905
rect 1398 6831 1454 6840
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 5846 1440 6734
rect 1400 5840 1452 5846
rect 1400 5782 1452 5788
rect 1308 5772 1360 5778
rect 1308 5714 1360 5720
rect 1320 3097 1348 5714
rect 1398 4992 1454 5001
rect 1398 4927 1454 4936
rect 1412 4826 1440 4927
rect 1400 4820 1452 4826
rect 1400 4762 1452 4768
rect 1400 3936 1452 3942
rect 1400 3878 1452 3884
rect 1306 3088 1362 3097
rect 1306 3023 1362 3032
rect 1412 480 1440 3878
rect 1504 1057 1532 9318
rect 1596 7177 1624 13670
rect 1780 10810 1808 15263
rect 2412 14408 2464 14414
rect 2042 14376 2098 14385
rect 2412 14350 2464 14356
rect 2042 14311 2098 14320
rect 1952 14272 2004 14278
rect 1952 14214 2004 14220
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1676 10464 1728 10470
rect 1676 10406 1728 10412
rect 1688 9518 1716 10406
rect 1768 10192 1820 10198
rect 1768 10134 1820 10140
rect 1780 9761 1808 10134
rect 1766 9752 1822 9761
rect 1766 9687 1822 9696
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1780 9382 1808 9687
rect 1768 9376 1820 9382
rect 1768 9318 1820 9324
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1780 8430 1808 8774
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1780 8090 1808 8366
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 1674 7576 1730 7585
rect 1674 7511 1730 7520
rect 1582 7168 1638 7177
rect 1582 7103 1638 7112
rect 1584 6248 1636 6254
rect 1584 6190 1636 6196
rect 1596 2378 1624 6190
rect 1688 4078 1716 7511
rect 1780 7410 1808 8026
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1872 5817 1900 13126
rect 1964 12442 1992 14214
rect 2056 14074 2084 14311
rect 2044 14068 2096 14074
rect 2044 14010 2096 14016
rect 2056 13870 2084 14010
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 2228 13864 2280 13870
rect 2228 13806 2280 13812
rect 2136 13796 2188 13802
rect 2136 13738 2188 13744
rect 2148 12850 2176 13738
rect 2136 12844 2188 12850
rect 2136 12786 2188 12792
rect 2044 12708 2096 12714
rect 2044 12650 2096 12656
rect 1952 12436 2004 12442
rect 1952 12378 2004 12384
rect 1964 9994 1992 12378
rect 2056 12170 2084 12650
rect 2044 12164 2096 12170
rect 2044 12106 2096 12112
rect 2148 11898 2176 12786
rect 2136 11892 2188 11898
rect 2136 11834 2188 11840
rect 2044 11620 2096 11626
rect 2044 11562 2096 11568
rect 2056 11286 2084 11562
rect 2044 11280 2096 11286
rect 2044 11222 2096 11228
rect 2044 10804 2096 10810
rect 2044 10746 2096 10752
rect 1952 9988 2004 9994
rect 1952 9930 2004 9936
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 1964 9178 1992 9318
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1858 5808 1914 5817
rect 1858 5743 1914 5752
rect 1964 5710 1992 6598
rect 2056 5914 2084 10746
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2148 9382 2176 9998
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 2148 7732 2176 9114
rect 2240 8362 2268 13806
rect 2320 13184 2372 13190
rect 2320 13126 2372 13132
rect 2332 12850 2360 13126
rect 2320 12844 2372 12850
rect 2320 12786 2372 12792
rect 2424 12442 2452 14350
rect 2872 13932 2924 13938
rect 2872 13874 2924 13880
rect 2596 13388 2648 13394
rect 2596 13330 2648 13336
rect 2504 13252 2556 13258
rect 2504 13194 2556 13200
rect 2516 12866 2544 13194
rect 2608 12986 2636 13330
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2516 12838 2636 12866
rect 2412 12436 2464 12442
rect 2412 12378 2464 12384
rect 2320 12300 2372 12306
rect 2320 12242 2372 12248
rect 2332 12209 2360 12242
rect 2318 12200 2374 12209
rect 2318 12135 2374 12144
rect 2424 11762 2452 12378
rect 2608 12345 2636 12838
rect 2594 12336 2650 12345
rect 2594 12271 2650 12280
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2320 10532 2372 10538
rect 2320 10474 2372 10480
rect 2332 10062 2360 10474
rect 2320 10056 2372 10062
rect 2320 9998 2372 10004
rect 2596 9648 2648 9654
rect 2594 9616 2596 9625
rect 2648 9616 2650 9625
rect 2594 9551 2650 9560
rect 2412 9512 2464 9518
rect 2700 9466 2728 13126
rect 2780 12844 2832 12850
rect 2780 12786 2832 12792
rect 2792 12442 2820 12786
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2792 10606 2820 11494
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2792 10266 2820 10542
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2884 9518 2912 13874
rect 2964 13252 3016 13258
rect 2964 13194 3016 13200
rect 2412 9454 2464 9460
rect 2228 8356 2280 8362
rect 2228 8298 2280 8304
rect 2240 7886 2268 8298
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2148 7704 2268 7732
rect 2134 7032 2190 7041
rect 2134 6967 2190 6976
rect 2044 5908 2096 5914
rect 2044 5850 2096 5856
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 1964 5250 1992 5646
rect 2056 5370 2084 5850
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 1964 5222 2084 5250
rect 2056 5098 2084 5222
rect 2044 5092 2096 5098
rect 2044 5034 2096 5040
rect 1950 4720 2006 4729
rect 1950 4655 2006 4664
rect 1676 4072 1728 4078
rect 1676 4014 1728 4020
rect 1688 3738 1716 4014
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 1584 2372 1636 2378
rect 1584 2314 1636 2320
rect 1490 1048 1546 1057
rect 1490 983 1546 992
rect 1964 480 1992 4655
rect 2056 2446 2084 5034
rect 2148 3058 2176 6967
rect 2240 4185 2268 7704
rect 2332 7546 2360 7890
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 2332 7002 2360 7346
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2332 6458 2360 6938
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 2332 5914 2360 6394
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2332 5098 2360 5850
rect 2320 5092 2372 5098
rect 2320 5034 2372 5040
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 2226 4176 2282 4185
rect 2226 4111 2282 4120
rect 2332 4010 2360 4422
rect 2320 4004 2372 4010
rect 2320 3946 2372 3952
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 2240 2650 2268 3470
rect 2332 3369 2360 3946
rect 2424 3890 2452 9454
rect 2608 9438 2728 9466
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2504 8356 2556 8362
rect 2504 8298 2556 8304
rect 2516 7342 2544 8298
rect 2608 7857 2636 9438
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2594 7848 2650 7857
rect 2594 7783 2650 7792
rect 2596 7744 2648 7750
rect 2596 7686 2648 7692
rect 2504 7336 2556 7342
rect 2504 7278 2556 7284
rect 2608 7154 2636 7686
rect 2516 7126 2636 7154
rect 2516 6254 2544 7126
rect 2700 6934 2728 9318
rect 2884 8634 2912 9454
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2870 8256 2926 8265
rect 2870 8191 2926 8200
rect 2688 6928 2740 6934
rect 2884 6882 2912 8191
rect 2976 7750 3004 13194
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 3068 12186 3096 12582
rect 3160 12374 3188 27503
rect 15752 26308 15804 26314
rect 15752 26250 15804 26256
rect 3514 26208 3570 26217
rect 3514 26143 3570 26152
rect 3422 25528 3478 25537
rect 3422 25463 3478 25472
rect 3436 24954 3464 25463
rect 3424 24948 3476 24954
rect 3424 24890 3476 24896
rect 3528 24886 3556 26143
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 13268 24948 13320 24954
rect 13268 24890 13320 24896
rect 3516 24880 3568 24886
rect 3516 24822 3568 24828
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 3422 24168 3478 24177
rect 3422 24103 3478 24112
rect 3238 23488 3294 23497
rect 3238 23423 3294 23432
rect 3252 17218 3280 23423
rect 3436 22273 3464 24103
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 10966 23760 11022 23769
rect 10966 23695 11022 23704
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5998 22672 6054 22681
rect 5998 22607 6054 22616
rect 3422 22264 3478 22273
rect 3422 22199 3478 22208
rect 3422 22128 3478 22137
rect 3422 22063 3478 22072
rect 3436 17649 3464 22063
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 4066 20768 4122 20777
rect 4066 20703 4122 20712
rect 3790 19408 3846 19417
rect 3790 19343 3846 19352
rect 3422 17640 3478 17649
rect 3422 17575 3478 17584
rect 3698 17368 3754 17377
rect 3698 17303 3754 17312
rect 3252 17190 3556 17218
rect 3238 16008 3294 16017
rect 3238 15943 3294 15952
rect 3148 12368 3200 12374
rect 3148 12310 3200 12316
rect 3068 12158 3188 12186
rect 3160 12102 3188 12158
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 3160 11626 3188 12038
rect 3148 11620 3200 11626
rect 3148 11562 3200 11568
rect 3160 10470 3188 11562
rect 3148 10464 3200 10470
rect 3148 10406 3200 10412
rect 3160 10266 3188 10406
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 3148 9444 3200 9450
rect 3148 9386 3200 9392
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 3068 7562 3096 9318
rect 3160 9042 3188 9386
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 3252 7886 3280 15943
rect 3330 14648 3386 14657
rect 3330 14583 3386 14592
rect 3344 12594 3372 14583
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 3436 12714 3464 13126
rect 3424 12708 3476 12714
rect 3424 12650 3476 12656
rect 3344 12566 3464 12594
rect 3332 12436 3384 12442
rect 3332 12378 3384 12384
rect 3344 11694 3372 12378
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 3344 11354 3372 11630
rect 3332 11348 3384 11354
rect 3332 11290 3384 11296
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 2688 6870 2740 6876
rect 2792 6854 2912 6882
rect 2976 7534 3096 7562
rect 2504 6248 2556 6254
rect 2504 6190 2556 6196
rect 2686 6216 2742 6225
rect 2686 6151 2742 6160
rect 2700 5642 2728 6151
rect 2688 5636 2740 5642
rect 2688 5578 2740 5584
rect 2792 4554 2820 6854
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 2884 4622 2912 6734
rect 2976 6662 3004 7534
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 3068 6798 3096 7278
rect 3252 7206 3280 7822
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2964 6180 3016 6186
rect 3148 6180 3200 6186
rect 3016 6140 3096 6168
rect 2964 6122 3016 6128
rect 2964 5840 3016 5846
rect 2962 5808 2964 5817
rect 3016 5808 3018 5817
rect 2962 5743 3018 5752
rect 3068 5681 3096 6140
rect 3148 6122 3200 6128
rect 3160 6089 3188 6122
rect 3146 6080 3202 6089
rect 3146 6015 3202 6024
rect 3054 5672 3110 5681
rect 3054 5607 3110 5616
rect 3160 5370 3188 6015
rect 3148 5364 3200 5370
rect 3148 5306 3200 5312
rect 3056 4752 3108 4758
rect 3056 4694 3108 4700
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 2780 4548 2832 4554
rect 2780 4490 2832 4496
rect 2596 4480 2648 4486
rect 2596 4422 2648 4428
rect 2424 3862 2544 3890
rect 2412 3732 2464 3738
rect 2412 3674 2464 3680
rect 2318 3360 2374 3369
rect 2424 3346 2452 3674
rect 2516 3618 2544 3862
rect 2608 3738 2636 4422
rect 2884 4214 2912 4558
rect 2872 4208 2924 4214
rect 2872 4150 2924 4156
rect 2976 4146 3004 4558
rect 3068 4214 3096 4694
rect 3146 4584 3202 4593
rect 3146 4519 3202 4528
rect 3056 4208 3108 4214
rect 3054 4176 3056 4185
rect 3108 4176 3110 4185
rect 2964 4140 3016 4146
rect 3054 4111 3110 4120
rect 2964 4082 3016 4088
rect 2780 4004 2832 4010
rect 2780 3946 2832 3952
rect 2792 3890 2820 3946
rect 2700 3862 2820 3890
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 2516 3590 2636 3618
rect 2502 3496 2558 3505
rect 2502 3431 2504 3440
rect 2556 3431 2558 3440
rect 2504 3402 2556 3408
rect 2424 3318 2544 3346
rect 2318 3295 2374 3304
rect 2228 2644 2280 2650
rect 2228 2586 2280 2592
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 2516 480 2544 3318
rect 2608 3233 2636 3590
rect 2594 3224 2650 3233
rect 2594 3159 2650 3168
rect 2700 2582 2728 3862
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 2688 2576 2740 2582
rect 2688 2518 2740 2524
rect 2688 2440 2740 2446
rect 2792 2394 2820 3538
rect 2884 3516 2912 3878
rect 2976 3754 3004 4082
rect 2976 3738 3096 3754
rect 2976 3732 3108 3738
rect 2976 3726 3056 3732
rect 3056 3674 3108 3680
rect 2964 3664 3016 3670
rect 2962 3632 2964 3641
rect 3016 3632 3018 3641
rect 2962 3567 3018 3576
rect 2964 3528 3016 3534
rect 2884 3488 2964 3516
rect 2964 3470 3016 3476
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2884 2922 2912 2994
rect 2872 2916 2924 2922
rect 2872 2858 2924 2864
rect 2740 2388 2820 2394
rect 2688 2382 2820 2388
rect 2700 2366 2820 2382
rect 2976 1465 3004 3470
rect 3056 3460 3108 3466
rect 3056 3402 3108 3408
rect 2962 1456 3018 1465
rect 2962 1391 3018 1400
rect 3068 480 3096 3402
rect 294 0 350 480
rect 846 0 902 480
rect 1398 0 1454 480
rect 1950 0 2006 480
rect 2502 0 2558 480
rect 3054 0 3110 480
rect 3160 377 3188 4519
rect 3344 4434 3372 9046
rect 3436 5409 3464 12566
rect 3528 11393 3556 17190
rect 3712 12986 3740 17303
rect 3700 12980 3752 12986
rect 3700 12922 3752 12928
rect 3712 12714 3740 12922
rect 3700 12708 3752 12714
rect 3700 12650 3752 12656
rect 3608 12368 3660 12374
rect 3608 12310 3660 12316
rect 3514 11384 3570 11393
rect 3514 11319 3570 11328
rect 3516 11008 3568 11014
rect 3516 10950 3568 10956
rect 3528 9926 3556 10950
rect 3516 9920 3568 9926
rect 3516 9862 3568 9868
rect 3528 9178 3556 9862
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 3620 9110 3648 12310
rect 3700 11348 3752 11354
rect 3700 11290 3752 11296
rect 3608 9104 3660 9110
rect 3608 9046 3660 9052
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3516 8356 3568 8362
rect 3516 8298 3568 8304
rect 3528 7954 3556 8298
rect 3620 8090 3648 8774
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3516 7948 3568 7954
rect 3516 7890 3568 7896
rect 3528 7818 3556 7890
rect 3516 7812 3568 7818
rect 3516 7754 3568 7760
rect 3620 7546 3648 8026
rect 3608 7540 3660 7546
rect 3608 7482 3660 7488
rect 3606 5944 3662 5953
rect 3606 5879 3662 5888
rect 3422 5400 3478 5409
rect 3422 5335 3478 5344
rect 3620 5137 3648 5879
rect 3606 5128 3662 5137
rect 3606 5063 3662 5072
rect 3712 4457 3740 11290
rect 3804 10169 3832 19343
rect 3974 18728 4030 18737
rect 3974 18663 4030 18672
rect 3882 18048 3938 18057
rect 3882 17983 3938 17992
rect 3896 12374 3924 17983
rect 3988 13569 4016 18663
rect 4080 16017 4108 20703
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 4066 16008 4122 16017
rect 4066 15943 4122 15952
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 3974 13560 4030 13569
rect 3974 13495 4030 13504
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 4160 13320 4212 13326
rect 5000 13297 5028 13330
rect 4160 13262 4212 13268
rect 4986 13288 5042 13297
rect 3974 12880 4030 12889
rect 3974 12815 4030 12824
rect 3988 12617 4016 12815
rect 3974 12608 4030 12617
rect 3974 12543 4030 12552
rect 3884 12368 3936 12374
rect 3884 12310 3936 12316
rect 4172 12288 4200 13262
rect 4986 13223 5042 13232
rect 4804 13184 4856 13190
rect 4804 13126 4856 13132
rect 4712 12912 4764 12918
rect 4712 12854 4764 12860
rect 4620 12708 4672 12714
rect 4620 12650 4672 12656
rect 3988 12260 4200 12288
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 3896 10470 3924 11154
rect 3884 10464 3936 10470
rect 3884 10406 3936 10412
rect 3790 10160 3846 10169
rect 3790 10095 3846 10104
rect 3988 9586 4016 12260
rect 4632 12238 4660 12650
rect 4724 12481 4752 12854
rect 4710 12472 4766 12481
rect 4710 12407 4766 12416
rect 4620 12232 4672 12238
rect 4158 12200 4214 12209
rect 4620 12174 4672 12180
rect 4158 12135 4214 12144
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 3804 8090 3832 9318
rect 3974 9208 4030 9217
rect 3974 9143 4030 9152
rect 3988 8537 4016 9143
rect 3974 8528 4030 8537
rect 3974 8463 4030 8472
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 3792 7948 3844 7954
rect 3792 7890 3844 7896
rect 3804 7750 3832 7890
rect 4080 7750 4108 12038
rect 4172 8906 4200 12135
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 4264 9450 4292 12038
rect 4632 11558 4660 12174
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4632 11082 4660 11494
rect 4620 11076 4672 11082
rect 4620 11018 4672 11024
rect 4632 10538 4660 11018
rect 4620 10532 4672 10538
rect 4620 10474 4672 10480
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 4356 10305 4384 10406
rect 4342 10296 4398 10305
rect 4342 10231 4398 10240
rect 4620 10192 4672 10198
rect 4620 10134 4672 10140
rect 4632 9722 4660 10134
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 4436 9648 4488 9654
rect 4436 9590 4488 9596
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 4252 9444 4304 9450
rect 4252 9386 4304 9392
rect 4160 8900 4212 8906
rect 4160 8842 4212 8848
rect 4356 8106 4384 9522
rect 4448 9489 4476 9590
rect 4434 9480 4490 9489
rect 4434 9415 4490 9424
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 4540 8566 4568 8910
rect 4528 8560 4580 8566
rect 4528 8502 4580 8508
rect 4436 8288 4488 8294
rect 4540 8265 4568 8502
rect 4436 8230 4488 8236
rect 4526 8256 4582 8265
rect 4172 8078 4384 8106
rect 3792 7744 3844 7750
rect 3792 7686 3844 7692
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 3804 6798 3832 7686
rect 4080 6934 4108 7686
rect 4068 6928 4120 6934
rect 4068 6870 4120 6876
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3804 4826 3832 6734
rect 4172 6730 4200 8078
rect 4344 8016 4396 8022
rect 4344 7958 4396 7964
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 3974 6488 4030 6497
rect 4264 6458 4292 6938
rect 3974 6423 4030 6432
rect 4252 6452 4304 6458
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3252 4406 3372 4434
rect 3698 4448 3754 4457
rect 3252 3670 3280 4406
rect 3698 4383 3754 4392
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3240 3664 3292 3670
rect 3240 3606 3292 3612
rect 3252 3126 3280 3606
rect 3606 3360 3662 3369
rect 3606 3295 3662 3304
rect 3240 3120 3292 3126
rect 3240 3062 3292 3068
rect 3330 3088 3386 3097
rect 3330 3023 3332 3032
rect 3384 3023 3386 3032
rect 3332 2994 3384 3000
rect 3240 2848 3292 2854
rect 3238 2816 3240 2825
rect 3292 2816 3294 2825
rect 3238 2751 3294 2760
rect 3620 480 3648 3295
rect 3712 2990 3740 3878
rect 3896 3466 3924 5510
rect 3988 5137 4016 6423
rect 4252 6394 4304 6400
rect 4264 5914 4292 6394
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4068 5636 4120 5642
rect 4068 5578 4120 5584
rect 3974 5128 4030 5137
rect 3974 5063 4030 5072
rect 4080 4826 4108 5578
rect 4172 5370 4200 5714
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4160 5092 4212 5098
rect 4264 5080 4292 5646
rect 4356 5302 4384 7958
rect 4448 7954 4476 8230
rect 4526 8191 4582 8200
rect 4632 8022 4660 9658
rect 4724 9518 4752 12407
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4620 8016 4672 8022
rect 4620 7958 4672 7964
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4528 7880 4580 7886
rect 4526 7848 4528 7857
rect 4580 7848 4582 7857
rect 4526 7783 4582 7792
rect 4540 7546 4568 7783
rect 4632 7546 4660 7958
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 4540 7313 4568 7482
rect 4526 7304 4582 7313
rect 4526 7239 4582 7248
rect 4724 6934 4752 7822
rect 4712 6928 4764 6934
rect 4712 6870 4764 6876
rect 4436 6860 4488 6866
rect 4436 6802 4488 6808
rect 4448 5574 4476 6802
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 4724 6118 4752 6734
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4618 5400 4674 5409
rect 4618 5335 4620 5344
rect 4672 5335 4674 5344
rect 4620 5306 4672 5312
rect 4344 5296 4396 5302
rect 4344 5238 4396 5244
rect 4212 5052 4292 5080
rect 4160 5034 4212 5040
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4172 4690 4200 5034
rect 4160 4684 4212 4690
rect 4160 4626 4212 4632
rect 4068 4004 4120 4010
rect 4068 3946 4120 3952
rect 3884 3460 3936 3466
rect 3884 3402 3936 3408
rect 4080 3194 4108 3946
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 3712 1329 3740 2926
rect 3988 2446 4016 2926
rect 4068 2576 4120 2582
rect 4172 2564 4200 3334
rect 4120 2536 4200 2564
rect 4068 2518 4120 2524
rect 3976 2440 4028 2446
rect 4172 2417 4200 2536
rect 3976 2382 4028 2388
rect 4158 2408 4214 2417
rect 4158 2343 4214 2352
rect 4356 2258 4384 5238
rect 4724 4729 4752 6054
rect 4710 4720 4766 4729
rect 4710 4655 4766 4664
rect 4816 4010 4844 13126
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5448 12844 5500 12850
rect 5500 12804 5580 12832
rect 5448 12786 5500 12792
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4908 9994 4936 12582
rect 5264 12368 5316 12374
rect 5264 12310 5316 12316
rect 5356 12368 5408 12374
rect 5356 12310 5408 12316
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 5000 11121 5028 12038
rect 5276 11898 5304 12310
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5368 11558 5396 12310
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5356 11552 5408 11558
rect 5356 11494 5408 11500
rect 5264 11144 5316 11150
rect 4986 11112 5042 11121
rect 5264 11086 5316 11092
rect 4986 11047 5042 11056
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 5092 10062 5120 10474
rect 5276 10470 5304 11086
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 4896 9988 4948 9994
rect 4896 9930 4948 9936
rect 4908 9450 4936 9930
rect 4896 9444 4948 9450
rect 4896 9386 4948 9392
rect 5092 9178 5120 9998
rect 5184 9382 5212 10066
rect 5368 9738 5396 11494
rect 5460 11354 5488 12174
rect 5552 11762 5580 12804
rect 5906 12472 5962 12481
rect 5906 12407 5962 12416
rect 5920 12374 5948 12407
rect 5908 12368 5960 12374
rect 5908 12310 5960 12316
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5540 11280 5592 11286
rect 5540 11222 5592 11228
rect 5552 10810 5580 11222
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5552 10266 5580 10746
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5446 9752 5502 9761
rect 5368 9710 5446 9738
rect 5552 9722 5580 10202
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5446 9687 5502 9696
rect 5540 9716 5592 9722
rect 5460 9602 5488 9687
rect 5540 9658 5592 9664
rect 5460 9586 5580 9602
rect 5460 9580 5592 9586
rect 5460 9574 5540 9580
rect 5540 9522 5592 9528
rect 5172 9376 5224 9382
rect 5170 9344 5172 9353
rect 5224 9344 5226 9353
rect 5170 9279 5226 9288
rect 5184 9253 5212 9279
rect 5538 9208 5594 9217
rect 5080 9172 5132 9178
rect 5538 9143 5540 9152
rect 5080 9114 5132 9120
rect 5592 9143 5594 9152
rect 5540 9114 5592 9120
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 5368 8362 5396 9046
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5368 7585 5396 8298
rect 5354 7576 5410 7585
rect 5354 7511 5410 7520
rect 5264 7472 5316 7478
rect 5262 7440 5264 7449
rect 5316 7440 5318 7449
rect 5262 7375 5318 7384
rect 5368 7177 5396 7511
rect 5354 7168 5410 7177
rect 5354 7103 5410 7112
rect 5170 6896 5226 6905
rect 5170 6831 5226 6840
rect 5184 6798 5212 6831
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 5184 6458 5212 6734
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5354 6352 5410 6361
rect 5354 6287 5410 6296
rect 5368 6254 5396 6287
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5264 5296 5316 5302
rect 5262 5264 5264 5273
rect 5316 5264 5318 5273
rect 5262 5199 5318 5208
rect 5368 4758 5396 5510
rect 5460 4865 5488 5714
rect 5446 4856 5502 4865
rect 5446 4791 5502 4800
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 5552 4078 5580 8366
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5736 6769 5764 7346
rect 5816 7268 5868 7274
rect 5816 7210 5868 7216
rect 5828 6934 5856 7210
rect 5816 6928 5868 6934
rect 5816 6870 5868 6876
rect 6012 6866 6040 22607
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 8758 22264 8814 22273
rect 10289 22256 10585 22276
rect 8758 22199 8814 22208
rect 7838 13560 7894 13569
rect 7838 13495 7840 13504
rect 7892 13495 7894 13504
rect 7840 13466 7892 13472
rect 6090 13016 6146 13025
rect 6090 12951 6092 12960
rect 6144 12951 6146 12960
rect 6092 12922 6144 12928
rect 7852 12714 7880 13466
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 7840 12708 7892 12714
rect 7840 12650 7892 12656
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6472 11558 6500 12174
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6274 11384 6330 11393
rect 6274 11319 6330 11328
rect 6288 10198 6316 11319
rect 6656 10810 6684 12582
rect 7472 12096 7524 12102
rect 7472 12038 7524 12044
rect 7484 11626 7512 12038
rect 8114 11656 8170 11665
rect 7472 11620 7524 11626
rect 8114 11591 8170 11600
rect 7472 11562 7524 11568
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6366 10568 6422 10577
rect 6366 10503 6422 10512
rect 6380 10266 6408 10503
rect 6748 10470 6776 11494
rect 7024 11354 7052 11494
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 7378 11112 7434 11121
rect 7378 11047 7434 11056
rect 7392 10470 7420 11047
rect 7484 11014 7512 11562
rect 8128 11082 8156 11591
rect 8312 11354 8340 12854
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8116 11076 8168 11082
rect 8116 11018 8168 11024
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7484 10538 7512 10950
rect 8220 10810 8248 11154
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8588 10810 8616 11086
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 7380 10464 7432 10470
rect 7380 10406 7432 10412
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6276 10192 6328 10198
rect 6276 10134 6328 10140
rect 6460 10192 6512 10198
rect 6460 10134 6512 10140
rect 6288 9722 6316 10134
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6472 9586 6500 10134
rect 6748 9654 6776 10406
rect 7378 10296 7434 10305
rect 7484 10266 7512 10474
rect 8484 10464 8536 10470
rect 8114 10432 8170 10441
rect 8484 10406 8536 10412
rect 8114 10367 8170 10376
rect 8022 10296 8078 10305
rect 7378 10231 7434 10240
rect 7472 10260 7524 10266
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6736 9648 6788 9654
rect 6736 9590 6788 9596
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 6182 9208 6238 9217
rect 6182 9143 6238 9152
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6104 8362 6132 8978
rect 6092 8356 6144 8362
rect 6092 8298 6144 8304
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 5722 6760 5778 6769
rect 5722 6695 5724 6704
rect 5776 6695 5778 6704
rect 5724 6666 5776 6672
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6012 6458 6040 6802
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6012 4593 6040 6054
rect 5998 4584 6054 4593
rect 5998 4519 6054 4528
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 4804 4004 4856 4010
rect 4804 3946 4856 3952
rect 5816 4004 5868 4010
rect 5816 3946 5868 3952
rect 5080 3936 5132 3942
rect 5264 3936 5316 3942
rect 5080 3878 5132 3884
rect 5262 3904 5264 3913
rect 5724 3936 5776 3942
rect 5316 3904 5318 3913
rect 4620 3664 4672 3670
rect 4620 3606 4672 3612
rect 4632 2854 4660 3606
rect 5092 3534 5120 3878
rect 5724 3878 5776 3884
rect 5262 3839 5318 3848
rect 5736 3777 5764 3878
rect 5722 3768 5778 3777
rect 5722 3703 5778 3712
rect 5828 3670 5856 3946
rect 5816 3664 5868 3670
rect 5816 3606 5868 3612
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 4724 2961 4752 3470
rect 5092 3398 5120 3470
rect 5080 3392 5132 3398
rect 5644 3380 5672 3538
rect 5080 3334 5132 3340
rect 5552 3352 5672 3380
rect 4802 3224 4858 3233
rect 4802 3159 4858 3168
rect 4710 2952 4766 2961
rect 4710 2887 4766 2896
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4724 2582 4752 2887
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 4816 2394 4844 3159
rect 5092 2990 5120 3334
rect 5552 3194 5580 3352
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5552 3097 5580 3130
rect 5538 3088 5594 3097
rect 5538 3023 5594 3032
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 5448 2916 5500 2922
rect 5448 2858 5500 2864
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 4172 2230 4384 2258
rect 4724 2366 4844 2394
rect 3698 1320 3754 1329
rect 3698 1255 3754 1264
rect 4172 480 4200 2230
rect 4724 480 4752 2366
rect 5276 480 5304 2790
rect 5460 2650 5488 2858
rect 6012 2650 6040 4422
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 6000 2644 6052 2650
rect 6000 2586 6052 2592
rect 5622 2204 5918 2224
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6104 1986 6132 8298
rect 6196 7342 6224 9143
rect 6748 9058 6776 9590
rect 6840 9194 6868 10066
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 6840 9166 6960 9194
rect 6932 9110 6960 9166
rect 6920 9104 6972 9110
rect 6748 9030 6868 9058
rect 6920 9046 6972 9052
rect 6840 8838 6868 9030
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6182 4312 6238 4321
rect 6182 4247 6184 4256
rect 6236 4247 6238 4256
rect 6184 4218 6236 4224
rect 6380 4060 6408 8774
rect 6656 8362 6684 8774
rect 6840 8430 6868 8774
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6564 8022 6592 8230
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 6564 7206 6592 7958
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6656 7721 6684 7890
rect 7012 7812 7064 7818
rect 7012 7754 7064 7760
rect 6920 7744 6972 7750
rect 6642 7712 6698 7721
rect 6920 7686 6972 7692
rect 6642 7647 6698 7656
rect 6656 7546 6684 7647
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6564 6118 6592 7142
rect 6656 7002 6684 7482
rect 6644 6996 6696 7002
rect 6644 6938 6696 6944
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6564 5234 6592 6054
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6748 5574 6776 5714
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6564 5030 6592 5170
rect 6748 5098 6776 5510
rect 6736 5092 6788 5098
rect 6736 5034 6788 5040
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6748 4826 6776 5034
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6380 4032 6500 4060
rect 6276 3664 6328 3670
rect 6276 3606 6328 3612
rect 6288 2922 6316 3606
rect 6276 2916 6328 2922
rect 6276 2858 6328 2864
rect 6288 2650 6316 2858
rect 6366 2816 6422 2825
rect 6366 2751 6422 2760
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 5828 1958 6132 1986
rect 5828 480 5856 1958
rect 6380 480 6408 2751
rect 6472 2553 6500 4032
rect 6840 3602 6868 5850
rect 6932 5642 6960 7686
rect 7024 5846 7052 7754
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7116 5914 7144 6598
rect 7208 5953 7236 9318
rect 7288 8356 7340 8362
rect 7288 8298 7340 8304
rect 7300 7750 7328 8298
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7300 7274 7328 7686
rect 7288 7268 7340 7274
rect 7288 7210 7340 7216
rect 7392 6934 7420 10231
rect 8128 10266 8156 10367
rect 8022 10231 8078 10240
rect 8116 10260 8168 10266
rect 7472 10202 7524 10208
rect 8036 10062 8064 10231
rect 8116 10202 8168 10208
rect 8024 10056 8076 10062
rect 7562 10024 7618 10033
rect 8024 9998 8076 10004
rect 7562 9959 7564 9968
rect 7616 9959 7618 9968
rect 7564 9930 7616 9936
rect 8036 9722 8064 9998
rect 8128 9926 8156 10202
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 8312 9500 8340 10066
rect 8496 9722 8524 10406
rect 8588 10266 8616 10746
rect 8668 10736 8720 10742
rect 8668 10678 8720 10684
rect 8680 10470 8708 10678
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8484 9716 8536 9722
rect 8484 9658 8536 9664
rect 8392 9512 8444 9518
rect 8312 9472 8392 9500
rect 7930 8120 7986 8129
rect 7930 8055 7986 8064
rect 7562 7848 7618 7857
rect 7562 7783 7618 7792
rect 7576 7410 7604 7783
rect 7944 7546 7972 8055
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 7748 7472 7800 7478
rect 7748 7414 7800 7420
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7760 7002 7788 7414
rect 7944 7206 7972 7482
rect 8036 7274 8064 7686
rect 8024 7268 8076 7274
rect 8024 7210 8076 7216
rect 7932 7200 7984 7206
rect 7932 7142 7984 7148
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7380 6928 7432 6934
rect 7380 6870 7432 6876
rect 7840 6928 7892 6934
rect 7840 6870 7892 6876
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7194 5944 7250 5953
rect 7104 5908 7156 5914
rect 7194 5879 7250 5888
rect 7104 5850 7156 5856
rect 7012 5840 7064 5846
rect 7012 5782 7064 5788
rect 7196 5704 7248 5710
rect 7300 5692 7328 6190
rect 7248 5664 7328 5692
rect 7196 5646 7248 5652
rect 6920 5636 6972 5642
rect 6920 5578 6972 5584
rect 6932 4758 6960 5578
rect 7300 5370 7328 5664
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 6920 4752 6972 4758
rect 6920 4694 6972 4700
rect 6920 4480 6972 4486
rect 6918 4448 6920 4457
rect 6972 4448 6974 4457
rect 6918 4383 6974 4392
rect 7300 4214 7328 5306
rect 7392 4826 7420 6598
rect 7668 5846 7696 6802
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7564 5840 7616 5846
rect 7562 5808 7564 5817
rect 7656 5840 7708 5846
rect 7616 5808 7618 5817
rect 7656 5782 7708 5788
rect 7562 5743 7618 5752
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7484 4865 7512 4966
rect 7470 4856 7526 4865
rect 7380 4820 7432 4826
rect 7576 4826 7604 5743
rect 7668 5273 7696 5782
rect 7654 5264 7710 5273
rect 7654 5199 7710 5208
rect 7470 4791 7526 4800
rect 7564 4820 7616 4826
rect 7380 4762 7432 4768
rect 7484 4758 7512 4791
rect 7564 4762 7616 4768
rect 7472 4752 7524 4758
rect 7378 4720 7434 4729
rect 7472 4694 7524 4700
rect 7378 4655 7434 4664
rect 7288 4208 7340 4214
rect 7288 4150 7340 4156
rect 7392 4146 7420 4655
rect 7484 4282 7512 4694
rect 7760 4282 7788 6734
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7116 3738 7144 4082
rect 7656 4004 7708 4010
rect 7656 3946 7708 3952
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 6748 2650 6776 2926
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 7116 2582 7144 3674
rect 7668 3398 7696 3946
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 7378 3088 7434 3097
rect 7378 3023 7434 3032
rect 7392 2990 7420 3023
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 7104 2576 7156 2582
rect 6458 2544 6514 2553
rect 7104 2518 7156 2524
rect 6458 2479 6514 2488
rect 7852 610 7880 6870
rect 8036 6254 8064 7210
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 8024 4208 8076 4214
rect 8024 4150 8076 4156
rect 8036 3738 8064 4150
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 6920 604 6972 610
rect 6920 546 6972 552
rect 7564 604 7616 610
rect 7564 546 7616 552
rect 7840 604 7892 610
rect 7840 546 7892 552
rect 6932 480 6960 546
rect 7576 480 7604 546
rect 8128 480 8156 9454
rect 8312 9178 8340 9472
rect 8392 9454 8444 9460
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8772 9110 8800 22199
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10289 21168 10585 21188
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10690 17640 10746 17649
rect 10690 17575 10746 17584
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 9954 14376 10010 14385
rect 9954 14311 10010 14320
rect 9586 13424 9642 13433
rect 9586 13359 9642 13368
rect 9600 13161 9628 13359
rect 9586 13152 9642 13161
rect 9586 13087 9642 13096
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8850 12336 8906 12345
rect 8850 12271 8906 12280
rect 8208 9104 8260 9110
rect 8760 9104 8812 9110
rect 8208 9046 8260 9052
rect 8390 9072 8446 9081
rect 8220 8634 8248 9046
rect 8760 9046 8812 9052
rect 8390 9007 8446 9016
rect 8208 8628 8260 8634
rect 8260 8588 8340 8616
rect 8208 8570 8260 8576
rect 8312 8090 8340 8588
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8404 7954 8432 9007
rect 8772 8634 8800 9046
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8220 6662 8248 7278
rect 8404 7041 8432 7890
rect 8496 7410 8524 8502
rect 8666 7576 8722 7585
rect 8666 7511 8722 7520
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8390 7032 8446 7041
rect 8390 6967 8446 6976
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8404 6118 8432 6734
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8404 5778 8432 6054
rect 8392 5772 8444 5778
rect 8392 5714 8444 5720
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8392 4684 8444 4690
rect 8392 4626 8444 4632
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8206 4040 8262 4049
rect 8206 3975 8262 3984
rect 8220 3602 8248 3975
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8312 2650 8340 4422
rect 8404 4010 8432 4626
rect 8392 4004 8444 4010
rect 8392 3946 8444 3952
rect 8496 2961 8524 5510
rect 8574 5128 8630 5137
rect 8574 5063 8630 5072
rect 8588 4826 8616 5063
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 8680 3670 8708 7511
rect 8760 7200 8812 7206
rect 8760 7142 8812 7148
rect 8772 4185 8800 7142
rect 8758 4176 8814 4185
rect 8758 4111 8814 4120
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 8864 3210 8892 12271
rect 8956 11898 8984 12718
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 8944 11892 8996 11898
rect 8944 11834 8996 11840
rect 8956 10606 8984 11834
rect 9036 11144 9088 11150
rect 9034 11112 9036 11121
rect 9088 11112 9090 11121
rect 9034 11047 9090 11056
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 8956 10266 8984 10542
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 9140 8974 9168 12582
rect 9402 10704 9458 10713
rect 9402 10639 9458 10648
rect 9416 10470 9444 10639
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9402 10160 9458 10169
rect 9402 10095 9458 10104
rect 9416 9178 9444 10095
rect 9496 9376 9548 9382
rect 9496 9318 9548 9324
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9508 9042 9536 9318
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9140 8634 9168 8910
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9036 8356 9088 8362
rect 9036 8298 9088 8304
rect 9048 7750 9076 8298
rect 9324 7750 9352 8366
rect 9508 8362 9536 8978
rect 9496 8356 9548 8362
rect 9600 8344 9628 12582
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9784 11558 9812 12174
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 9784 11150 9812 11494
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9692 10441 9720 11018
rect 9784 10538 9812 11086
rect 9772 10532 9824 10538
rect 9772 10474 9824 10480
rect 9678 10432 9734 10441
rect 9678 10367 9734 10376
rect 9680 10192 9732 10198
rect 9678 10160 9680 10169
rect 9732 10160 9734 10169
rect 9678 10095 9734 10104
rect 9862 10160 9918 10169
rect 9862 10095 9918 10104
rect 9876 9994 9904 10095
rect 9864 9988 9916 9994
rect 9864 9930 9916 9936
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9692 9217 9720 9590
rect 9772 9444 9824 9450
rect 9772 9386 9824 9392
rect 9784 9353 9812 9386
rect 9770 9344 9826 9353
rect 9770 9279 9826 9288
rect 9678 9208 9734 9217
rect 9678 9143 9734 9152
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9600 8316 9720 8344
rect 9496 8298 9548 8304
rect 9692 8022 9720 8316
rect 9680 8016 9732 8022
rect 9680 7958 9732 7964
rect 9784 7954 9812 8774
rect 9876 8129 9904 8842
rect 9862 8120 9918 8129
rect 9862 8055 9918 8064
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9770 7848 9826 7857
rect 9770 7783 9772 7792
rect 9824 7783 9826 7792
rect 9772 7754 9824 7760
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9048 7002 9076 7686
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 9036 6996 9088 7002
rect 9036 6938 9088 6944
rect 9036 5024 9088 5030
rect 9034 4992 9036 5001
rect 9088 4992 9090 5001
rect 9034 4927 9090 4936
rect 9140 4842 9168 7278
rect 9324 6730 9352 7686
rect 9772 7472 9824 7478
rect 9772 7414 9824 7420
rect 9496 7268 9548 7274
rect 9496 7210 9548 7216
rect 9312 6724 9364 6730
rect 9312 6666 9364 6672
rect 9324 6458 9352 6666
rect 9508 6474 9536 7210
rect 9678 6488 9734 6497
rect 9312 6452 9364 6458
rect 9508 6446 9678 6474
rect 9678 6423 9734 6432
rect 9312 6394 9364 6400
rect 9324 5778 9352 6394
rect 9678 6352 9734 6361
rect 9678 6287 9734 6296
rect 9312 5772 9364 5778
rect 9312 5714 9364 5720
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9310 5128 9366 5137
rect 9310 5063 9366 5072
rect 8680 3182 8892 3210
rect 9048 4814 9168 4842
rect 8482 2952 8538 2961
rect 8482 2887 8538 2896
rect 8496 2854 8524 2887
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8680 480 8708 3182
rect 9048 678 9076 4814
rect 9324 4282 9352 5063
rect 9416 4554 9444 5510
rect 9692 5386 9720 6287
rect 9784 6254 9812 7414
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9784 5914 9812 6190
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9692 5358 9812 5386
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9404 4548 9456 4554
rect 9404 4490 9456 4496
rect 9312 4276 9364 4282
rect 9312 4218 9364 4224
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 9126 3496 9182 3505
rect 9126 3431 9182 3440
rect 9140 3194 9168 3431
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9036 672 9088 678
rect 9036 614 9088 620
rect 9232 480 9260 3946
rect 9324 3777 9352 4218
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 9310 3768 9366 3777
rect 9416 3738 9444 3946
rect 9508 3890 9536 4762
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9600 4214 9628 4422
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 9692 4049 9720 5238
rect 9784 4078 9812 5358
rect 9876 4826 9904 6938
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9862 4720 9918 4729
rect 9862 4655 9918 4664
rect 9772 4072 9824 4078
rect 9678 4040 9734 4049
rect 9772 4014 9824 4020
rect 9678 3975 9734 3984
rect 9772 3936 9824 3942
rect 9508 3862 9720 3890
rect 9876 3913 9904 4655
rect 9772 3878 9824 3884
rect 9862 3904 9918 3913
rect 9310 3703 9366 3712
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9588 3392 9640 3398
rect 9692 3369 9720 3862
rect 9588 3334 9640 3340
rect 9678 3360 9734 3369
rect 9600 3210 9628 3334
rect 9678 3295 9734 3304
rect 9678 3224 9734 3233
rect 9600 3182 9678 3210
rect 9678 3159 9734 3168
rect 9784 3074 9812 3878
rect 9862 3839 9918 3848
rect 9876 3670 9904 3839
rect 9864 3664 9916 3670
rect 9864 3606 9916 3612
rect 9692 3046 9812 3074
rect 9496 2984 9548 2990
rect 9496 2926 9548 2932
rect 9508 2514 9536 2926
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9600 2650 9628 2790
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9692 2106 9720 3046
rect 9968 2802 9996 14311
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10140 12368 10192 12374
rect 10140 12310 10192 12316
rect 10152 11558 10180 12310
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 10060 10305 10088 11494
rect 10152 10810 10180 11494
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10046 10296 10102 10305
rect 10289 10288 10585 10308
rect 10046 10231 10102 10240
rect 10232 10192 10284 10198
rect 10232 10134 10284 10140
rect 10244 9586 10272 10134
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10046 8256 10102 8265
rect 10046 8191 10102 8200
rect 10060 7410 10088 8191
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10140 8016 10192 8022
rect 10140 7958 10192 7964
rect 10324 8016 10376 8022
rect 10324 7958 10376 7964
rect 10152 7546 10180 7958
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10336 7478 10364 7958
rect 10324 7472 10376 7478
rect 10324 7414 10376 7420
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 10704 7342 10732 17575
rect 10782 13288 10838 13297
rect 10782 13223 10838 13232
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10289 7100 10585 7120
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10289 7024 10585 7044
rect 10704 6866 10732 7278
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10060 6633 10088 6802
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10046 6624 10102 6633
rect 10046 6559 10102 6568
rect 10060 6225 10088 6559
rect 10046 6216 10102 6225
rect 10046 6151 10102 6160
rect 10152 6089 10180 6734
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10138 6080 10194 6089
rect 10138 6015 10194 6024
rect 10152 5914 10180 6015
rect 10289 6012 10585 6032
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 10060 5370 10088 5714
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 10704 5250 10732 6598
rect 10796 5370 10824 13223
rect 10980 12594 11008 23695
rect 11702 19816 11758 19825
rect 11702 19751 11758 19760
rect 11242 13016 11298 13025
rect 11242 12951 11298 12960
rect 10980 12566 11100 12594
rect 11072 12356 11100 12566
rect 10980 12328 11100 12356
rect 10876 8288 10928 8294
rect 10876 8230 10928 8236
rect 10888 8022 10916 8230
rect 10876 8016 10928 8022
rect 10876 7958 10928 7964
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 10888 6905 10916 7822
rect 10980 7562 11008 12328
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 11164 11286 11192 12038
rect 11256 11898 11284 12951
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 11164 10266 11192 11222
rect 11152 10260 11204 10266
rect 11152 10202 11204 10208
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 11164 9081 11192 9862
rect 11426 9616 11482 9625
rect 11426 9551 11482 9560
rect 11244 9444 11296 9450
rect 11244 9386 11296 9392
rect 11150 9072 11206 9081
rect 11150 9007 11206 9016
rect 11256 8838 11284 9386
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11348 8906 11376 9318
rect 11336 8900 11388 8906
rect 11336 8842 11388 8848
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 11256 7721 11284 8774
rect 11336 7744 11388 7750
rect 11242 7712 11298 7721
rect 11336 7686 11388 7692
rect 11242 7647 11298 7656
rect 10980 7534 11284 7562
rect 10968 7472 11020 7478
rect 10968 7414 11020 7420
rect 10874 6896 10930 6905
rect 10874 6831 10930 6840
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10888 5846 10916 6054
rect 10876 5840 10928 5846
rect 10876 5782 10928 5788
rect 10980 5409 11008 7414
rect 11060 6792 11112 6798
rect 11058 6760 11060 6769
rect 11112 6760 11114 6769
rect 11058 6695 11114 6704
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 11256 5794 11284 7534
rect 11348 7410 11376 7686
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 11348 7313 11376 7346
rect 11334 7304 11390 7313
rect 11334 7239 11390 7248
rect 11348 6934 11376 7239
rect 11336 6928 11388 6934
rect 11336 6870 11388 6876
rect 11348 6458 11376 6870
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 10966 5400 11022 5409
rect 10784 5364 10836 5370
rect 11072 5370 11100 5782
rect 11256 5766 11376 5794
rect 11242 5672 11298 5681
rect 11242 5607 11298 5616
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 10966 5335 11022 5344
rect 11060 5364 11112 5370
rect 10784 5306 10836 5312
rect 11060 5306 11112 5312
rect 10704 5222 10916 5250
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10784 5160 10836 5166
rect 10784 5102 10836 5108
rect 10140 5092 10192 5098
rect 10140 5034 10192 5040
rect 10152 4486 10180 5034
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10232 4752 10284 4758
rect 10232 4694 10284 4700
rect 10140 4480 10192 4486
rect 10140 4422 10192 4428
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 9876 2774 9996 2802
rect 9876 2666 9904 2774
rect 9784 2638 9904 2666
rect 9680 2100 9732 2106
rect 9680 2042 9732 2048
rect 9784 480 9812 2638
rect 10060 2582 10088 4082
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 10152 3670 10180 4014
rect 10244 4010 10272 4694
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 10428 4282 10456 4626
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10232 4004 10284 4010
rect 10232 3946 10284 3952
rect 10289 3836 10585 3856
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10140 3664 10192 3670
rect 10140 3606 10192 3612
rect 10704 3194 10732 5102
rect 10692 3188 10744 3194
rect 10692 3130 10744 3136
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10289 2672 10585 2692
rect 10796 2632 10824 5102
rect 10888 4298 10916 5222
rect 11164 4826 11192 5510
rect 11256 5166 11284 5607
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 10888 4270 11008 4298
rect 10876 4208 10928 4214
rect 10874 4176 10876 4185
rect 10928 4176 10930 4185
rect 10874 4111 10930 4120
rect 10876 4004 10928 4010
rect 10876 3946 10928 3952
rect 10336 2604 10824 2632
rect 10048 2576 10100 2582
rect 10046 2544 10048 2553
rect 10100 2544 10102 2553
rect 10046 2479 10102 2488
rect 10336 480 10364 2604
rect 10888 480 10916 3946
rect 10980 3346 11008 4270
rect 11164 4146 11192 4762
rect 11348 4758 11376 5766
rect 11440 5114 11468 9551
rect 11532 9518 11560 9998
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11532 7206 11560 7822
rect 11624 7392 11652 9522
rect 11716 9110 11744 19751
rect 11794 13832 11850 13841
rect 11794 13767 11850 13776
rect 11704 9104 11756 9110
rect 11704 9046 11756 9052
rect 11716 8634 11744 9046
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11624 7364 11744 7392
rect 11612 7268 11664 7274
rect 11612 7210 11664 7216
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 11532 6662 11560 7142
rect 11520 6656 11572 6662
rect 11520 6598 11572 6604
rect 11532 6254 11560 6598
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11520 5908 11572 5914
rect 11520 5850 11572 5856
rect 11532 5234 11560 5850
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11440 5086 11560 5114
rect 11428 5024 11480 5030
rect 11428 4966 11480 4972
rect 11336 4752 11388 4758
rect 11256 4712 11336 4740
rect 11256 4282 11284 4712
rect 11336 4694 11388 4700
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11244 4276 11296 4282
rect 11244 4218 11296 4224
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11348 4049 11376 4422
rect 11334 4040 11390 4049
rect 11334 3975 11336 3984
rect 11388 3975 11390 3984
rect 11336 3946 11388 3952
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 11072 3738 11100 3878
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 10980 3318 11100 3346
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 10980 1737 11008 3130
rect 11072 2689 11100 3318
rect 11150 3088 11206 3097
rect 11150 3023 11206 3032
rect 11058 2680 11114 2689
rect 11164 2650 11192 3023
rect 11058 2615 11114 2624
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11440 2009 11468 4966
rect 11532 2446 11560 5086
rect 11624 3670 11652 7210
rect 11716 4826 11744 7364
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 11716 4321 11744 4762
rect 11702 4312 11758 4321
rect 11702 4247 11704 4256
rect 11756 4247 11758 4256
rect 11704 4218 11756 4224
rect 11716 4187 11744 4218
rect 11808 3738 11836 13767
rect 12622 11792 12678 11801
rect 12622 11727 12678 11736
rect 12164 11552 12216 11558
rect 12164 11494 12216 11500
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 12084 10606 12112 10950
rect 12072 10600 12124 10606
rect 12072 10542 12124 10548
rect 12084 10198 12112 10542
rect 12072 10192 12124 10198
rect 12072 10134 12124 10140
rect 12084 9722 12112 10134
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 11980 9444 12032 9450
rect 11980 9386 12032 9392
rect 11888 9104 11940 9110
rect 11888 9046 11940 9052
rect 11900 8362 11928 9046
rect 11992 8974 12020 9386
rect 11980 8968 12032 8974
rect 11980 8910 12032 8916
rect 11888 8356 11940 8362
rect 11888 8298 11940 8304
rect 11900 7426 11928 8298
rect 11992 8090 12020 8910
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 11900 7398 12112 7426
rect 12084 5846 12112 7398
rect 12072 5840 12124 5846
rect 12072 5782 12124 5788
rect 11980 5636 12032 5642
rect 11980 5578 12032 5584
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11900 4758 11928 5306
rect 11888 4752 11940 4758
rect 11888 4694 11940 4700
rect 11796 3732 11848 3738
rect 11848 3692 11928 3720
rect 11796 3674 11848 3680
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11624 3194 11652 3606
rect 11796 3528 11848 3534
rect 11794 3496 11796 3505
rect 11848 3496 11850 3505
rect 11794 3431 11850 3440
rect 11900 3194 11928 3692
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 11888 3188 11940 3194
rect 11888 3130 11940 3136
rect 11520 2440 11572 2446
rect 11520 2382 11572 2388
rect 11426 2000 11482 2009
rect 11426 1935 11482 1944
rect 11426 1864 11482 1873
rect 11426 1799 11482 1808
rect 10966 1728 11022 1737
rect 10966 1663 11022 1672
rect 11440 480 11468 1799
rect 11992 480 12020 5578
rect 12084 5030 12112 5782
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 12084 4593 12112 4966
rect 12070 4584 12126 4593
rect 12070 4519 12126 4528
rect 12176 4146 12204 11494
rect 12348 11076 12400 11082
rect 12348 11018 12400 11024
rect 12360 10849 12388 11018
rect 12346 10840 12402 10849
rect 12346 10775 12402 10784
rect 12532 10736 12584 10742
rect 12532 10678 12584 10684
rect 12544 9625 12572 10678
rect 12530 9616 12586 9625
rect 12530 9551 12586 9560
rect 12256 8900 12308 8906
rect 12256 8842 12308 8848
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 12268 610 12296 8842
rect 12636 8634 12664 11727
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12622 7984 12678 7993
rect 12348 7948 12400 7954
rect 12622 7919 12678 7928
rect 12348 7890 12400 7896
rect 12360 7206 12388 7890
rect 12438 7576 12494 7585
rect 12636 7546 12664 7919
rect 12438 7511 12494 7520
rect 12624 7540 12676 7546
rect 12452 7342 12480 7511
rect 12624 7482 12676 7488
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12348 7200 12400 7206
rect 12348 7142 12400 7148
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12636 6662 12664 7142
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12348 5160 12400 5166
rect 12544 5148 12572 6190
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12400 5120 12572 5148
rect 12348 5102 12400 5108
rect 12544 4826 12572 5120
rect 12636 5030 12664 5510
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12544 3738 12572 4762
rect 12728 3942 12756 11494
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 13004 10470 13032 10950
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 13004 10169 13032 10406
rect 12990 10160 13046 10169
rect 12990 10095 13046 10104
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 13004 9518 13032 9862
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12992 9512 13044 9518
rect 12992 9454 13044 9460
rect 12820 8906 12848 9454
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 13004 8401 13032 8774
rect 12990 8392 13046 8401
rect 12990 8327 13046 8336
rect 12900 7744 12952 7750
rect 12898 7712 12900 7721
rect 12952 7712 12954 7721
rect 12898 7647 12954 7656
rect 13174 6896 13230 6905
rect 13174 6831 13176 6840
rect 13228 6831 13230 6840
rect 13176 6802 13228 6808
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 12820 6254 12848 6394
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12806 6080 12862 6089
rect 12806 6015 12862 6024
rect 12820 4282 12848 6015
rect 12990 5400 13046 5409
rect 12990 5335 13046 5344
rect 13004 4593 13032 5335
rect 12990 4584 13046 4593
rect 12990 4519 13046 4528
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 13004 4010 13032 4519
rect 13096 4486 13124 6598
rect 13280 5778 13308 24890
rect 14004 24880 14056 24886
rect 14004 24822 14056 24828
rect 13818 16008 13874 16017
rect 13818 15943 13874 15952
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13372 9110 13400 11086
rect 13360 9104 13412 9110
rect 13360 9046 13412 9052
rect 13372 8566 13400 9046
rect 13544 8900 13596 8906
rect 13544 8842 13596 8848
rect 13360 8560 13412 8566
rect 13360 8502 13412 8508
rect 13556 8294 13584 8842
rect 13636 8356 13688 8362
rect 13636 8298 13688 8304
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13556 7954 13584 8230
rect 13544 7948 13596 7954
rect 13464 7908 13544 7936
rect 13464 6458 13492 7908
rect 13544 7890 13596 7896
rect 13544 7200 13596 7206
rect 13542 7168 13544 7177
rect 13596 7168 13598 7177
rect 13542 7103 13598 7112
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13544 6248 13596 6254
rect 13544 6190 13596 6196
rect 13556 5846 13584 6190
rect 13544 5840 13596 5846
rect 13358 5808 13414 5817
rect 13268 5772 13320 5778
rect 13544 5782 13596 5788
rect 13358 5743 13414 5752
rect 13268 5714 13320 5720
rect 13266 4992 13322 5001
rect 13266 4927 13322 4936
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 13096 4146 13124 4422
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 12992 4004 13044 4010
rect 12992 3946 13044 3952
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 13280 3738 13308 4927
rect 13372 4622 13400 5743
rect 13452 5568 13504 5574
rect 13452 5510 13504 5516
rect 13464 4758 13492 5510
rect 13452 4752 13504 4758
rect 13452 4694 13504 4700
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13372 4282 13400 4558
rect 13360 4276 13412 4282
rect 13360 4218 13412 4224
rect 13464 3913 13492 4694
rect 13450 3904 13506 3913
rect 13450 3839 13506 3848
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 12544 2990 12572 3674
rect 12716 3528 12768 3534
rect 12622 3496 12678 3505
rect 12716 3470 12768 3476
rect 12622 3431 12678 3440
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 12544 2650 12572 2926
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12544 2514 12572 2586
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 12636 1578 12664 3431
rect 12728 2990 12756 3470
rect 13280 3466 13308 3674
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13268 3460 13320 3466
rect 13268 3402 13320 3408
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12820 1601 12848 3334
rect 13372 3194 13400 3470
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13082 2000 13138 2009
rect 13082 1935 13138 1944
rect 12544 1550 12664 1578
rect 12806 1592 12862 1601
rect 12256 604 12308 610
rect 12256 546 12308 552
rect 12544 480 12572 1550
rect 12806 1527 12862 1536
rect 13096 480 13124 1935
rect 13648 480 13676 8298
rect 13832 8090 13860 15943
rect 13910 10568 13966 10577
rect 13910 10503 13966 10512
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13832 7274 13860 8026
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13924 7002 13952 10503
rect 13912 6996 13964 7002
rect 13912 6938 13964 6944
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13740 5642 13768 6802
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 13728 5636 13780 5642
rect 13728 5578 13780 5584
rect 13832 5370 13860 5782
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 13924 5370 13952 5714
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 13726 5264 13782 5273
rect 13726 5199 13782 5208
rect 13740 4554 13768 5199
rect 13728 4548 13780 4554
rect 13728 4490 13780 4496
rect 14016 4078 14044 24822
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15382 20904 15438 20913
rect 15382 20839 15438 20848
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14108 9042 14136 9318
rect 14832 9172 14884 9178
rect 14832 9114 14884 9120
rect 14096 9036 14148 9042
rect 14096 8978 14148 8984
rect 14108 8362 14136 8978
rect 14096 8356 14148 8362
rect 14096 8298 14148 8304
rect 14740 8288 14792 8294
rect 14740 8230 14792 8236
rect 14752 8022 14780 8230
rect 14740 8016 14792 8022
rect 14740 7958 14792 7964
rect 14372 7880 14424 7886
rect 14372 7822 14424 7828
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14200 4146 14228 7142
rect 14280 6656 14332 6662
rect 14278 6624 14280 6633
rect 14332 6624 14334 6633
rect 14278 6559 14334 6568
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 14016 3738 14044 4014
rect 14188 3936 14240 3942
rect 14188 3878 14240 3884
rect 14200 3777 14228 3878
rect 14186 3768 14242 3777
rect 14004 3732 14056 3738
rect 14186 3703 14242 3712
rect 14004 3674 14056 3680
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13832 2582 13860 3130
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 13820 2576 13872 2582
rect 14016 2553 14044 2586
rect 13820 2518 13872 2524
rect 14002 2544 14058 2553
rect 14002 2479 14058 2488
rect 14292 480 14320 6054
rect 14384 3602 14412 7822
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14476 7342 14504 7686
rect 14752 7410 14780 7958
rect 14844 7546 14872 9114
rect 15304 9110 15332 9998
rect 15292 9104 15344 9110
rect 15292 9046 15344 9052
rect 15396 8922 15424 20839
rect 15474 12880 15530 12889
rect 15474 12815 15530 12824
rect 15304 8894 15424 8922
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14832 7540 14884 7546
rect 14832 7482 14884 7488
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 15028 7002 15056 7346
rect 15016 6996 15068 7002
rect 15016 6938 15068 6944
rect 14832 6860 14884 6866
rect 14832 6802 14884 6808
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14660 6225 14688 6598
rect 14646 6216 14702 6225
rect 14646 6151 14702 6160
rect 14844 6118 14872 6802
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15304 6474 15332 8894
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15396 7993 15424 8774
rect 15382 7984 15438 7993
rect 15382 7919 15438 7928
rect 15488 6730 15516 12815
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15580 10985 15608 11018
rect 15566 10976 15622 10985
rect 15566 10911 15622 10920
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15476 6724 15528 6730
rect 15476 6666 15528 6672
rect 15304 6458 15424 6474
rect 15304 6452 15436 6458
rect 15304 6446 15384 6452
rect 15384 6394 15436 6400
rect 15292 6384 15344 6390
rect 15292 6326 15344 6332
rect 14832 6112 14884 6118
rect 14832 6054 14884 6060
rect 15304 5846 15332 6326
rect 15384 6112 15436 6118
rect 15384 6054 15436 6060
rect 15292 5840 15344 5846
rect 15292 5782 15344 5788
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 14844 5370 14872 5646
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 14832 5364 14884 5370
rect 14832 5306 14884 5312
rect 15304 5114 15332 5782
rect 15120 5086 15332 5114
rect 15120 4826 15148 5086
rect 15108 4820 15160 4826
rect 15108 4762 15160 4768
rect 14648 4616 14700 4622
rect 14646 4584 14648 4593
rect 14700 4584 14702 4593
rect 14646 4519 14702 4528
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14476 3738 14504 4082
rect 15396 3942 15424 6054
rect 15580 5817 15608 9318
rect 15660 9104 15712 9110
rect 15660 9046 15712 9052
rect 15672 8634 15700 9046
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15566 5808 15622 5817
rect 15566 5743 15622 5752
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15488 5166 15516 5510
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15488 4214 15516 5102
rect 15764 4826 15792 26250
rect 19622 25596 19918 25616
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 19622 22332 19918 22352
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 24122 21040 24178 21049
rect 24122 20975 24178 20984
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19522 13424 19578 13433
rect 19522 13359 19578 13368
rect 16396 11892 16448 11898
rect 16396 11834 16448 11840
rect 16212 11212 16264 11218
rect 16212 11154 16264 11160
rect 16224 10742 16252 11154
rect 16212 10736 16264 10742
rect 16210 10704 16212 10713
rect 16264 10704 16266 10713
rect 16210 10639 16266 10648
rect 16408 9654 16436 11834
rect 16670 11656 16726 11665
rect 16670 11591 16726 11600
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 16396 9648 16448 9654
rect 16500 9636 16528 11086
rect 16684 10606 16712 11591
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16948 10532 17000 10538
rect 16948 10474 17000 10480
rect 16500 9608 16712 9636
rect 16396 9590 16448 9596
rect 16684 9382 16712 9608
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 15948 8634 15976 8910
rect 16684 8634 16712 9114
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 15948 8090 15976 8570
rect 16212 8356 16264 8362
rect 16212 8298 16264 8304
rect 15936 8084 15988 8090
rect 15936 8026 15988 8032
rect 15948 7274 15976 8026
rect 16028 7948 16080 7954
rect 16028 7890 16080 7896
rect 16040 7342 16068 7890
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 15936 7268 15988 7274
rect 15936 7210 15988 7216
rect 15948 7002 15976 7210
rect 16224 7041 16252 8298
rect 16396 7268 16448 7274
rect 16396 7210 16448 7216
rect 16210 7032 16266 7041
rect 15936 6996 15988 7002
rect 16210 6967 16266 6976
rect 15936 6938 15988 6944
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 16316 6322 16344 6802
rect 16408 6798 16436 7210
rect 16856 7200 16908 7206
rect 16856 7142 16908 7148
rect 16868 6934 16896 7142
rect 16856 6928 16908 6934
rect 16856 6870 16908 6876
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 16408 6458 16436 6734
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16408 5778 16436 6394
rect 15936 5772 15988 5778
rect 15936 5714 15988 5720
rect 16396 5772 16448 5778
rect 16396 5714 16448 5720
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 15476 4208 15528 4214
rect 15476 4150 15528 4156
rect 15764 4078 15792 4762
rect 15752 4072 15804 4078
rect 15752 4014 15804 4020
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 14384 3194 14412 3538
rect 14660 3233 14688 3878
rect 14740 3664 14792 3670
rect 14738 3632 14740 3641
rect 14792 3632 14794 3641
rect 15856 3602 15884 4762
rect 15948 4690 15976 5714
rect 16408 5370 16436 5714
rect 16960 5409 16988 10474
rect 17868 9648 17920 9654
rect 17868 9590 17920 9596
rect 18050 9616 18106 9625
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17788 6458 17816 8910
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17788 6186 17816 6394
rect 17776 6180 17828 6186
rect 17776 6122 17828 6128
rect 17592 5704 17644 5710
rect 17590 5672 17592 5681
rect 17644 5672 17646 5681
rect 17590 5607 17646 5616
rect 17682 5536 17738 5545
rect 17682 5471 17738 5480
rect 16946 5400 17002 5409
rect 16396 5364 16448 5370
rect 16946 5335 17002 5344
rect 16396 5306 16448 5312
rect 17592 5160 17644 5166
rect 17590 5128 17592 5137
rect 17644 5128 17646 5137
rect 17590 5063 17646 5072
rect 16212 5024 16264 5030
rect 17224 5024 17276 5030
rect 16212 4966 16264 4972
rect 17222 4992 17224 5001
rect 17276 4992 17278 5001
rect 16224 4690 16252 4966
rect 17222 4927 17278 4936
rect 16394 4856 16450 4865
rect 16394 4791 16450 4800
rect 15936 4684 15988 4690
rect 15936 4626 15988 4632
rect 16212 4684 16264 4690
rect 16212 4626 16264 4632
rect 15948 4282 15976 4626
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 15936 4004 15988 4010
rect 15936 3946 15988 3952
rect 14738 3567 14794 3576
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 15568 3528 15620 3534
rect 15382 3496 15438 3505
rect 15568 3470 15620 3476
rect 15382 3431 15438 3440
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14646 3224 14702 3233
rect 14372 3188 14424 3194
rect 14956 3216 15252 3236
rect 14646 3159 14702 3168
rect 14372 3130 14424 3136
rect 14738 3088 14794 3097
rect 15396 3058 15424 3431
rect 15580 3097 15608 3470
rect 15658 3360 15714 3369
rect 15658 3295 15714 3304
rect 15566 3088 15622 3097
rect 14738 3023 14740 3032
rect 14792 3023 14794 3032
rect 15384 3052 15436 3058
rect 14740 2994 14792 3000
rect 15566 3023 15622 3032
rect 15384 2994 15436 3000
rect 14832 2984 14884 2990
rect 14830 2952 14832 2961
rect 14884 2952 14886 2961
rect 14830 2887 14886 2896
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 14648 2304 14700 2310
rect 14648 2246 14700 2252
rect 14660 1465 14688 2246
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15384 2100 15436 2106
rect 15384 2042 15436 2048
rect 14646 1456 14702 1465
rect 14646 1391 14702 1400
rect 14832 1148 14884 1154
rect 14832 1090 14884 1096
rect 14844 480 14872 1090
rect 15396 480 15424 2042
rect 15488 1465 15516 2450
rect 15474 1456 15530 1465
rect 15474 1391 15530 1400
rect 15672 1154 15700 3295
rect 15948 3194 15976 3946
rect 16224 3738 16252 4626
rect 16302 3904 16358 3913
rect 16302 3839 16358 3848
rect 16316 3738 16344 3839
rect 16212 3732 16264 3738
rect 16212 3674 16264 3680
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 15764 2145 15792 2382
rect 15750 2136 15806 2145
rect 15750 2071 15806 2080
rect 16408 1714 16436 4791
rect 17316 4480 17368 4486
rect 16486 4448 16542 4457
rect 17316 4422 17368 4428
rect 16486 4383 16542 4392
rect 16500 3194 16528 4383
rect 16764 4276 16816 4282
rect 16764 4218 16816 4224
rect 16776 3602 16804 4218
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 16960 3738 16988 4082
rect 17132 4072 17184 4078
rect 17130 4040 17132 4049
rect 17184 4040 17186 4049
rect 17328 4010 17356 4422
rect 17130 3975 17186 3984
rect 17316 4004 17368 4010
rect 17316 3946 17368 3952
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 16764 3596 16816 3602
rect 16764 3538 16816 3544
rect 16776 3194 16804 3538
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 16580 2984 16632 2990
rect 16580 2926 16632 2932
rect 16592 2650 16620 2926
rect 16960 2922 16988 3674
rect 17328 3670 17356 3946
rect 17316 3664 17368 3670
rect 17316 3606 17368 3612
rect 17590 3224 17646 3233
rect 17590 3159 17646 3168
rect 16948 2916 17000 2922
rect 16948 2858 17000 2864
rect 16762 2680 16818 2689
rect 16580 2644 16632 2650
rect 16762 2615 16818 2624
rect 16580 2586 16632 2592
rect 16776 2514 16804 2615
rect 17040 2576 17092 2582
rect 17038 2544 17040 2553
rect 17092 2544 17094 2553
rect 16764 2508 16816 2514
rect 17038 2479 17094 2488
rect 16764 2450 16816 2456
rect 16670 2136 16726 2145
rect 16670 2071 16672 2080
rect 16724 2071 16726 2080
rect 16854 2136 16910 2145
rect 16854 2071 16910 2080
rect 16672 2042 16724 2048
rect 16408 1686 16528 1714
rect 15660 1148 15712 1154
rect 15660 1090 15712 1096
rect 15936 604 15988 610
rect 15936 546 15988 552
rect 15948 480 15976 546
rect 16500 480 16528 1686
rect 16868 1601 16896 2071
rect 16854 1592 16910 1601
rect 16854 1527 16910 1536
rect 17038 1592 17094 1601
rect 17038 1527 17094 1536
rect 17052 480 17080 1527
rect 17604 480 17632 3159
rect 17696 3058 17724 5471
rect 17880 4826 17908 9590
rect 18050 9551 18106 9560
rect 18064 9518 18092 9551
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 18328 9444 18380 9450
rect 18328 9386 18380 9392
rect 18340 9042 18368 9386
rect 18696 9376 18748 9382
rect 18696 9318 18748 9324
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 18340 8634 18368 8978
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 17958 8392 18014 8401
rect 17958 8327 18014 8336
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 17774 4584 17830 4593
rect 17972 4570 18000 8327
rect 18326 7984 18382 7993
rect 18326 7919 18328 7928
rect 18380 7919 18382 7928
rect 18328 7890 18380 7896
rect 18144 7744 18196 7750
rect 18144 7686 18196 7692
rect 18050 7576 18106 7585
rect 18050 7511 18106 7520
rect 18064 7410 18092 7511
rect 18052 7404 18104 7410
rect 18052 7346 18104 7352
rect 18156 7342 18184 7686
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 18156 6730 18184 7278
rect 18340 7002 18368 7890
rect 18328 6996 18380 7002
rect 18328 6938 18380 6944
rect 18144 6724 18196 6730
rect 18144 6666 18196 6672
rect 18156 6474 18184 6666
rect 18156 6446 18276 6474
rect 18144 6384 18196 6390
rect 18144 6326 18196 6332
rect 18156 5778 18184 6326
rect 18248 6322 18276 6446
rect 18236 6316 18288 6322
rect 18236 6258 18288 6264
rect 18248 5914 18276 6258
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 18144 5772 18196 5778
rect 18144 5714 18196 5720
rect 18708 5166 18736 9318
rect 19156 8832 19208 8838
rect 19156 8774 19208 8780
rect 18878 7032 18934 7041
rect 18878 6967 18934 6976
rect 18788 5704 18840 5710
rect 18786 5672 18788 5681
rect 18840 5672 18842 5681
rect 18786 5607 18842 5616
rect 18328 5160 18380 5166
rect 18328 5102 18380 5108
rect 18696 5160 18748 5166
rect 18696 5102 18748 5108
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18248 4865 18276 4966
rect 18234 4856 18290 4865
rect 18234 4791 18290 4800
rect 18236 4752 18288 4758
rect 18234 4720 18236 4729
rect 18288 4720 18290 4729
rect 18234 4655 18290 4664
rect 17972 4542 18276 4570
rect 17774 4519 17830 4528
rect 17788 4146 17816 4519
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 17684 3052 17736 3058
rect 17684 2994 17736 3000
rect 17972 2990 18000 3334
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 18142 2952 18198 2961
rect 17972 2650 18000 2926
rect 18142 2887 18198 2896
rect 17960 2644 18012 2650
rect 17960 2586 18012 2592
rect 18156 480 18184 2887
rect 18248 2514 18276 4542
rect 18340 4146 18368 5102
rect 18604 4752 18656 4758
rect 18604 4694 18656 4700
rect 18512 4480 18564 4486
rect 18512 4422 18564 4428
rect 18524 4321 18552 4422
rect 18510 4312 18566 4321
rect 18510 4247 18566 4256
rect 18328 4140 18380 4146
rect 18328 4082 18380 4088
rect 18510 3768 18566 3777
rect 18616 3754 18644 4694
rect 18892 4622 18920 6967
rect 18972 5772 19024 5778
rect 18972 5714 19024 5720
rect 18984 5370 19012 5714
rect 18972 5364 19024 5370
rect 18972 5306 19024 5312
rect 18880 4616 18932 4622
rect 18880 4558 18932 4564
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 18892 4282 18920 4558
rect 19076 4282 19104 4558
rect 18880 4276 18932 4282
rect 18880 4218 18932 4224
rect 19064 4276 19116 4282
rect 19064 4218 19116 4224
rect 19168 4049 19196 8774
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19352 6866 19380 7822
rect 19430 7304 19486 7313
rect 19430 7239 19486 7248
rect 19444 7206 19472 7239
rect 19432 7200 19484 7206
rect 19432 7142 19484 7148
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 19352 6458 19380 6802
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 19444 6089 19472 6190
rect 19430 6080 19486 6089
rect 19430 6015 19486 6024
rect 19248 5024 19300 5030
rect 19248 4966 19300 4972
rect 19154 4040 19210 4049
rect 18696 4004 18748 4010
rect 19154 3975 19210 3984
rect 18696 3946 18748 3952
rect 18566 3726 18644 3754
rect 18510 3703 18566 3712
rect 18524 3670 18552 3703
rect 18512 3664 18564 3670
rect 18418 3632 18474 3641
rect 18512 3606 18564 3612
rect 18602 3632 18658 3641
rect 18418 3567 18420 3576
rect 18472 3567 18474 3576
rect 18602 3567 18658 3576
rect 18420 3538 18472 3544
rect 18616 2582 18644 3567
rect 18604 2576 18656 2582
rect 18604 2518 18656 2524
rect 18236 2508 18288 2514
rect 18236 2450 18288 2456
rect 18708 480 18736 3946
rect 19260 480 19288 4966
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 19352 3369 19380 4014
rect 19536 3942 19564 13359
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 20810 11248 20866 11257
rect 20810 11183 20866 11192
rect 19982 10976 20038 10985
rect 19982 10911 20038 10920
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19800 5704 19852 5710
rect 19800 5646 19852 5652
rect 19812 5545 19840 5646
rect 19798 5536 19854 5545
rect 19798 5471 19854 5480
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19430 3768 19486 3777
rect 19622 3760 19918 3780
rect 19996 3738 20024 10911
rect 20442 8528 20498 8537
rect 20442 8463 20498 8472
rect 20258 5400 20314 5409
rect 20258 5335 20314 5344
rect 20272 5166 20300 5335
rect 20260 5160 20312 5166
rect 20260 5102 20312 5108
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 19430 3703 19432 3712
rect 19484 3703 19486 3712
rect 19984 3732 20036 3738
rect 19432 3674 19484 3680
rect 19984 3674 20036 3680
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 19338 3360 19394 3369
rect 19338 3295 19394 3304
rect 19996 3194 20024 3538
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 19984 3052 20036 3058
rect 19984 2994 20036 3000
rect 19432 2848 19484 2854
rect 19430 2816 19432 2825
rect 19484 2816 19486 2825
rect 19430 2751 19486 2760
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19996 2650 20024 2994
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 20088 2530 20116 4966
rect 20260 4072 20312 4078
rect 20260 4014 20312 4020
rect 20350 4040 20406 4049
rect 20272 3942 20300 4014
rect 20350 3975 20406 3984
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 20272 3505 20300 3878
rect 20258 3496 20314 3505
rect 20258 3431 20314 3440
rect 20168 3392 20220 3398
rect 20168 3334 20220 3340
rect 19616 2508 19668 2514
rect 19616 2450 19668 2456
rect 19812 2502 20116 2530
rect 19432 2304 19484 2310
rect 19432 2246 19484 2252
rect 19444 1465 19472 2246
rect 19628 1873 19656 2450
rect 19614 1864 19670 1873
rect 19614 1799 19670 1808
rect 19430 1456 19486 1465
rect 19430 1391 19486 1400
rect 19812 480 19840 2502
rect 20180 1329 20208 3334
rect 20166 1320 20222 1329
rect 20166 1255 20222 1264
rect 20364 480 20392 3975
rect 20456 3058 20484 8463
rect 20534 7440 20590 7449
rect 20534 7375 20590 7384
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 20548 2990 20576 7375
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20640 3913 20668 6598
rect 20626 3904 20682 3913
rect 20626 3839 20682 3848
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 20536 2984 20588 2990
rect 20536 2926 20588 2932
rect 20536 2440 20588 2446
rect 20534 2408 20536 2417
rect 20588 2408 20590 2417
rect 20534 2343 20590 2352
rect 20732 2106 20760 3538
rect 20824 3534 20852 11183
rect 20902 10024 20958 10033
rect 20902 9959 20958 9968
rect 20916 7954 20944 9959
rect 20904 7948 20956 7954
rect 20904 7890 20956 7896
rect 20916 7546 20944 7890
rect 22008 7880 22060 7886
rect 21362 7848 21418 7857
rect 22008 7822 22060 7828
rect 21362 7783 21418 7792
rect 20904 7540 20956 7546
rect 20904 7482 20956 7488
rect 21376 7342 21404 7783
rect 21364 7336 21416 7342
rect 21364 7278 21416 7284
rect 21640 7268 21692 7274
rect 21640 7210 21692 7216
rect 20904 6180 20956 6186
rect 20904 6122 20956 6128
rect 20916 5778 20944 6122
rect 20904 5772 20956 5778
rect 20904 5714 20956 5720
rect 20916 5370 20944 5714
rect 21362 5672 21418 5681
rect 21362 5607 21418 5616
rect 21088 5568 21140 5574
rect 21088 5510 21140 5516
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 20996 4684 21048 4690
rect 20996 4626 21048 4632
rect 20904 4480 20956 4486
rect 20904 4422 20956 4428
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 20812 3392 20864 3398
rect 20812 3334 20864 3340
rect 20824 3233 20852 3334
rect 20810 3224 20866 3233
rect 20810 3159 20866 3168
rect 20720 2100 20772 2106
rect 20720 2042 20772 2048
rect 20916 480 20944 4422
rect 21008 3942 21036 4626
rect 20996 3936 21048 3942
rect 20996 3878 21048 3884
rect 21008 3641 21036 3878
rect 20994 3632 21050 3641
rect 20994 3567 21050 3576
rect 20996 3528 21048 3534
rect 20996 3470 21048 3476
rect 21008 2650 21036 3470
rect 21100 2825 21128 5510
rect 21376 5166 21404 5607
rect 21364 5160 21416 5166
rect 21364 5102 21416 5108
rect 21652 4049 21680 7210
rect 22020 5250 22048 7822
rect 24136 7585 24164 20975
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24289 11920 24585 11940
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24289 8732 24585 8752
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24122 7576 24178 7585
rect 24289 7568 24585 7588
rect 24122 7511 24178 7520
rect 24136 6254 24164 7511
rect 24766 7032 24822 7041
rect 24766 6967 24822 6976
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24780 6254 24808 6967
rect 25504 6384 25556 6390
rect 25502 6352 25504 6361
rect 25556 6352 25558 6361
rect 25502 6287 25558 6296
rect 24124 6248 24176 6254
rect 24124 6190 24176 6196
rect 24768 6248 24820 6254
rect 24768 6190 24820 6196
rect 24136 5914 24164 6190
rect 24124 5908 24176 5914
rect 24124 5850 24176 5856
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 22466 5264 22522 5273
rect 22020 5222 22140 5250
rect 22112 5166 22140 5222
rect 22466 5199 22522 5208
rect 22100 5160 22152 5166
rect 22100 5102 22152 5108
rect 22008 5092 22060 5098
rect 22008 5034 22060 5040
rect 21730 4176 21786 4185
rect 22020 4162 22048 5034
rect 22480 4690 22508 5199
rect 23572 5024 23624 5030
rect 23572 4966 23624 4972
rect 22468 4684 22520 4690
rect 22468 4626 22520 4632
rect 22480 4282 22508 4626
rect 23478 4448 23534 4457
rect 23478 4383 23534 4392
rect 22742 4312 22798 4321
rect 22468 4276 22520 4282
rect 22742 4247 22798 4256
rect 22468 4218 22520 4224
rect 22020 4134 22140 4162
rect 21730 4111 21786 4120
rect 21744 4078 21772 4111
rect 21732 4072 21784 4078
rect 21638 4040 21694 4049
rect 21732 4014 21784 4020
rect 21638 3975 21694 3984
rect 22008 4004 22060 4010
rect 22008 3946 22060 3952
rect 21546 3904 21602 3913
rect 21546 3839 21602 3848
rect 21086 2816 21142 2825
rect 21086 2751 21142 2760
rect 20996 2644 21048 2650
rect 20996 2586 21048 2592
rect 21180 2508 21232 2514
rect 21180 2450 21232 2456
rect 21192 2009 21220 2450
rect 21178 2000 21234 2009
rect 21178 1935 21234 1944
rect 21560 480 21588 3839
rect 22020 3641 22048 3946
rect 22006 3632 22062 3641
rect 21640 3596 21692 3602
rect 22006 3567 22062 3576
rect 21640 3538 21692 3544
rect 21652 3194 21680 3538
rect 21640 3188 21692 3194
rect 21640 3130 21692 3136
rect 21822 3088 21878 3097
rect 21822 3023 21878 3032
rect 21836 2990 21864 3023
rect 21824 2984 21876 2990
rect 21824 2926 21876 2932
rect 22006 2952 22062 2961
rect 22006 2887 22062 2896
rect 22020 2854 22048 2887
rect 22008 2848 22060 2854
rect 22008 2790 22060 2796
rect 22112 480 22140 4134
rect 22756 3602 22784 4247
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 22756 3194 22784 3538
rect 23204 3392 23256 3398
rect 23204 3334 23256 3340
rect 22744 3188 22796 3194
rect 22744 3130 22796 3136
rect 22650 2816 22706 2825
rect 22650 2751 22706 2760
rect 22282 2544 22338 2553
rect 22282 2479 22284 2488
rect 22336 2479 22338 2488
rect 22284 2450 22336 2456
rect 22468 2304 22520 2310
rect 22468 2246 22520 2252
rect 22480 1601 22508 2246
rect 22466 1592 22522 1601
rect 22466 1527 22522 1536
rect 22664 480 22692 2751
rect 23216 480 23244 3334
rect 23492 3194 23520 4383
rect 23584 3890 23612 4966
rect 23756 4684 23808 4690
rect 23756 4626 23808 4632
rect 23768 4282 23796 4626
rect 25412 4480 25464 4486
rect 25412 4422 25464 4428
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 23756 4276 23808 4282
rect 23756 4218 23808 4224
rect 23664 4072 23716 4078
rect 23662 4040 23664 4049
rect 24768 4072 24820 4078
rect 23716 4040 23718 4049
rect 24768 4014 24820 4020
rect 23662 3975 23718 3984
rect 24124 3936 24176 3942
rect 23584 3862 23704 3890
rect 24124 3878 24176 3884
rect 23480 3188 23532 3194
rect 23480 3130 23532 3136
rect 23492 2990 23520 3130
rect 23480 2984 23532 2990
rect 23480 2926 23532 2932
rect 23676 2530 23704 3862
rect 24032 3596 24084 3602
rect 24032 3538 24084 3544
rect 24044 2990 24072 3538
rect 24032 2984 24084 2990
rect 24032 2926 24084 2932
rect 23676 2502 23796 2530
rect 23768 480 23796 2502
rect 24032 2508 24084 2514
rect 24032 2450 24084 2456
rect 24044 2145 24072 2450
rect 24030 2136 24086 2145
rect 24030 2071 24086 2080
rect 24136 1986 24164 3878
rect 24780 3670 24808 4014
rect 24768 3664 24820 3670
rect 24768 3606 24820 3612
rect 25134 3632 25190 3641
rect 25134 3567 25136 3576
rect 25188 3567 25190 3576
rect 25136 3538 25188 3544
rect 24952 3392 25004 3398
rect 24952 3334 25004 3340
rect 24289 3292 24585 3312
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24768 2984 24820 2990
rect 24768 2926 24820 2932
rect 24780 2582 24808 2926
rect 24768 2576 24820 2582
rect 24768 2518 24820 2524
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24136 1958 24348 1986
rect 24320 480 24348 1958
rect 24964 1714 24992 3334
rect 25148 3194 25176 3538
rect 25136 3188 25188 3194
rect 25136 3130 25188 3136
rect 25044 2916 25096 2922
rect 25044 2858 25096 2864
rect 25056 2514 25084 2858
rect 25136 2848 25188 2854
rect 25134 2816 25136 2825
rect 25188 2816 25190 2825
rect 25134 2751 25190 2760
rect 25044 2508 25096 2514
rect 25044 2450 25096 2456
rect 24872 1686 24992 1714
rect 24872 480 24900 1686
rect 25424 480 25452 4422
rect 25964 3936 26016 3942
rect 25964 3878 26016 3884
rect 25976 480 26004 3878
rect 27066 2816 27122 2825
rect 27066 2751 27122 2760
rect 26516 2372 26568 2378
rect 26516 2314 26568 2320
rect 26528 480 26556 2314
rect 27080 480 27108 2751
rect 27618 1728 27674 1737
rect 27618 1663 27674 1672
rect 27632 480 27660 1663
rect 3146 368 3202 377
rect 3146 303 3202 312
rect 3606 0 3662 480
rect 4158 0 4214 480
rect 4710 0 4766 480
rect 5262 0 5318 480
rect 5814 0 5870 480
rect 6366 0 6422 480
rect 6918 0 6974 480
rect 7562 0 7618 480
rect 8114 0 8170 480
rect 8666 0 8722 480
rect 9218 0 9274 480
rect 9770 0 9826 480
rect 10322 0 10378 480
rect 10874 0 10930 480
rect 11426 0 11482 480
rect 11978 0 12034 480
rect 12530 0 12586 480
rect 13082 0 13138 480
rect 13634 0 13690 480
rect 14278 0 14334 480
rect 14830 0 14886 480
rect 15382 0 15438 480
rect 15934 0 15990 480
rect 16486 0 16542 480
rect 17038 0 17094 480
rect 17590 0 17646 480
rect 18142 0 18198 480
rect 18694 0 18750 480
rect 19246 0 19302 480
rect 19798 0 19854 480
rect 20350 0 20406 480
rect 20902 0 20958 480
rect 21546 0 21602 480
rect 22098 0 22154 480
rect 22650 0 22706 480
rect 23202 0 23258 480
rect 23754 0 23810 480
rect 24306 0 24362 480
rect 24858 0 24914 480
rect 25410 0 25466 480
rect 25962 0 26018 480
rect 26514 0 26570 480
rect 27066 0 27122 480
rect 27618 0 27674 480
<< via2 >>
rect 3146 27512 3202 27568
rect 2962 26832 3018 26888
rect 570 24792 626 24848
rect 570 23704 626 23760
rect 1490 16632 1546 16688
rect 1766 15272 1822 15328
rect 570 9832 626 9888
rect 846 7248 902 7304
rect 294 4120 350 4176
rect 1398 6840 1454 6896
rect 1398 4936 1454 4992
rect 1306 3032 1362 3088
rect 2042 14320 2098 14376
rect 1766 9696 1822 9752
rect 1674 7520 1730 7576
rect 1582 7112 1638 7168
rect 1858 5752 1914 5808
rect 2318 12144 2374 12200
rect 2594 12280 2650 12336
rect 2594 9596 2596 9616
rect 2596 9596 2648 9616
rect 2648 9596 2650 9616
rect 2594 9560 2650 9596
rect 2134 6976 2190 7032
rect 1950 4664 2006 4720
rect 1490 992 1546 1048
rect 2226 4120 2282 4176
rect 2594 7792 2650 7848
rect 2870 8200 2926 8256
rect 3514 26152 3570 26208
rect 3422 25472 3478 25528
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 3422 24112 3478 24168
rect 3238 23432 3294 23488
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 10966 23704 11022 23760
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5998 22616 6054 22672
rect 3422 22208 3478 22264
rect 3422 22072 3478 22128
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 4066 20712 4122 20768
rect 3790 19352 3846 19408
rect 3422 17584 3478 17640
rect 3698 17312 3754 17368
rect 3238 15952 3294 16008
rect 3330 14592 3386 14648
rect 2686 6160 2742 6216
rect 2962 5788 2964 5808
rect 2964 5788 3016 5808
rect 3016 5788 3018 5808
rect 2962 5752 3018 5788
rect 3146 6024 3202 6080
rect 3054 5616 3110 5672
rect 2318 3304 2374 3360
rect 3146 4528 3202 4584
rect 3054 4156 3056 4176
rect 3056 4156 3108 4176
rect 3108 4156 3110 4176
rect 3054 4120 3110 4156
rect 2502 3460 2558 3496
rect 2502 3440 2504 3460
rect 2504 3440 2556 3460
rect 2556 3440 2558 3460
rect 2594 3168 2650 3224
rect 2962 3612 2964 3632
rect 2964 3612 3016 3632
rect 3016 3612 3018 3632
rect 2962 3576 3018 3612
rect 2962 1400 3018 1456
rect 3514 11328 3570 11384
rect 3606 5888 3662 5944
rect 3422 5344 3478 5400
rect 3606 5072 3662 5128
rect 3974 18672 4030 18728
rect 3882 17992 3938 18048
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 4066 15952 4122 16008
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 3974 13504 4030 13560
rect 3974 12824 4030 12880
rect 3974 12552 4030 12608
rect 4986 13232 5042 13288
rect 3790 10104 3846 10160
rect 4710 12416 4766 12472
rect 4158 12144 4214 12200
rect 3974 9152 4030 9208
rect 3974 8472 4030 8528
rect 4342 10240 4398 10296
rect 4434 9424 4490 9480
rect 3974 6432 4030 6488
rect 3698 4392 3754 4448
rect 3606 3304 3662 3360
rect 3330 3052 3386 3088
rect 3330 3032 3332 3052
rect 3332 3032 3384 3052
rect 3384 3032 3386 3052
rect 3238 2796 3240 2816
rect 3240 2796 3292 2816
rect 3292 2796 3294 2816
rect 3238 2760 3294 2796
rect 3974 5072 4030 5128
rect 4526 8200 4582 8256
rect 4526 7828 4528 7848
rect 4528 7828 4580 7848
rect 4580 7828 4582 7848
rect 4526 7792 4582 7828
rect 4526 7248 4582 7304
rect 4618 5364 4674 5400
rect 4618 5344 4620 5364
rect 4620 5344 4672 5364
rect 4672 5344 4674 5364
rect 4158 2352 4214 2408
rect 4710 4664 4766 4720
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 4986 11056 5042 11112
rect 5906 12416 5962 12472
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5446 9696 5502 9752
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5170 9324 5172 9344
rect 5172 9324 5224 9344
rect 5224 9324 5226 9344
rect 5170 9288 5226 9324
rect 5538 9172 5594 9208
rect 5538 9152 5540 9172
rect 5540 9152 5592 9172
rect 5592 9152 5594 9172
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5354 7520 5410 7576
rect 5262 7420 5264 7440
rect 5264 7420 5316 7440
rect 5316 7420 5318 7440
rect 5262 7384 5318 7420
rect 5354 7112 5410 7168
rect 5170 6840 5226 6896
rect 5354 6296 5410 6352
rect 5262 5244 5264 5264
rect 5264 5244 5316 5264
rect 5316 5244 5318 5264
rect 5262 5208 5318 5244
rect 5446 4800 5502 4856
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 8758 22208 8814 22264
rect 7838 13524 7894 13560
rect 7838 13504 7840 13524
rect 7840 13504 7892 13524
rect 7892 13504 7894 13524
rect 6090 12980 6146 13016
rect 6090 12960 6092 12980
rect 6092 12960 6144 12980
rect 6144 12960 6146 12980
rect 6274 11328 6330 11384
rect 8114 11600 8170 11656
rect 6366 10512 6422 10568
rect 7378 11056 7434 11112
rect 7378 10240 7434 10296
rect 8114 10376 8170 10432
rect 6182 9152 6238 9208
rect 5722 6724 5778 6760
rect 5722 6704 5724 6724
rect 5724 6704 5776 6724
rect 5776 6704 5778 6724
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 5998 4528 6054 4584
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5262 3884 5264 3904
rect 5264 3884 5316 3904
rect 5316 3884 5318 3904
rect 5262 3848 5318 3884
rect 5722 3712 5778 3768
rect 4802 3168 4858 3224
rect 4710 2896 4766 2952
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 5538 3032 5594 3088
rect 3698 1264 3754 1320
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6182 4276 6238 4312
rect 6182 4256 6184 4276
rect 6184 4256 6236 4276
rect 6236 4256 6238 4276
rect 6642 7656 6698 7712
rect 6366 2760 6422 2816
rect 8022 10240 8078 10296
rect 7562 9988 7618 10024
rect 7562 9968 7564 9988
rect 7564 9968 7616 9988
rect 7616 9968 7618 9988
rect 7930 8064 7986 8120
rect 7562 7792 7618 7848
rect 7194 5888 7250 5944
rect 6918 4428 6920 4448
rect 6920 4428 6972 4448
rect 6972 4428 6974 4448
rect 6918 4392 6974 4428
rect 7562 5788 7564 5808
rect 7564 5788 7616 5808
rect 7616 5788 7618 5808
rect 7562 5752 7618 5788
rect 7470 4800 7526 4856
rect 7654 5208 7710 5264
rect 7378 4664 7434 4720
rect 7378 3032 7434 3088
rect 6458 2488 6514 2544
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10690 17584 10746 17640
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 9954 14320 10010 14376
rect 9586 13368 9642 13424
rect 9586 13096 9642 13152
rect 8850 12280 8906 12336
rect 8390 9016 8446 9072
rect 8666 7520 8722 7576
rect 8390 6976 8446 7032
rect 8206 3984 8262 4040
rect 8574 5072 8630 5128
rect 8758 4120 8814 4176
rect 9034 11092 9036 11112
rect 9036 11092 9088 11112
rect 9088 11092 9090 11112
rect 9034 11056 9090 11092
rect 9402 10648 9458 10704
rect 9402 10104 9458 10160
rect 9678 10376 9734 10432
rect 9678 10140 9680 10160
rect 9680 10140 9732 10160
rect 9732 10140 9734 10160
rect 9678 10104 9734 10140
rect 9862 10104 9918 10160
rect 9770 9288 9826 9344
rect 9678 9152 9734 9208
rect 9862 8064 9918 8120
rect 9770 7812 9826 7848
rect 9770 7792 9772 7812
rect 9772 7792 9824 7812
rect 9824 7792 9826 7812
rect 9034 4972 9036 4992
rect 9036 4972 9088 4992
rect 9088 4972 9090 4992
rect 9034 4936 9090 4972
rect 9678 6432 9734 6488
rect 9678 6296 9734 6352
rect 9310 5072 9366 5128
rect 8482 2896 8538 2952
rect 9126 3440 9182 3496
rect 9310 3712 9366 3768
rect 9862 4664 9918 4720
rect 9678 3984 9734 4040
rect 9678 3304 9734 3360
rect 9678 3168 9734 3224
rect 9862 3848 9918 3904
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10046 10240 10102 10296
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10046 8200 10102 8256
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 10782 13232 10838 13288
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10046 6568 10102 6624
rect 10046 6160 10102 6216
rect 10138 6024 10194 6080
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 11702 19760 11758 19816
rect 11242 12960 11298 13016
rect 11426 9560 11482 9616
rect 11150 9016 11206 9072
rect 11242 7656 11298 7712
rect 10874 6840 10930 6896
rect 11058 6740 11060 6760
rect 11060 6740 11112 6760
rect 11112 6740 11114 6760
rect 11058 6704 11114 6740
rect 11334 7248 11390 7304
rect 10966 5344 11022 5400
rect 11242 5616 11298 5672
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10874 4156 10876 4176
rect 10876 4156 10928 4176
rect 10928 4156 10930 4176
rect 10874 4120 10930 4156
rect 10046 2524 10048 2544
rect 10048 2524 10100 2544
rect 10100 2524 10102 2544
rect 10046 2488 10102 2524
rect 11794 13776 11850 13832
rect 11334 4004 11390 4040
rect 11334 3984 11336 4004
rect 11336 3984 11388 4004
rect 11388 3984 11390 4004
rect 11150 3032 11206 3088
rect 11058 2624 11114 2680
rect 11702 4276 11758 4312
rect 11702 4256 11704 4276
rect 11704 4256 11756 4276
rect 11756 4256 11758 4276
rect 12622 11736 12678 11792
rect 11794 3476 11796 3496
rect 11796 3476 11848 3496
rect 11848 3476 11850 3496
rect 11794 3440 11850 3476
rect 11426 1944 11482 2000
rect 11426 1808 11482 1864
rect 10966 1672 11022 1728
rect 12070 4528 12126 4584
rect 12346 10784 12402 10840
rect 12530 9560 12586 9616
rect 12622 7928 12678 7984
rect 12438 7520 12494 7576
rect 12990 10104 13046 10160
rect 12990 8336 13046 8392
rect 12898 7692 12900 7712
rect 12900 7692 12952 7712
rect 12952 7692 12954 7712
rect 12898 7656 12954 7692
rect 13174 6860 13230 6896
rect 13174 6840 13176 6860
rect 13176 6840 13228 6860
rect 13228 6840 13230 6860
rect 12806 6024 12862 6080
rect 12990 5344 13046 5400
rect 12990 4528 13046 4584
rect 13818 15952 13874 16008
rect 13542 7148 13544 7168
rect 13544 7148 13596 7168
rect 13596 7148 13598 7168
rect 13542 7112 13598 7148
rect 13358 5752 13414 5808
rect 13266 4936 13322 4992
rect 13450 3848 13506 3904
rect 12622 3440 12678 3496
rect 13082 1944 13138 2000
rect 12806 1536 12862 1592
rect 13910 10512 13966 10568
rect 13726 5208 13782 5264
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 15382 20848 15438 20904
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 14278 6604 14280 6624
rect 14280 6604 14332 6624
rect 14332 6604 14334 6624
rect 14278 6568 14334 6604
rect 14186 3712 14242 3768
rect 14002 2488 14058 2544
rect 15474 12824 15530 12880
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14646 6160 14702 6216
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 15382 7928 15438 7984
rect 15566 10920 15622 10976
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14646 4564 14648 4584
rect 14648 4564 14700 4584
rect 14700 4564 14702 4584
rect 14646 4528 14702 4564
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 15566 5752 15622 5808
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 24122 20984 24178 21040
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 19522 13368 19578 13424
rect 16210 10684 16212 10704
rect 16212 10684 16264 10704
rect 16264 10684 16266 10704
rect 16210 10648 16266 10684
rect 16670 11600 16726 11656
rect 16210 6976 16266 7032
rect 14738 3612 14740 3632
rect 14740 3612 14792 3632
rect 14792 3612 14794 3632
rect 14738 3576 14794 3612
rect 17590 5652 17592 5672
rect 17592 5652 17644 5672
rect 17644 5652 17646 5672
rect 17590 5616 17646 5652
rect 17682 5480 17738 5536
rect 16946 5344 17002 5400
rect 17590 5108 17592 5128
rect 17592 5108 17644 5128
rect 17644 5108 17646 5128
rect 17590 5072 17646 5108
rect 17222 4972 17224 4992
rect 17224 4972 17276 4992
rect 17276 4972 17278 4992
rect 17222 4936 17278 4972
rect 16394 4800 16450 4856
rect 15382 3440 15438 3496
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 14646 3168 14702 3224
rect 14738 3052 14794 3088
rect 15658 3304 15714 3360
rect 14738 3032 14740 3052
rect 14740 3032 14792 3052
rect 14792 3032 14794 3052
rect 15566 3032 15622 3088
rect 14830 2932 14832 2952
rect 14832 2932 14884 2952
rect 14884 2932 14886 2952
rect 14830 2896 14886 2932
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 14646 1400 14702 1456
rect 15474 1400 15530 1456
rect 16302 3848 16358 3904
rect 15750 2080 15806 2136
rect 16486 4392 16542 4448
rect 17130 4020 17132 4040
rect 17132 4020 17184 4040
rect 17184 4020 17186 4040
rect 17130 3984 17186 4020
rect 17590 3168 17646 3224
rect 16762 2624 16818 2680
rect 17038 2524 17040 2544
rect 17040 2524 17092 2544
rect 17092 2524 17094 2544
rect 17038 2488 17094 2524
rect 16670 2100 16726 2136
rect 16670 2080 16672 2100
rect 16672 2080 16724 2100
rect 16724 2080 16726 2100
rect 16854 2080 16910 2136
rect 16854 1536 16910 1592
rect 17038 1536 17094 1592
rect 18050 9560 18106 9616
rect 17958 8336 18014 8392
rect 17774 4528 17830 4584
rect 18326 7948 18382 7984
rect 18326 7928 18328 7948
rect 18328 7928 18380 7948
rect 18380 7928 18382 7948
rect 18050 7520 18106 7576
rect 18878 6976 18934 7032
rect 18786 5652 18788 5672
rect 18788 5652 18840 5672
rect 18840 5652 18842 5672
rect 18786 5616 18842 5652
rect 18234 4800 18290 4856
rect 18234 4700 18236 4720
rect 18236 4700 18288 4720
rect 18288 4700 18290 4720
rect 18234 4664 18290 4700
rect 18142 2896 18198 2952
rect 18510 4256 18566 4312
rect 18510 3712 18566 3768
rect 19430 7248 19486 7304
rect 19430 6024 19486 6080
rect 19154 3984 19210 4040
rect 18418 3596 18474 3632
rect 18418 3576 18420 3596
rect 18420 3576 18472 3596
rect 18472 3576 18474 3596
rect 18602 3576 18658 3632
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 20810 11192 20866 11248
rect 19982 10920 20038 10976
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19798 5480 19854 5536
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19430 3732 19486 3768
rect 20442 8472 20498 8528
rect 20258 5344 20314 5400
rect 19430 3712 19432 3732
rect 19432 3712 19484 3732
rect 19484 3712 19486 3732
rect 19338 3304 19394 3360
rect 19430 2796 19432 2816
rect 19432 2796 19484 2816
rect 19484 2796 19486 2816
rect 19430 2760 19486 2796
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 20350 3984 20406 4040
rect 20258 3440 20314 3496
rect 19614 1808 19670 1864
rect 19430 1400 19486 1456
rect 20166 1264 20222 1320
rect 20534 7384 20590 7440
rect 20626 3848 20682 3904
rect 20534 2388 20536 2408
rect 20536 2388 20588 2408
rect 20588 2388 20590 2408
rect 20534 2352 20590 2388
rect 20902 9968 20958 10024
rect 21362 7792 21418 7848
rect 21362 5616 21418 5672
rect 20810 3168 20866 3224
rect 20994 3576 21050 3632
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 24122 7520 24178 7576
rect 24766 6976 24822 7032
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 25502 6332 25504 6352
rect 25504 6332 25556 6352
rect 25556 6332 25558 6352
rect 25502 6296 25558 6332
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 22466 5208 22522 5264
rect 21730 4120 21786 4176
rect 23478 4392 23534 4448
rect 22742 4256 22798 4312
rect 21638 3984 21694 4040
rect 21546 3848 21602 3904
rect 21086 2760 21142 2816
rect 21178 1944 21234 2000
rect 22006 3576 22062 3632
rect 21822 3032 21878 3088
rect 22006 2896 22062 2952
rect 22650 2760 22706 2816
rect 22282 2508 22338 2544
rect 22282 2488 22284 2508
rect 22284 2488 22336 2508
rect 22336 2488 22338 2508
rect 22466 1536 22522 1592
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 23662 4020 23664 4040
rect 23664 4020 23716 4040
rect 23716 4020 23718 4040
rect 23662 3984 23718 4020
rect 24030 2080 24086 2136
rect 25134 3596 25190 3632
rect 25134 3576 25136 3596
rect 25136 3576 25188 3596
rect 25188 3576 25190 3596
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 25134 2796 25136 2816
rect 25136 2796 25188 2816
rect 25188 2796 25190 2816
rect 25134 2760 25190 2796
rect 27066 2760 27122 2816
rect 27618 1672 27674 1728
rect 3146 312 3202 368
<< metal3 >>
rect 0 27570 480 27600
rect 3141 27570 3207 27573
rect 0 27568 3207 27570
rect 0 27512 3146 27568
rect 3202 27512 3207 27568
rect 0 27510 3207 27512
rect 0 27480 480 27510
rect 3141 27507 3207 27510
rect 0 26890 480 26920
rect 2957 26890 3023 26893
rect 0 26888 3023 26890
rect 0 26832 2962 26888
rect 3018 26832 3023 26888
rect 0 26830 3023 26832
rect 0 26800 480 26830
rect 2957 26827 3023 26830
rect 0 26210 480 26240
rect 3509 26210 3575 26213
rect 0 26208 3575 26210
rect 0 26152 3514 26208
rect 3570 26152 3575 26208
rect 0 26150 3575 26152
rect 0 26120 480 26150
rect 3509 26147 3575 26150
rect 10277 25600 10597 25601
rect 0 25530 480 25560
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 3417 25530 3483 25533
rect 0 25528 3483 25530
rect 0 25472 3422 25528
rect 3478 25472 3483 25528
rect 0 25470 3483 25472
rect 0 25440 480 25470
rect 3417 25467 3483 25470
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 0 24850 480 24880
rect 565 24850 631 24853
rect 0 24848 631 24850
rect 0 24792 570 24848
rect 626 24792 631 24848
rect 0 24790 631 24792
rect 0 24760 480 24790
rect 565 24787 631 24790
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 0 24170 480 24200
rect 3417 24170 3483 24173
rect 0 24168 3483 24170
rect 0 24112 3422 24168
rect 3478 24112 3483 24168
rect 0 24110 3483 24112
rect 0 24080 480 24110
rect 3417 24107 3483 24110
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 565 23762 631 23765
rect 10961 23762 11027 23765
rect 565 23760 11027 23762
rect 565 23704 570 23760
rect 626 23704 10966 23760
rect 11022 23704 11027 23760
rect 565 23702 11027 23704
rect 565 23699 631 23702
rect 10961 23699 11027 23702
rect 0 23490 480 23520
rect 3233 23490 3299 23493
rect 0 23488 3299 23490
rect 0 23432 3238 23488
rect 3294 23432 3299 23488
rect 0 23430 3299 23432
rect 0 23400 480 23430
rect 3233 23427 3299 23430
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 5610 22880 5930 22881
rect 0 22810 480 22840
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 0 22750 5458 22810
rect 0 22720 480 22750
rect 5398 22674 5458 22750
rect 5993 22674 6059 22677
rect 5398 22672 6059 22674
rect 5398 22616 5998 22672
rect 6054 22616 6059 22672
rect 5398 22614 6059 22616
rect 5993 22611 6059 22614
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 3417 22266 3483 22269
rect 8753 22266 8819 22269
rect 3417 22264 8819 22266
rect 3417 22208 3422 22264
rect 3478 22208 8758 22264
rect 8814 22208 8819 22264
rect 3417 22206 8819 22208
rect 3417 22203 3483 22206
rect 8753 22203 8819 22206
rect 0 22130 480 22160
rect 3417 22130 3483 22133
rect 0 22128 3483 22130
rect 0 22072 3422 22128
rect 3478 22072 3483 22128
rect 0 22070 3483 22072
rect 0 22040 480 22070
rect 3417 22067 3483 22070
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 21727 24597 21728
rect 0 21450 480 21480
rect 0 21390 674 21450
rect 0 21360 480 21390
rect 614 20906 674 21390
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 21183 19930 21184
rect 24117 21042 24183 21045
rect 27520 21042 28000 21072
rect 24117 21040 28000 21042
rect 24117 20984 24122 21040
rect 24178 20984 28000 21040
rect 24117 20982 28000 20984
rect 24117 20979 24183 20982
rect 27520 20952 28000 20982
rect 15377 20906 15443 20909
rect 614 20904 15443 20906
rect 614 20848 15382 20904
rect 15438 20848 15443 20904
rect 614 20846 15443 20848
rect 15377 20843 15443 20846
rect 0 20770 480 20800
rect 4061 20770 4127 20773
rect 0 20768 4127 20770
rect 0 20712 4066 20768
rect 4122 20712 4127 20768
rect 0 20710 4127 20712
rect 0 20680 480 20710
rect 4061 20707 4127 20710
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 20639 24597 20640
rect 10277 20160 10597 20161
rect 0 20090 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 0 20030 674 20090
rect 0 20000 480 20030
rect 614 19818 674 20030
rect 11697 19818 11763 19821
rect 614 19816 11763 19818
rect 614 19760 11702 19816
rect 11758 19760 11763 19816
rect 614 19758 11763 19760
rect 11697 19755 11763 19758
rect 5610 19616 5930 19617
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 0 19410 480 19440
rect 3785 19410 3851 19413
rect 0 19408 3851 19410
rect 0 19352 3790 19408
rect 3846 19352 3851 19408
rect 0 19350 3851 19352
rect 0 19320 480 19350
rect 3785 19347 3851 19350
rect 10277 19072 10597 19073
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 0 18730 480 18760
rect 3969 18730 4035 18733
rect 0 18728 4035 18730
rect 0 18672 3974 18728
rect 4030 18672 4035 18728
rect 0 18670 4035 18672
rect 0 18640 480 18670
rect 3969 18667 4035 18670
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 0 18050 480 18080
rect 3877 18050 3943 18053
rect 0 18048 3943 18050
rect 0 17992 3882 18048
rect 3938 17992 3943 18048
rect 0 17990 3943 17992
rect 0 17960 480 17990
rect 3877 17987 3943 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 3417 17642 3483 17645
rect 10685 17642 10751 17645
rect 3417 17640 10751 17642
rect 3417 17584 3422 17640
rect 3478 17584 10690 17640
rect 10746 17584 10751 17640
rect 3417 17582 10751 17584
rect 3417 17579 3483 17582
rect 10685 17579 10751 17582
rect 5610 17440 5930 17441
rect 0 17370 480 17400
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 3693 17370 3759 17373
rect 0 17368 3759 17370
rect 0 17312 3698 17368
rect 3754 17312 3759 17368
rect 0 17310 3759 17312
rect 0 17280 480 17310
rect 3693 17307 3759 17310
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 0 16690 480 16720
rect 1485 16690 1551 16693
rect 0 16688 1551 16690
rect 0 16632 1490 16688
rect 1546 16632 1551 16688
rect 0 16630 1551 16632
rect 0 16600 480 16630
rect 1485 16627 1551 16630
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 0 16010 480 16040
rect 3233 16010 3299 16013
rect 0 16008 3299 16010
rect 0 15952 3238 16008
rect 3294 15952 3299 16008
rect 0 15950 3299 15952
rect 0 15920 480 15950
rect 3233 15947 3299 15950
rect 4061 16010 4127 16013
rect 13813 16010 13879 16013
rect 4061 16008 13879 16010
rect 4061 15952 4066 16008
rect 4122 15952 13818 16008
rect 13874 15952 13879 16008
rect 4061 15950 13879 15952
rect 4061 15947 4127 15950
rect 13813 15947 13879 15950
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 0 15330 480 15360
rect 1761 15330 1827 15333
rect 0 15328 1827 15330
rect 0 15272 1766 15328
rect 1822 15272 1827 15328
rect 0 15270 1827 15272
rect 0 15240 480 15270
rect 1761 15267 1827 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 10277 14720 10597 14721
rect 0 14650 480 14680
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 3325 14650 3391 14653
rect 0 14648 3391 14650
rect 0 14592 3330 14648
rect 3386 14592 3391 14648
rect 0 14590 3391 14592
rect 0 14560 480 14590
rect 3325 14587 3391 14590
rect 2037 14378 2103 14381
rect 9949 14378 10015 14381
rect 2037 14376 10015 14378
rect 2037 14320 2042 14376
rect 2098 14320 9954 14376
rect 10010 14320 10015 14376
rect 2037 14318 10015 14320
rect 2037 14315 2103 14318
rect 9949 14315 10015 14318
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 0 13970 480 14000
rect 0 13910 1410 13970
rect 0 13880 480 13910
rect 1350 13834 1410 13910
rect 11789 13834 11855 13837
rect 1350 13832 11855 13834
rect 1350 13776 11794 13832
rect 11850 13776 11855 13832
rect 1350 13774 11855 13776
rect 11789 13771 11855 13774
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 3969 13562 4035 13565
rect 7833 13562 7899 13565
rect 3969 13560 7899 13562
rect 3969 13504 3974 13560
rect 4030 13504 7838 13560
rect 7894 13504 7899 13560
rect 3969 13502 7899 13504
rect 3969 13499 4035 13502
rect 7833 13499 7899 13502
rect 9581 13426 9647 13429
rect 19517 13426 19583 13429
rect 4846 13424 9647 13426
rect 4846 13368 9586 13424
rect 9642 13368 9647 13424
rect 4846 13366 9647 13368
rect 0 13290 480 13320
rect 4846 13290 4906 13366
rect 9581 13363 9647 13366
rect 12022 13424 19583 13426
rect 12022 13368 19522 13424
rect 19578 13368 19583 13424
rect 12022 13366 19583 13368
rect 0 13230 4906 13290
rect 4981 13290 5047 13293
rect 10777 13290 10843 13293
rect 4981 13288 10843 13290
rect 4981 13232 4986 13288
rect 5042 13232 10782 13288
rect 10838 13232 10843 13288
rect 4981 13230 10843 13232
rect 0 13200 480 13230
rect 4981 13227 5047 13230
rect 10777 13227 10843 13230
rect 9581 13154 9647 13157
rect 12022 13154 12082 13366
rect 19517 13363 19583 13366
rect 9581 13152 12082 13154
rect 9581 13096 9586 13152
rect 9642 13096 12082 13152
rect 9581 13094 12082 13096
rect 9581 13091 9647 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 13023 24597 13024
rect 6085 13018 6151 13021
rect 11237 13018 11303 13021
rect 6085 13016 11303 13018
rect 6085 12960 6090 13016
rect 6146 12960 11242 13016
rect 11298 12960 11303 13016
rect 6085 12958 11303 12960
rect 6085 12955 6151 12958
rect 11237 12955 11303 12958
rect 3969 12882 4035 12885
rect 15469 12882 15535 12885
rect 3969 12880 15535 12882
rect 3969 12824 3974 12880
rect 4030 12824 15474 12880
rect 15530 12824 15535 12880
rect 3969 12822 15535 12824
rect 3969 12819 4035 12822
rect 15469 12819 15535 12822
rect 0 12610 480 12640
rect 3969 12610 4035 12613
rect 0 12608 4035 12610
rect 0 12552 3974 12608
rect 4030 12552 4035 12608
rect 0 12550 4035 12552
rect 0 12520 480 12550
rect 3969 12547 4035 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 4705 12474 4771 12477
rect 5901 12474 5967 12477
rect 4705 12472 5967 12474
rect 4705 12416 4710 12472
rect 4766 12416 5906 12472
rect 5962 12416 5967 12472
rect 4705 12414 5967 12416
rect 4705 12411 4771 12414
rect 5901 12411 5967 12414
rect 2589 12338 2655 12341
rect 8845 12338 8911 12341
rect 2589 12336 8911 12338
rect 2589 12280 2594 12336
rect 2650 12280 8850 12336
rect 8906 12280 8911 12336
rect 2589 12278 8911 12280
rect 2589 12275 2655 12278
rect 8845 12275 8911 12278
rect 2313 12202 2379 12205
rect 4153 12202 4219 12205
rect 2313 12200 4219 12202
rect 2313 12144 2318 12200
rect 2374 12144 4158 12200
rect 4214 12144 4219 12200
rect 2313 12142 4219 12144
rect 2313 12139 2379 12142
rect 4153 12139 4219 12142
rect 5610 12000 5930 12001
rect 0 11930 480 11960
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 0 11896 2698 11930
rect 0 11870 2882 11896
rect 0 11840 480 11870
rect 2638 11836 2882 11870
rect 2822 11794 2882 11836
rect 12617 11794 12683 11797
rect 2822 11792 12683 11794
rect 2822 11736 12622 11792
rect 12678 11736 12683 11792
rect 2822 11734 12683 11736
rect 12617 11731 12683 11734
rect 8109 11658 8175 11661
rect 16665 11658 16731 11661
rect 8109 11656 16731 11658
rect 8109 11600 8114 11656
rect 8170 11600 16670 11656
rect 16726 11600 16731 11656
rect 8109 11598 16731 11600
rect 8109 11595 8175 11598
rect 16665 11595 16731 11598
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 3509 11386 3575 11389
rect 6269 11386 6335 11389
rect 3509 11384 6335 11386
rect 3509 11328 3514 11384
rect 3570 11328 6274 11384
rect 6330 11328 6335 11384
rect 3509 11326 6335 11328
rect 3509 11323 3575 11326
rect 6269 11323 6335 11326
rect 0 11250 480 11280
rect 20805 11250 20871 11253
rect 0 11248 20871 11250
rect 0 11192 20810 11248
rect 20866 11192 20871 11248
rect 0 11190 20871 11192
rect 0 11160 480 11190
rect 20805 11187 20871 11190
rect 4981 11114 5047 11117
rect 7373 11114 7439 11117
rect 9029 11114 9095 11117
rect 4981 11112 9095 11114
rect 4981 11056 4986 11112
rect 5042 11056 7378 11112
rect 7434 11056 9034 11112
rect 9090 11056 9095 11112
rect 4981 11054 9095 11056
rect 4981 11051 5047 11054
rect 7373 11051 7439 11054
rect 9029 11051 9095 11054
rect 15561 10978 15627 10981
rect 19977 10978 20043 10981
rect 15561 10976 20043 10978
rect 15561 10920 15566 10976
rect 15622 10920 19982 10976
rect 20038 10920 20043 10976
rect 15561 10918 20043 10920
rect 15561 10915 15627 10918
rect 19977 10915 20043 10918
rect 5610 10912 5930 10913
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 12341 10842 12407 10845
rect 6088 10840 12407 10842
rect 6088 10784 12346 10840
rect 12402 10784 12407 10840
rect 6088 10782 12407 10784
rect 0 10570 480 10600
rect 6088 10570 6148 10782
rect 12341 10779 12407 10782
rect 9397 10706 9463 10709
rect 16205 10706 16271 10709
rect 9397 10704 16271 10706
rect 9397 10648 9402 10704
rect 9458 10648 16210 10704
rect 16266 10648 16271 10704
rect 9397 10646 16271 10648
rect 9397 10643 9463 10646
rect 16205 10643 16271 10646
rect 0 10510 6148 10570
rect 6361 10570 6427 10573
rect 13905 10570 13971 10573
rect 6361 10568 13971 10570
rect 6361 10512 6366 10568
rect 6422 10512 13910 10568
rect 13966 10512 13971 10568
rect 6361 10510 13971 10512
rect 0 10480 480 10510
rect 6361 10507 6427 10510
rect 13905 10507 13971 10510
rect 8109 10434 8175 10437
rect 9673 10434 9739 10437
rect 8109 10432 9739 10434
rect 8109 10376 8114 10432
rect 8170 10376 9678 10432
rect 9734 10376 9739 10432
rect 8109 10374 9739 10376
rect 8109 10371 8175 10374
rect 9673 10371 9739 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 4337 10298 4403 10301
rect 7373 10298 7439 10301
rect 4337 10296 7439 10298
rect 4337 10240 4342 10296
rect 4398 10240 7378 10296
rect 7434 10240 7439 10296
rect 4337 10238 7439 10240
rect 4337 10235 4403 10238
rect 7373 10235 7439 10238
rect 8017 10298 8083 10301
rect 10041 10298 10107 10301
rect 8017 10296 10107 10298
rect 8017 10240 8022 10296
rect 8078 10240 10046 10296
rect 10102 10240 10107 10296
rect 8017 10238 10107 10240
rect 8017 10235 8083 10238
rect 10041 10235 10107 10238
rect 3785 10162 3851 10165
rect 9397 10162 9463 10165
rect 9673 10162 9739 10165
rect 3785 10160 9739 10162
rect 3785 10104 3790 10160
rect 3846 10104 9402 10160
rect 9458 10104 9678 10160
rect 9734 10104 9739 10160
rect 3785 10102 9739 10104
rect 3785 10099 3851 10102
rect 9397 10099 9463 10102
rect 9673 10099 9739 10102
rect 9857 10162 9923 10165
rect 12985 10162 13051 10165
rect 9857 10160 13051 10162
rect 9857 10104 9862 10160
rect 9918 10104 12990 10160
rect 13046 10104 13051 10160
rect 9857 10102 13051 10104
rect 9857 10099 9923 10102
rect 12985 10099 13051 10102
rect 7557 10026 7623 10029
rect 20897 10026 20963 10029
rect 7557 10024 20963 10026
rect 7557 9968 7562 10024
rect 7618 9968 20902 10024
rect 20958 9968 20963 10024
rect 7557 9966 20963 9968
rect 7557 9963 7623 9966
rect 20897 9963 20963 9966
rect 0 9890 480 9920
rect 565 9890 631 9893
rect 0 9888 631 9890
rect 0 9832 570 9888
rect 626 9832 631 9888
rect 0 9830 631 9832
rect 0 9800 480 9830
rect 565 9827 631 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 1761 9754 1827 9757
rect 5441 9754 5507 9757
rect 1761 9752 5507 9754
rect 1761 9696 1766 9752
rect 1822 9696 5446 9752
rect 5502 9696 5507 9752
rect 1761 9694 5507 9696
rect 1761 9691 1827 9694
rect 5441 9691 5507 9694
rect 2589 9618 2655 9621
rect 11421 9618 11487 9621
rect 2589 9616 11487 9618
rect 2589 9560 2594 9616
rect 2650 9560 11426 9616
rect 11482 9560 11487 9616
rect 2589 9558 11487 9560
rect 2589 9555 2655 9558
rect 11421 9555 11487 9558
rect 12525 9618 12591 9621
rect 18045 9618 18111 9621
rect 12525 9616 18111 9618
rect 12525 9560 12530 9616
rect 12586 9560 18050 9616
rect 18106 9560 18111 9616
rect 12525 9558 18111 9560
rect 12525 9555 12591 9558
rect 18045 9555 18111 9558
rect 4429 9482 4495 9485
rect 14590 9482 14596 9484
rect 4429 9480 14596 9482
rect 4429 9424 4434 9480
rect 4490 9424 14596 9480
rect 4429 9422 14596 9424
rect 4429 9419 4495 9422
rect 14590 9420 14596 9422
rect 14660 9420 14666 9484
rect 5165 9346 5231 9349
rect 9765 9346 9831 9349
rect 5165 9344 9831 9346
rect 5165 9288 5170 9344
rect 5226 9288 9770 9344
rect 9826 9288 9831 9344
rect 5165 9286 9831 9288
rect 5165 9283 5231 9286
rect 9765 9283 9831 9286
rect 10277 9280 10597 9281
rect 0 9210 480 9240
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 3969 9210 4035 9213
rect 0 9208 4035 9210
rect 0 9152 3974 9208
rect 4030 9152 4035 9208
rect 0 9150 4035 9152
rect 0 9120 480 9150
rect 3969 9147 4035 9150
rect 5533 9210 5599 9213
rect 6177 9210 6243 9213
rect 9673 9210 9739 9213
rect 5533 9208 9739 9210
rect 5533 9152 5538 9208
rect 5594 9152 6182 9208
rect 6238 9152 9678 9208
rect 9734 9152 9739 9208
rect 5533 9150 9739 9152
rect 5533 9147 5599 9150
rect 6177 9147 6243 9150
rect 9673 9147 9739 9150
rect 8385 9074 8451 9077
rect 11145 9074 11211 9077
rect 8385 9072 11211 9074
rect 8385 9016 8390 9072
rect 8446 9016 11150 9072
rect 11206 9016 11211 9072
rect 8385 9014 11211 9016
rect 8385 9011 8451 9014
rect 11145 9011 11211 9014
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 0 8530 480 8560
rect 3969 8530 4035 8533
rect 20437 8530 20503 8533
rect 0 8470 2698 8530
rect 0 8440 480 8470
rect 2638 8122 2698 8470
rect 3969 8528 20503 8530
rect 3969 8472 3974 8528
rect 4030 8472 20442 8528
rect 20498 8472 20503 8528
rect 3969 8470 20503 8472
rect 3969 8467 4035 8470
rect 20437 8467 20503 8470
rect 12985 8394 13051 8397
rect 17953 8394 18019 8397
rect 12985 8392 18019 8394
rect 12985 8336 12990 8392
rect 13046 8336 17958 8392
rect 18014 8336 18019 8392
rect 12985 8334 18019 8336
rect 12985 8331 13051 8334
rect 17953 8331 18019 8334
rect 2865 8258 2931 8261
rect 4521 8258 4587 8261
rect 10041 8258 10107 8261
rect 2865 8256 10107 8258
rect 2865 8200 2870 8256
rect 2926 8200 4526 8256
rect 4582 8200 10046 8256
rect 10102 8200 10107 8256
rect 2865 8198 10107 8200
rect 2865 8195 2931 8198
rect 4521 8195 4587 8198
rect 10041 8195 10107 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 7925 8122 7991 8125
rect 9857 8122 9923 8125
rect 2638 8062 2928 8122
rect 2868 7986 2928 8062
rect 7925 8120 9923 8122
rect 7925 8064 7930 8120
rect 7986 8064 9862 8120
rect 9918 8064 9923 8120
rect 7925 8062 9923 8064
rect 7925 8059 7991 8062
rect 9857 8059 9923 8062
rect 12617 7986 12683 7989
rect 2868 7984 12683 7986
rect 2868 7928 12622 7984
rect 12678 7928 12683 7984
rect 2868 7926 12683 7928
rect 12617 7923 12683 7926
rect 15377 7986 15443 7989
rect 18321 7986 18387 7989
rect 15377 7984 18387 7986
rect 15377 7928 15382 7984
rect 15438 7928 18326 7984
rect 18382 7928 18387 7984
rect 15377 7926 18387 7928
rect 15377 7923 15443 7926
rect 18321 7923 18387 7926
rect 0 7850 480 7880
rect 2589 7850 2655 7853
rect 0 7848 2655 7850
rect 0 7792 2594 7848
rect 2650 7792 2655 7848
rect 0 7790 2655 7792
rect 0 7760 480 7790
rect 2589 7787 2655 7790
rect 4521 7850 4587 7853
rect 7557 7850 7623 7853
rect 4521 7848 7623 7850
rect 4521 7792 4526 7848
rect 4582 7792 7562 7848
rect 7618 7792 7623 7848
rect 4521 7790 7623 7792
rect 4521 7787 4587 7790
rect 7557 7787 7623 7790
rect 9765 7850 9831 7853
rect 21357 7850 21423 7853
rect 9765 7848 21423 7850
rect 9765 7792 9770 7848
rect 9826 7792 21362 7848
rect 21418 7792 21423 7848
rect 9765 7790 21423 7792
rect 9765 7787 9831 7790
rect 21357 7787 21423 7790
rect 6637 7714 6703 7717
rect 11237 7714 11303 7717
rect 12893 7714 12959 7717
rect 6637 7712 12959 7714
rect 6637 7656 6642 7712
rect 6698 7656 11242 7712
rect 11298 7656 12898 7712
rect 12954 7656 12959 7712
rect 6637 7654 12959 7656
rect 6637 7651 6703 7654
rect 11237 7651 11303 7654
rect 12893 7651 12959 7654
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 1669 7578 1735 7581
rect 5349 7578 5415 7581
rect 1669 7576 5415 7578
rect 1669 7520 1674 7576
rect 1730 7520 5354 7576
rect 5410 7520 5415 7576
rect 1669 7518 5415 7520
rect 1669 7515 1735 7518
rect 5349 7515 5415 7518
rect 8661 7578 8727 7581
rect 12433 7578 12499 7581
rect 8661 7576 12499 7578
rect 8661 7520 8666 7576
rect 8722 7520 12438 7576
rect 12494 7520 12499 7576
rect 8661 7518 12499 7520
rect 8661 7515 8727 7518
rect 12433 7515 12499 7518
rect 18045 7578 18111 7581
rect 24117 7578 24183 7581
rect 18045 7576 24183 7578
rect 18045 7520 18050 7576
rect 18106 7520 24122 7576
rect 24178 7520 24183 7576
rect 18045 7518 24183 7520
rect 18045 7515 18111 7518
rect 24117 7515 24183 7518
rect 5257 7442 5323 7445
rect 20529 7442 20595 7445
rect 5257 7440 20595 7442
rect 5257 7384 5262 7440
rect 5318 7384 20534 7440
rect 20590 7384 20595 7440
rect 5257 7382 20595 7384
rect 5257 7379 5323 7382
rect 20529 7379 20595 7382
rect 841 7306 907 7309
rect 4521 7306 4587 7309
rect 11329 7306 11395 7309
rect 19425 7306 19491 7309
rect 841 7304 4587 7306
rect 841 7248 846 7304
rect 902 7248 4526 7304
rect 4582 7248 4587 7304
rect 841 7246 4587 7248
rect 841 7243 907 7246
rect 4521 7243 4587 7246
rect 9446 7246 10794 7306
rect 0 7170 480 7200
rect 1577 7170 1643 7173
rect 0 7168 1643 7170
rect 0 7112 1582 7168
rect 1638 7112 1643 7168
rect 0 7110 1643 7112
rect 0 7080 480 7110
rect 1577 7107 1643 7110
rect 5349 7170 5415 7173
rect 9446 7170 9506 7246
rect 5349 7168 9506 7170
rect 5349 7112 5354 7168
rect 5410 7112 9506 7168
rect 5349 7110 9506 7112
rect 10734 7170 10794 7246
rect 11329 7304 19491 7306
rect 11329 7248 11334 7304
rect 11390 7248 19430 7304
rect 19486 7248 19491 7304
rect 11329 7246 19491 7248
rect 11329 7243 11395 7246
rect 19425 7243 19491 7246
rect 13537 7170 13603 7173
rect 10734 7168 13603 7170
rect 10734 7112 13542 7168
rect 13598 7112 13603 7168
rect 10734 7110 13603 7112
rect 5349 7107 5415 7110
rect 13537 7107 13603 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 2129 7034 2195 7037
rect 8385 7034 8451 7037
rect 2129 7032 8451 7034
rect 2129 6976 2134 7032
rect 2190 6976 8390 7032
rect 8446 6976 8451 7032
rect 2129 6974 8451 6976
rect 2129 6971 2195 6974
rect 8385 6971 8451 6974
rect 16205 7034 16271 7037
rect 18873 7034 18939 7037
rect 16205 7032 18939 7034
rect 16205 6976 16210 7032
rect 16266 6976 18878 7032
rect 18934 6976 18939 7032
rect 16205 6974 18939 6976
rect 16205 6971 16271 6974
rect 18873 6971 18939 6974
rect 24761 7034 24827 7037
rect 27520 7034 28000 7064
rect 24761 7032 28000 7034
rect 24761 6976 24766 7032
rect 24822 6976 28000 7032
rect 24761 6974 28000 6976
rect 24761 6971 24827 6974
rect 27520 6944 28000 6974
rect 1393 6898 1459 6901
rect 5165 6898 5231 6901
rect 1393 6896 5231 6898
rect 1393 6840 1398 6896
rect 1454 6840 5170 6896
rect 5226 6840 5231 6896
rect 1393 6838 5231 6840
rect 1393 6835 1459 6838
rect 5165 6835 5231 6838
rect 10869 6898 10935 6901
rect 13169 6898 13235 6901
rect 10869 6896 13235 6898
rect 10869 6840 10874 6896
rect 10930 6840 13174 6896
rect 13230 6840 13235 6896
rect 10869 6838 13235 6840
rect 10869 6835 10935 6838
rect 13169 6835 13235 6838
rect 5717 6762 5783 6765
rect 11053 6762 11119 6765
rect 5717 6760 11119 6762
rect 5717 6704 5722 6760
rect 5778 6704 11058 6760
rect 11114 6704 11119 6760
rect 5717 6702 11119 6704
rect 5717 6699 5783 6702
rect 11053 6699 11119 6702
rect 10041 6626 10107 6629
rect 14273 6626 14339 6629
rect 10041 6624 14339 6626
rect 10041 6568 10046 6624
rect 10102 6568 14278 6624
rect 14334 6568 14339 6624
rect 10041 6566 14339 6568
rect 10041 6563 10107 6566
rect 14273 6563 14339 6566
rect 5610 6560 5930 6561
rect 0 6490 480 6520
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 3969 6490 4035 6493
rect 0 6488 4035 6490
rect 0 6432 3974 6488
rect 4030 6432 4035 6488
rect 0 6430 4035 6432
rect 0 6400 480 6430
rect 3969 6427 4035 6430
rect 9673 6490 9739 6493
rect 9673 6488 14474 6490
rect 9673 6432 9678 6488
rect 9734 6432 14474 6488
rect 9673 6430 14474 6432
rect 9673 6427 9739 6430
rect 5349 6354 5415 6357
rect 9673 6354 9739 6357
rect 14414 6354 14474 6430
rect 25497 6354 25563 6357
rect 5349 6352 10242 6354
rect 5349 6296 5354 6352
rect 5410 6296 9678 6352
rect 9734 6296 10242 6352
rect 5349 6294 10242 6296
rect 14414 6352 25563 6354
rect 14414 6296 25502 6352
rect 25558 6296 25563 6352
rect 14414 6294 25563 6296
rect 5349 6291 5415 6294
rect 9673 6291 9739 6294
rect 2681 6218 2747 6221
rect 10041 6218 10107 6221
rect 2681 6216 10107 6218
rect 2681 6160 2686 6216
rect 2742 6160 10046 6216
rect 10102 6160 10107 6216
rect 2681 6158 10107 6160
rect 10182 6218 10242 6294
rect 25497 6291 25563 6294
rect 14641 6218 14707 6221
rect 10182 6216 14707 6218
rect 10182 6160 14646 6216
rect 14702 6160 14707 6216
rect 10182 6158 14707 6160
rect 2681 6155 2747 6158
rect 10041 6155 10107 6158
rect 14641 6155 14707 6158
rect 3141 6082 3207 6085
rect 10133 6082 10199 6085
rect 3141 6080 10199 6082
rect 3141 6024 3146 6080
rect 3202 6024 10138 6080
rect 10194 6024 10199 6080
rect 3141 6022 10199 6024
rect 3141 6019 3207 6022
rect 10133 6019 10199 6022
rect 12801 6082 12867 6085
rect 19425 6082 19491 6085
rect 12801 6080 19491 6082
rect 12801 6024 12806 6080
rect 12862 6024 19430 6080
rect 19486 6024 19491 6080
rect 12801 6022 19491 6024
rect 12801 6019 12867 6022
rect 19425 6019 19491 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 5951 19930 5952
rect 3601 5946 3667 5949
rect 7189 5946 7255 5949
rect 3601 5944 7255 5946
rect 3601 5888 3606 5944
rect 3662 5888 7194 5944
rect 7250 5888 7255 5944
rect 3601 5886 7255 5888
rect 3601 5883 3667 5886
rect 7189 5883 7255 5886
rect 0 5810 480 5840
rect 1853 5810 1919 5813
rect 0 5808 1919 5810
rect 0 5752 1858 5808
rect 1914 5752 1919 5808
rect 0 5750 1919 5752
rect 0 5720 480 5750
rect 1853 5747 1919 5750
rect 2957 5810 3023 5813
rect 7557 5810 7623 5813
rect 2957 5808 7623 5810
rect 2957 5752 2962 5808
rect 3018 5752 7562 5808
rect 7618 5752 7623 5808
rect 2957 5750 7623 5752
rect 2957 5747 3023 5750
rect 7557 5747 7623 5750
rect 13353 5810 13419 5813
rect 15561 5810 15627 5813
rect 13353 5808 15627 5810
rect 13353 5752 13358 5808
rect 13414 5752 15566 5808
rect 15622 5752 15627 5808
rect 13353 5750 15627 5752
rect 13353 5747 13419 5750
rect 15561 5747 15627 5750
rect 3049 5674 3115 5677
rect 11237 5674 11303 5677
rect 17585 5674 17651 5677
rect 3049 5672 17651 5674
rect 3049 5616 3054 5672
rect 3110 5616 11242 5672
rect 11298 5616 17590 5672
rect 17646 5616 17651 5672
rect 3049 5614 17651 5616
rect 3049 5611 3115 5614
rect 11237 5611 11303 5614
rect 17585 5611 17651 5614
rect 18781 5674 18847 5677
rect 21357 5674 21423 5677
rect 18781 5672 21423 5674
rect 18781 5616 18786 5672
rect 18842 5616 21362 5672
rect 21418 5616 21423 5672
rect 18781 5614 21423 5616
rect 18781 5611 18847 5614
rect 21357 5611 21423 5614
rect 17677 5538 17743 5541
rect 19793 5538 19859 5541
rect 17677 5536 19859 5538
rect 17677 5480 17682 5536
rect 17738 5480 19798 5536
rect 19854 5480 19859 5536
rect 17677 5478 19859 5480
rect 17677 5475 17743 5478
rect 19793 5475 19859 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 3417 5402 3483 5405
rect 4613 5402 4679 5405
rect 3417 5400 4679 5402
rect 3417 5344 3422 5400
rect 3478 5344 4618 5400
rect 4674 5344 4679 5400
rect 3417 5342 4679 5344
rect 3417 5339 3483 5342
rect 4613 5339 4679 5342
rect 10961 5402 11027 5405
rect 12985 5402 13051 5405
rect 10961 5400 13051 5402
rect 10961 5344 10966 5400
rect 11022 5344 12990 5400
rect 13046 5344 13051 5400
rect 10961 5342 13051 5344
rect 10961 5339 11027 5342
rect 12985 5339 13051 5342
rect 16941 5402 17007 5405
rect 20253 5402 20319 5405
rect 16941 5400 20319 5402
rect 16941 5344 16946 5400
rect 17002 5344 20258 5400
rect 20314 5344 20319 5400
rect 16941 5342 20319 5344
rect 16941 5339 17007 5342
rect 20253 5339 20319 5342
rect 5257 5266 5323 5269
rect 7649 5266 7715 5269
rect 5257 5264 7715 5266
rect 5257 5208 5262 5264
rect 5318 5208 7654 5264
rect 7710 5208 7715 5264
rect 5257 5206 7715 5208
rect 5257 5203 5323 5206
rect 7649 5203 7715 5206
rect 13721 5266 13787 5269
rect 22461 5266 22527 5269
rect 13721 5264 22527 5266
rect 13721 5208 13726 5264
rect 13782 5208 22466 5264
rect 22522 5208 22527 5264
rect 13721 5206 22527 5208
rect 13721 5203 13787 5206
rect 22461 5203 22527 5206
rect 0 5130 480 5160
rect 3601 5130 3667 5133
rect 0 5128 3667 5130
rect 0 5072 3606 5128
rect 3662 5072 3667 5128
rect 0 5070 3667 5072
rect 0 5040 480 5070
rect 3601 5067 3667 5070
rect 3969 5130 4035 5133
rect 8569 5130 8635 5133
rect 3969 5128 8635 5130
rect 3969 5072 3974 5128
rect 4030 5072 8574 5128
rect 8630 5072 8635 5128
rect 3969 5070 8635 5072
rect 3969 5067 4035 5070
rect 8569 5067 8635 5070
rect 9305 5130 9371 5133
rect 17585 5130 17651 5133
rect 9305 5128 17651 5130
rect 9305 5072 9310 5128
rect 9366 5072 17590 5128
rect 17646 5072 17651 5128
rect 9305 5070 17651 5072
rect 9305 5067 9371 5070
rect 17585 5067 17651 5070
rect 1393 4994 1459 4997
rect 9029 4994 9095 4997
rect 1393 4992 9095 4994
rect 1393 4936 1398 4992
rect 1454 4936 9034 4992
rect 9090 4936 9095 4992
rect 1393 4934 9095 4936
rect 1393 4931 1459 4934
rect 9029 4931 9095 4934
rect 13261 4994 13327 4997
rect 17217 4994 17283 4997
rect 13261 4992 17283 4994
rect 13261 4936 13266 4992
rect 13322 4936 17222 4992
rect 17278 4936 17283 4992
rect 13261 4934 17283 4936
rect 13261 4931 13327 4934
rect 17217 4931 17283 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 4863 19930 4864
rect 5441 4858 5507 4861
rect 7465 4858 7531 4861
rect 5441 4856 7531 4858
rect 5441 4800 5446 4856
rect 5502 4800 7470 4856
rect 7526 4800 7531 4856
rect 5441 4798 7531 4800
rect 5441 4795 5507 4798
rect 7465 4795 7531 4798
rect 16389 4858 16455 4861
rect 18229 4858 18295 4861
rect 16389 4856 18295 4858
rect 16389 4800 16394 4856
rect 16450 4800 18234 4856
rect 18290 4800 18295 4856
rect 16389 4798 18295 4800
rect 16389 4795 16455 4798
rect 18229 4795 18295 4798
rect 1945 4722 2011 4725
rect 4705 4722 4771 4725
rect 7373 4722 7439 4725
rect 9857 4722 9923 4725
rect 18229 4722 18295 4725
rect 1945 4720 9690 4722
rect 1945 4664 1950 4720
rect 2006 4664 4710 4720
rect 4766 4664 7378 4720
rect 7434 4664 9690 4720
rect 1945 4662 9690 4664
rect 1945 4659 2011 4662
rect 4705 4659 4771 4662
rect 7373 4659 7439 4662
rect 3141 4586 3207 4589
rect 5993 4586 6059 4589
rect 3141 4584 6059 4586
rect 3141 4528 3146 4584
rect 3202 4528 5998 4584
rect 6054 4528 6059 4584
rect 3141 4526 6059 4528
rect 9630 4586 9690 4662
rect 9857 4720 18295 4722
rect 9857 4664 9862 4720
rect 9918 4664 18234 4720
rect 18290 4664 18295 4720
rect 9857 4662 18295 4664
rect 9857 4659 9923 4662
rect 18229 4659 18295 4662
rect 12065 4586 12131 4589
rect 9630 4584 12131 4586
rect 9630 4528 12070 4584
rect 12126 4528 12131 4584
rect 9630 4526 12131 4528
rect 3141 4523 3207 4526
rect 5993 4523 6059 4526
rect 12065 4523 12131 4526
rect 12985 4586 13051 4589
rect 14641 4586 14707 4589
rect 17769 4586 17835 4589
rect 12985 4584 14707 4586
rect 12985 4528 12990 4584
rect 13046 4528 14646 4584
rect 14702 4528 14707 4584
rect 12985 4526 14707 4528
rect 12985 4523 13051 4526
rect 14641 4523 14707 4526
rect 14782 4584 17835 4586
rect 14782 4528 17774 4584
rect 17830 4528 17835 4584
rect 14782 4526 17835 4528
rect 0 4450 480 4480
rect 3693 4450 3759 4453
rect 0 4448 3759 4450
rect 0 4392 3698 4448
rect 3754 4392 3759 4448
rect 0 4390 3759 4392
rect 0 4360 480 4390
rect 3693 4387 3759 4390
rect 6913 4450 6979 4453
rect 14782 4450 14842 4526
rect 17769 4523 17835 4526
rect 6913 4448 14842 4450
rect 6913 4392 6918 4448
rect 6974 4392 14842 4448
rect 6913 4390 14842 4392
rect 16481 4450 16547 4453
rect 23473 4450 23539 4453
rect 16481 4448 23539 4450
rect 16481 4392 16486 4448
rect 16542 4392 23478 4448
rect 23534 4392 23539 4448
rect 16481 4390 23539 4392
rect 6913 4387 6979 4390
rect 16481 4387 16547 4390
rect 23473 4387 23539 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 4319 24597 4320
rect 6177 4314 6243 4317
rect 11697 4314 11763 4317
rect 6177 4312 11763 4314
rect 6177 4256 6182 4312
rect 6238 4256 11702 4312
rect 11758 4256 11763 4312
rect 6177 4254 11763 4256
rect 6177 4251 6243 4254
rect 11697 4251 11763 4254
rect 18505 4314 18571 4317
rect 22737 4314 22803 4317
rect 18505 4312 22803 4314
rect 18505 4256 18510 4312
rect 18566 4256 22742 4312
rect 22798 4256 22803 4312
rect 18505 4254 22803 4256
rect 18505 4251 18571 4254
rect 22737 4251 22803 4254
rect 289 4178 355 4181
rect 2221 4178 2287 4181
rect 3049 4178 3115 4181
rect 8753 4178 8819 4181
rect 289 4176 3115 4178
rect 289 4120 294 4176
rect 350 4120 2226 4176
rect 2282 4120 3054 4176
rect 3110 4120 3115 4176
rect 289 4118 3115 4120
rect 289 4115 355 4118
rect 2221 4115 2287 4118
rect 3049 4115 3115 4118
rect 3972 4176 8819 4178
rect 3972 4120 8758 4176
rect 8814 4120 8819 4176
rect 3972 4118 8819 4120
rect 0 3770 480 3800
rect 3972 3770 4032 4118
rect 8753 4115 8819 4118
rect 10869 4178 10935 4181
rect 21725 4178 21791 4181
rect 10869 4176 21791 4178
rect 10869 4120 10874 4176
rect 10930 4120 21730 4176
rect 21786 4120 21791 4176
rect 10869 4118 21791 4120
rect 10869 4115 10935 4118
rect 21725 4115 21791 4118
rect 8201 4042 8267 4045
rect 9673 4042 9739 4045
rect 11094 4042 11100 4044
rect 8201 4040 11100 4042
rect 8201 3984 8206 4040
rect 8262 3984 9678 4040
rect 9734 3984 11100 4040
rect 8201 3982 11100 3984
rect 8201 3979 8267 3982
rect 9673 3979 9739 3982
rect 11094 3980 11100 3982
rect 11164 3980 11170 4044
rect 11329 4042 11395 4045
rect 17125 4042 17191 4045
rect 11329 4040 17191 4042
rect 11329 3984 11334 4040
rect 11390 3984 17130 4040
rect 17186 3984 17191 4040
rect 11329 3982 17191 3984
rect 11329 3979 11395 3982
rect 17125 3979 17191 3982
rect 19149 4042 19215 4045
rect 20345 4042 20411 4045
rect 19149 4040 20411 4042
rect 19149 3984 19154 4040
rect 19210 3984 20350 4040
rect 20406 3984 20411 4040
rect 19149 3982 20411 3984
rect 19149 3979 19215 3982
rect 20345 3979 20411 3982
rect 21633 4042 21699 4045
rect 23657 4042 23723 4045
rect 21633 4040 23723 4042
rect 21633 3984 21638 4040
rect 21694 3984 23662 4040
rect 23718 3984 23723 4040
rect 21633 3982 23723 3984
rect 21633 3979 21699 3982
rect 23657 3979 23723 3982
rect 5257 3906 5323 3909
rect 9857 3906 9923 3909
rect 5257 3904 9923 3906
rect 5257 3848 5262 3904
rect 5318 3848 9862 3904
rect 9918 3848 9923 3904
rect 5257 3846 9923 3848
rect 5257 3843 5323 3846
rect 9857 3843 9923 3846
rect 13445 3906 13511 3909
rect 16297 3906 16363 3909
rect 13445 3904 16363 3906
rect 13445 3848 13450 3904
rect 13506 3848 16302 3904
rect 16358 3848 16363 3904
rect 13445 3846 16363 3848
rect 13445 3843 13511 3846
rect 16297 3843 16363 3846
rect 20621 3906 20687 3909
rect 21541 3906 21607 3909
rect 20621 3904 21607 3906
rect 20621 3848 20626 3904
rect 20682 3848 21546 3904
rect 21602 3848 21607 3904
rect 20621 3846 21607 3848
rect 20621 3843 20687 3846
rect 21541 3843 21607 3846
rect 10277 3840 10597 3841
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 0 3710 4032 3770
rect 5717 3770 5783 3773
rect 9305 3770 9371 3773
rect 5717 3768 9371 3770
rect 5717 3712 5722 3768
rect 5778 3712 9310 3768
rect 9366 3712 9371 3768
rect 5717 3710 9371 3712
rect 0 3680 480 3710
rect 5717 3707 5783 3710
rect 9305 3707 9371 3710
rect 14181 3770 14247 3773
rect 18505 3770 18571 3773
rect 19425 3772 19491 3773
rect 19374 3770 19380 3772
rect 14181 3768 18571 3770
rect 14181 3712 14186 3768
rect 14242 3712 18510 3768
rect 18566 3712 18571 3768
rect 14181 3710 18571 3712
rect 19334 3710 19380 3770
rect 19444 3768 19491 3772
rect 19486 3712 19491 3768
rect 14181 3707 14247 3710
rect 18505 3707 18571 3710
rect 19374 3708 19380 3710
rect 19444 3708 19491 3712
rect 19425 3707 19491 3708
rect 2957 3634 3023 3637
rect 14733 3634 14799 3637
rect 18413 3634 18479 3637
rect 2957 3632 14799 3634
rect 2957 3576 2962 3632
rect 3018 3576 14738 3632
rect 14794 3576 14799 3632
rect 2957 3574 14799 3576
rect 2957 3571 3023 3574
rect 14733 3571 14799 3574
rect 15150 3632 18479 3634
rect 15150 3576 18418 3632
rect 18474 3576 18479 3632
rect 15150 3574 18479 3576
rect 2497 3498 2563 3501
rect 9121 3498 9187 3501
rect 11789 3498 11855 3501
rect 2497 3496 8954 3498
rect 2497 3440 2502 3496
rect 2558 3440 8954 3496
rect 2497 3438 8954 3440
rect 2497 3435 2563 3438
rect 2313 3362 2379 3365
rect 3601 3362 3667 3365
rect 2313 3360 3667 3362
rect 2313 3304 2318 3360
rect 2374 3304 3606 3360
rect 3662 3304 3667 3360
rect 2313 3302 3667 3304
rect 8894 3362 8954 3438
rect 9121 3496 11855 3498
rect 9121 3440 9126 3496
rect 9182 3440 11794 3496
rect 11850 3440 11855 3496
rect 9121 3438 11855 3440
rect 9121 3435 9187 3438
rect 11789 3435 11855 3438
rect 12617 3498 12683 3501
rect 15150 3498 15210 3574
rect 18413 3571 18479 3574
rect 18597 3634 18663 3637
rect 20989 3634 21055 3637
rect 18597 3632 21055 3634
rect 18597 3576 18602 3632
rect 18658 3576 20994 3632
rect 21050 3576 21055 3632
rect 18597 3574 21055 3576
rect 18597 3571 18663 3574
rect 20989 3571 21055 3574
rect 22001 3634 22067 3637
rect 25129 3634 25195 3637
rect 22001 3632 25195 3634
rect 22001 3576 22006 3632
rect 22062 3576 25134 3632
rect 25190 3576 25195 3632
rect 22001 3574 25195 3576
rect 22001 3571 22067 3574
rect 25129 3571 25195 3574
rect 12617 3496 15210 3498
rect 12617 3440 12622 3496
rect 12678 3440 15210 3496
rect 12617 3438 15210 3440
rect 15377 3498 15443 3501
rect 20253 3498 20319 3501
rect 15377 3496 20319 3498
rect 15377 3440 15382 3496
rect 15438 3440 20258 3496
rect 20314 3440 20319 3496
rect 15377 3438 20319 3440
rect 12617 3435 12683 3438
rect 15377 3435 15443 3438
rect 20253 3435 20319 3438
rect 9673 3362 9739 3365
rect 8894 3360 9739 3362
rect 8894 3304 9678 3360
rect 9734 3304 9739 3360
rect 8894 3302 9739 3304
rect 2313 3299 2379 3302
rect 3601 3299 3667 3302
rect 9673 3299 9739 3302
rect 15653 3362 15719 3365
rect 19333 3362 19399 3365
rect 15653 3360 19399 3362
rect 15653 3304 15658 3360
rect 15714 3304 19338 3360
rect 19394 3304 19399 3360
rect 15653 3302 19399 3304
rect 15653 3299 15719 3302
rect 19333 3299 19399 3302
rect 5610 3296 5930 3297
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 2589 3226 2655 3229
rect 4797 3226 4863 3229
rect 2589 3224 4863 3226
rect 2589 3168 2594 3224
rect 2650 3168 4802 3224
rect 4858 3168 4863 3224
rect 2589 3166 4863 3168
rect 2589 3163 2655 3166
rect 4797 3163 4863 3166
rect 9673 3226 9739 3229
rect 14641 3226 14707 3229
rect 9673 3224 14707 3226
rect 9673 3168 9678 3224
rect 9734 3168 14646 3224
rect 14702 3168 14707 3224
rect 9673 3166 14707 3168
rect 9673 3163 9739 3166
rect 14641 3163 14707 3166
rect 17585 3226 17651 3229
rect 20805 3226 20871 3229
rect 17585 3224 20871 3226
rect 17585 3168 17590 3224
rect 17646 3168 20810 3224
rect 20866 3168 20871 3224
rect 17585 3166 20871 3168
rect 17585 3163 17651 3166
rect 20805 3163 20871 3166
rect 0 3090 480 3120
rect 1301 3090 1367 3093
rect 0 3088 1367 3090
rect 0 3032 1306 3088
rect 1362 3032 1367 3088
rect 0 3030 1367 3032
rect 0 3000 480 3030
rect 1301 3027 1367 3030
rect 3325 3090 3391 3093
rect 5533 3090 5599 3093
rect 3325 3088 5599 3090
rect 3325 3032 3330 3088
rect 3386 3032 5538 3088
rect 5594 3032 5599 3088
rect 3325 3030 5599 3032
rect 3325 3027 3391 3030
rect 5533 3027 5599 3030
rect 7373 3090 7439 3093
rect 11145 3090 11211 3093
rect 7373 3088 11211 3090
rect 7373 3032 7378 3088
rect 7434 3032 11150 3088
rect 11206 3032 11211 3088
rect 7373 3030 11211 3032
rect 7373 3027 7439 3030
rect 11145 3027 11211 3030
rect 14590 3028 14596 3092
rect 14660 3090 14666 3092
rect 14733 3090 14799 3093
rect 14660 3088 14799 3090
rect 14660 3032 14738 3088
rect 14794 3032 14799 3088
rect 14660 3030 14799 3032
rect 14660 3028 14666 3030
rect 14733 3027 14799 3030
rect 15561 3090 15627 3093
rect 21817 3090 21883 3093
rect 15561 3088 21883 3090
rect 15561 3032 15566 3088
rect 15622 3032 21822 3088
rect 21878 3032 21883 3088
rect 15561 3030 21883 3032
rect 15561 3027 15627 3030
rect 21817 3027 21883 3030
rect 4705 2954 4771 2957
rect 8477 2954 8543 2957
rect 4705 2952 8543 2954
rect 4705 2896 4710 2952
rect 4766 2896 8482 2952
rect 8538 2896 8543 2952
rect 4705 2894 8543 2896
rect 4705 2891 4771 2894
rect 8477 2891 8543 2894
rect 14825 2954 14891 2957
rect 18137 2954 18203 2957
rect 22001 2954 22067 2957
rect 14825 2952 15578 2954
rect 14825 2896 14830 2952
rect 14886 2896 15578 2952
rect 14825 2894 15578 2896
rect 14825 2891 14891 2894
rect 3233 2818 3299 2821
rect 6361 2818 6427 2821
rect 3233 2816 6427 2818
rect 3233 2760 3238 2816
rect 3294 2760 6366 2816
rect 6422 2760 6427 2816
rect 3233 2758 6427 2760
rect 15518 2818 15578 2894
rect 18137 2952 22067 2954
rect 18137 2896 18142 2952
rect 18198 2896 22006 2952
rect 22062 2896 22067 2952
rect 18137 2894 22067 2896
rect 18137 2891 18203 2894
rect 22001 2891 22067 2894
rect 19425 2818 19491 2821
rect 15518 2816 19491 2818
rect 15518 2760 19430 2816
rect 19486 2760 19491 2816
rect 15518 2758 19491 2760
rect 3233 2755 3299 2758
rect 6361 2755 6427 2758
rect 19425 2755 19491 2758
rect 21081 2818 21147 2821
rect 22645 2818 22711 2821
rect 21081 2816 22711 2818
rect 21081 2760 21086 2816
rect 21142 2760 22650 2816
rect 22706 2760 22711 2816
rect 21081 2758 22711 2760
rect 21081 2755 21147 2758
rect 22645 2755 22711 2758
rect 25129 2818 25195 2821
rect 27061 2818 27127 2821
rect 25129 2816 27127 2818
rect 25129 2760 25134 2816
rect 25190 2760 27066 2816
rect 27122 2760 27127 2816
rect 25129 2758 27127 2760
rect 25129 2755 25195 2758
rect 27061 2755 27127 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 11053 2682 11119 2685
rect 16757 2682 16823 2685
rect 11053 2680 16823 2682
rect 11053 2624 11058 2680
rect 11114 2624 16762 2680
rect 16818 2624 16823 2680
rect 11053 2622 16823 2624
rect 11053 2619 11119 2622
rect 16757 2619 16823 2622
rect 6453 2546 6519 2549
rect 3190 2544 6519 2546
rect 3190 2488 6458 2544
rect 6514 2488 6519 2544
rect 3190 2486 6519 2488
rect 0 2410 480 2440
rect 3190 2410 3250 2486
rect 6453 2483 6519 2486
rect 10041 2546 10107 2549
rect 13997 2546 14063 2549
rect 10041 2544 14063 2546
rect 10041 2488 10046 2544
rect 10102 2488 14002 2544
rect 14058 2488 14063 2544
rect 10041 2486 14063 2488
rect 10041 2483 10107 2486
rect 13997 2483 14063 2486
rect 17033 2546 17099 2549
rect 22277 2546 22343 2549
rect 17033 2544 22343 2546
rect 17033 2488 17038 2544
rect 17094 2488 22282 2544
rect 22338 2488 22343 2544
rect 17033 2486 22343 2488
rect 17033 2483 17099 2486
rect 22277 2483 22343 2486
rect 0 2350 3250 2410
rect 4153 2410 4219 2413
rect 20529 2410 20595 2413
rect 4153 2408 20595 2410
rect 4153 2352 4158 2408
rect 4214 2352 20534 2408
rect 20590 2352 20595 2408
rect 4153 2350 20595 2352
rect 0 2320 480 2350
rect 4153 2347 4219 2350
rect 20529 2347 20595 2350
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 15745 2138 15811 2141
rect 16665 2138 16731 2141
rect 15745 2136 16731 2138
rect 15745 2080 15750 2136
rect 15806 2080 16670 2136
rect 16726 2080 16731 2136
rect 15745 2078 16731 2080
rect 15745 2075 15811 2078
rect 16665 2075 16731 2078
rect 16849 2138 16915 2141
rect 24025 2138 24091 2141
rect 16849 2136 24091 2138
rect 16849 2080 16854 2136
rect 16910 2080 24030 2136
rect 24086 2080 24091 2136
rect 16849 2078 24091 2080
rect 16849 2075 16915 2078
rect 24025 2075 24091 2078
rect 11421 2002 11487 2005
rect 3374 2000 11487 2002
rect 3374 1944 11426 2000
rect 11482 1944 11487 2000
rect 3374 1942 11487 1944
rect 0 1730 480 1760
rect 3374 1730 3434 1942
rect 11421 1939 11487 1942
rect 13077 2002 13143 2005
rect 21173 2002 21239 2005
rect 13077 2000 21239 2002
rect 13077 1944 13082 2000
rect 13138 1944 21178 2000
rect 21234 1944 21239 2000
rect 13077 1942 21239 1944
rect 13077 1939 13143 1942
rect 21173 1939 21239 1942
rect 11421 1866 11487 1869
rect 19609 1866 19675 1869
rect 11421 1864 19675 1866
rect 11421 1808 11426 1864
rect 11482 1808 19614 1864
rect 19670 1808 19675 1864
rect 11421 1806 19675 1808
rect 11421 1803 11487 1806
rect 19609 1803 19675 1806
rect 0 1670 3434 1730
rect 10961 1730 11027 1733
rect 27613 1730 27679 1733
rect 10961 1728 27679 1730
rect 10961 1672 10966 1728
rect 11022 1672 27618 1728
rect 27674 1672 27679 1728
rect 10961 1670 27679 1672
rect 0 1640 480 1670
rect 10961 1667 11027 1670
rect 27613 1667 27679 1670
rect 12801 1594 12867 1597
rect 16849 1594 16915 1597
rect 12801 1592 16915 1594
rect 12801 1536 12806 1592
rect 12862 1536 16854 1592
rect 16910 1536 16915 1592
rect 12801 1534 16915 1536
rect 12801 1531 12867 1534
rect 16849 1531 16915 1534
rect 17033 1594 17099 1597
rect 22461 1594 22527 1597
rect 17033 1592 22527 1594
rect 17033 1536 17038 1592
rect 17094 1536 22466 1592
rect 22522 1536 22527 1592
rect 17033 1534 22527 1536
rect 17033 1531 17099 1534
rect 22461 1531 22527 1534
rect 2957 1458 3023 1461
rect 14641 1458 14707 1461
rect 2957 1456 14707 1458
rect 2957 1400 2962 1456
rect 3018 1400 14646 1456
rect 14702 1400 14707 1456
rect 2957 1398 14707 1400
rect 2957 1395 3023 1398
rect 14641 1395 14707 1398
rect 15469 1458 15535 1461
rect 19425 1458 19491 1461
rect 15469 1456 19491 1458
rect 15469 1400 15474 1456
rect 15530 1400 19430 1456
rect 19486 1400 19491 1456
rect 15469 1398 19491 1400
rect 15469 1395 15535 1398
rect 19425 1395 19491 1398
rect 3693 1322 3759 1325
rect 20161 1322 20227 1325
rect 3693 1320 20227 1322
rect 3693 1264 3698 1320
rect 3754 1264 20166 1320
rect 20222 1264 20227 1320
rect 3693 1262 20227 1264
rect 3693 1259 3759 1262
rect 20161 1259 20227 1262
rect 0 1050 480 1080
rect 1485 1050 1551 1053
rect 0 1048 1551 1050
rect 0 992 1490 1048
rect 1546 992 1551 1048
rect 0 990 1551 992
rect 0 960 480 990
rect 1485 987 1551 990
rect 0 370 480 400
rect 3141 370 3207 373
rect 0 368 3207 370
rect 0 312 3146 368
rect 3202 312 3207 368
rect 0 310 3207 312
rect 0 280 480 310
rect 3141 307 3207 310
<< via3 >>
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 14596 9420 14660 9484
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 11100 3980 11164 4044
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 19380 3768 19444 3772
rect 19380 3712 19430 3768
rect 19430 3712 19444 3768
rect 19380 3708 19444 3712
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 14596 3028 14660 3092
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
<< metal4 >>
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 5610 9824 5931 10848
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 5610 3296 5931 4320
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 19072 10597 20096
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 19616 15264 20640
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 18528 15264 19552
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 12000 15264 13024
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 10912 15264 11936
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14595 9484 14661 9485
rect 14595 9420 14596 9484
rect 14660 9420 14661 9484
rect 14595 9419 14661 9420
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 6016 10597 7040
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 3840 10597 4864
rect 11099 4044 11165 4045
rect 11099 3980 11100 4044
rect 11164 3980 11165 4044
rect 11099 3979 11165 3980
rect 11102 3858 11162 3979
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 2752 10597 3776
rect 14598 3093 14658 9419
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 3296 15264 4320
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 19072 19930 20096
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 12544 19930 13568
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 19610 3840 19930 4864
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14595 3092 14661 3093
rect 14595 3028 14596 3092
rect 14660 3028 14661 3092
rect 14595 3027 14661 3028
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 19610 2752 19930 3776
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2128 19930 2688
rect 24277 25056 24597 25616
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
<< via4 >>
rect 11014 3622 11250 3858
rect 19294 3772 19530 3858
rect 19294 3708 19380 3772
rect 19380 3708 19444 3772
rect 19444 3708 19530 3772
rect 19294 3622 19530 3708
<< metal5 >>
rect 10972 3858 19572 3900
rect 10972 3622 11014 3858
rect 11250 3622 19294 3858
rect 19530 3622 19572 3858
rect 10972 3580 19572 3622
use scs8hd_fill_2  FILLER_1_9 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_6
timestamp 1586364061
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_buf_4  mux_left_track_9.scs8hd_buf_4_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 590 592
use scs8hd_conb_1  _34_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_13
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_10
timestamp 1586364061
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_9.mux_l1_in_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2668 0 1 2720
box -38 -48 866 592
use scs8hd_mux2_2  mux_left_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_26
timestamp 1586364061
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_30
timestamp 1586364061
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_86 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_0_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 4232 0 1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_51 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5796 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_55 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 6164 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 7176 0 -1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_left_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 7084 0 1 2720
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  FILLER_1_62
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_88
timestamp 1586364061
transform 1 0 9200 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_84
timestamp 1586364061
transform 1 0 8832 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_89
timestamp 1586364061
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_85
timestamp 1586364061
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9016 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_left_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11868 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_113
timestamp 1586364061
transform 1 0 11500 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_117
timestamp 1586364061
transform 1 0 11868 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_111
timestamp 1586364061
transform 1 0 11316 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_115
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_119
timestamp 1586364061
transform 1 0 12052 0 1 2720
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_39.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_left_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_142
timestamp 1586364061
transform 1 0 14168 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_144
timestamp 1586364061
transform 1 0 14352 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_150
timestamp 1586364061
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_146
timestamp 1586364061
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_152
timestamp 1586364061
transform 1 0 15088 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_0_148
timestamp 1586364061
transform 1 0 14720 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 14904 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_9.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15088 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_158
timestamp 1586364061
transform 1 0 15640 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_4  mux_bottom_track_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_162
timestamp 1586364061
transform 1 0 16008 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_168
timestamp 1586364061
transform 1 0 16560 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_162
timestamp 1586364061
transform 1 0 16008 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 15824 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16376 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_37.mux_l2_in_0_
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_176
timestamp 1586364061
transform 1 0 17296 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_3.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16744 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_180
timestamp 1586364061
transform 1 0 17664 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_4  mux_bottom_track_17.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_197
timestamp 1586364061
transform 1 0 19228 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_193
timestamp 1586364061
transform 1 0 18860 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 19044 0 -1 2720
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_39.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_1_203
timestamp 1586364061
transform 1 0 19780 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_205
timestamp 1586364061
transform 1 0 19964 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 19412 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__52__A
timestamp 1586364061
transform 1 0 19964 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _54_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 19596 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_207
timestamp 1586364061
transform 1 0 20148 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_209
timestamp 1586364061
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__54__A
timestamp 1586364061
transform 1 0 20148 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_4  mux_bottom_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20516 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_217
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_213
timestamp 1586364061
transform 1 0 20700 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _51_
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_221
timestamp 1586364061
transform 1 0 21436 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_226
timestamp 1586364061
transform 1 0 21896 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_222
timestamp 1586364061
transform 1 0 21528 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__85__A
timestamp 1586364061
transform 1 0 21620 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 21252 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__51__A
timestamp 1586364061
transform 1 0 21712 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _84_
timestamp 1586364061
transform 1 0 21804 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_233
timestamp 1586364061
transform 1 0 22540 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_229
timestamp 1586364061
transform 1 0 22172 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_234
timestamp 1586364061
transform 1 0 22632 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__84__A
timestamp 1586364061
transform 1 0 22356 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22724 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _86_
timestamp 1586364061
transform 1 0 22264 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_4  FILLER_1_237
timestamp 1586364061
transform 1 0 22908 0 1 2720
box -38 -48 406 592
use scs8hd_decap_8  FILLER_0_238 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 23000 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__86__A
timestamp 1586364061
transform 1 0 22816 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_241
timestamp 1586364061
transform 1 0 23276 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_251
timestamp 1586364061
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_246
timestamp 1586364061
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_4  mux_bottom_track_39.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 590 592
use scs8hd_buf_4  mux_bottom_track_37.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_255
timestamp 1586364061
transform 1 0 24564 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_255
timestamp 1586364061
transform 1 0 24564 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 24748 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__68__A
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__75__A
timestamp 1586364061
transform 1 0 24380 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_263
timestamp 1586364061
transform 1 0 25300 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_259
timestamp 1586364061
transform 1 0 24932 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__72__A
timestamp 1586364061
transform 1 0 25484 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _69_
timestamp 1586364061
transform 1 0 25300 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _68_
timestamp 1586364061
transform 1 0 24932 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_275
timestamp 1586364061
transform 1 0 26404 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_1_267
timestamp 1586364061
transform 1 0 25668 0 1 2720
box -38 -48 774 592
use scs8hd_decap_6  FILLER_0_271 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 26036 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_267
timestamp 1586364061
transform 1 0 25668 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__69__A
timestamp 1586364061
transform 1 0 25852 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use scs8hd_conb_1  _33_
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_6
timestamp 1586364061
transform 1 0 1656 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_2_12
timestamp 1586364061
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_23
timestamp 1586364061
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_27
timestamp 1586364061
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_left_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5704 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5428 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_41
timestamp 1586364061
transform 1 0 4876 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_45
timestamp 1586364061
transform 1 0 5244 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_49
timestamp 1586364061
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use scs8hd_buf_4  mux_left_track_25.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 8188 0 -1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 7636 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 8004 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_69
timestamp 1586364061
transform 1 0 7452 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_73
timestamp 1586364061
transform 1 0 7820 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_4  mux_left_track_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_83
timestamp 1586364061
transform 1 0 8740 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_87
timestamp 1586364061
transform 1 0 9108 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_90
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_99
timestamp 1586364061
transform 1 0 10212 0 -1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_39.mux_l1_in_0_
timestamp 1586364061
transform 1 0 11132 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10396 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_103
timestamp 1586364061
transform 1 0 10580 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_107
timestamp 1586364061
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_118
timestamp 1586364061
transform 1 0 11960 0 -1 3808
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_39.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12696 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_39.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_122
timestamp 1586364061
transform 1 0 12328 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_125
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_4  FILLER_2_135
timestamp 1586364061
transform 1 0 13524 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_4  mux_bottom_track_7.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14720 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_139
timestamp 1586364061
transform 1 0 13892 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_142
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_146
timestamp 1586364061
transform 1 0 14536 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_150
timestamp 1586364061
transform 1 0 14904 0 -1 3808
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_37.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16744 0 -1 3808
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 16008 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 16376 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_160
timestamp 1586364061
transform 1 0 15824 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_164
timestamp 1586364061
transform 1 0 16192 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_168
timestamp 1586364061
transform 1 0 16560 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _52_
timestamp 1586364061
transform 1 0 19228 0 -1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 18676 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_189
timestamp 1586364061
transform 1 0 18492 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_193
timestamp 1586364061
transform 1 0 18860 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _85_
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20148 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_201
timestamp 1586364061
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_205
timestamp 1586364061
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_209
timestamp 1586364061
transform 1 0 20332 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_213
timestamp 1586364061
transform 1 0 20700 0 -1 3808
box -38 -48 130 592
use scs8hd_buf_4  mux_bottom_track_35.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22724 0 -1 3808
box -38 -48 590 592
use scs8hd_decap_12  FILLER_2_219 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 21252 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_2_231
timestamp 1586364061
transform 1 0 22356 0 -1 3808
box -38 -48 406 592
use scs8hd_buf_2  _75_
timestamp 1586364061
transform 1 0 24012 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_8  FILLER_2_241
timestamp 1586364061
transform 1 0 23276 0 -1 3808
box -38 -48 774 592
use scs8hd_decap_8  FILLER_2_253
timestamp 1586364061
transform 1 0 24380 0 -1 3808
box -38 -48 774 592
use scs8hd_buf_2  _72_
timestamp 1586364061
transform 1 0 25116 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_265
timestamp 1586364061
transform 1 0 25484 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_2_273
timestamp 1586364061
transform 1 0 26220 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_276
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l1_in_1_
timestamp 1586364061
transform 1 0 2024 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_3_7
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_19
timestamp 1586364061
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 3588 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_23
timestamp 1586364061
transform 1 0 3220 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_36
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_40
timestamp 1586364061
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l1_in_1_
timestamp 1586364061
transform 1 0 7636 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 7452 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 6992 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_62
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_66
timestamp 1586364061
transform 1 0 7176 0 1 3808
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__58__A
timestamp 1586364061
transform 1 0 8648 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_80
timestamp 1586364061
transform 1 0 8464 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_84
timestamp 1586364061
transform 1 0 8832 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_97
timestamp 1586364061
transform 1 0 10028 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_31.mux_l2_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_101
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_23.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_132
timestamp 1586364061
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_136
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_35.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 15180 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_149
timestamp 1586364061
transform 1 0 14812 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_155
timestamp 1586364061
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_37.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_37.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16744 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_168
timestamp 1586364061
transform 1 0 16560 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_172
timestamp 1586364061
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_176
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 406 592
use scs8hd_buf_2  _48_
timestamp 1586364061
transform 1 0 19320 0 1 3808
box -38 -48 406 592
use scs8hd_buf_4  mux_bottom_track_1.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 18768 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_35.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_180
timestamp 1586364061
transform 1 0 17664 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_190
timestamp 1586364061
transform 1 0 18584 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_194
timestamp 1586364061
transform 1 0 18952 0 1 3808
box -38 -48 222 592
use scs8hd_buf_2  _83_
timestamp 1586364061
transform 1 0 20424 0 1 3808
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__48__A
timestamp 1586364061
transform 1 0 19872 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__79__A
timestamp 1586364061
transform 1 0 20976 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__83__A
timestamp 1586364061
transform 1 0 20240 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_202
timestamp 1586364061
transform 1 0 19688 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_206
timestamp 1586364061
transform 1 0 20056 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_214
timestamp 1586364061
transform 1 0 20792 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_218
timestamp 1586364061
transform 1 0 21160 0 1 3808
box -38 -48 590 592
use scs8hd_buf_4  mux_bottom_track_31.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 21712 0 1 3808
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_230
timestamp 1586364061
transform 1 0 22264 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_234
timestamp 1586364061
transform 1 0 22632 0 1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_3_238
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 590 592
use scs8hd_buf_2  _70_
timestamp 1586364061
transform 1 0 24748 0 1 3808
box -38 -48 406 592
use scs8hd_buf_2  _73_
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__73__A
timestamp 1586364061
transform 1 0 24196 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__71__A
timestamp 1586364061
transform 1 0 24564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_249
timestamp 1586364061
transform 1 0 24012 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_253
timestamp 1586364061
transform 1 0 24380 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__70__A
timestamp 1586364061
transform 1 0 25300 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_261
timestamp 1586364061
transform 1 0 25116 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_265
timestamp 1586364061
transform 1 0 25484 0 1 3808
box -38 -48 1142 592
use scs8hd_conb_1  _32_
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l1_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_6
timestamp 1586364061
transform 1 0 1656 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_12
timestamp 1586364061
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_23
timestamp 1586364061
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5980 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_51
timestamp 1586364061
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_55
timestamp 1586364061
transform 1 0 6164 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_59
timestamp 1586364061
transform 1 0 6532 0 -1 4896
box -38 -48 130 592
use scs8hd_buf_2  _58_
timestamp 1586364061
transform 1 0 8372 0 -1 4896
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l3_in_0_
timestamp 1586364061
transform 1 0 6808 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_71
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_75
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_left_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_83
timestamp 1586364061
transform 1 0 8740 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_87
timestamp 1586364061
transform 1 0 9108 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_90
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_31.mux_l1_in_0_
timestamp 1586364061
transform 1 0 11224 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_102
timestamp 1586364061
transform 1 0 10488 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_3  FILLER_4_107
timestamp 1586364061
transform 1 0 10948 0 -1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_4_119
timestamp 1586364061
transform 1 0 12052 0 -1 4896
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_33.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12880 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 12420 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_125
timestamp 1586364061
transform 1 0 12604 0 -1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_4_137
timestamp 1586364061
transform 1 0 13708 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_141
timestamp 1586364061
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 14260 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 13892 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_158
timestamp 1586364061
transform 1 0 15640 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_154
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_37.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15916 0 -1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_37.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15732 0 -1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_35.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18400 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17848 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_180
timestamp 1586364061
transform 1 0 17664 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_184
timestamp 1586364061
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_4_197
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 1142 592
use scs8hd_buf_2  _79_
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_4_209
timestamp 1586364061
transform 1 0 20332 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_213
timestamp 1586364061
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use scs8hd_buf_4  mux_bottom_track_33.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 22448 0 -1 4896
box -38 -48 590 592
use scs8hd_decap_12  FILLER_4_219
timestamp 1586364061
transform 1 0 21252 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_231
timestamp 1586364061
transform 1 0 22356 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_238
timestamp 1586364061
transform 1 0 23000 0 -1 4896
box -38 -48 774 592
use scs8hd_buf_2  _71_
timestamp 1586364061
transform 1 0 23736 0 -1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_4_250
timestamp 1586364061
transform 1 0 24104 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_262
timestamp 1586364061
transform 1 0 25208 0 -1 4896
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_4_274
timestamp 1586364061
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 1840 0 1 4896
box -38 -48 1786 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 1564 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_7
timestamp 1586364061
transform 1 0 1748 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3864 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_32
timestamp 1586364061
transform 1 0 4048 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_36
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l1_in_2_
timestamp 1586364061
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_40
timestamp 1586364061
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 7084 0 1 4896
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_decap_3  FILLER_5_62
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use scs8hd_mux2_2  mux_left_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9568 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_84
timestamp 1586364061
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_88
timestamp 1586364061
transform 1 0 9200 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _65_
timestamp 1586364061
transform 1 0 11132 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_31.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11684 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_101
timestamp 1586364061
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_105
timestamp 1586364061
transform 1 0 10764 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_113
timestamp 1586364061
transform 1 0 11500 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_117
timestamp 1586364061
transform 1 0 11868 0 1 4896
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_35.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 14904 0 1 4896
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 14352 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14720 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_142
timestamp 1586364061
transform 1 0 14168 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_146
timestamp 1586364061
transform 1 0 14536 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 16836 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_39.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_169
timestamp 1586364061
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_173
timestamp 1586364061
transform 1 0 17020 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_177
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _82_
timestamp 1586364061
transform 1 0 19136 0 1 4896
box -38 -48 406 592
use scs8hd_buf_2  _87_
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__87__A
timestamp 1586364061
transform 1 0 18584 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18952 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_181
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_188
timestamp 1586364061
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_192
timestamp 1586364061
transform 1 0 18768 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _81_
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__82__A
timestamp 1586364061
transform 1 0 19688 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__81__A
timestamp 1586364061
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__76__A
timestamp 1586364061
transform 1 0 21160 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_200
timestamp 1586364061
transform 1 0 19504 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_204
timestamp 1586364061
transform 1 0 19872 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_212
timestamp 1586364061
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_216
timestamp 1586364061
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use scs8hd_buf_2  _74_
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 406 592
use scs8hd_buf_2  _77_
timestamp 1586364061
transform 1 0 21344 0 1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__77__A
timestamp 1586364061
transform 1 0 21896 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__74__A
timestamp 1586364061
transform 1 0 23000 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_224
timestamp 1586364061
transform 1 0 21712 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_228
timestamp 1586364061
transform 1 0 22080 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_decap_4  FILLER_5_240
timestamp 1586364061
transform 1 0 23184 0 1 4896
box -38 -48 406 592
use scs8hd_decap_12  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_257
timestamp 1586364061
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use scs8hd_decap_8  FILLER_5_269
timestamp 1586364061
transform 1 0 25852 0 1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_3
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_4  mux_left_track_5.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 1564 0 1 5984
box -38 -48 590 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l2_in_1_
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_11
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_16
timestamp 1586364061
transform 1 0 2576 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_12
timestamp 1586364061
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2760 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 2668 0 1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 2852 0 1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_6_27
timestamp 1586364061
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_23
timestamp 1586364061
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_3.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use scs8hd_conb_1  _35_
timestamp 1586364061
transform 1 0 2944 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_38
timestamp 1586364061
transform 1 0 4600 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_36
timestamp 1586364061
transform 1 0 4416 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 4232 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_3.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 4692 0 -1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_7_42
timestamp 1586364061
transform 1 0 4968 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 5152 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 4784 0 1 5984
box -38 -48 222 592
use scs8hd_buf_2  _67_
timestamp 1586364061
transform 1 0 5336 0 1 5984
box -38 -48 406 592
use scs8hd_decap_4  FILLER_7_54
timestamp 1586364061
transform 1 0 6072 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_50
timestamp 1586364061
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_58
timestamp 1586364061
transform 1 0 6440 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_58
timestamp 1586364061
transform 1 0 6440 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_62
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_62
timestamp 1586364061
transform 1 0 6808 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6992 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l2_in_1_
timestamp 1586364061
transform 1 0 7176 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_79
timestamp 1586364061
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_75
timestamp 1586364061
transform 1 0 8004 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8188 0 -1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6992 0 1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_7_87
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_83
timestamp 1586364061
transform 1 0 8740 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_87
timestamp 1586364061
transform 1 0 9108 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_83
timestamp 1586364061
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8556 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_97
timestamp 1586364061
transform 1 0 10028 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_left_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 10212 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_31.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_31.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9476 0 1 5984
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_31.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10396 0 -1 5984
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 11408 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_110
timestamp 1586364061
transform 1 0 11224 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_123
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_125
timestamp 1586364061
transform 1 0 12604 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_120
timestamp 1586364061
transform 1 0 12144 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12420 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_33.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12604 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_33.mux_l1_in_0_
timestamp 1586364061
transform 1 0 12880 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_6_137
timestamp 1586364061
transform 1 0 13708 0 -1 5984
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_33.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12788 0 1 5984
box -38 -48 1786 592
use scs8hd_fill_2  FILLER_7_146
timestamp 1586364061
transform 1 0 14536 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 14260 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__49__A
timestamp 1586364061
transform 1 0 14720 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__53__A
timestamp 1586364061
transform 1 0 13892 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_154
timestamp 1586364061
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_150
timestamp 1586364061
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_152
timestamp 1586364061
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_1  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_35.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14904 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 15088 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_21.mux_l1_in_0_
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 866 592
use scs8hd_dfxbp_1  mem_bottom_track_35.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 16652 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 17020 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 17204 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_173
timestamp 1586364061
transform 1 0 17020 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_177
timestamp 1586364061
transform 1 0 17388 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_167
timestamp 1586364061
transform 1 0 16468 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_171
timestamp 1586364061
transform 1 0 16836 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_175
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_179
timestamp 1586364061
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_186
timestamp 1586364061
transform 1 0 18216 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  FILLER_6_181
timestamp 1586364061
transform 1 0 17756 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__65__A
timestamp 1586364061
transform 1 0 17572 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_21.mux_l2_in_0_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use scs8hd_decap_6  FILLER_7_193
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 590 592
use scs8hd_decap_8  FILLER_6_195
timestamp 1586364061
transform 1 0 19044 0 -1 5984
box -38 -48 774 592
use scs8hd_buf_4  mux_bottom_track_21.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18492 0 -1 5984
box -38 -48 590 592
use scs8hd_conb_1  _26_
timestamp 1586364061
transform 1 0 19780 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_2  _76_
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use scs8hd_buf_4  mux_bottom_track_23.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__78__A
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20332 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_206
timestamp 1586364061
transform 1 0 20056 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_207
timestamp 1586364061
transform 1 0 20148 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_7_211
timestamp 1586364061
transform 1 0 20516 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_219
timestamp 1586364061
transform 1 0 21252 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_231
timestamp 1586364061
transform 1 0 22356 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_223
timestamp 1586364061
transform 1 0 21620 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_235
timestamp 1586364061
transform 1 0 22724 0 1 5984
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_bottom_track_1.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 24104 0 1 5984
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 23920 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_1.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 24104 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_6_243
timestamp 1586364061
transform 1 0 23460 0 -1 5984
box -38 -48 590 592
use scs8hd_fill_1  FILLER_6_249
timestamp 1586364061
transform 1 0 24012 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_252
timestamp 1586364061
transform 1 0 24288 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_7_243
timestamp 1586364061
transform 1 0 23460 0 1 5984
box -38 -48 130 592
use scs8hd_decap_3  FILLER_7_245
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_264
timestamp 1586364061
transform 1 0 25392 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_272
timestamp 1586364061
transform 1 0 26128 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_276
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_7_269
timestamp 1586364061
transform 1 0 25852 0 1 5984
box -38 -48 774 592
use scs8hd_conb_1  _46_
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l2_in_0_
timestamp 1586364061
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 1840 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_10
timestamp 1586364061
transform 1 0 2024 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l1_in_1_
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__S
timestamp 1586364061
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_23
timestamp 1586364061
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_27
timestamp 1586364061
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l1_in_1_
timestamp 1586364061
transform 1 0 5612 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_41
timestamp 1586364061
transform 1 0 4876 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  FILLER_8_46
timestamp 1586364061
transform 1 0 5336 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_8_58
timestamp 1586364061
transform 1 0 6440 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7176 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 6624 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 8188 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_62
timestamp 1586364061
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_75
timestamp 1586364061
transform 1 0 8004 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_79
timestamp 1586364061
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_3.mux_l3_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 9292 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8556 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 8924 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_83
timestamp 1586364061
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_87
timestamp 1586364061
transform 1 0 9108 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_91
timestamp 1586364061
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_23.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 11224 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_102
timestamp 1586364061
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_106
timestamp 1586364061
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_2  _53_
timestamp 1586364061
transform 1 0 13708 0 -1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 13156 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 13524 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_129
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_133
timestamp 1586364061
transform 1 0 13340 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_2  _49_
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 14260 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__67__A
timestamp 1586364061
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_141
timestamp 1586364061
transform 1 0 14076 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_145
timestamp 1586364061
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_149
timestamp 1586364061
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_158
timestamp 1586364061
transform 1 0 15640 0 -1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_21.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 16376 0 -1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 15824 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 16192 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_162
timestamp 1586364061
transform 1 0 16008 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18308 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_185
timestamp 1586364061
transform 1 0 18124 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_8_189
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_8_197
timestamp 1586364061
transform 1 0 19228 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_2  _78_
timestamp 1586364061
transform 1 0 19412 0 -1 7072
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_203
timestamp 1586364061
transform 1 0 19780 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_211
timestamp 1586364061
transform 1 0 20516 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_215
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_227
timestamp 1586364061
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_239
timestamp 1586364061
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_251
timestamp 1586364061
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_263
timestamp 1586364061
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use scs8hd_conb_1  _43_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 2392 0 1 7072
box -38 -48 1786 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1586364061
transform 1 0 2208 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_6
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_10
timestamp 1586364061
transform 1 0 2024 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_33
timestamp 1586364061
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_37
timestamp 1586364061
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l2_in_0_
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_41
timestamp 1586364061
transform 1 0 4876 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_1.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7636 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7084 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_62
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_67
timestamp 1586364061
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _62_
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__62__A
timestamp 1586364061
transform 1 0 9752 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 8648 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_80
timestamp 1586364061
transform 1 0 8464 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_84
timestamp 1586364061
transform 1 0 8832 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_92
timestamp 1586364061
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_96
timestamp 1586364061
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_23.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10672 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10488 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_25.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12052 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_100
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_113
timestamp 1586364061
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_117
timestamp 1586364061
transform 1 0 11868 0 1 7072
box -38 -48 222 592
use scs8hd_buf_2  _55_
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use scs8hd_mux2_2  mux_bottom_track_19.mux_l1_in_0_
timestamp 1586364061
transform 1 0 13708 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_121
timestamp 1586364061
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use scs8hd_decap_4  FILLER_9_127
timestamp 1586364061
transform 1 0 12788 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_133
timestamp 1586364061
transform 1 0 13340 0 1 7072
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_21.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_21.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_146
timestamp 1586364061
transform 1 0 14536 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_152
timestamp 1586364061
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_175
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 590 592
use scs8hd_dfxbp_1  mem_bottom_track_23.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_203
timestamp 1586364061
transform 1 0 19780 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  FILLER_9_217
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 314 592
use scs8hd_buf_4  mux_bottom_track_29.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 21344 0 1 7072
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 22080 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_226
timestamp 1586364061
transform 1 0 21896 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_230
timestamp 1586364061
transform 1 0 22264 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_242
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_257
timestamp 1586364061
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_269
timestamp 1586364061
transform 1 0 25852 0 1 7072
box -38 -48 774 592
use scs8hd_conb_1  _28_
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l1_in_2_
timestamp 1586364061
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_6
timestamp 1586364061
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_10
timestamp 1586364061
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_23
timestamp 1586364061
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_27
timestamp 1586364061
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 5888 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_41
timestamp 1586364061
transform 1 0 4876 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_45
timestamp 1586364061
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_49
timestamp 1586364061
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use scs8hd_buf_2  _63_
timestamp 1586364061
transform 1 0 8372 0 -1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8188 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_71
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_75
timestamp 1586364061
transform 1 0 8004 0 -1 8160
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_29.mux_l2_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 9292 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 8924 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_83
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_87
timestamp 1586364061
transform 1 0 9108 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_25.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 11500 0 -1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11316 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 10672 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_102
timestamp 1586364061
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_106
timestamp 1586364061
transform 1 0 10856 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_110
timestamp 1586364061
transform 1 0 11224 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 13708 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_132
timestamp 1586364061
transform 1 0 13248 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_136
timestamp 1586364061
transform 1 0 13616 0 -1 8160
box -38 -48 130 592
use scs8hd_conb_1  _27_
timestamp 1586364061
transform 1 0 13984 0 -1 8160
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_19.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__55__A
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_10_139
timestamp 1586364061
transform 1 0 13892 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_10_143
timestamp 1586364061
transform 1 0 14260 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_147
timestamp 1586364061
transform 1 0 14628 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_8  FILLER_10_173
timestamp 1586364061
transform 1 0 17020 0 -1 8160
box -38 -48 774 592
use scs8hd_buf_4  mux_bottom_track_19.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18308 0 -1 8160
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_23.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 18032 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_181
timestamp 1586364061
transform 1 0 17756 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_1  FILLER_10_186
timestamp 1586364061
transform 1 0 18216 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_193
timestamp 1586364061
transform 1 0 18860 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_4  mux_bottom_track_27.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_205
timestamp 1586364061
transform 1 0 19964 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_213
timestamp 1586364061
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_221
timestamp 1586364061
transform 1 0 21436 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_233
timestamp 1586364061
transform 1 0 22540 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_245
timestamp 1586364061
transform 1 0 23644 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_257
timestamp 1586364061
transform 1 0 24748 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_6  FILLER_10_269
timestamp 1586364061
transform 1 0 25852 0 -1 8160
box -38 -48 590 592
use scs8hd_fill_1  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l2_in_1_
timestamp 1586364061
transform 1 0 1656 0 1 8160
box -38 -48 866 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2668 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_3
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_15
timestamp 1586364061
transform 1 0 2484 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_19
timestamp 1586364061
transform 1 0 2852 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_5.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 3220 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_5.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use scs8hd_conb_1  _31_
timestamp 1586364061
transform 1 0 5704 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 5152 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__64__A
timestamp 1586364061
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_42
timestamp 1586364061
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_46
timestamp 1586364061
transform 1 0 5336 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_53
timestamp 1586364061
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_57
timestamp 1586364061
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_27.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_29.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 9292 0 1 8160
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_29.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 8740 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_81
timestamp 1586364061
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_85
timestamp 1586364061
transform 1 0 8924 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 11316 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_108
timestamp 1586364061
transform 1 0 11040 0 1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_11_113
timestamp 1586364061
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_117
timestamp 1586364061
transform 1 0 11868 0 1 8160
box -38 -48 314 592
use scs8hd_buf_2  _50_
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_19.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 13708 0 1 8160
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__50__A
timestamp 1586364061
transform 1 0 12972 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_127
timestamp 1586364061
transform 1 0 12788 0 1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_11_131
timestamp 1586364061
transform 1 0 13156 0 1 8160
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 15640 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_156
timestamp 1586364061
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use scs8hd_conb_1  _25_
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 16008 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_19.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 16652 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_160
timestamp 1586364061
transform 1 0 15824 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_167
timestamp 1586364061
transform 1 0 16468 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_171
timestamp 1586364061
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__80__A
timestamp 1586364061
transform 1 0 18308 0 1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_11_189
timestamp 1586364061
transform 1 0 18492 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_201
timestamp 1586364061
transform 1 0 19596 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_213
timestamp 1586364061
transform 1 0 20700 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_225
timestamp 1586364061
transform 1 0 21804 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_11_237
timestamp 1586364061
transform 1 0 22908 0 1 8160
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_11_243
timestamp 1586364061
transform 1 0 23460 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_bottom_track_7.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 1472 0 -1 9248
box -38 -48 1786 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_1  FILLER_12_3
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_7.mux_l1_in_1_
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_23
timestamp 1586364061
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_27
timestamp 1586364061
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use scs8hd_buf_2  _64_
timestamp 1586364061
transform 1 0 5612 0 -1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5060 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 5428 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_41
timestamp 1586364061
transform 1 0 4876 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_45
timestamp 1586364061
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_4  FILLER_12_53
timestamp 1586364061
transform 1 0 5980 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_57
timestamp 1586364061
transform 1 0 6348 0 -1 9248
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_27.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 7084 0 -1 9248
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_27.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_60
timestamp 1586364061
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_1  FILLER_12_64
timestamp 1586364061
transform 1 0 6992 0 -1 9248
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_29.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_84
timestamp 1586364061
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_88
timestamp 1586364061
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l1_in_0_
timestamp 1586364061
transform 1 0 11316 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 11132 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_12_102
timestamp 1586364061
transform 1 0 10488 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_107
timestamp 1586364061
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_17.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12880 0 -1 9248
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 12696 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 12328 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_120
timestamp 1586364061
transform 1 0 12144 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_124
timestamp 1586364061
transform 1 0 12512 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_137
timestamp 1586364061
transform 1 0 13708 0 -1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_19.mux_l2_in_0_
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_19.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 13892 0 -1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 14260 0 -1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_8  FILLER_12_145
timestamp 1586364061
transform 1 0 14444 0 -1 9248
box -38 -48 774 592
use scs8hd_conb_1  _41_
timestamp 1586364061
transform 1 0 16836 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_8  FILLER_12_163
timestamp 1586364061
transform 1 0 16100 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_12_174
timestamp 1586364061
transform 1 0 17112 0 -1 9248
box -38 -48 1142 592
use scs8hd_buf_2  _80_
timestamp 1586364061
transform 1 0 18308 0 -1 9248
box -38 -48 406 592
use scs8hd_fill_1  FILLER_12_186
timestamp 1586364061
transform 1 0 18216 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_191
timestamp 1586364061
transform 1 0 18676 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_203
timestamp 1586364061
transform 1 0 19780 0 -1 9248
box -38 -48 774 592
use scs8hd_decap_3  FILLER_12_211
timestamp 1586364061
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_7
timestamp 1586364061
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_7.mux_l1_in_0_
timestamp 1586364061
transform 1 0 1656 0 -1 10336
box -38 -48 866 592
use scs8hd_buf_2  _66_
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_19
timestamp 1586364061
transform 1 0 2852 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_11
timestamp 1586364061
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_2__CLK
timestamp 1586364061
transform 1 0 2668 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_5.mux_l3_in_0_
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_23
timestamp 1586364061
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_13_28
timestamp 1586364061
transform 1 0 3680 0 1 9248
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_24
timestamp 1586364061
transform 1 0 3312 0 1 9248
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_2__D
timestamp 1586364061
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3036 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_31
timestamp 1586364061
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 4140 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l2_in_0_
timestamp 1586364061
transform 1 0 4324 0 1 9248
box -38 -48 866 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4324 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_48
timestamp 1586364061
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_13_48
timestamp 1586364061
transform 1 0 5520 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_44
timestamp 1586364061
transform 1 0 5152 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 5336 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_58
timestamp 1586364061
transform 1 0 6440 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_54
timestamp 1586364061
transform 1 0 6072 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 5704 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 6256 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 5888 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_27.mux_l1_in_0_
timestamp 1586364061
transform 1 0 5888 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_65
timestamp 1586364061
transform 1 0 7084 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_14_61
timestamp 1586364061
transform 1 0 6716 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_66
timestamp 1586364061
transform 1 0 7176 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__60__A
timestamp 1586364061
transform 1 0 7360 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_27.mux_l2_in_0_
timestamp 1586364061
transform 1 0 7452 0 -1 10336
box -38 -48 866 592
use scs8hd_buf_2  _60_
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_78
timestamp 1586364061
transform 1 0 8280 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_70
timestamp 1586364061
transform 1 0 7544 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 7728 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_29.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_29.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 8280 0 1 9248
box -38 -48 1786 592
use scs8hd_decap_4  FILLER_14_86
timestamp 1586364061
transform 1 0 9016 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_14_82
timestamp 1586364061
transform 1 0 8648 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 222 592
use scs8hd_fill_1  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_97
timestamp 1586364061
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_15.mux_l1_in_0_
timestamp 1586364061
transform 1 0 9752 0 -1 10336
box -38 -48 866 592
use scs8hd_fill_2  FILLER_14_108
timestamp 1586364061
transform 1 0 11040 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_14_103
timestamp 1586364061
transform 1 0 10580 0 -1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_101
timestamp 1586364061
transform 1 0 10396 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 10580 0 1 9248
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_25.mux_l1_in_0_
timestamp 1586364061
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use scs8hd_decap_4  FILLER_14_112
timestamp 1586364061
transform 1 0 11408 0 -1 10336
box -38 -48 406 592
use scs8hd_fill_2  FILLER_13_118
timestamp 1586364061
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use scs8hd_fill_2  FILLER_13_114
timestamp 1586364061
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__63__A
timestamp 1586364061
transform 1 0 11224 0 -1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 11776 0 -1 10336
box -38 -48 1786 592
use scs8hd_dfxbp_1  mem_bottom_track_17.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 12696 0 1 9248
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_17.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 13708 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_14_135
timestamp 1586364061
transform 1 0 13524 0 -1 10336
box -38 -48 222 592
use scs8hd_conb_1  _24_
timestamp 1586364061
transform 1 0 15180 0 1 9248
box -38 -48 314 592
use scs8hd_conb_1  _40_
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_145
timestamp 1586364061
transform 1 0 14444 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_13_156
timestamp 1586364061
transform 1 0 15456 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_139
timestamp 1586364061
transform 1 0 13892 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_14_151
timestamp 1586364061
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_14_157
timestamp 1586364061
transform 1 0 15548 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_168
timestamp 1586364061
transform 1 0 16560 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_169
timestamp 1586364061
transform 1 0 16652 0 -1 10336
box -38 -48 1142 592
use scs8hd_buf_4  mux_bottom_track_15.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 18768 0 1 9248
box -38 -48 222 592
use scs8hd_decap_3  FILLER_13_180
timestamp 1586364061
transform 1 0 17664 0 1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_13_190
timestamp 1586364061
transform 1 0 18584 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_194
timestamp 1586364061
transform 1 0 18952 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_181
timestamp 1586364061
transform 1 0 17756 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_193
timestamp 1586364061
transform 1 0 18860 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_206
timestamp 1586364061
transform 1 0 20056 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_218
timestamp 1586364061
transform 1 0 21160 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_14_205
timestamp 1586364061
transform 1 0 19964 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_213
timestamp 1586364061
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_230
timestamp 1586364061
transform 1 0 22264 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_242
timestamp 1586364061
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_8  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_7.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 1748 0 1 10336
box -38 -48 1786 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__66__A
timestamp 1586364061
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 4232 0 1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA__61__A
timestamp 1586364061
transform 1 0 4048 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 3680 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_26
timestamp 1586364061
transform 1 0 3496 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_30
timestamp 1586364061
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_53
timestamp 1586364061
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use scs8hd_fill_2  FILLER_15_57
timestamp 1586364061
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_11.mux_l2_in_0_
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 8004 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_71
timestamp 1586364061
transform 1 0 7636 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  FILLER_15_77
timestamp 1586364061
transform 1 0 8188 0 1 10336
box -38 -48 314 592
use scs8hd_dfxbp_1  mem_bottom_track_13.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 8648 0 1 10336
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use scs8hd_conb_1  _38_
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 10856 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use scs8hd_decap_4  FILLER_15_101
timestamp 1586364061
transform 1 0 10396 0 1 10336
box -38 -48 406 592
use scs8hd_fill_1  FILLER_15_105
timestamp 1586364061
transform 1 0 10764 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_108
timestamp 1586364061
transform 1 0 11040 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_113
timestamp 1586364061
transform 1 0 11500 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_118
timestamp 1586364061
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_15.mux_l2_in_0_
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_132
timestamp 1586364061
transform 1 0 13248 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_144
timestamp 1586364061
transform 1 0 14352 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_156
timestamp 1586364061
transform 1 0 15456 0 1 10336
box -38 -48 774 592
use scs8hd_buf_4  mux_bottom_track_13.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16652 0 1 10336
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use scs8hd_decap_3  FILLER_15_166
timestamp 1586364061
transform 1 0 16376 0 1 10336
box -38 -48 314 592
use scs8hd_fill_2  FILLER_15_175
timestamp 1586364061
transform 1 0 17204 0 1 10336
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_15_179
timestamp 1586364061
transform 1 0 17572 0 1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use scs8hd_decap_8  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 774 592
use scs8hd_dfxbp_1  mem_bottom_track_7.scs8hd_dfxbp_1_2_
timestamp 1586364061
transform 1 0 1472 0 -1 11424
box -38 -48 1786 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_fill_1  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 130 592
use scs8hd_buf_2  _61_
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_7.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_23
timestamp 1586364061
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_36
timestamp 1586364061
transform 1 0 4416 0 -1 11424
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_11.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 5336 0 -1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 4876 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_16_40
timestamp 1586364061
transform 1 0 4784 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_43
timestamp 1586364061
transform 1 0 5060 0 -1 11424
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_13.mux_l2_in_0_
timestamp 1586364061
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_65
timestamp 1586364061
transform 1 0 7084 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_69
timestamp 1586364061
transform 1 0 7452 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  FILLER_16_72
timestamp 1586364061
transform 1 0 7728 0 -1 11424
box -38 -48 314 592
use scs8hd_conb_1  _37_
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9016 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_27.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 10120 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_84
timestamp 1586364061
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_88
timestamp 1586364061
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_96
timestamp 1586364061
transform 1 0 9936 0 -1 11424
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_15.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 10856 0 -1 11424
box -38 -48 1786 592
use scs8hd_decap_6  FILLER_16_100
timestamp 1586364061
transform 1 0 10304 0 -1 11424
box -38 -48 590 592
use scs8hd_conb_1  _39_
timestamp 1586364061
transform 1 0 13340 0 -1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_15.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_16_125
timestamp 1586364061
transform 1 0 12604 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_136
timestamp 1586364061
transform 1 0 13616 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_148
timestamp 1586364061
transform 1 0 14720 0 -1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_16_152
timestamp 1586364061
transform 1 0 15088 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 774 592
use scs8hd_buf_4  mux_bottom_track_11.scs8hd_buf_4_0_
timestamp 1586364061
transform 1 0 16192 0 -1 11424
box -38 -48 590 592
use scs8hd_fill_2  FILLER_16_162
timestamp 1586364061
transform 1 0 16008 0 -1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_16_170
timestamp 1586364061
transform 1 0 16744 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_182
timestamp 1586364061
transform 1 0 17848 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_194
timestamp 1586364061
transform 1 0 18952 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_206
timestamp 1586364061
transform 1 0 20056 0 -1 11424
box -38 -48 774 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_7.mux_l2_in_1_
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 866 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 2392 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_12
timestamp 1586364061
transform 1 0 2208 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_16
timestamp 1586364061
transform 1 0 2576 0 1 11424
box -38 -48 406 592
use scs8hd_dfxbp_1  mem_bottom_track_9.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 3220 0 1 11424
box -38 -48 1786 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 3036 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_20
timestamp 1586364061
transform 1 0 2944 0 1 11424
box -38 -48 130 592
use scs8hd_conb_1  _30_
timestamp 1586364061
transform 1 0 5704 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 5152 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_1__CLK
timestamp 1586364061
transform 1 0 6440 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_42
timestamp 1586364061
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_46
timestamp 1586364061
transform 1 0 5336 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_53
timestamp 1586364061
transform 1 0 5980 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_57
timestamp 1586364061
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use scs8hd_dfxbp_1  mem_bottom_track_13.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 7544 0 1 11424
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_13.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 7360 0 1 11424
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_11.scs8hd_dfxbp_1_1__D
timestamp 1586364061
transform 1 0 6992 0 1 11424
box -38 -48 222 592
use scs8hd_fill_1  FILLER_17_60
timestamp 1586364061
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_66
timestamp 1586364061
transform 1 0 7176 0 1 11424
box -38 -48 222 592
use scs8hd_conb_1  _44_
timestamp 1586364061
transform 1 0 10028 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_0__CLK
timestamp 1586364061
transform 1 0 9752 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_89
timestamp 1586364061
transform 1 0 9292 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_93
timestamp 1586364061
transform 1 0 9660 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_96
timestamp 1586364061
transform 1 0 9936 0 1 11424
box -38 -48 130 592
use scs8hd_conb_1  _42_
timestamp 1586364061
transform 1 0 11132 0 1 11424
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_15.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 10488 0 1 11424
box -38 -48 222 592
use scs8hd_fill_2  FILLER_17_100
timestamp 1586364061
transform 1 0 10304 0 1 11424
box -38 -48 222 592
use scs8hd_decap_4  FILLER_17_104
timestamp 1586364061
transform 1 0 10672 0 1 11424
box -38 -48 406 592
use scs8hd_fill_1  FILLER_17_108
timestamp 1586364061
transform 1 0 11040 0 1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_17_112
timestamp 1586364061
transform 1 0 11408 0 1 11424
box -38 -48 774 592
use scs8hd_conb_1  _47_
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_120
timestamp 1586364061
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_126
timestamp 1586364061
transform 1 0 12696 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_138
timestamp 1586364061
transform 1 0 13800 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_150
timestamp 1586364061
transform 1 0 14904 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_162
timestamp 1586364061
transform 1 0 16008 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_174
timestamp 1586364061
transform 1 0 17112 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_fill_1  FILLER_17_182
timestamp 1586364061
transform 1 0 17848 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use scs8hd_decap_8  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 774 592
use scs8hd_mux2_2  mux_bottom_track_7.mux_l2_in_0_
timestamp 1586364061
transform 1 0 1472 0 -1 12512
box -38 -48 866 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__A0
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_1__S
timestamp 1586364061
transform 1 0 2852 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_13
timestamp 1586364061
transform 1 0 2300 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_17
timestamp 1586364061
transform 1 0 2668 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_21
timestamp 1586364061
transform 1 0 3036 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_25
timestamp 1586364061
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_track_9.scs8hd_dfxbp_1_0__D
timestamp 1586364061
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_29
timestamp 1586364061
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__S
timestamp 1586364061
transform 1 0 4232 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_18_36
timestamp 1586364061
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use scs8hd_dfxbp_1  mem_bottom_track_11.scs8hd_dfxbp_1_1_
timestamp 1586364061
transform 1 0 6440 0 -1 12512
box -38 -48 1786 592
use scs8hd_mux2_2  mux_bottom_track_11.mux_l1_in_0_
timestamp 1586364061
transform 1 0 4876 0 -1 12512
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 5888 0 -1 12512
box -38 -48 222 592
use scs8hd_fill_1  FILLER_18_40
timestamp 1586364061
transform 1 0 4784 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_18_50
timestamp 1586364061
transform 1 0 5704 0 -1 12512
box -38 -48 222 592
use scs8hd_decap_4  FILLER_18_54
timestamp 1586364061
transform 1 0 6072 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_77
timestamp 1586364061
transform 1 0 8188 0 -1 12512
box -38 -48 1142 592
use scs8hd_dfxbp_1  mem_bottom_track_15.scs8hd_dfxbp_1_0_
timestamp 1586364061
transform 1 0 9752 0 -1 12512
box -38 -48 1786 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  FILLER_18_89
timestamp 1586364061
transform 1 0 9292 0 -1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_113
timestamp 1586364061
transform 1 0 11500 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_125
timestamp 1586364061
transform 1 0 12604 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_137
timestamp 1586364061
transform 1 0 13708 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_149
timestamp 1586364061
transform 1 0 14812 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use scs8hd_fill_2  FILLER_20_7
timestamp 1586364061
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__59__A
timestamp 1586364061
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_mux2_2  mux_bottom_track_7.mux_l3_in_0_
timestamp 1586364061
transform 1 0 1564 0 1 12512
box -38 -48 866 592
use scs8hd_buf_2  _59_
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_2  FILLER_20_19
timestamp 1586364061
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_11
timestamp 1586364061
transform 1 0 2116 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_18
timestamp 1586364061
transform 1 0 2760 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_14
timestamp 1586364061
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__S
timestamp 1586364061
transform 1 0 2300 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__56__A
timestamp 1586364061
transform 1 0 2576 0 1 12512
box -38 -48 222 592
use scs8hd_buf_2  _56_
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__S
timestamp 1586364061
transform 1 0 2944 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_22
timestamp 1586364061
transform 1 0 3128 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0
timestamp 1586364061
transform 1 0 3312 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A1
timestamp 1586364061
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_23
timestamp 1586364061
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1
timestamp 1586364061
transform 1 0 3680 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_26
timestamp 1586364061
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_5.scs8hd_buf_4_0__A
timestamp 1586364061
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 4232 0 -1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_mux2_2  mux_bottom_track_9.mux_l1_in_1_
timestamp 1586364061
transform 1 0 3864 0 1 12512
box -38 -48 866 592
use scs8hd_decap_12  FILLER_20_36
timestamp 1586364061
transform 1 0 4416 0 -1 13600
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 4876 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_43
timestamp 1586364061
transform 1 0 5060 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_19_55
timestamp 1586364061
transform 1 0 6164 0 1 12512
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_48
timestamp 1586364061
transform 1 0 5520 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_19_69
timestamp 1586364061
transform 1 0 7452 0 1 12512
box -38 -48 222 592
use scs8hd_fill_2  FILLER_19_65
timestamp 1586364061
transform 1 0 7084 0 1 12512
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__S
timestamp 1586364061
transform 1 0 7268 0 1 12512
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_conb_1  _36_
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use scs8hd_fill_1  FILLER_20_72
timestamp 1586364061
transform 1 0 7728 0 -1 13600
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A0
timestamp 1586364061
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1586364061
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use scs8hd_mux2_2  mux_bottom_track_13.mux_l1_in_0_
timestamp 1586364061
transform 1 0 7820 0 1 12512
box -38 -48 866 592
use scs8hd_decap_12  FILLER_20_75
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_60
timestamp 1586364061
transform 1 0 6624 0 -1 13600
box -38 -48 1142 592
use scs8hd_conb_1  _45_
timestamp 1586364061
transform 1 0 9384 0 1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_82
timestamp 1586364061
transform 1 0 8648 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_19_93
timestamp 1586364061
transform 1 0 9660 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 406 592
use scs8hd_fill_1  FILLER_20_91
timestamp 1586364061
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_20_93
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_105
timestamp 1586364061
transform 1 0 10764 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_19_117
timestamp 1586364061
transform 1 0 11868 0 1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_105
timestamp 1586364061
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_117
timestamp 1586364061
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_fill_1  FILLER_19_121
timestamp 1586364061
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_129
timestamp 1586364061
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_141
timestamp 1586364061
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_154
timestamp 1586364061
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_166
timestamp 1586364061
transform 1 0 16376 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_178
timestamp 1586364061
transform 1 0 17480 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_190
timestamp 1586364061
transform 1 0 18584 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_202
timestamp 1586364061
transform 1 0 19688 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_215
timestamp 1586364061
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_227
timestamp 1586364061
transform 1 0 21988 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_239
timestamp 1586364061
transform 1 0 23092 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_251
timestamp 1586364061
transform 1 0 24196 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_8  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_263
timestamp 1586364061
transform 1 0 25300 0 -1 13600
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_20_276
timestamp 1586364061
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use scs8hd_buf_2  _57_
timestamp 1586364061
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use scs8hd_decap_3  PHY_42
timestamp 1586364061
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__57__A
timestamp 1586364061
transform 1 0 1932 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1586364061
transform 1 0 2300 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_7
timestamp 1586364061
transform 1 0 1748 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_11
timestamp 1586364061
transform 1 0 2116 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_15
timestamp 1586364061
transform 1 0 2484 0 1 13600
box -38 -48 222 592
use scs8hd_fill_2  FILLER_21_19
timestamp 1586364061
transform 1 0 2852 0 1 13600
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l3_in_0__A0
timestamp 1586364061
transform 1 0 3036 0 1 13600
box -38 -48 222 592
use scs8hd_decap_12  FILLER_21_23
timestamp 1586364061
transform 1 0 3220 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_35
timestamp 1586364061
transform 1 0 4324 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_47
timestamp 1586364061
transform 1 0 5428 0 1 13600
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_21_59
timestamp 1586364061
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_62
timestamp 1586364061
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_74
timestamp 1586364061
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_86
timestamp 1586364061
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_98
timestamp 1586364061
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_110
timestamp 1586364061
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_123
timestamp 1586364061
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_135
timestamp 1586364061
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_147
timestamp 1586364061
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_159
timestamp 1586364061
transform 1 0 15732 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_171
timestamp 1586364061
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_184
timestamp 1586364061
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_196
timestamp 1586364061
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_208
timestamp 1586364061
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_220
timestamp 1586364061
transform 1 0 21344 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_232
timestamp 1586364061
transform 1 0 22448 0 1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_21_245
timestamp 1586364061
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_21_257
timestamp 1586364061
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_43
timestamp 1586364061
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use scs8hd_decap_8  FILLER_21_269
timestamp 1586364061
transform 1 0 25852 0 1 13600
box -38 -48 774 592
use scs8hd_conb_1  _29_
timestamp 1586364061
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use scs8hd_decap_3  PHY_44
timestamp 1586364061
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A1
timestamp 1586364061
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_track_7.mux_l2_in_0__A0
timestamp 1586364061
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_6
timestamp 1586364061
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use scs8hd_fill_2  FILLER_22_10
timestamp 1586364061
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use scs8hd_decap_12  FILLER_22_14
timestamp 1586364061
transform 1 0 2392 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_4  FILLER_22_26
timestamp 1586364061
transform 1 0 3496 0 -1 14688
box -38 -48 406 592
use scs8hd_fill_1  FILLER_22_30
timestamp 1586364061
transform 1 0 3864 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_32
timestamp 1586364061
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_44
timestamp 1586364061
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_56
timestamp 1586364061
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_68
timestamp 1586364061
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_80
timestamp 1586364061
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_93
timestamp 1586364061
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_105
timestamp 1586364061
transform 1 0 10764 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_117
timestamp 1586364061
transform 1 0 11868 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_129
timestamp 1586364061
transform 1 0 12972 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_141
timestamp 1586364061
transform 1 0 14076 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_154
timestamp 1586364061
transform 1 0 15272 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_166
timestamp 1586364061
transform 1 0 16376 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_178
timestamp 1586364061
transform 1 0 17480 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_190
timestamp 1586364061
transform 1 0 18584 0 -1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_191
timestamp 1586364061
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_202
timestamp 1586364061
transform 1 0 19688 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_215
timestamp 1586364061
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_227
timestamp 1586364061
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_239
timestamp 1586364061
transform 1 0 23092 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_22_251
timestamp 1586364061
transform 1 0 24196 0 -1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_45
timestamp 1586364061
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_192
timestamp 1586364061
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_22_263
timestamp 1586364061
transform 1 0 25300 0 -1 14688
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_22_276
timestamp 1586364061
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use scs8hd_decap_3  PHY_46
timestamp 1586364061
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use scs8hd_decap_12  FILLER_23_3
timestamp 1586364061
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_15
timestamp 1586364061
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_27
timestamp 1586364061
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_39
timestamp 1586364061
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_23_51
timestamp 1586364061
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use scs8hd_fill_2  FILLER_23_59
timestamp 1586364061
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_193
timestamp 1586364061
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_62
timestamp 1586364061
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_74
timestamp 1586364061
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_86
timestamp 1586364061
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_98
timestamp 1586364061
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_110
timestamp 1586364061
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_194
timestamp 1586364061
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_123
timestamp 1586364061
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_135
timestamp 1586364061
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_147
timestamp 1586364061
transform 1 0 14628 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_159
timestamp 1586364061
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_171
timestamp 1586364061
transform 1 0 16836 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_195
timestamp 1586364061
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_184
timestamp 1586364061
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_196
timestamp 1586364061
transform 1 0 19136 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_208
timestamp 1586364061
transform 1 0 20240 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_220
timestamp 1586364061
transform 1 0 21344 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_232
timestamp 1586364061
transform 1 0 22448 0 1 14688
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_196
timestamp 1586364061
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use scs8hd_decap_12  FILLER_23_245
timestamp 1586364061
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_23_257
timestamp 1586364061
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use scs8hd_decap_3  PHY_47
timestamp 1586364061
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use scs8hd_decap_8  FILLER_23_269
timestamp 1586364061
transform 1 0 25852 0 1 14688
box -38 -48 774 592
use scs8hd_decap_3  PHY_48
timestamp 1586364061
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_24_3
timestamp 1586364061
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_15
timestamp 1586364061
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_197
timestamp 1586364061
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_4  FILLER_24_27
timestamp 1586364061
transform 1 0 3588 0 -1 15776
box -38 -48 406 592
use scs8hd_decap_12  FILLER_24_32
timestamp 1586364061
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_44
timestamp 1586364061
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_56
timestamp 1586364061
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_68
timestamp 1586364061
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_198
timestamp 1586364061
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_80
timestamp 1586364061
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_93
timestamp 1586364061
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_105
timestamp 1586364061
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_117
timestamp 1586364061
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_129
timestamp 1586364061
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_199
timestamp 1586364061
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_141
timestamp 1586364061
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_154
timestamp 1586364061
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_166
timestamp 1586364061
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_178
timestamp 1586364061
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_190
timestamp 1586364061
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_200
timestamp 1586364061
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_202
timestamp 1586364061
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_215
timestamp 1586364061
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_227
timestamp 1586364061
transform 1 0 21988 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_239
timestamp 1586364061
transform 1 0 23092 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_24_251
timestamp 1586364061
transform 1 0 24196 0 -1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_49
timestamp 1586364061
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_201
timestamp 1586364061
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_24_263
timestamp 1586364061
transform 1 0 25300 0 -1 15776
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_24_276
timestamp 1586364061
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use scs8hd_decap_3  PHY_50
timestamp 1586364061
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use scs8hd_decap_12  FILLER_25_3
timestamp 1586364061
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_15
timestamp 1586364061
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_27
timestamp 1586364061
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_39
timestamp 1586364061
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_25_51
timestamp 1586364061
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use scs8hd_fill_2  FILLER_25_59
timestamp 1586364061
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_202
timestamp 1586364061
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_62
timestamp 1586364061
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_74
timestamp 1586364061
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_86
timestamp 1586364061
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_98
timestamp 1586364061
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_110
timestamp 1586364061
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_203
timestamp 1586364061
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_123
timestamp 1586364061
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_135
timestamp 1586364061
transform 1 0 13524 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_147
timestamp 1586364061
transform 1 0 14628 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_159
timestamp 1586364061
transform 1 0 15732 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_171
timestamp 1586364061
transform 1 0 16836 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_204
timestamp 1586364061
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_184
timestamp 1586364061
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_196
timestamp 1586364061
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_208
timestamp 1586364061
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_220
timestamp 1586364061
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_232
timestamp 1586364061
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_205
timestamp 1586364061
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use scs8hd_decap_12  FILLER_25_245
timestamp 1586364061
transform 1 0 23644 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_25_257
timestamp 1586364061
transform 1 0 24748 0 1 15776
box -38 -48 1142 592
use scs8hd_decap_3  PHY_51
timestamp 1586364061
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use scs8hd_decap_8  FILLER_25_269
timestamp 1586364061
transform 1 0 25852 0 1 15776
box -38 -48 774 592
use scs8hd_decap_3  PHY_52
timestamp 1586364061
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_54
timestamp 1586364061
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use scs8hd_decap_12  FILLER_26_3
timestamp 1586364061
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_15
timestamp 1586364061
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_3
timestamp 1586364061
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_15
timestamp 1586364061
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_206
timestamp 1586364061
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_4  FILLER_26_27
timestamp 1586364061
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use scs8hd_decap_12  FILLER_26_32
timestamp 1586364061
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_27
timestamp 1586364061
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_39
timestamp 1586364061
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_44
timestamp 1586364061
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_56
timestamp 1586364061
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_27_51
timestamp 1586364061
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use scs8hd_fill_2  FILLER_27_59
timestamp 1586364061
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_211
timestamp 1586364061
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_68
timestamp 1586364061
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_62
timestamp 1586364061
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_74
timestamp 1586364061
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_207
timestamp 1586364061
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_80
timestamp 1586364061
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_93
timestamp 1586364061
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_86
timestamp 1586364061
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_98
timestamp 1586364061
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_105
timestamp 1586364061
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_117
timestamp 1586364061
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_110
timestamp 1586364061
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_212
timestamp 1586364061
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_129
timestamp 1586364061
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_123
timestamp 1586364061
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_135
timestamp 1586364061
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_208
timestamp 1586364061
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_141
timestamp 1586364061
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_154
timestamp 1586364061
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_147
timestamp 1586364061
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_166
timestamp 1586364061
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_178
timestamp 1586364061
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_159
timestamp 1586364061
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_171
timestamp 1586364061
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_213
timestamp 1586364061
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_190
timestamp 1586364061
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_184
timestamp 1586364061
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_196
timestamp 1586364061
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_209
timestamp 1586364061
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_202
timestamp 1586364061
transform 1 0 19688 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_215
timestamp 1586364061
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_208
timestamp 1586364061
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_227
timestamp 1586364061
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_220
timestamp 1586364061
transform 1 0 21344 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_232
timestamp 1586364061
transform 1 0 22448 0 1 16864
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_214
timestamp 1586364061
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_239
timestamp 1586364061
transform 1 0 23092 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_26_251
timestamp 1586364061
transform 1 0 24196 0 -1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_245
timestamp 1586364061
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_27_257
timestamp 1586364061
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use scs8hd_decap_3  PHY_53
timestamp 1586364061
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use scs8hd_decap_3  PHY_55
timestamp 1586364061
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_210
timestamp 1586364061
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_12  FILLER_26_263
timestamp 1586364061
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_26_276
timestamp 1586364061
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use scs8hd_decap_8  FILLER_27_269
timestamp 1586364061
transform 1 0 25852 0 1 16864
box -38 -48 774 592
use scs8hd_decap_3  PHY_56
timestamp 1586364061
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_28_3
timestamp 1586364061
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_15
timestamp 1586364061
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_215
timestamp 1586364061
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_4  FILLER_28_27
timestamp 1586364061
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use scs8hd_decap_12  FILLER_28_32
timestamp 1586364061
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_44
timestamp 1586364061
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_56
timestamp 1586364061
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_68
timestamp 1586364061
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_216
timestamp 1586364061
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_80
timestamp 1586364061
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_93
timestamp 1586364061
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_105
timestamp 1586364061
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_117
timestamp 1586364061
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_129
timestamp 1586364061
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_217
timestamp 1586364061
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_141
timestamp 1586364061
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_154
timestamp 1586364061
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_166
timestamp 1586364061
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_178
timestamp 1586364061
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_190
timestamp 1586364061
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_218
timestamp 1586364061
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_202
timestamp 1586364061
transform 1 0 19688 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_215
timestamp 1586364061
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_227
timestamp 1586364061
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_239
timestamp 1586364061
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_28_251
timestamp 1586364061
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_57
timestamp 1586364061
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_219
timestamp 1586364061
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_28_263
timestamp 1586364061
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_28_276
timestamp 1586364061
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use scs8hd_decap_3  PHY_58
timestamp 1586364061
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use scs8hd_decap_12  FILLER_29_3
timestamp 1586364061
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_15
timestamp 1586364061
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_27
timestamp 1586364061
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_39
timestamp 1586364061
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_29_51
timestamp 1586364061
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use scs8hd_fill_2  FILLER_29_59
timestamp 1586364061
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_220
timestamp 1586364061
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_62
timestamp 1586364061
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_74
timestamp 1586364061
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_86
timestamp 1586364061
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_98
timestamp 1586364061
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_110
timestamp 1586364061
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_221
timestamp 1586364061
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_123
timestamp 1586364061
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_135
timestamp 1586364061
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_147
timestamp 1586364061
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_159
timestamp 1586364061
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_171
timestamp 1586364061
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_222
timestamp 1586364061
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_184
timestamp 1586364061
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_196
timestamp 1586364061
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_208
timestamp 1586364061
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_220
timestamp 1586364061
transform 1 0 21344 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_232
timestamp 1586364061
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_223
timestamp 1586364061
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use scs8hd_decap_12  FILLER_29_245
timestamp 1586364061
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_29_257
timestamp 1586364061
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use scs8hd_decap_3  PHY_59
timestamp 1586364061
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use scs8hd_decap_8  FILLER_29_269
timestamp 1586364061
transform 1 0 25852 0 1 17952
box -38 -48 774 592
use scs8hd_decap_3  PHY_60
timestamp 1586364061
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_30_3
timestamp 1586364061
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_15
timestamp 1586364061
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_224
timestamp 1586364061
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_4  FILLER_30_27
timestamp 1586364061
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use scs8hd_decap_12  FILLER_30_32
timestamp 1586364061
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_44
timestamp 1586364061
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_56
timestamp 1586364061
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_68
timestamp 1586364061
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_225
timestamp 1586364061
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_80
timestamp 1586364061
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_93
timestamp 1586364061
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_105
timestamp 1586364061
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_117
timestamp 1586364061
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_129
timestamp 1586364061
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_226
timestamp 1586364061
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_141
timestamp 1586364061
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_154
timestamp 1586364061
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_166
timestamp 1586364061
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_178
timestamp 1586364061
transform 1 0 17480 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_190
timestamp 1586364061
transform 1 0 18584 0 -1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_227
timestamp 1586364061
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_202
timestamp 1586364061
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_215
timestamp 1586364061
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_227
timestamp 1586364061
transform 1 0 21988 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_239
timestamp 1586364061
transform 1 0 23092 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_30_251
timestamp 1586364061
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_61
timestamp 1586364061
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_228
timestamp 1586364061
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_30_263
timestamp 1586364061
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_30_276
timestamp 1586364061
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use scs8hd_decap_3  PHY_62
timestamp 1586364061
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use scs8hd_decap_12  FILLER_31_3
timestamp 1586364061
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_15
timestamp 1586364061
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_27
timestamp 1586364061
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_39
timestamp 1586364061
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_31_51
timestamp 1586364061
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use scs8hd_fill_2  FILLER_31_59
timestamp 1586364061
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_229
timestamp 1586364061
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_62
timestamp 1586364061
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_74
timestamp 1586364061
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_86
timestamp 1586364061
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_98
timestamp 1586364061
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_110
timestamp 1586364061
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_230
timestamp 1586364061
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_123
timestamp 1586364061
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_135
timestamp 1586364061
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_147
timestamp 1586364061
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_159
timestamp 1586364061
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_171
timestamp 1586364061
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_231
timestamp 1586364061
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_184
timestamp 1586364061
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_196
timestamp 1586364061
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_208
timestamp 1586364061
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_220
timestamp 1586364061
transform 1 0 21344 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_232
timestamp 1586364061
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_232
timestamp 1586364061
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use scs8hd_decap_12  FILLER_31_245
timestamp 1586364061
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_31_257
timestamp 1586364061
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use scs8hd_decap_3  PHY_63
timestamp 1586364061
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use scs8hd_decap_8  FILLER_31_269
timestamp 1586364061
transform 1 0 25852 0 1 19040
box -38 -48 774 592
use scs8hd_decap_3  PHY_64
timestamp 1586364061
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use scs8hd_decap_12  FILLER_32_3
timestamp 1586364061
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_15
timestamp 1586364061
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_233
timestamp 1586364061
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_4  FILLER_32_27
timestamp 1586364061
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use scs8hd_decap_12  FILLER_32_32
timestamp 1586364061
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_44
timestamp 1586364061
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_56
timestamp 1586364061
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_68
timestamp 1586364061
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_234
timestamp 1586364061
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_80
timestamp 1586364061
transform 1 0 8464 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_93
timestamp 1586364061
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_105
timestamp 1586364061
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_117
timestamp 1586364061
transform 1 0 11868 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_129
timestamp 1586364061
transform 1 0 12972 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_235
timestamp 1586364061
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_141
timestamp 1586364061
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_154
timestamp 1586364061
transform 1 0 15272 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_166
timestamp 1586364061
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_178
timestamp 1586364061
transform 1 0 17480 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_190
timestamp 1586364061
transform 1 0 18584 0 -1 20128
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_236
timestamp 1586364061
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_202
timestamp 1586364061
transform 1 0 19688 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_215
timestamp 1586364061
transform 1 0 20884 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_227
timestamp 1586364061
transform 1 0 21988 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_239
timestamp 1586364061
transform 1 0 23092 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_32_251
timestamp 1586364061
transform 1 0 24196 0 -1 20128
box -38 -48 1142 592
use scs8hd_decap_3  PHY_65
timestamp 1586364061
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_237
timestamp 1586364061
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_32_263
timestamp 1586364061
transform 1 0 25300 0 -1 20128
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_32_276
timestamp 1586364061
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use scs8hd_decap_3  PHY_66
timestamp 1586364061
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_68
timestamp 1586364061
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_33_3
timestamp 1586364061
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_15
timestamp 1586364061
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_3
timestamp 1586364061
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_15
timestamp 1586364061
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_242
timestamp 1586364061
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_27
timestamp 1586364061
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_39
timestamp 1586364061
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_34_27
timestamp 1586364061
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use scs8hd_decap_12  FILLER_34_32
timestamp 1586364061
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_33_51
timestamp 1586364061
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use scs8hd_fill_2  FILLER_33_59
timestamp 1586364061
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use scs8hd_decap_12  FILLER_34_44
timestamp 1586364061
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_56
timestamp 1586364061
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_238
timestamp 1586364061
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_62
timestamp 1586364061
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_74
timestamp 1586364061
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_68
timestamp 1586364061
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_243
timestamp 1586364061
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_86
timestamp 1586364061
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_98
timestamp 1586364061
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_80
timestamp 1586364061
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_93
timestamp 1586364061
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_110
timestamp 1586364061
transform 1 0 11224 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_105
timestamp 1586364061
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_117
timestamp 1586364061
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_239
timestamp 1586364061
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_123
timestamp 1586364061
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_135
timestamp 1586364061
transform 1 0 13524 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_129
timestamp 1586364061
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_244
timestamp 1586364061
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_147
timestamp 1586364061
transform 1 0 14628 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_141
timestamp 1586364061
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_154
timestamp 1586364061
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_159
timestamp 1586364061
transform 1 0 15732 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_171
timestamp 1586364061
transform 1 0 16836 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_166
timestamp 1586364061
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_178
timestamp 1586364061
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_240
timestamp 1586364061
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_184
timestamp 1586364061
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_196
timestamp 1586364061
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_190
timestamp 1586364061
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_245
timestamp 1586364061
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_208
timestamp 1586364061
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_202
timestamp 1586364061
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_215
timestamp 1586364061
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_220
timestamp 1586364061
transform 1 0 21344 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_232
timestamp 1586364061
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_227
timestamp 1586364061
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_241
timestamp 1586364061
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use scs8hd_decap_12  FILLER_33_245
timestamp 1586364061
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_33_257
timestamp 1586364061
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_239
timestamp 1586364061
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_34_251
timestamp 1586364061
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_67
timestamp 1586364061
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use scs8hd_decap_3  PHY_69
timestamp 1586364061
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_246
timestamp 1586364061
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_8  FILLER_33_269
timestamp 1586364061
transform 1 0 25852 0 1 20128
box -38 -48 774 592
use scs8hd_decap_12  FILLER_34_263
timestamp 1586364061
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_34_276
timestamp 1586364061
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use scs8hd_decap_3  PHY_70
timestamp 1586364061
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use scs8hd_decap_12  FILLER_35_3
timestamp 1586364061
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_15
timestamp 1586364061
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_27
timestamp 1586364061
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_39
timestamp 1586364061
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_35_51
timestamp 1586364061
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use scs8hd_fill_2  FILLER_35_59
timestamp 1586364061
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_247
timestamp 1586364061
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_62
timestamp 1586364061
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_74
timestamp 1586364061
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_86
timestamp 1586364061
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_98
timestamp 1586364061
transform 1 0 10120 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_110
timestamp 1586364061
transform 1 0 11224 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_248
timestamp 1586364061
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_123
timestamp 1586364061
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_135
timestamp 1586364061
transform 1 0 13524 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_147
timestamp 1586364061
transform 1 0 14628 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_159
timestamp 1586364061
transform 1 0 15732 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_171
timestamp 1586364061
transform 1 0 16836 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_249
timestamp 1586364061
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_184
timestamp 1586364061
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_196
timestamp 1586364061
transform 1 0 19136 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_208
timestamp 1586364061
transform 1 0 20240 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_220
timestamp 1586364061
transform 1 0 21344 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_232
timestamp 1586364061
transform 1 0 22448 0 1 21216
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_250
timestamp 1586364061
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use scs8hd_decap_12  FILLER_35_245
timestamp 1586364061
transform 1 0 23644 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_35_257
timestamp 1586364061
transform 1 0 24748 0 1 21216
box -38 -48 1142 592
use scs8hd_decap_3  PHY_71
timestamp 1586364061
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use scs8hd_decap_8  FILLER_35_269
timestamp 1586364061
transform 1 0 25852 0 1 21216
box -38 -48 774 592
use scs8hd_decap_3  PHY_72
timestamp 1586364061
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_36_3
timestamp 1586364061
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_15
timestamp 1586364061
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_251
timestamp 1586364061
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_4  FILLER_36_27
timestamp 1586364061
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use scs8hd_decap_12  FILLER_36_32
timestamp 1586364061
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_44
timestamp 1586364061
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_56
timestamp 1586364061
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_68
timestamp 1586364061
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_252
timestamp 1586364061
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_80
timestamp 1586364061
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_93
timestamp 1586364061
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_105
timestamp 1586364061
transform 1 0 10764 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_117
timestamp 1586364061
transform 1 0 11868 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_129
timestamp 1586364061
transform 1 0 12972 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_253
timestamp 1586364061
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_141
timestamp 1586364061
transform 1 0 14076 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_154
timestamp 1586364061
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_166
timestamp 1586364061
transform 1 0 16376 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_178
timestamp 1586364061
transform 1 0 17480 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_190
timestamp 1586364061
transform 1 0 18584 0 -1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_254
timestamp 1586364061
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_202
timestamp 1586364061
transform 1 0 19688 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_215
timestamp 1586364061
transform 1 0 20884 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_227
timestamp 1586364061
transform 1 0 21988 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_239
timestamp 1586364061
transform 1 0 23092 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_36_251
timestamp 1586364061
transform 1 0 24196 0 -1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_73
timestamp 1586364061
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_255
timestamp 1586364061
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_36_263
timestamp 1586364061
transform 1 0 25300 0 -1 22304
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_36_276
timestamp 1586364061
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use scs8hd_decap_3  PHY_74
timestamp 1586364061
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use scs8hd_decap_12  FILLER_37_3
timestamp 1586364061
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_15
timestamp 1586364061
transform 1 0 2484 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_27
timestamp 1586364061
transform 1 0 3588 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_39
timestamp 1586364061
transform 1 0 4692 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_37_51
timestamp 1586364061
transform 1 0 5796 0 1 22304
box -38 -48 774 592
use scs8hd_fill_2  FILLER_37_59
timestamp 1586364061
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_256
timestamp 1586364061
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_62
timestamp 1586364061
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_74
timestamp 1586364061
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_86
timestamp 1586364061
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_98
timestamp 1586364061
transform 1 0 10120 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_110
timestamp 1586364061
transform 1 0 11224 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_257
timestamp 1586364061
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_123
timestamp 1586364061
transform 1 0 12420 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_135
timestamp 1586364061
transform 1 0 13524 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_147
timestamp 1586364061
transform 1 0 14628 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_159
timestamp 1586364061
transform 1 0 15732 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_171
timestamp 1586364061
transform 1 0 16836 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_258
timestamp 1586364061
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_184
timestamp 1586364061
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_196
timestamp 1586364061
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_208
timestamp 1586364061
transform 1 0 20240 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_220
timestamp 1586364061
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_232
timestamp 1586364061
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_259
timestamp 1586364061
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use scs8hd_decap_12  FILLER_37_245
timestamp 1586364061
transform 1 0 23644 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_37_257
timestamp 1586364061
transform 1 0 24748 0 1 22304
box -38 -48 1142 592
use scs8hd_decap_3  PHY_75
timestamp 1586364061
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use scs8hd_decap_8  FILLER_37_269
timestamp 1586364061
transform 1 0 25852 0 1 22304
box -38 -48 774 592
use scs8hd_decap_3  PHY_76
timestamp 1586364061
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use scs8hd_decap_12  FILLER_38_3
timestamp 1586364061
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_15
timestamp 1586364061
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_260
timestamp 1586364061
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_4  FILLER_38_27
timestamp 1586364061
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use scs8hd_decap_12  FILLER_38_32
timestamp 1586364061
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_44
timestamp 1586364061
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_56
timestamp 1586364061
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_68
timestamp 1586364061
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_261
timestamp 1586364061
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_80
timestamp 1586364061
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_93
timestamp 1586364061
transform 1 0 9660 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_105
timestamp 1586364061
transform 1 0 10764 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_117
timestamp 1586364061
transform 1 0 11868 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_129
timestamp 1586364061
transform 1 0 12972 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_262
timestamp 1586364061
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_141
timestamp 1586364061
transform 1 0 14076 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_154
timestamp 1586364061
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_166
timestamp 1586364061
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_178
timestamp 1586364061
transform 1 0 17480 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_190
timestamp 1586364061
transform 1 0 18584 0 -1 23392
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_263
timestamp 1586364061
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_202
timestamp 1586364061
transform 1 0 19688 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_215
timestamp 1586364061
transform 1 0 20884 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_227
timestamp 1586364061
transform 1 0 21988 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_239
timestamp 1586364061
transform 1 0 23092 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_38_251
timestamp 1586364061
transform 1 0 24196 0 -1 23392
box -38 -48 1142 592
use scs8hd_decap_3  PHY_77
timestamp 1586364061
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_264
timestamp 1586364061
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_38_263
timestamp 1586364061
transform 1 0 25300 0 -1 23392
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_38_276
timestamp 1586364061
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use scs8hd_decap_3  PHY_78
timestamp 1586364061
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_80
timestamp 1586364061
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_39_3
timestamp 1586364061
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_15
timestamp 1586364061
transform 1 0 2484 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_3
timestamp 1586364061
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_15
timestamp 1586364061
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_269
timestamp 1586364061
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_27
timestamp 1586364061
transform 1 0 3588 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_39
timestamp 1586364061
transform 1 0 4692 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_40_27
timestamp 1586364061
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use scs8hd_decap_12  FILLER_40_32
timestamp 1586364061
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_39_51
timestamp 1586364061
transform 1 0 5796 0 1 23392
box -38 -48 774 592
use scs8hd_fill_2  FILLER_39_59
timestamp 1586364061
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use scs8hd_decap_12  FILLER_40_44
timestamp 1586364061
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_56
timestamp 1586364061
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_265
timestamp 1586364061
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_62
timestamp 1586364061
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_74
timestamp 1586364061
transform 1 0 7912 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_68
timestamp 1586364061
transform 1 0 7360 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_270
timestamp 1586364061
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_86
timestamp 1586364061
transform 1 0 9016 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_98
timestamp 1586364061
transform 1 0 10120 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_80
timestamp 1586364061
transform 1 0 8464 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_93
timestamp 1586364061
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_110
timestamp 1586364061
transform 1 0 11224 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_105
timestamp 1586364061
transform 1 0 10764 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_117
timestamp 1586364061
transform 1 0 11868 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_266
timestamp 1586364061
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_123
timestamp 1586364061
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_135
timestamp 1586364061
transform 1 0 13524 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_129
timestamp 1586364061
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_271
timestamp 1586364061
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_147
timestamp 1586364061
transform 1 0 14628 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_141
timestamp 1586364061
transform 1 0 14076 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_154
timestamp 1586364061
transform 1 0 15272 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_159
timestamp 1586364061
transform 1 0 15732 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_171
timestamp 1586364061
transform 1 0 16836 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_166
timestamp 1586364061
transform 1 0 16376 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_178
timestamp 1586364061
transform 1 0 17480 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_267
timestamp 1586364061
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_184
timestamp 1586364061
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_196
timestamp 1586364061
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_190
timestamp 1586364061
transform 1 0 18584 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_272
timestamp 1586364061
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_208
timestamp 1586364061
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_202
timestamp 1586364061
transform 1 0 19688 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_215
timestamp 1586364061
transform 1 0 20884 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_220
timestamp 1586364061
transform 1 0 21344 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_232
timestamp 1586364061
transform 1 0 22448 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_227
timestamp 1586364061
transform 1 0 21988 0 -1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_268
timestamp 1586364061
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use scs8hd_decap_12  FILLER_39_245
timestamp 1586364061
transform 1 0 23644 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_39_257
timestamp 1586364061
transform 1 0 24748 0 1 23392
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_239
timestamp 1586364061
transform 1 0 23092 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_40_251
timestamp 1586364061
transform 1 0 24196 0 -1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_79
timestamp 1586364061
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use scs8hd_decap_3  PHY_81
timestamp 1586364061
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_273
timestamp 1586364061
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_8  FILLER_39_269
timestamp 1586364061
transform 1 0 25852 0 1 23392
box -38 -48 774 592
use scs8hd_decap_12  FILLER_40_263
timestamp 1586364061
transform 1 0 25300 0 -1 24480
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_40_276
timestamp 1586364061
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use scs8hd_decap_3  PHY_82
timestamp 1586364061
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use scs8hd_decap_12  FILLER_41_3
timestamp 1586364061
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_15
timestamp 1586364061
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_27
timestamp 1586364061
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_39
timestamp 1586364061
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_41_51
timestamp 1586364061
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use scs8hd_fill_2  FILLER_41_59
timestamp 1586364061
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_274
timestamp 1586364061
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_62
timestamp 1586364061
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_74
timestamp 1586364061
transform 1 0 7912 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_86
timestamp 1586364061
transform 1 0 9016 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_98
timestamp 1586364061
transform 1 0 10120 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_110
timestamp 1586364061
transform 1 0 11224 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_275
timestamp 1586364061
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_123
timestamp 1586364061
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_135
timestamp 1586364061
transform 1 0 13524 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_147
timestamp 1586364061
transform 1 0 14628 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_159
timestamp 1586364061
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_171
timestamp 1586364061
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_276
timestamp 1586364061
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_184
timestamp 1586364061
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_196
timestamp 1586364061
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_208
timestamp 1586364061
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_220
timestamp 1586364061
transform 1 0 21344 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_232
timestamp 1586364061
transform 1 0 22448 0 1 24480
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_277
timestamp 1586364061
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use scs8hd_decap_12  FILLER_41_245
timestamp 1586364061
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_41_257
timestamp 1586364061
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use scs8hd_decap_3  PHY_83
timestamp 1586364061
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use scs8hd_decap_8  FILLER_41_269
timestamp 1586364061
transform 1 0 25852 0 1 24480
box -38 -48 774 592
use scs8hd_decap_3  PHY_84
timestamp 1586364061
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_3
timestamp 1586364061
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_15
timestamp 1586364061
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_278
timestamp 1586364061
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_4  FILLER_42_27
timestamp 1586364061
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use scs8hd_decap_12  FILLER_42_32
timestamp 1586364061
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_44
timestamp 1586364061
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_56
timestamp 1586364061
transform 1 0 6256 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_279
timestamp 1586364061
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_63
timestamp 1586364061
transform 1 0 6900 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_75
timestamp 1586364061
transform 1 0 8004 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_280
timestamp 1586364061
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_87
timestamp 1586364061
transform 1 0 9108 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_94
timestamp 1586364061
transform 1 0 9752 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_106
timestamp 1586364061
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_118
timestamp 1586364061
transform 1 0 11960 0 -1 25568
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_281
timestamp 1586364061
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_125
timestamp 1586364061
transform 1 0 12604 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_137
timestamp 1586364061
transform 1 0 13708 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_282
timestamp 1586364061
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_149
timestamp 1586364061
transform 1 0 14812 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_156
timestamp 1586364061
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_168
timestamp 1586364061
transform 1 0 16560 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_283
timestamp 1586364061
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_180
timestamp 1586364061
transform 1 0 17664 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_187
timestamp 1586364061
transform 1 0 18308 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_284
timestamp 1586364061
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_12  FILLER_42_199
timestamp 1586364061
transform 1 0 19412 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_42_211
timestamp 1586364061
transform 1 0 20516 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_218
timestamp 1586364061
transform 1 0 21160 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_42_230
timestamp 1586364061
transform 1 0 22264 0 -1 25568
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_285
timestamp 1586364061
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use scs8hd_decap_6  FILLER_42_242
timestamp 1586364061
transform 1 0 23368 0 -1 25568
box -38 -48 590 592
use scs8hd_decap_12  FILLER_42_249
timestamp 1586364061
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_3  PHY_85
timestamp 1586364061
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use scs8hd_decap_12  FILLER_42_261
timestamp 1586364061
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_42_273
timestamp 1586364061
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 294 0 350 480 6 bottom_left_grid_pin_34_
port 0 nsew default input
rlabel metal2 s 846 0 902 480 6 bottom_left_grid_pin_35_
port 1 nsew default input
rlabel metal2 s 1398 0 1454 480 6 bottom_left_grid_pin_36_
port 2 nsew default input
rlabel metal2 s 1950 0 2006 480 6 bottom_left_grid_pin_37_
port 3 nsew default input
rlabel metal2 s 2502 0 2558 480 6 bottom_left_grid_pin_38_
port 4 nsew default input
rlabel metal2 s 3054 0 3110 480 6 bottom_left_grid_pin_39_
port 5 nsew default input
rlabel metal2 s 3606 0 3662 480 6 bottom_left_grid_pin_40_
port 6 nsew default input
rlabel metal2 s 4158 0 4214 480 6 bottom_left_grid_pin_41_
port 7 nsew default input
rlabel metal2 s 15934 0 15990 480 6 bottom_right_grid_pin_1_
port 8 nsew default input
rlabel metal3 s 27520 6944 28000 7064 6 ccff_head
port 9 nsew default input
rlabel metal2 s 27618 0 27674 480 6 ccff_tail
port 10 nsew default tristate
rlabel metal3 s 0 13880 480 14000 6 chanx_left_in[0]
port 11 nsew default input
rlabel metal3 s 0 20680 480 20800 6 chanx_left_in[10]
port 12 nsew default input
rlabel metal3 s 0 21360 480 21480 6 chanx_left_in[11]
port 13 nsew default input
rlabel metal3 s 0 22040 480 22160 6 chanx_left_in[12]
port 14 nsew default input
rlabel metal3 s 0 22720 480 22840 6 chanx_left_in[13]
port 15 nsew default input
rlabel metal3 s 0 23400 480 23520 6 chanx_left_in[14]
port 16 nsew default input
rlabel metal3 s 0 24080 480 24200 6 chanx_left_in[15]
port 17 nsew default input
rlabel metal3 s 0 24760 480 24880 6 chanx_left_in[16]
port 18 nsew default input
rlabel metal3 s 0 25440 480 25560 6 chanx_left_in[17]
port 19 nsew default input
rlabel metal3 s 0 26120 480 26240 6 chanx_left_in[18]
port 20 nsew default input
rlabel metal3 s 0 26800 480 26920 6 chanx_left_in[19]
port 21 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[1]
port 22 nsew default input
rlabel metal3 s 0 15240 480 15360 6 chanx_left_in[2]
port 23 nsew default input
rlabel metal3 s 0 15920 480 16040 6 chanx_left_in[3]
port 24 nsew default input
rlabel metal3 s 0 16600 480 16720 6 chanx_left_in[4]
port 25 nsew default input
rlabel metal3 s 0 17280 480 17400 6 chanx_left_in[5]
port 26 nsew default input
rlabel metal3 s 0 17960 480 18080 6 chanx_left_in[6]
port 27 nsew default input
rlabel metal3 s 0 18640 480 18760 6 chanx_left_in[7]
port 28 nsew default input
rlabel metal3 s 0 19320 480 19440 6 chanx_left_in[8]
port 29 nsew default input
rlabel metal3 s 0 20000 480 20120 6 chanx_left_in[9]
port 30 nsew default input
rlabel metal3 s 0 280 480 400 6 chanx_left_out[0]
port 31 nsew default tristate
rlabel metal3 s 0 7080 480 7200 6 chanx_left_out[10]
port 32 nsew default tristate
rlabel metal3 s 0 7760 480 7880 6 chanx_left_out[11]
port 33 nsew default tristate
rlabel metal3 s 0 8440 480 8560 6 chanx_left_out[12]
port 34 nsew default tristate
rlabel metal3 s 0 9120 480 9240 6 chanx_left_out[13]
port 35 nsew default tristate
rlabel metal3 s 0 9800 480 9920 6 chanx_left_out[14]
port 36 nsew default tristate
rlabel metal3 s 0 10480 480 10600 6 chanx_left_out[15]
port 37 nsew default tristate
rlabel metal3 s 0 11160 480 11280 6 chanx_left_out[16]
port 38 nsew default tristate
rlabel metal3 s 0 11840 480 11960 6 chanx_left_out[17]
port 39 nsew default tristate
rlabel metal3 s 0 12520 480 12640 6 chanx_left_out[18]
port 40 nsew default tristate
rlabel metal3 s 0 13200 480 13320 6 chanx_left_out[19]
port 41 nsew default tristate
rlabel metal3 s 0 960 480 1080 6 chanx_left_out[1]
port 42 nsew default tristate
rlabel metal3 s 0 1640 480 1760 6 chanx_left_out[2]
port 43 nsew default tristate
rlabel metal3 s 0 2320 480 2440 6 chanx_left_out[3]
port 44 nsew default tristate
rlabel metal3 s 0 3000 480 3120 6 chanx_left_out[4]
port 45 nsew default tristate
rlabel metal3 s 0 3680 480 3800 6 chanx_left_out[5]
port 46 nsew default tristate
rlabel metal3 s 0 4360 480 4480 6 chanx_left_out[6]
port 47 nsew default tristate
rlabel metal3 s 0 5040 480 5160 6 chanx_left_out[7]
port 48 nsew default tristate
rlabel metal3 s 0 5720 480 5840 6 chanx_left_out[8]
port 49 nsew default tristate
rlabel metal3 s 0 6400 480 6520 6 chanx_left_out[9]
port 50 nsew default tristate
rlabel metal2 s 4710 0 4766 480 6 chany_bottom_in[0]
port 51 nsew default input
rlabel metal2 s 10322 0 10378 480 6 chany_bottom_in[10]
port 52 nsew default input
rlabel metal2 s 10874 0 10930 480 6 chany_bottom_in[11]
port 53 nsew default input
rlabel metal2 s 11426 0 11482 480 6 chany_bottom_in[12]
port 54 nsew default input
rlabel metal2 s 11978 0 12034 480 6 chany_bottom_in[13]
port 55 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[14]
port 56 nsew default input
rlabel metal2 s 13082 0 13138 480 6 chany_bottom_in[15]
port 57 nsew default input
rlabel metal2 s 13634 0 13690 480 6 chany_bottom_in[16]
port 58 nsew default input
rlabel metal2 s 14278 0 14334 480 6 chany_bottom_in[17]
port 59 nsew default input
rlabel metal2 s 14830 0 14886 480 6 chany_bottom_in[18]
port 60 nsew default input
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_in[19]
port 61 nsew default input
rlabel metal2 s 5262 0 5318 480 6 chany_bottom_in[1]
port 62 nsew default input
rlabel metal2 s 5814 0 5870 480 6 chany_bottom_in[2]
port 63 nsew default input
rlabel metal2 s 6366 0 6422 480 6 chany_bottom_in[3]
port 64 nsew default input
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_in[4]
port 65 nsew default input
rlabel metal2 s 7562 0 7618 480 6 chany_bottom_in[5]
port 66 nsew default input
rlabel metal2 s 8114 0 8170 480 6 chany_bottom_in[6]
port 67 nsew default input
rlabel metal2 s 8666 0 8722 480 6 chany_bottom_in[7]
port 68 nsew default input
rlabel metal2 s 9218 0 9274 480 6 chany_bottom_in[8]
port 69 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[9]
port 70 nsew default input
rlabel metal2 s 16486 0 16542 480 6 chany_bottom_out[0]
port 71 nsew default tristate
rlabel metal2 s 22098 0 22154 480 6 chany_bottom_out[10]
port 72 nsew default tristate
rlabel metal2 s 22650 0 22706 480 6 chany_bottom_out[11]
port 73 nsew default tristate
rlabel metal2 s 23202 0 23258 480 6 chany_bottom_out[12]
port 74 nsew default tristate
rlabel metal2 s 23754 0 23810 480 6 chany_bottom_out[13]
port 75 nsew default tristate
rlabel metal2 s 24306 0 24362 480 6 chany_bottom_out[14]
port 76 nsew default tristate
rlabel metal2 s 24858 0 24914 480 6 chany_bottom_out[15]
port 77 nsew default tristate
rlabel metal2 s 25410 0 25466 480 6 chany_bottom_out[16]
port 78 nsew default tristate
rlabel metal2 s 25962 0 26018 480 6 chany_bottom_out[17]
port 79 nsew default tristate
rlabel metal2 s 26514 0 26570 480 6 chany_bottom_out[18]
port 80 nsew default tristate
rlabel metal2 s 27066 0 27122 480 6 chany_bottom_out[19]
port 81 nsew default tristate
rlabel metal2 s 17038 0 17094 480 6 chany_bottom_out[1]
port 82 nsew default tristate
rlabel metal2 s 17590 0 17646 480 6 chany_bottom_out[2]
port 83 nsew default tristate
rlabel metal2 s 18142 0 18198 480 6 chany_bottom_out[3]
port 84 nsew default tristate
rlabel metal2 s 18694 0 18750 480 6 chany_bottom_out[4]
port 85 nsew default tristate
rlabel metal2 s 19246 0 19302 480 6 chany_bottom_out[5]
port 86 nsew default tristate
rlabel metal2 s 19798 0 19854 480 6 chany_bottom_out[6]
port 87 nsew default tristate
rlabel metal2 s 20350 0 20406 480 6 chany_bottom_out[7]
port 88 nsew default tristate
rlabel metal2 s 20902 0 20958 480 6 chany_bottom_out[8]
port 89 nsew default tristate
rlabel metal2 s 21546 0 21602 480 6 chany_bottom_out[9]
port 90 nsew default tristate
rlabel metal3 s 0 27480 480 27600 6 left_top_grid_pin_1_
port 91 nsew default input
rlabel metal3 s 27520 20952 28000 21072 6 prog_clk
port 92 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 vpwr
port 93 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 vgnd
port 94 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 27600
<< end >>
