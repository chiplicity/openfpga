* NGSPICE file created from grid_io_top.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_1 abstract view
.subckt scs8hd_ebufn_1 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_and4_4 abstract view
.subckt scs8hd_and4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_1 abstract view
.subckt scs8hd_buf_1 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor4_4 abstract view
.subckt scs8hd_nor4_4 A B C D Y vgnd vpwr
.ends

.subckt grid_io_top address[0] address[1] address[2] address[3] bottom_width_0_height_0__pin_0_
+ bottom_width_0_height_0__pin_10_ bottom_width_0_height_0__pin_11_ bottom_width_0_height_0__pin_12_
+ bottom_width_0_height_0__pin_13_ bottom_width_0_height_0__pin_14_ bottom_width_0_height_0__pin_15_
+ bottom_width_0_height_0__pin_1_ bottom_width_0_height_0__pin_2_ bottom_width_0_height_0__pin_3_
+ bottom_width_0_height_0__pin_4_ bottom_width_0_height_0__pin_5_ bottom_width_0_height_0__pin_6_
+ bottom_width_0_height_0__pin_7_ bottom_width_0_height_0__pin_8_ bottom_width_0_height_0__pin_9_
+ data_in enable gfpga_pad_GPIO_PAD[0] gfpga_pad_GPIO_PAD[1] gfpga_pad_GPIO_PAD[2]
+ gfpga_pad_GPIO_PAD[3] gfpga_pad_GPIO_PAD[4] gfpga_pad_GPIO_PAD[5] gfpga_pad_GPIO_PAD[6]
+ gfpga_pad_GPIO_PAD[7] vpwr vgnd
XFILLER_18_406 vgnd vpwr scs8hd_fill_1
XFILLER_9_159 vgnd vpwr scs8hd_decap_12
XFILLER_3_45 vgnd vpwr scs8hd_decap_3
XFILLER_5_354 vgnd vpwr scs8hd_decap_12
XFILLER_12_98 vgnd vpwr scs8hd_decap_12
XFILLER_12_32 vgnd vpwr scs8hd_decap_12
XFILLER_6_129 vgnd vpwr scs8hd_decap_12
XFILLER_2_324 vgnd vpwr scs8hd_decap_12
XFILLER_5_184 vgnd vpwr scs8hd_decap_12
XFILLER_2_154 vgnd vpwr scs8hd_decap_12
XFILLER_2_198 vgnd vpwr scs8hd_decap_12
XFILLER_20_242 vgnd vpwr scs8hd_decap_6
XFILLER_11_220 vgnd vpwr scs8hd_decap_12
XFILLER_7_235 vpwr vgnd scs8hd_fill_2
XFILLER_7_213 vpwr vgnd scs8hd_fill_2
XFILLER_19_342 vgnd vpwr scs8hd_decap_12
XFILLER_20_87 vgnd vpwr scs8hd_decap_6
XFILLER_20_32 vgnd vpwr scs8hd_decap_12
XFILLER_16_312 vgnd vpwr scs8hd_decap_12
XFILLER_4_227 vgnd vpwr scs8hd_decap_12
XFILLER_13_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_56 vgnd vpwr scs8hd_decap_12
XFILLER_15_98 vgnd vpwr scs8hd_decap_12
XFILLER_1_208 vgnd vpwr scs8hd_decap_12
XPHY_181 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_170 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_385 vgnd vpwr scs8hd_decap_12
XFILLER_13_123 vgnd vpwr scs8hd_decap_12
XFILLER_9_116 vpwr vgnd scs8hd_fill_2
XFILLER_18_215 vgnd vpwr scs8hd_decap_12
XFILLER_12_44 vgnd vpwr scs8hd_decap_12
XFILLER_17_281 vgnd vpwr scs8hd_decap_12
XFILLER_1_391 vgnd vpwr scs8hd_decap_12
XFILLER_5_196 vgnd vpwr scs8hd_decap_12
XFILLER_14_251 vgnd vpwr scs8hd_decap_12
XFILLER_0_36 vgnd vpwr scs8hd_fill_1
XFILLER_2_166 vgnd vpwr scs8hd_decap_12
XFILLER_18_32 vgnd vpwr scs8hd_decap_12
XFILLER_11_243 vgnd vpwr scs8hd_fill_1
XFILLER_7_225 vgnd vpwr scs8hd_decap_4
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _10_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_354 vgnd vpwr scs8hd_decap_12
XFILLER_20_44 vgnd vpwr scs8hd_decap_12
XFILLER_4_239 vgnd vpwr scs8hd_decap_12
XFILLER_19_184 vgnd vpwr scs8hd_decap_12
XFILLER_16_324 vgnd vpwr scs8hd_decap_12
XFILLER_6_68 vgnd vpwr scs8hd_decap_12
XPHY_182 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_160 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_154 vgnd vpwr scs8hd_decap_12
XFILLER_0_275 vgnd vpwr scs8hd_decap_4
XFILLER_13_135 vgnd vpwr scs8hd_decap_12
XFILLER_5_367 vgnd vpwr scs8hd_decap_12
XFILLER_12_56 vgnd vpwr scs8hd_decap_12
XFILLER_2_337 vgnd vpwr scs8hd_decap_12
XFILLER_18_227 vgnd vpwr scs8hd_decap_12
XFILLER_17_293 vgnd vpwr scs8hd_decap_12
XFILLER_15_208 vgnd vpwr scs8hd_decap_12
XFILLER_14_263 vgnd vpwr scs8hd_decap_12
XFILLER_11_403 vgnd vpwr scs8hd_decap_4
XFILLER_0_59 vgnd vpwr scs8hd_decap_3
XFILLER_0_15 vpwr vgnd scs8hd_fill_2
XFILLER_2_178 vgnd vpwr scs8hd_decap_6
XFILLER_3_3 vgnd vpwr scs8hd_decap_12
XFILLER_20_211 vgnd vpwr scs8hd_decap_6
XFILLER_18_44 vgnd vpwr scs8hd_decap_12
XFILLER_6_270 vgnd vpwr scs8hd_decap_4
XFILLER_20_56 vgnd vpwr scs8hd_decap_6
XFILLER_3_273 vgnd vpwr scs8hd_decap_12
XFILLER_19_196 vgnd vpwr scs8hd_decap_12
XFILLER_15_391 vgnd vpwr scs8hd_decap_12
XFILLER_16_166 vgnd vpwr scs8hd_decap_12
XFILLER_13_306 vgnd vpwr scs8hd_decap_12
XANTENNA__04__A address[3] vgnd vpwr scs8hd_diode_2
XPHY_183 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_361 vgnd vpwr scs8hd_decap_12
XFILLER_8_398 vgnd vpwr scs8hd_decap_8
XFILLER_13_147 vgnd vpwr scs8hd_decap_12
XFILLER_3_15 vgnd vpwr scs8hd_decap_4
XFILLER_5_379 vgnd vpwr scs8hd_decap_12
XFILLER_12_68 vgnd vpwr scs8hd_decap_12
XFILLER_18_239 vgnd vpwr scs8hd_decap_12
XFILLER_2_349 vgnd vpwr scs8hd_decap_12
XFILLER_5_110 vgnd vpwr scs8hd_decap_12
XFILLER_20_404 vgnd vpwr scs8hd_decap_3
Xlogical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ bottom_width_0_height_0__pin_8_ logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[4] vgnd vpwr scs8hd_ebufn_1
XFILLER_4_91 vgnd vpwr scs8hd_fill_1
XANTENNA__12__A _06_/Y vgnd vpwr scs8hd_diode_2
XFILLER_0_27 vgnd vpwr scs8hd_decap_4
XFILLER_18_56 vgnd vpwr scs8hd_decap_12
XANTENNA__07__A _04_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_367 vgnd vpwr scs8hd_decap_12
XFILLER_11_245 vgnd vpwr scs8hd_decap_12
XFILLER_7_249 vgnd vpwr scs8hd_fill_1
XFILLER_16_337 vgnd vpwr scs8hd_decap_12
XFILLER_6_15 vgnd vpwr scs8hd_decap_12
XFILLER_3_285 vgnd vpwr scs8hd_decap_12
XFILLER_13_318 vgnd vpwr scs8hd_decap_12
XANTENNA__20__A gfpga_pad_GPIO_PAD[1] vgnd vpwr scs8hd_diode_2
XFILLER_0_255 vpwr vgnd scs8hd_fill_2
XFILLER_0_288 vgnd vpwr scs8hd_decap_12
XPHY_184 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_178 vgnd vpwr scs8hd_decap_12
XPHY_151 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_373 vgnd vpwr scs8hd_decap_12
XFILLER_11_3 vgnd vpwr scs8hd_decap_12
XFILLER_8_300 vgnd vpwr scs8hd_decap_12
XFILLER_7_91 vpwr vgnd scs8hd_fill_2
XFILLER_13_159 vgnd vpwr scs8hd_decap_12
XFILLER_9_108 vpwr vgnd scs8hd_fill_2
XANTENNA__15__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_8_152 vgnd vpwr scs8hd_fill_1
XANTENNA__12__B _11_/Y vgnd vpwr scs8hd_diode_2
Xlogical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _12_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_14_276 vgnd vpwr scs8hd_decap_12
XFILLER_9_59 vpwr vgnd scs8hd_fill_2
XFILLER_9_15 vgnd vpwr scs8hd_decap_12
XFILLER_0_39 vpwr vgnd scs8hd_fill_2
XFILLER_18_68 vgnd vpwr scs8hd_decap_12
XFILLER_19_379 vgnd vpwr scs8hd_decap_12
XFILLER_11_257 vgnd vpwr scs8hd_decap_12
XFILLER_11_235 vpwr vgnd scs8hd_fill_2
XFILLER_7_239 vpwr vgnd scs8hd_fill_2
XANTENNA__07__B address[2] vgnd vpwr scs8hd_diode_2
XFILLER_7_217 vpwr vgnd scs8hd_fill_2
XANTENNA__23__A gfpga_pad_GPIO_PAD[4] vgnd vpwr scs8hd_diode_2
XFILLER_16_349 vgnd vpwr scs8hd_decap_12
XANTENNA__18__A gfpga_pad_GPIO_PAD[7] vgnd vpwr scs8hd_diode_2
XFILLER_0_404 vgnd vpwr scs8hd_decap_3
XFILLER_19_110 vgnd vpwr scs8hd_decap_12
XFILLER_10_80 vgnd vpwr scs8hd_decap_12
XFILLER_3_297 vgnd vpwr scs8hd_decap_8
XFILLER_6_27 vgnd vpwr scs8hd_decap_4
XPHY_185 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_152 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_385 vgnd vpwr scs8hd_decap_12
XPHY_130 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_312 vgnd vpwr scs8hd_decap_12
XANTENNA__15__B _11_/Y vgnd vpwr scs8hd_diode_2
XFILLER_12_15 vgnd vpwr scs8hd_decap_12
XFILLER_10_119 vgnd vpwr scs8hd_decap_12
XFILLER_5_123 vgnd vpwr scs8hd_decap_12
XANTENNA__12__C _04_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_71 vgnd vpwr scs8hd_decap_12
XFILLER_4_93 vgnd vpwr scs8hd_decap_12
XFILLER_14_288 vgnd vpwr scs8hd_decap_12
XFILLER_9_27 vgnd vpwr scs8hd_decap_12
XFILLER_9_281 vgnd vpwr scs8hd_decap_12
XFILLER_11_269 vgnd vpwr scs8hd_decap_12
XANTENNA__07__C _06_/Y vgnd vpwr scs8hd_diode_2
XFILLER_6_251 vgnd vpwr scs8hd_fill_1
XFILLER_20_15 vgnd vpwr scs8hd_decap_12
XFILLER_3_243 vgnd vpwr scs8hd_fill_1
XFILLER_15_59 vpwr vgnd scs8hd_fill_2
XFILLER_15_15 vgnd vpwr scs8hd_decap_12
XPHY_186 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_175 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_153 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_142 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_324 vgnd vpwr scs8hd_decap_12
XFILLER_0_246 vpwr vgnd scs8hd_fill_2
XFILLER_0_213 vpwr vgnd scs8hd_fill_2
XPHY_0 vgnd vpwr scs8hd_decap_3
XANTENNA__15__C _04_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_80 vgnd vpwr scs8hd_decap_12
XFILLER_8_154 vgnd vpwr scs8hd_decap_12
XFILLER_8_110 vgnd vpwr scs8hd_decap_12
XFILLER_12_27 vgnd vpwr scs8hd_decap_4
XFILLER_17_220 vgnd vpwr scs8hd_decap_12
XFILLER_1_330 vgnd vpwr scs8hd_decap_12
XFILLER_5_135 vgnd vpwr scs8hd_decap_12
XFILLER_4_83 vgnd vpwr scs8hd_decap_8
XFILLER_4_190 vgnd vpwr scs8hd_decap_12
XANTENNA__12__D _08_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_39 vgnd vpwr scs8hd_decap_12
XFILLER_2_105 vgnd vpwr scs8hd_decap_12
XFILLER_9_293 vgnd vpwr scs8hd_decap_12
XFILLER_1_171 vpwr vgnd scs8hd_fill_2
XFILLER_18_15 vgnd vpwr scs8hd_decap_12
XANTENNA__07__D enable vgnd vpwr scs8hd_diode_2
XFILLER_7_208 vgnd vpwr scs8hd_decap_3
XFILLER_3_403 vgnd vpwr scs8hd_decap_4
XFILLER_6_274 vgnd vpwr scs8hd_fill_1
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_20_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_62 vgnd vpwr scs8hd_decap_12
XFILLER_19_123 vgnd vpwr scs8hd_decap_12
XFILLER_10_93 vgnd vpwr scs8hd_decap_3
XFILLER_15_27 vgnd vpwr scs8hd_decap_12
X_09_ address[1] enable address[3] _08_/Y _09_/X vgnd vpwr scs8hd_and4_4
XPHY_187 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_398 vgnd vpwr scs8hd_decap_8
XPHY_1 vgnd vpwr scs8hd_decap_3
XFILLER_7_391 vgnd vpwr scs8hd_decap_12
XANTENNA__15__D address[2] vgnd vpwr scs8hd_diode_2
XFILLER_5_306 vgnd vpwr scs8hd_decap_12
XFILLER_8_166 vgnd vpwr scs8hd_decap_12
XFILLER_8_122 vgnd vpwr scs8hd_decap_12
XFILLER_3_19 vgnd vpwr scs8hd_fill_1
XFILLER_4_361 vgnd vpwr scs8hd_decap_12
XFILLER_1_342 vgnd vpwr scs8hd_decap_12
XFILLER_5_147 vgnd vpwr scs8hd_decap_12
XFILLER_17_232 vgnd vpwr scs8hd_decap_12
XFILLER_14_202 vgnd vpwr scs8hd_decap_12
XFILLER_2_117 vgnd vpwr scs8hd_decap_12
XFILLER_20_249 vgnd vpwr scs8hd_decap_12
XFILLER_18_27 vgnd vpwr scs8hd_decap_4
XFILLER_1_74 vgnd vpwr scs8hd_decap_12
XFILLER_3_212 vpwr vgnd scs8hd_fill_2
XFILLER_3_245 vgnd vpwr scs8hd_decap_12
XFILLER_19_135 vgnd vpwr scs8hd_decap_12
XFILLER_15_330 vgnd vpwr scs8hd_decap_12
X_08_ address[2] _08_/Y vgnd vpwr scs8hd_inv_8
Xlogical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ bottom_width_0_height_0__pin_10_ logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[5] vgnd vpwr scs8hd_ebufn_1
XFILLER_18_190 vgnd vpwr scs8hd_decap_12
XFILLER_16_105 vgnd vpwr scs8hd_decap_12
XFILLER_15_39 vgnd vpwr scs8hd_decap_12
XPHY_100 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_0_226 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ bottom_width_0_height_0__pin_14_ vgnd vpwr scs8hd_diode_2
XFILLER_0_259 vpwr vgnd scs8hd_fill_2
XPHY_177 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_171 vgnd vpwr scs8hd_decap_12
XPHY_144 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_300 vgnd vpwr scs8hd_decap_12
XPHY_122 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_111 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_337 vgnd vpwr scs8hd_decap_12
XPHY_2 vgnd vpwr scs8hd_decap_3
XFILLER_7_95 vpwr vgnd scs8hd_fill_2
XFILLER_7_51 vgnd vpwr scs8hd_decap_8
XFILLER_7_62 vgnd vpwr scs8hd_decap_12
XFILLER_17_403 vgnd vpwr scs8hd_decap_4
XFILLER_16_93 vgnd vpwr scs8hd_decap_12
XFILLER_12_152 vgnd vpwr scs8hd_fill_1
XFILLER_8_178 vgnd vpwr scs8hd_decap_12
XFILLER_8_134 vgnd vpwr scs8hd_decap_12
XFILLER_5_318 vgnd vpwr scs8hd_decap_12
XFILLER_4_373 vgnd vpwr scs8hd_decap_12
XFILLER_14_406 vgnd vpwr scs8hd_fill_1
XFILLER_1_354 vgnd vpwr scs8hd_decap_12
XFILLER_5_159 vgnd vpwr scs8hd_decap_12
XFILLER_2_129 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ bottom_width_0_height_0__pin_10_ vgnd vpwr scs8hd_diode_2
XFILLER_1_184 vgnd vpwr scs8hd_decap_12
XFILLER_11_239 vpwr vgnd scs8hd_fill_2
XFILLER_19_306 vgnd vpwr scs8hd_decap_12
XFILLER_18_361 vgnd vpwr scs8hd_decap_12
XFILLER_6_276 vgnd vpwr scs8hd_decap_12
XFILLER_6_254 vpwr vgnd scs8hd_fill_2
XFILLER_1_86 vgnd vpwr scs8hd_decap_12
XFILLER_1_31 vgnd vpwr scs8hd_decap_12
XFILLER_3_257 vgnd vpwr scs8hd_decap_3
XFILLER_19_147 vgnd vpwr scs8hd_decap_12
XFILLER_15_342 vgnd vpwr scs8hd_decap_12
X_07_ _04_/X address[2] _06_/Y enable _07_/X vgnd vpwr scs8hd_and4_4
XFILLER_0_249 vpwr vgnd scs8hd_fill_2
XFILLER_0_238 vgnd vpwr scs8hd_decap_8
XPHY_189 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_117 vgnd vpwr scs8hd_decap_12
XPHY_145 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_312 vgnd vpwr scs8hd_decap_12
XPHY_123 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_349 vgnd vpwr scs8hd_decap_12
XPHY_101 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ bottom_width_0_height_0__pin_6_ vgnd vpwr scs8hd_diode_2
XPHY_3 vgnd vpwr scs8hd_decap_3
XFILLER_7_74 vgnd vpwr scs8hd_decap_12
XFILLER_12_175 vgnd vpwr scs8hd_decap_12
XFILLER_8_146 vgnd vpwr scs8hd_decap_6
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_4_385 vgnd vpwr scs8hd_decap_12
XFILLER_17_245 vgnd vpwr scs8hd_decap_12
XFILLER_14_215 vgnd vpwr scs8hd_decap_12
XFILLER_13_62 vgnd vpwr scs8hd_decap_12
XFILLER_13_51 vgnd vpwr scs8hd_decap_8
XFILLER_1_196 vgnd vpwr scs8hd_decap_12
XFILLER_20_218 vgnd vpwr scs8hd_decap_12
XFILLER_13_281 vgnd vpwr scs8hd_decap_12
XFILLER_19_318 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ bottom_width_0_height_0__pin_2_ vgnd vpwr scs8hd_diode_2
XFILLER_18_373 vgnd vpwr scs8hd_decap_12
XFILLER_10_251 vgnd vpwr scs8hd_decap_12
XFILLER_6_288 vgnd vpwr scs8hd_decap_12
X_23_ gfpga_pad_GPIO_PAD[4] bottom_width_0_height_0__pin_9_ vgnd vpwr scs8hd_buf_2
XFILLER_1_98 vgnd vpwr scs8hd_decap_12
XFILLER_1_43 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _12_/Y vgnd vpwr scs8hd_diode_2
XFILLER_19_159 vgnd vpwr scs8hd_decap_12
XFILLER_15_354 vgnd vpwr scs8hd_decap_12
X_06_ address[1] _06_/Y vgnd vpwr scs8hd_inv_8
XPHY_179 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_157 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_129 vgnd vpwr scs8hd_decap_12
XPHY_146 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_324 vgnd vpwr scs8hd_decap_12
XPHY_124 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_184 vgnd vpwr scs8hd_decap_12
XFILLER_7_86 vgnd vpwr scs8hd_decap_3
XPHY_4 vgnd vpwr scs8hd_decap_3
XFILLER_12_187 vgnd vpwr scs8hd_decap_12
XFILLER_12_154 vgnd vpwr scs8hd_decap_12
XFILLER_12_110 vgnd vpwr scs8hd_decap_12
XFILLER_17_257 vgnd vpwr scs8hd_decap_12
XFILLER_1_367 vgnd vpwr scs8hd_decap_12
XFILLER_4_32 vgnd vpwr scs8hd_decap_12
XFILLER_14_227 vgnd vpwr scs8hd_decap_12
XFILLER_13_74 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_13_293 vgnd vpwr scs8hd_decap_12
XFILLER_1_175 vgnd vpwr scs8hd_decap_8
Xlogical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _05_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_208 vgnd vpwr scs8hd_decap_12
XFILLER_18_385 vgnd vpwr scs8hd_decap_12
XFILLER_10_263 vgnd vpwr scs8hd_decap_12
X_22_ gfpga_pad_GPIO_PAD[3] bottom_width_0_height_0__pin_7_ vgnd vpwr scs8hd_buf_2
XFILLER_1_55 vgnd vpwr scs8hd_decap_6
XFILLER_1_11 vpwr vgnd scs8hd_fill_2
XFILLER_19_62 vgnd vpwr scs8hd_decap_12
XFILLER_19_51 vgnd vpwr scs8hd_decap_8
XFILLER_18_3 vgnd vpwr scs8hd_decap_12
X_05_ _04_/X address[2] address[1] enable _05_/X vgnd vpwr scs8hd_and4_4
XPHY_169 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_158 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_196 vgnd vpwr scs8hd_decap_12
XFILLER_11_391 vgnd vpwr scs8hd_decap_12
XPHY_5 vgnd vpwr scs8hd_decap_3
XFILLER_12_199 vgnd vpwr scs8hd_decap_12
XFILLER_12_122 vgnd vpwr scs8hd_decap_12
XFILLER_4_398 vgnd vpwr scs8hd_decap_8
XFILLER_17_269 vgnd vpwr scs8hd_decap_12
XFILLER_1_379 vgnd vpwr scs8hd_decap_12
XFILLER_4_44 vgnd vpwr scs8hd_decap_4
XFILLER_14_239 vgnd vpwr scs8hd_decap_12
XFILLER_13_86 vgnd vpwr scs8hd_decap_12
XFILLER_9_243 vgnd vpwr scs8hd_fill_1
XFILLER_1_110 vgnd vpwr scs8hd_decap_12
XFILLER_6_202 vgnd vpwr scs8hd_decap_12
X_21_ gfpga_pad_GPIO_PAD[2] bottom_width_0_height_0__pin_5_ vgnd vpwr scs8hd_buf_2
XFILLER_19_74 vgnd vpwr scs8hd_decap_12
XFILLER_10_98 vpwr vgnd scs8hd_fill_2
XFILLER_10_32 vgnd vpwr scs8hd_decap_12
XFILLER_3_227 vgnd vpwr scs8hd_decap_12
XFILLER_15_367 vgnd vpwr scs8hd_decap_12
X_04_ address[3] _04_/X vgnd vpwr scs8hd_buf_1
XFILLER_2_260 vpwr vgnd scs8hd_fill_2
Xlogical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _13_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XPHY_159 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_337 vgnd vpwr scs8hd_decap_12
XPHY_126 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_7_330 vgnd vpwr scs8hd_decap_12
XPHY_6 vgnd vpwr scs8hd_decap_3
XFILLER_7_99 vpwr vgnd scs8hd_fill_2
XFILLER_12_134 vgnd vpwr scs8hd_decap_12
XFILLER_4_300 vgnd vpwr scs8hd_decap_12
XFILLER_7_171 vgnd vpwr scs8hd_decap_12
XFILLER_9_403 vgnd vpwr scs8hd_decap_4
Xlogical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ bottom_width_0_height_0__pin_12_ logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[6] vgnd vpwr scs8hd_ebufn_1
XFILLER_4_23 vgnd vpwr scs8hd_decap_8
XFILLER_4_141 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_98 vgnd vpwr scs8hd_decap_12
XFILLER_9_211 vgnd vpwr scs8hd_decap_12
XFILLER_8_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_406 vgnd vpwr scs8hd_fill_1
XFILLER_10_276 vgnd vpwr scs8hd_decap_12
XFILLER_6_258 vgnd vpwr scs8hd_decap_12
XFILLER_18_398 vgnd vpwr scs8hd_decap_8
X_20_ gfpga_pad_GPIO_PAD[1] bottom_width_0_height_0__pin_3_ vgnd vpwr scs8hd_buf_2
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_10_44 vgnd vpwr scs8hd_decap_12
XFILLER_3_239 vgnd vpwr scs8hd_decap_4
XFILLER_19_86 vgnd vpwr scs8hd_decap_12
XFILLER_15_379 vgnd vpwr scs8hd_decap_12
XFILLER_2_272 vgnd vpwr scs8hd_decap_3
XPHY_116 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_105 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_110 vgnd vpwr scs8hd_decap_12
XPHY_138 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_12_349 vgnd vpwr scs8hd_decap_12
XPHY_127 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XPHY_7 vgnd vpwr scs8hd_decap_3
XFILLER_7_342 vgnd vpwr scs8hd_decap_12
XFILLER_16_32 vgnd vpwr scs8hd_decap_12
XFILLER_12_146 vgnd vpwr scs8hd_decap_6
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _05_/X vgnd vpwr scs8hd_diode_2
XFILLER_4_312 vgnd vpwr scs8hd_decap_12
XFILLER_1_304 vgnd vpwr scs8hd_fill_1
XANTENNA_logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_1_123 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_13_230 vgnd vpwr scs8hd_decap_12
XFILLER_9_245 vgnd vpwr scs8hd_decap_12
XFILLER_9_223 vgnd vpwr scs8hd_decap_12
XFILLER_6_215 vgnd vpwr scs8hd_decap_12
XFILLER_18_300 vgnd vpwr scs8hd_decap_12
XFILLER_10_288 vgnd vpwr scs8hd_decap_12
XFILLER_10_56 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_3_207 vgnd vpwr scs8hd_decap_3
XFILLER_5_281 vgnd vpwr scs8hd_decap_12
XFILLER_19_98 vgnd vpwr scs8hd_decap_12
XFILLER_18_141 vgnd vpwr scs8hd_decap_12
XPHY_139 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_106 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_3 vgnd vpwr scs8hd_decap_12
XFILLER_7_354 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XPHY_8 vgnd vpwr scs8hd_decap_3
XFILLER_16_44 vgnd vpwr scs8hd_decap_12
XFILLER_20_180 vgnd vpwr scs8hd_decap_6
XFILLER_11_180 vgnd vpwr scs8hd_decap_3
XFILLER_4_324 vgnd vpwr scs8hd_decap_12
XFILLER_7_184 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_D
+ data_in vgnd vpwr scs8hd_diode_2
XFILLER_4_154 vgnd vpwr scs8hd_decap_12
XFILLER_1_135 vgnd vpwr scs8hd_decap_12
XFILLER_13_242 vpwr vgnd scs8hd_fill_2
XFILLER_9_257 vgnd vpwr scs8hd_decap_12
XFILLER_9_235 vgnd vpwr scs8hd_decap_8
XFILLER_18_312 vgnd vpwr scs8hd_decap_12
XFILLER_10_212 vpwr vgnd scs8hd_fill_2
XFILLER_6_227 vgnd vpwr scs8hd_decap_12
XFILLER_1_15 vpwr vgnd scs8hd_fill_2
XFILLER_5_293 vgnd vpwr scs8hd_decap_12
XFILLER_10_68 vgnd vpwr scs8hd_decap_12
XFILLER_20_373 vgnd vpwr scs8hd_decap_12
XPHY_129 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA__10__A _06_/Y vgnd vpwr scs8hd_diode_2
XPHY_107 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_80 vgnd vpwr scs8hd_decap_6
XFILLER_15_123 vgnd vpwr scs8hd_decap_12
XPHY_9 vgnd vpwr scs8hd_decap_3
XFILLER_16_56 vgnd vpwr scs8hd_decap_12
XANTENNA__05__A _04_/X vgnd vpwr scs8hd_diode_2
XFILLER_19_281 vgnd vpwr scs8hd_decap_12
XFILLER_7_196 vgnd vpwr scs8hd_decap_12
XFILLER_3_391 vgnd vpwr scs8hd_decap_12
XFILLER_1_306 vgnd vpwr scs8hd_decap_12
XFILLER_16_251 vgnd vpwr scs8hd_decap_12
XFILLER_4_15 vgnd vpwr scs8hd_decap_6
XFILLER_4_59 vgnd vpwr scs8hd_decap_12
XFILLER_4_166 vgnd vpwr scs8hd_decap_12
XFILLER_1_147 vgnd vpwr scs8hd_decap_12
XFILLER_9_269 vgnd vpwr scs8hd_decap_12
XFILLER_18_324 vgnd vpwr scs8hd_decap_12
XANTENNA__13__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_6_239 vgnd vpwr scs8hd_decap_12
XFILLER_6_3 vgnd vpwr scs8hd_decap_12
XANTENNA__08__A address[2] vgnd vpwr scs8hd_diode_2
XFILLER_18_154 vgnd vpwr scs8hd_decap_12
XFILLER_2_264 vgnd vpwr scs8hd_decap_8
XFILLER_20_385 vgnd vpwr scs8hd_decap_12
XPHY_119 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_108 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_15_135 vgnd vpwr scs8hd_decap_12
XFILLER_11_330 vgnd vpwr scs8hd_decap_12
XANTENNA__10__B enable vgnd vpwr scs8hd_diode_2
XFILLER_7_367 vgnd vpwr scs8hd_decap_12
XFILLER_7_15 vgnd vpwr scs8hd_decap_12
XFILLER_7_59 vpwr vgnd scs8hd_fill_2
XFILLER_14_190 vgnd vpwr scs8hd_decap_12
XFILLER_16_68 vgnd vpwr scs8hd_decap_12
XANTENNA__05__B address[2] vgnd vpwr scs8hd_diode_2
XANTENNA__21__A gfpga_pad_GPIO_PAD[2] vgnd vpwr scs8hd_diode_2
XFILLER_4_337 vgnd vpwr scs8hd_decap_12
XFILLER_19_293 vgnd vpwr scs8hd_decap_12
XFILLER_17_208 vgnd vpwr scs8hd_decap_12
XFILLER_13_403 vgnd vpwr scs8hd_decap_4
XFILLER_8_80 vgnd vpwr scs8hd_decap_12
XANTENNA__16__A gfpga_pad_GPIO_PAD[5] vgnd vpwr scs8hd_diode_2
XFILLER_1_318 vgnd vpwr scs8hd_decap_12
XFILLER_16_263 vgnd vpwr scs8hd_decap_12
XFILLER_0_373 vgnd vpwr scs8hd_decap_12
XFILLER_4_178 vgnd vpwr scs8hd_decap_12
XFILLER_10_406 vgnd vpwr scs8hd_fill_1
XFILLER_1_159 vgnd vpwr scs8hd_decap_8
XANTENNA__13__B _11_/Y vgnd vpwr scs8hd_diode_2
XFILLER_17_391 vgnd vpwr scs8hd_decap_12
XFILLER_15_306 vgnd vpwr scs8hd_decap_12
XFILLER_10_15 vgnd vpwr scs8hd_decap_12
XFILLER_18_166 vgnd vpwr scs8hd_decap_12
XFILLER_14_361 vgnd vpwr scs8hd_decap_12
XFILLER_2_210 vgnd vpwr scs8hd_decap_4
XFILLER_2_276 vgnd vpwr scs8hd_decap_12
XFILLER_20_342 vgnd vpwr scs8hd_decap_12
XPHY_109 vgnd vpwr scs8hd_tapvpwrvgnd_1
Xlogical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ bottom_width_0_height_0__pin_14_ logical_tile_io_mode_io__7.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[7] vgnd vpwr scs8hd_ebufn_1
XFILLER_2_93 vgnd vpwr scs8hd_decap_12
XFILLER_20_397 vgnd vpwr scs8hd_decap_6
XFILLER_15_147 vgnd vpwr scs8hd_decap_12
XFILLER_11_342 vgnd vpwr scs8hd_decap_12
XANTENNA__10__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_7_379 vgnd vpwr scs8hd_decap_12
XANTENNA__19__A gfpga_pad_GPIO_PAD[0] vgnd vpwr scs8hd_diode_2
XFILLER_7_27 vgnd vpwr scs8hd_decap_12
XANTENNA__05__C address[1] vgnd vpwr scs8hd_diode_2
XFILLER_4_349 vgnd vpwr scs8hd_decap_12
XFILLER_14_3 vgnd vpwr scs8hd_decap_12
XFILLER_0_385 vgnd vpwr scs8hd_decap_12
XFILLER_13_15 vgnd vpwr scs8hd_decap_12
XFILLER_13_245 vgnd vpwr scs8hd_decap_12
XFILLER_13_59 vpwr vgnd scs8hd_fill_2
XFILLER_0_171 vgnd vpwr scs8hd_decap_12
XFILLER_0_160 vgnd vpwr scs8hd_fill_1
XFILLER_10_215 vgnd vpwr scs8hd_decap_12
XFILLER_10_204 vgnd vpwr scs8hd_decap_8
XANTENNA__13__C _04_/X vgnd vpwr scs8hd_diode_2
XFILLER_5_60 vgnd vpwr scs8hd_fill_1
XFILLER_18_337 vgnd vpwr scs8hd_decap_12
XFILLER_14_80 vgnd vpwr scs8hd_decap_12
XFILLER_10_27 vgnd vpwr scs8hd_decap_4
XFILLER_15_318 vgnd vpwr scs8hd_decap_12
XFILLER_2_288 vgnd vpwr scs8hd_decap_12
XFILLER_18_178 vgnd vpwr scs8hd_decap_12
XFILLER_14_373 vgnd vpwr scs8hd_decap_12
XPHY_90 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _13_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_354 vgnd vpwr scs8hd_decap_12
XFILLER_15_159 vgnd vpwr scs8hd_decap_12
XANTENNA__10__D _08_/Y vgnd vpwr scs8hd_diode_2
Xlogical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _07_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_11_354 vgnd vpwr scs8hd_decap_12
XFILLER_11_92 vpwr vgnd scs8hd_fill_2
XFILLER_7_39 vgnd vpwr scs8hd_decap_12
XFILLER_16_15 vgnd vpwr scs8hd_decap_12
XANTENNA__05__D enable vgnd vpwr scs8hd_diode_2
XFILLER_11_184 vgnd vpwr scs8hd_decap_12
XFILLER_0_342 vgnd vpwr scs8hd_decap_12
XFILLER_0_397 vgnd vpwr scs8hd_decap_6
XFILLER_16_276 vgnd vpwr scs8hd_decap_12
XFILLER_13_27 vgnd vpwr scs8hd_decap_12
XFILLER_13_257 vgnd vpwr scs8hd_decap_12
XFILLER_0_183 vgnd vpwr scs8hd_decap_3
XFILLER_10_227 vgnd vpwr scs8hd_decap_12
XANTENNA__13__D _08_/Y vgnd vpwr scs8hd_diode_2
XFILLER_8_250 vpwr vgnd scs8hd_fill_2
XFILLER_18_349 vgnd vpwr scs8hd_decap_12
XFILLER_1_19 vgnd vpwr scs8hd_decap_12
XFILLER_5_220 vgnd vpwr scs8hd_decap_12
XFILLER_19_59 vpwr vgnd scs8hd_fill_2
XFILLER_19_15 vgnd vpwr scs8hd_decap_12
XFILLER_4_3 vgnd vpwr scs8hd_decap_12
XFILLER_14_385 vgnd vpwr scs8hd_decap_12
XPHY_91 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_80 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_20_366 vgnd vpwr scs8hd_decap_6
XFILLER_20_311 vgnd vpwr scs8hd_decap_12
XFILLER_16_27 vgnd vpwr scs8hd_decap_4
XFILLER_11_196 vgnd vpwr scs8hd_decap_12
XFILLER_7_123 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _14_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_16_288 vgnd vpwr scs8hd_decap_12
XFILLER_0_354 vgnd vpwr scs8hd_decap_12
XFILLER_13_39 vgnd vpwr scs8hd_decap_12
XFILLER_13_269 vgnd vpwr scs8hd_decap_12
XFILLER_5_62 vgnd vpwr scs8hd_decap_12
XFILLER_10_239 vgnd vpwr scs8hd_decap_12
XFILLER_14_93 vgnd vpwr scs8hd_decap_12
XFILLER_5_232 vgnd vpwr scs8hd_decap_12
XFILLER_19_27 vgnd vpwr scs8hd_decap_12
XPHY_92 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_70 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_81 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_20_323 vgnd vpwr scs8hd_decap_12
XFILLER_2_30 vgnd vpwr scs8hd_fill_1
XFILLER_11_367 vgnd vpwr scs8hd_decap_12
XFILLER_19_220 vgnd vpwr scs8hd_decap_12
XFILLER_7_135 vgnd vpwr scs8hd_decap_12
XFILLER_3_330 vgnd vpwr scs8hd_decap_12
XFILLER_6_190 vgnd vpwr scs8hd_decap_12
XFILLER_4_105 vgnd vpwr scs8hd_decap_12
XFILLER_0_300 vgnd vpwr scs8hd_decap_8
XFILLER_0_311 vgnd vpwr scs8hd_decap_12
XFILLER_0_366 vgnd vpwr scs8hd_decap_6
XFILLER_12_3 vgnd vpwr scs8hd_decap_12
XFILLER_3_171 vgnd vpwr scs8hd_decap_8
XFILLER_13_204 vgnd vpwr scs8hd_decap_3
XFILLER_5_403 vgnd vpwr scs8hd_decap_4
XFILLER_8_274 vgnd vpwr scs8hd_fill_1
XFILLER_5_74 vgnd vpwr scs8hd_decap_12
XFILLER_2_406 vgnd vpwr scs8hd_fill_1
XFILLER_19_39 vgnd vpwr scs8hd_decap_12
XFILLER_14_398 vgnd vpwr scs8hd_decap_8
XPHY_93 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_60 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_247 vpwr vgnd scs8hd_fill_2
XPHY_71 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_82 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_20_335 vgnd vpwr scs8hd_decap_6
XFILLER_9_391 vgnd vpwr scs8hd_decap_12
XFILLER_1_280 vgnd vpwr scs8hd_decap_12
XFILLER_2_86 vgnd vpwr scs8hd_fill_1
XFILLER_11_379 vgnd vpwr scs8hd_decap_12
XFILLER_11_62 vgnd vpwr scs8hd_decap_12
XFILLER_11_51 vgnd vpwr scs8hd_decap_8
XFILLER_7_306 vgnd vpwr scs8hd_decap_12
XFILLER_6_361 vgnd vpwr scs8hd_decap_12
XFILLER_20_187 vgnd vpwr scs8hd_decap_12
XFILLER_19_232 vgnd vpwr scs8hd_decap_12
XFILLER_11_165 vgnd vpwr scs8hd_fill_1
XFILLER_11_121 vgnd vpwr scs8hd_fill_1
XFILLER_7_147 vgnd vpwr scs8hd_decap_12
XFILLER_7_103 vpwr vgnd scs8hd_fill_2
XFILLER_3_342 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ bottom_width_0_height_0__pin_0_ logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[0] vgnd vpwr scs8hd_ebufn_1
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _07_/X vgnd vpwr scs8hd_diode_2
XFILLER_16_202 vgnd vpwr scs8hd_decap_12
XFILLER_0_323 vgnd vpwr scs8hd_decap_12
XFILLER_4_117 vgnd vpwr scs8hd_decap_12
XFILLER_8_242 vgnd vpwr scs8hd_decap_8
XFILLER_5_86 vgnd vpwr scs8hd_decap_12
XFILLER_17_330 vgnd vpwr scs8hd_decap_12
XFILLER_5_245 vgnd vpwr scs8hd_decap_12
XFILLER_18_105 vgnd vpwr scs8hd_decap_12
XFILLER_14_300 vgnd vpwr scs8hd_decap_12
XPHY_50 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_61 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_215 vgnd vpwr scs8hd_decap_12
XPHY_72 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_83 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_94 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_171 vgnd vpwr scs8hd_decap_12
XFILLER_1_292 vgnd vpwr scs8hd_decap_12
XFILLER_2_32 vgnd vpwr scs8hd_decap_12
XFILLER_7_318 vgnd vpwr scs8hd_decap_12
XFILLER_19_403 vgnd vpwr scs8hd_decap_4
XFILLER_14_141 vgnd vpwr scs8hd_decap_12
XFILLER_11_74 vgnd vpwr scs8hd_decap_12
XFILLER_6_373 vgnd vpwr scs8hd_decap_12
XFILLER_20_199 vgnd vpwr scs8hd_decap_12
XFILLER_16_406 vgnd vpwr scs8hd_fill_1
XFILLER_7_159 vgnd vpwr scs8hd_decap_12
XFILLER_3_354 vgnd vpwr scs8hd_decap_12
XFILLER_17_62 vgnd vpwr scs8hd_decap_12
XFILLER_17_51 vgnd vpwr scs8hd_decap_8
XFILLER_0_335 vgnd vpwr scs8hd_decap_6
XFILLER_4_129 vgnd vpwr scs8hd_decap_12
XFILLER_3_195 vgnd vpwr scs8hd_decap_12
XFILLER_12_272 vgnd vpwr scs8hd_decap_3
XFILLER_8_276 vgnd vpwr scs8hd_decap_12
XFILLER_8_254 vgnd vpwr scs8hd_decap_12
XFILLER_8_232 vgnd vpwr scs8hd_fill_1
XFILLER_0_187 vgnd vpwr scs8hd_decap_12
XFILLER_5_32 vgnd vpwr scs8hd_decap_12
XFILLER_5_98 vgnd vpwr scs8hd_decap_12
XFILLER_5_257 vgnd vpwr scs8hd_decap_12
XFILLER_17_342 vgnd vpwr scs8hd_decap_12
XFILLER_18_117 vgnd vpwr scs8hd_decap_12
XFILLER_2_227 vgnd vpwr scs8hd_decap_12
XPHY_40 vgnd vpwr scs8hd_decap_3
XFILLER_14_312 vgnd vpwr scs8hd_decap_12
XPHY_95 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_51 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_11 vgnd vpwr scs8hd_decap_8
XFILLER_2_44 vgnd vpwr scs8hd_decap_12
XPHY_62 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_73 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_84 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_20_304 vgnd vpwr scs8hd_decap_6
XFILLER_11_86 vgnd vpwr scs8hd_decap_4
XFILLER_20_156 vgnd vpwr scs8hd_decap_12
XFILLER_6_385 vgnd vpwr scs8hd_decap_12
XFILLER_11_123 vgnd vpwr scs8hd_decap_12
XFILLER_19_245 vgnd vpwr scs8hd_decap_12
XFILLER_8_32 vgnd vpwr scs8hd_decap_12
X_19_ gfpga_pad_GPIO_PAD[0] bottom_width_0_height_0__pin_1_ vgnd vpwr scs8hd_buf_2
XFILLER_17_74 vgnd vpwr scs8hd_decap_12
XFILLER_16_215 vgnd vpwr scs8hd_decap_12
XFILLER_15_281 vgnd vpwr scs8hd_decap_12
XFILLER_13_218 vgnd vpwr scs8hd_decap_12
XFILLER_12_240 vgnd vpwr scs8hd_decap_12
XFILLER_0_199 vgnd vpwr scs8hd_decap_12
XFILLER_10_3 vgnd vpwr scs8hd_decap_12
XFILLER_8_288 vgnd vpwr scs8hd_decap_12
XFILLER_8_266 vgnd vpwr scs8hd_decap_8
XFILLER_5_44 vgnd vpwr scs8hd_decap_12
XFILLER_5_269 vgnd vpwr scs8hd_decap_12
XFILLER_17_354 vgnd vpwr scs8hd_decap_12
XFILLER_2_239 vgnd vpwr scs8hd_decap_8
XPHY_41 vgnd vpwr scs8hd_decap_3
XFILLER_18_129 vgnd vpwr scs8hd_decap_12
XPHY_30 vgnd vpwr scs8hd_decap_3
XFILLER_14_324 vgnd vpwr scs8hd_decap_12
XPHY_96 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_52 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_2_56 vgnd vpwr scs8hd_decap_12
XFILLER_2_89 vgnd vpwr scs8hd_decap_3
XPHY_63 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_74 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_85 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_184 vgnd vpwr scs8hd_decap_12
XFILLER_14_154 vgnd vpwr scs8hd_decap_12
XFILLER_20_168 vgnd vpwr scs8hd_decap_12
XFILLER_11_168 vgnd vpwr scs8hd_decap_12
XFILLER_11_135 vgnd vpwr scs8hd_decap_12
XFILLER_11_113 vgnd vpwr scs8hd_decap_8
XFILLER_19_257 vgnd vpwr scs8hd_decap_12
XFILLER_10_190 vgnd vpwr scs8hd_decap_12
XFILLER_8_44 vgnd vpwr scs8hd_decap_12
XFILLER_3_367 vgnd vpwr scs8hd_decap_12
X_18_ gfpga_pad_GPIO_PAD[7] bottom_width_0_height_0__pin_15_ vgnd vpwr scs8hd_buf_2
XFILLER_17_86 vgnd vpwr scs8hd_decap_12
XFILLER_16_227 vgnd vpwr scs8hd_decap_12
XFILLER_15_293 vgnd vpwr scs8hd_decap_12
XFILLER_0_156 vgnd vpwr scs8hd_decap_4
XFILLER_12_252 vgnd vpwr scs8hd_decap_12
XFILLER_8_212 vpwr vgnd scs8hd_fill_2
XFILLER_5_56 vgnd vpwr scs8hd_decap_4
XFILLER_14_32 vgnd vpwr scs8hd_decap_12
XPHY_31 vgnd vpwr scs8hd_decap_3
XPHY_20 vgnd vpwr scs8hd_decap_3
XPHY_97 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_42 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_1_251 vpwr vgnd scs8hd_fill_2
XPHY_53 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_64 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_75 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_86 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_196 vgnd vpwr scs8hd_decap_12
XFILLER_13_391 vgnd vpwr scs8hd_decap_12
XFILLER_2_24 vgnd vpwr scs8hd_decap_6
XFILLER_2_68 vgnd vpwr scs8hd_decap_12
XFILLER_11_306 vgnd vpwr scs8hd_decap_12
XFILLER_14_166 vgnd vpwr scs8hd_decap_12
XFILLER_10_361 vgnd vpwr scs8hd_decap_12
XFILLER_6_398 vgnd vpwr scs8hd_decap_8
XFILLER_20_125 vgnd vpwr scs8hd_decap_12
XFILLER_19_269 vgnd vpwr scs8hd_decap_12
XFILLER_11_147 vgnd vpwr scs8hd_decap_12
XFILLER_8_56 vgnd vpwr scs8hd_decap_12
XFILLER_7_107 vgnd vpwr scs8hd_decap_12
XFILLER_3_379 vgnd vpwr scs8hd_decap_12
X_17_ gfpga_pad_GPIO_PAD[6] bottom_width_0_height_0__pin_13_ vgnd vpwr scs8hd_buf_2
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_17_98 vgnd vpwr scs8hd_decap_12
XFILLER_16_239 vgnd vpwr scs8hd_decap_12
XFILLER_3_110 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _09_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_0_102 vgnd vpwr scs8hd_decap_8
XFILLER_12_264 vgnd vpwr scs8hd_decap_8
XFILLER_8_224 vgnd vpwr scs8hd_decap_8
XFILLER_17_367 vgnd vpwr scs8hd_decap_12
XFILLER_14_44 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ bottom_width_0_height_0__pin_2_ logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[1] vgnd vpwr scs8hd_ebufn_1
XPHY_32 vgnd vpwr scs8hd_decap_3
XFILLER_14_337 vgnd vpwr scs8hd_decap_12
XPHY_21 vgnd vpwr scs8hd_decap_3
XPHY_98 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_43 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_54 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_65 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_76 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_10 vgnd vpwr scs8hd_decap_3
XPHY_87 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_330 vgnd vpwr scs8hd_decap_12
XFILLER_1_230 vgnd vpwr scs8hd_decap_12
XFILLER_11_318 vgnd vpwr scs8hd_decap_12
XFILLER_2_7 vpwr vgnd scs8hd_fill_2
XFILLER_14_178 vgnd vpwr scs8hd_decap_12
XFILLER_10_373 vgnd vpwr scs8hd_decap_12
XFILLER_6_300 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _14_/Y vgnd vpwr scs8hd_diode_2
XFILLER_20_137 vgnd vpwr scs8hd_decap_12
XFILLER_9_171 vgnd vpwr scs8hd_decap_12
XFILLER_11_159 vgnd vpwr scs8hd_decap_6
XFILLER_7_119 vgnd vpwr scs8hd_decap_3
XANTENNA_logical_tile_io_mode_io__6.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ bottom_width_0_height_0__pin_12_ vgnd vpwr scs8hd_diode_2
XFILLER_8_68 vgnd vpwr scs8hd_decap_12
XFILLER_6_141 vgnd vpwr scs8hd_decap_12
X_16_ gfpga_pad_GPIO_PAD[5] bottom_width_0_height_0__pin_11_ vgnd vpwr scs8hd_buf_2
XFILLER_8_406 vgnd vpwr scs8hd_fill_1
XFILLER_12_276 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_0_125 vgnd vpwr scs8hd_decap_12
XFILLER_0_114 vpwr vgnd scs8hd_fill_2
XFILLER_14_56 vgnd vpwr scs8hd_decap_12
XFILLER_17_379 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ bottom_width_0_height_0__pin_8_ vgnd vpwr scs8hd_diode_2
Xlogical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _15_/Y vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_4_272 vgnd vpwr scs8hd_decap_3
XPHY_33 vgnd vpwr scs8hd_decap_3
XFILLER_14_349 vgnd vpwr scs8hd_decap_12
XPHY_22 vgnd vpwr scs8hd_decap_3
XPHY_99 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_88 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_44 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_55 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_66 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_77 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vpwr scs8hd_decap_3
XFILLER_17_110 vgnd vpwr scs8hd_decap_12
XFILLER_9_342 vgnd vpwr scs8hd_decap_12
XFILLER_1_242 vpwr vgnd scs8hd_fill_2
XFILLER_1_220 vpwr vgnd scs8hd_fill_2
XFILLER_10_385 vgnd vpwr scs8hd_decap_12
XFILLER_6_312 vgnd vpwr scs8hd_decap_12
XFILLER_20_149 vgnd vpwr scs8hd_decap_6
XANTENNA__11__A enable vgnd vpwr scs8hd_diode_2
XFILLER_19_3 vgnd vpwr scs8hd_decap_12
X_15_ address[1] _11_/Y _04_/X address[2] _15_/Y vgnd vpwr scs8hd_nor4_4
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ bottom_width_0_height_0__pin_4_ vgnd vpwr scs8hd_diode_2
XANTENNA__06__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_3_123 vgnd vpwr scs8hd_decap_12
XFILLER_12_288 vgnd vpwr scs8hd_decap_12
XFILLER_12_211 vgnd vpwr scs8hd_decap_3
XFILLER_8_204 vgnd vpwr scs8hd_decap_8
XFILLER_0_137 vgnd vpwr scs8hd_decap_12
XFILLER_5_15 vgnd vpwr scs8hd_decap_4
XFILLER_14_68 vgnd vpwr scs8hd_decap_12
XFILLER_4_251 vgnd vpwr scs8hd_decap_8
XANTENNA_logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XPHY_12 vgnd vpwr scs8hd_decap_3
XFILLER_6_80 vgnd vpwr scs8hd_decap_12
XPHY_34 vgnd vpwr scs8hd_decap_3
XANTENNA__14__A _06_/Y vgnd vpwr scs8hd_diode_2
XPHY_23 vgnd vpwr scs8hd_decap_3
XPHY_89 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_56 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_45 vgnd vpwr scs8hd_tapvpwrvgnd_1
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_A
+ bottom_width_0_height_0__pin_0_ vgnd vpwr scs8hd_diode_2
XPHY_67 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_78 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_9_354 vgnd vpwr scs8hd_decap_12
XFILLER_6_324 vgnd vpwr scs8hd_decap_12
XANTENNA__09__A address[1] vgnd vpwr scs8hd_diode_2
XFILLER_20_106 vgnd vpwr scs8hd_decap_12
XFILLER_9_184 vgnd vpwr scs8hd_decap_12
XFILLER_8_15 vgnd vpwr scs8hd_decap_12
XFILLER_6_154 vgnd vpwr scs8hd_decap_12
X_14_ _06_/Y _11_/Y _04_/X address[2] _14_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_0_308 vpwr vgnd scs8hd_fill_2
XFILLER_15_220 vgnd vpwr scs8hd_decap_12
XANTENNA__22__A gfpga_pad_GPIO_PAD[3] vgnd vpwr scs8hd_diode_2
XFILLER_3_135 vgnd vpwr scs8hd_decap_12
XFILLER_3_179 vpwr vgnd scs8hd_fill_2
XFILLER_0_71 vgnd vpwr scs8hd_decap_12
XFILLER_9_80 vgnd vpwr scs8hd_fill_1
XFILLER_0_149 vgnd vpwr scs8hd_decap_4
XANTENNA__17__A gfpga_pad_GPIO_PAD[6] vgnd vpwr scs8hd_diode_2
XFILLER_5_208 vgnd vpwr scs8hd_decap_12
XFILLER_1_403 vgnd vpwr scs8hd_decap_4
XPHY_35 vgnd vpwr scs8hd_decap_3
XPHY_24 vgnd vpwr scs8hd_decap_3
XANTENNA__14__B _11_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_3 vgnd vpwr scs8hd_decap_12
XPHY_13 vgnd vpwr scs8hd_decap_3
XPHY_57 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_46 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_1_255 vgnd vpwr scs8hd_decap_3
XPHY_68 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_79 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_123 vgnd vpwr scs8hd_decap_12
XFILLER_11_59 vpwr vgnd scs8hd_fill_2
XFILLER_11_15 vgnd vpwr scs8hd_decap_12
XANTENNA__09__B enable vgnd vpwr scs8hd_diode_2
XFILLER_20_118 vgnd vpwr scs8hd_decap_6
XFILLER_10_398 vgnd vpwr scs8hd_decap_8
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer_TEB
+ logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ vgnd vpwr scs8hd_diode_2
XFILLER_3_60 vgnd vpwr scs8hd_fill_1
XFILLER_3_82 vgnd vpwr scs8hd_decap_3
XFILLER_5_391 vgnd vpwr scs8hd_decap_12
XFILLER_12_80 vgnd vpwr scs8hd_decap_12
XFILLER_10_151 vpwr vgnd scs8hd_fill_2
XFILLER_8_27 vgnd vpwr scs8hd_decap_4
XFILLER_6_166 vgnd vpwr scs8hd_decap_12
XFILLER_3_306 vgnd vpwr scs8hd_decap_12
XFILLER_18_251 vgnd vpwr scs8hd_decap_12
X_13_ address[1] _11_/Y _04_/X _08_/Y _13_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_2_361 vgnd vpwr scs8hd_decap_12
XFILLER_3_147 vgnd vpwr scs8hd_decap_12
XFILLER_15_232 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__5.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _09_/X vgnd vpwr scs8hd_diode_2
XFILLER_0_83 vgnd vpwr scs8hd_decap_4
XFILLER_14_15 vgnd vpwr scs8hd_decap_12
XFILLER_7_261 vgnd vpwr scs8hd_decap_12
XFILLER_6_93 vgnd vpwr scs8hd_decap_12
XFILLER_4_264 vgnd vpwr scs8hd_decap_8
XPHY_36 vgnd vpwr scs8hd_decap_3
XPHY_25 vgnd vpwr scs8hd_decap_3
XANTENNA__14__C _04_/X vgnd vpwr scs8hd_diode_2
XPHY_58 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_1_245 vgnd vpwr scs8hd_decap_4
XPHY_47 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_69 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_14 vgnd vpwr scs8hd_decap_3
XFILLER_17_135 vgnd vpwr scs8hd_decap_12
XFILLER_13_330 vgnd vpwr scs8hd_decap_12
XFILLER_9_367 vgnd vpwr scs8hd_decap_12
XFILLER_16_190 vgnd vpwr scs8hd_decap_12
XFILLER_11_27 vgnd vpwr scs8hd_decap_12
XANTENNA__09__C address[3] vgnd vpwr scs8hd_diode_2
XFILLER_14_105 vgnd vpwr scs8hd_decap_12
XFILLER_10_300 vgnd vpwr scs8hd_decap_12
XFILLER_6_337 vgnd vpwr scs8hd_decap_12
XFILLER_13_171 vgnd vpwr scs8hd_decap_12
XFILLER_9_120 vpwr vgnd scs8hd_fill_2
XFILLER_3_50 vpwr vgnd scs8hd_fill_2
XFILLER_19_208 vgnd vpwr scs8hd_decap_12
XFILLER_15_403 vgnd vpwr scs8hd_decap_4
XFILLER_3_318 vgnd vpwr scs8hd_decap_12
XFILLER_18_263 vgnd vpwr scs8hd_decap_12
X_12_ _06_/Y _11_/Y _04_/X _08_/Y _12_/Y vgnd vpwr scs8hd_nor4_4
XFILLER_6_178 vgnd vpwr scs8hd_decap_12
Xlogical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ bottom_width_0_height_0__pin_4_ logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[2] vgnd vpwr scs8hd_ebufn_1
XFILLER_2_373 vgnd vpwr scs8hd_decap_12
XFILLER_17_59 vpwr vgnd scs8hd_fill_2
XFILLER_17_15 vgnd vpwr scs8hd_decap_12
XFILLER_12_406 vgnd vpwr scs8hd_fill_1
XFILLER_3_159 vgnd vpwr scs8hd_decap_12
XFILLER_17_3 vgnd vpwr scs8hd_decap_12
XFILLER_0_118 vgnd vpwr scs8hd_decap_6
XFILLER_0_51 vgnd vpwr scs8hd_decap_8
XFILLER_20_280 vgnd vpwr scs8hd_decap_12
XFILLER_18_80 vgnd vpwr scs8hd_decap_12
XFILLER_19_391 vgnd vpwr scs8hd_decap_12
XFILLER_7_273 vgnd vpwr scs8hd_decap_12
XFILLER_17_306 vgnd vpwr scs8hd_decap_12
XFILLER_14_27 vgnd vpwr scs8hd_decap_4
XFILLER_16_361 vgnd vpwr scs8hd_decap_12
XFILLER_4_276 vgnd vpwr scs8hd_decap_12
XPHY_37 vgnd vpwr scs8hd_decap_3
XPHY_26 vgnd vpwr scs8hd_decap_3
XANTENNA__14__D address[2] vgnd vpwr scs8hd_diode_2
XPHY_15 vgnd vpwr scs8hd_decap_3
XPHY_48 vgnd vpwr scs8hd_tapvpwrvgnd_1
XPHY_59 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_147 vgnd vpwr scs8hd_decap_12
XFILLER_13_342 vgnd vpwr scs8hd_decap_12
XFILLER_9_379 vgnd vpwr scs8hd_decap_12
XFILLER_1_268 vgnd vpwr scs8hd_decap_12
XFILLER_2_19 vgnd vpwr scs8hd_decap_3
XFILLER_11_39 vgnd vpwr scs8hd_decap_12
XFILLER_14_117 vgnd vpwr scs8hd_decap_12
XFILLER_10_312 vgnd vpwr scs8hd_decap_12
XFILLER_6_349 vgnd vpwr scs8hd_decap_12
XANTENNA__09__D _08_/Y vgnd vpwr scs8hd_diode_2
XFILLER_9_198 vpwr vgnd scs8hd_fill_2
XFILLER_3_62 vgnd vpwr scs8hd_decap_12
X_11_ enable _11_/Y vgnd vpwr scs8hd_inv_8
XFILLER_12_93 vgnd vpwr scs8hd_decap_3
XFILLER_10_131 vgnd vpwr scs8hd_decap_12
XFILLER_2_385 vgnd vpwr scs8hd_decap_12
XFILLER_17_27 vgnd vpwr scs8hd_decap_12
XFILLER_15_245 vgnd vpwr scs8hd_decap_12
XFILLER_9_83 vpwr vgnd scs8hd_fill_2
XFILLER_20_292 vgnd vpwr scs8hd_decap_12
XFILLER_12_215 vgnd vpwr scs8hd_decap_12
XFILLER_11_281 vgnd vpwr scs8hd_decap_12
XFILLER_7_285 vgnd vpwr scs8hd_decap_12
XFILLER_17_318 vgnd vpwr scs8hd_decap_12
XFILLER_16_373 vgnd vpwr scs8hd_decap_12
XFILLER_4_288 vgnd vpwr scs8hd_decap_12
XPHY_38 vgnd vpwr scs8hd_decap_3
XPHY_27 vgnd vpwr scs8hd_decap_3
XPHY_16 vgnd vpwr scs8hd_decap_3
XPHY_49 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_17_159 vgnd vpwr scs8hd_decap_12
XFILLER_13_354 vgnd vpwr scs8hd_decap_12
XFILLER_14_129 vgnd vpwr scs8hd_decap_12
XFILLER_10_324 vgnd vpwr scs8hd_decap_12
XFILLER_7_3 vgnd vpwr scs8hd_decap_12
XFILLER_13_184 vgnd vpwr scs8hd_decap_12
XFILLER_3_74 vgnd vpwr scs8hd_decap_8
XFILLER_18_276 vgnd vpwr scs8hd_decap_12
XFILLER_10_154 vgnd vpwr scs8hd_decap_12
XFILLER_10_143 vgnd vpwr scs8hd_decap_8
X_10_ _06_/Y enable address[3] _08_/Y _10_/X vgnd vpwr scs8hd_and4_4
XFILLER_17_39 vgnd vpwr scs8hd_decap_12
XFILLER_15_257 vgnd vpwr scs8hd_decap_12
XFILLER_9_62 vgnd vpwr scs8hd_decap_12
XFILLER_9_51 vgnd vpwr scs8hd_decap_8
XFILLER_12_227 vgnd vpwr scs8hd_decap_4
XFILLER_18_93 vgnd vpwr scs8hd_decap_12
XFILLER_11_293 vgnd vpwr scs8hd_decap_12
XFILLER_7_297 vgnd vpwr scs8hd_decap_8
XFILLER_7_231 vpwr vgnd scs8hd_fill_2
XFILLER_20_94 vgnd vpwr scs8hd_decap_12
XFILLER_16_385 vgnd vpwr scs8hd_decap_12
XPHY_28 vgnd vpwr scs8hd_decap_3
XPHY_17 vgnd vpwr scs8hd_decap_3
XPHY_39 vgnd vpwr scs8hd_decap_3
XFILLER_1_226 vpwr vgnd scs8hd_fill_2
Xlogical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch
+ data_in logical_tile_io_mode_io__4.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ _10_/X vgnd vpwr scs8hd_lpflow_inputisolatch_1
XFILLER_13_196 vgnd vpwr scs8hd_decap_8
XFILLER_9_123 vgnd vpwr scs8hd_decap_12
XFILLER_9_112 vpwr vgnd scs8hd_fill_2
XFILLER_10_166 vgnd vpwr scs8hd_decap_12
XFILLER_2_398 vgnd vpwr scs8hd_decap_8
XFILLER_18_288 vgnd vpwr scs8hd_decap_12
XFILLER_15_269 vgnd vpwr scs8hd_decap_12
XFILLER_0_32 vgnd vpwr scs8hd_decap_4
XFILLER_9_74 vgnd vpwr scs8hd_decap_6
XFILLER_20_261 vgnd vpwr scs8hd_decap_12
XFILLER_7_243 vgnd vpwr scs8hd_fill_1
XFILLER_7_221 vpwr vgnd scs8hd_fill_2
XFILLER_15_3 vgnd vpwr scs8hd_decap_12
XFILLER_4_202 vgnd vpwr scs8hd_decap_12
XPHY_29 vgnd vpwr scs8hd_decap_3
XPHY_18 vgnd vpwr scs8hd_decap_3
XFILLER_15_62 vgnd vpwr scs8hd_decap_12
XFILLER_15_51 vgnd vpwr scs8hd_decap_8
XFILLER_13_367 vgnd vpwr scs8hd_decap_12
XFILLER_0_271 vpwr vgnd scs8hd_fill_2
XFILLER_10_337 vgnd vpwr scs8hd_decap_12
XFILLER_9_135 vgnd vpwr scs8hd_decap_12
XFILLER_8_190 vgnd vpwr scs8hd_decap_12
XFILLER_3_54 vgnd vpwr scs8hd_decap_6
XFILLER_3_98 vgnd vpwr scs8hd_decap_12
XFILLER_5_330 vgnd vpwr scs8hd_decap_12
XFILLER_10_178 vgnd vpwr scs8hd_decap_12
XFILLER_6_105 vgnd vpwr scs8hd_decap_12
XANTENNA_logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.GPIO_LATCH_mem.LATCH_0_.latch_SLEEPB
+ _15_/Y vgnd vpwr scs8hd_diode_2
XFILLER_2_300 vgnd vpwr scs8hd_decap_12
XFILLER_5_171 vgnd vpwr scs8hd_decap_12
XFILLER_7_403 vgnd vpwr scs8hd_decap_4
XFILLER_0_11 vpwr vgnd scs8hd_fill_2
XFILLER_2_141 vgnd vpwr scs8hd_decap_12
XFILLER_20_273 vgnd vpwr scs8hd_decap_6
XFILLER_4_406 vgnd vpwr scs8hd_fill_1
XFILLER_20_63 vgnd vpwr scs8hd_decap_12
XFILLER_16_398 vgnd vpwr scs8hd_decap_8
Xlogical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer
+ bottom_width_0_height_0__pin_6_ logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.GPIO_0_.buffer/TEB
+ gfpga_pad_GPIO_PAD[3] vgnd vpwr scs8hd_ebufn_1
XFILLER_6_32 vgnd vpwr scs8hd_decap_12
XPHY_19 vgnd vpwr scs8hd_decap_3
XFILLER_15_74 vgnd vpwr scs8hd_decap_12
XFILLER_13_379 vgnd vpwr scs8hd_decap_12
XFILLER_9_306 vgnd vpwr scs8hd_decap_12
XPHY_190 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_8_361 vgnd vpwr scs8hd_decap_12
XFILLER_10_349 vgnd vpwr scs8hd_decap_12
XFILLER_13_110 vgnd vpwr scs8hd_decap_12
XFILLER_9_147 vgnd vpwr scs8hd_decap_12
XFILLER_3_33 vgnd vpwr scs8hd_decap_12
XFILLER_5_342 vgnd vpwr scs8hd_decap_12
XFILLER_6_117 vgnd vpwr scs8hd_decap_12
XFILLER_18_202 vgnd vpwr scs8hd_decap_12
XFILLER_2_312 vgnd vpwr scs8hd_decap_12
XFILLER_5_3 vgnd vpwr scs8hd_decap_12
XFILLER_2_186 vgnd vpwr scs8hd_decap_12
XFILLER_9_87 vpwr vgnd scs8hd_fill_2
XFILLER_0_89 vpwr vgnd scs8hd_fill_2
XFILLER_0_67 vpwr vgnd scs8hd_fill_2
XFILLER_0_23 vpwr vgnd scs8hd_fill_2
XFILLER_20_230 vgnd vpwr scs8hd_decap_12
XFILLER_19_330 vgnd vpwr scs8hd_decap_12
XFILLER_7_245 vgnd vpwr scs8hd_decap_4
XFILLER_20_75 vgnd vpwr scs8hd_decap_12
XFILLER_16_300 vgnd vpwr scs8hd_decap_12
XFILLER_4_215 vgnd vpwr scs8hd_decap_12
XFILLER_4_259 vgnd vpwr scs8hd_decap_3
XFILLER_19_171 vgnd vpwr scs8hd_decap_12
XFILLER_20_3 vgnd vpwr scs8hd_decap_12
XFILLER_6_44 vgnd vpwr scs8hd_decap_12
XFILLER_15_86 vgnd vpwr scs8hd_decap_12
XFILLER_9_318 vgnd vpwr scs8hd_decap_12
XPHY_180 vgnd vpwr scs8hd_tapvpwrvgnd_1
XFILLER_16_141 vgnd vpwr scs8hd_decap_12
XFILLER_8_373 vgnd vpwr scs8hd_decap_12
XFILLER_0_284 vpwr vgnd scs8hd_fill_2
.ends

